

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6545, n6547, n6548, n6549, n6550, n6551, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15310;

  AND2_X1 U7293 ( .A1(n7102), .A2(n9103), .ZN(n13015) );
  OR2_X1 U7294 ( .A1(n12253), .A2(n12261), .ZN(n11566) );
  OR2_X1 U7295 ( .A1(n11557), .A2(n11556), .ZN(n12275) );
  NAND2_X2 U7296 ( .A1(n8095), .A2(n8094), .ZN(n13144) );
  XNOR2_X1 U7297 ( .A(n7977), .B(SI_20_), .ZN(n7976) );
  BUF_X1 U7298 ( .A(n10895), .Z(n6569) );
  INV_X1 U7299 ( .A(n11882), .ZN(n11930) );
  CLKBUF_X2 U7302 ( .A(n6620), .Z(n6825) );
  CLKBUF_X2 U7303 ( .A(n11940), .Z(n6565) );
  INV_X2 U7304 ( .A(n12673), .ZN(n12663) );
  INV_X1 U7305 ( .A(n9124), .ZN(n14748) );
  NAND2_X1 U7307 ( .A1(n6549), .A2(n7712), .ZN(n9765) );
  OAI211_X1 U7308 ( .C1(n8529), .C2(n9264), .A(n8292), .B(n6614), .ZN(n10298)
         );
  CLKBUF_X2 U7309 ( .A(n8288), .Z(n8529) );
  CLKBUF_X2 U7310 ( .A(n9653), .Z(n10364) );
  CLKBUF_X2 U7311 ( .A(n7691), .Z(n6563) );
  INV_X2 U7312 ( .A(n10252), .ZN(n13448) );
  XNOR2_X1 U7313 ( .A(n8250), .B(n8249), .ZN(n8746) );
  INV_X2 U7314 ( .A(n9251), .ZN(n9020) );
  INV_X1 U7315 ( .A(n8276), .ZN(n9251) );
  AND3_X2 U7316 ( .A1(n6612), .A2(n7471), .A3(n9200), .ZN(n9217) );
  AND3_X1 U7317 ( .A1(n9143), .A2(n9196), .A3(n9144), .ZN(n6612) );
  CLKBUF_X1 U7318 ( .A(n12088), .Z(n6545) );
  OAI21_X1 U7319 ( .B1(n9984), .B2(n9983), .A(n14934), .ZN(n12088) );
  INV_X1 U7321 ( .A(n15310), .ZN(n6547) );
  OAI22_X1 U7322 ( .A1(n8947), .A2(n7498), .B1(n8948), .B2(n7499), .ZN(n8953)
         );
  NAND2_X1 U7323 ( .A1(n12277), .A2(n12260), .ZN(n11423) );
  AND2_X2 U7324 ( .A1(n9653), .A2(n9652), .ZN(n11821) );
  NOR2_X1 U7325 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9147) );
  OR2_X1 U7326 ( .A1(n8639), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7327 ( .A1(n8613), .A2(n8612), .ZN(n12333) );
  NAND2_X1 U7328 ( .A1(n8746), .A2(n12610), .ZN(n9579) );
  AND2_X2 U7329 ( .A1(n14808), .A2(n9409), .ZN(n12673) );
  OR2_X1 U7330 ( .A1(n9953), .A2(n10060), .ZN(n10057) );
  OR2_X1 U7331 ( .A1(n13039), .A2(n7103), .ZN(n7102) );
  INV_X2 U7332 ( .A(n11884), .ZN(n11931) );
  INV_X1 U7333 ( .A(n10244), .ZN(n10252) );
  INV_X2 U7334 ( .A(n11063), .ZN(n13455) );
  INV_X1 U7335 ( .A(n12309), .ZN(n12054) );
  INV_X1 U7337 ( .A(n8682), .ZN(n8311) );
  INV_X1 U7338 ( .A(n7690), .ZN(n9029) );
  OAI21_X1 U7339 ( .B1(n12991), .B2(n12826), .A(n12983), .ZN(n8210) );
  AND2_X1 U7340 ( .A1(n6941), .A2(n6939), .ZN(n13029) );
  AND2_X1 U7341 ( .A1(n7141), .A2(n7142), .ZN(n13087) );
  NAND2_X1 U7342 ( .A1(n12860), .A2(n7678), .ZN(n7725) );
  NAND2_X1 U7343 ( .A1(n10798), .A2(n7488), .ZN(n7487) );
  AND2_X1 U7344 ( .A1(n10388), .A2(n10524), .ZN(n14554) );
  CLKBUF_X3 U7345 ( .A(n14557), .Z(n6570) );
  NAND2_X2 U7347 ( .A1(n7953), .A2(n7952), .ZN(n13078) );
  OAI21_X1 U7348 ( .B1(n13070), .B2(n8205), .A(n8206), .ZN(n13059) );
  AND2_X1 U7349 ( .A1(n8846), .A2(n12710), .ZN(n13146) );
  AOI21_X1 U7350 ( .B1(n11777), .B2(n14571), .A(n11776), .ZN(n14032) );
  NAND2_X1 U7351 ( .A1(n14134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9397) );
  AND2_X1 U7352 ( .A1(n9440), .A2(n9439), .ZN(n13952) );
  AND4_X1 U7353 ( .A1(n9150), .A2(n10094), .A3(n9149), .A4(n9148), .ZN(n6548)
         );
  AND2_X1 U7354 ( .A1(n7713), .A2(n6619), .ZN(n6549) );
  OR2_X1 U7355 ( .A1(n6945), .A2(n7314), .ZN(n6550) );
  NAND2_X2 U7356 ( .A1(n8199), .A2(n8198), .ZN(n11357) );
  NAND2_X2 U7358 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  INV_X1 U7359 ( .A(n11063), .ZN(n6551) );
  NAND2_X1 U7360 ( .A1(n11671), .A2(n9020), .ZN(n11063) );
  NOR2_X2 U7361 ( .A1(n8751), .A2(n10100), .ZN(n14930) );
  OAI21_X2 U7362 ( .B1(n14684), .B2(n14681), .A(n14680), .ZN(n12613) );
  NAND2_X2 U7363 ( .A1(n11115), .A2(n11114), .ZN(n14684) );
  CLKBUF_X2 U7365 ( .A(n8281), .Z(n6553) );
  NAND4_X1 U7366 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8281)
         );
  NAND2_X2 U7367 ( .A1(n7467), .A2(n7465), .ZN(n13306) );
  NAND2_X1 U7368 ( .A1(n11821), .A2(n6570), .ZN(n9656) );
  INV_X1 U7369 ( .A(n9656), .ZN(n11940) );
  NAND2_X2 U7370 ( .A1(n6966), .A2(n6967), .ZN(n7590) );
  NAND2_X2 U7372 ( .A1(n6594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9224) );
  NAND2_X2 U7373 ( .A1(n8603), .A2(n8602), .ZN(n8615) );
  INV_X1 U7374 ( .A(n14596), .ZN(n10348) );
  NAND2_X2 U7375 ( .A1(n8140), .A2(n8131), .ZN(n9173) );
  AND2_X2 U7376 ( .A1(n8240), .A2(n8239), .ZN(n8312) );
  BUF_X4 U7377 ( .A(n8312), .Z(n8710) );
  NAND2_X2 U7378 ( .A1(n11737), .A2(n11736), .ZN(n14045) );
  XNOR2_X2 U7379 ( .A(n8246), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U7380 ( .A1(n6759), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8246) );
  INV_X2 U7381 ( .A(n12673), .ZN(n6554) );
  NAND2_X1 U7382 ( .A1(n7574), .A2(n13259), .ZN(n8135) );
  XNOR2_X2 U7383 ( .A(n7566), .B(n7562), .ZN(n13259) );
  XNOR2_X2 U7384 ( .A(n13937), .B(n13582), .ZN(n13930) );
  AND2_X2 U7385 ( .A1(n9142), .A2(n9141), .ZN(n7471) );
  OAI21_X2 U7386 ( .B1(n12321), .B2(n8645), .A(n8646), .ZN(n12308) );
  XNOR2_X1 U7387 ( .A(n8346), .B(P3_IR_REG_6__SCAN_IN), .ZN(n9926) );
  NOR3_X2 U7388 ( .A1(n9123), .A2(n9122), .A3(n9121), .ZN(n9125) );
  AOI22_X2 U7389 ( .A1(n13007), .A2(n13006), .B1(n12724), .B2(n13168), .ZN(
        n12997) );
  NAND2_X1 U7390 ( .A1(n8746), .A2(n12610), .ZN(n6556) );
  NAND2_X1 U7391 ( .A1(n8746), .A2(n12610), .ZN(n6557) );
  XNOR2_X2 U7392 ( .A(n8589), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12222) );
  NAND2_X2 U7393 ( .A1(n7487), .A2(n7486), .ZN(n11333) );
  XNOR2_X2 U7394 ( .A(n12655), .B(n12654), .ZN(n12775) );
  NAND2_X2 U7395 ( .A1(n12714), .A2(n7319), .ZN(n12655) );
  AOI21_X2 U7396 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(n14229), .A(n14498), .ZN(
        n14232) );
  XNOR2_X1 U7397 ( .A(n8251), .B(n8237), .ZN(n12610) );
  NAND2_X2 U7398 ( .A1(n13301), .A2(n11868), .ZN(n13359) );
  OAI21_X2 U7399 ( .B1(n12333), .B2(n8629), .A(n8630), .ZN(n12321) );
  XNOR2_X2 U7400 ( .A(n13078), .B(n12788), .ZN(n13071) );
  XNOR2_X2 U7401 ( .A(n9397), .B(n9396), .ZN(n11808) );
  OR2_X2 U7403 ( .A1(n12138), .A2(n10298), .ZN(n11446) );
  XNOR2_X2 U7404 ( .A(n9398), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9399) );
  XNOR2_X2 U7405 ( .A(n6727), .B(n6714), .ZN(n11726) );
  OR2_X2 U7406 ( .A1(n8459), .A2(n8458), .ZN(n8468) );
  OAI21_X2 U7407 ( .B1(n8455), .B2(n8454), .A(n8456), .ZN(n8459) );
  NAND2_X2 U7408 ( .A1(n8725), .A2(n8724), .ZN(n12253) );
  NOR2_X2 U7409 ( .A1(n14200), .A2(n15303), .ZN(n14250) );
  NAND2_X1 U7410 ( .A1(n8817), .A2(n8816), .ZN(n11959) );
  NAND2_X1 U7411 ( .A1(n13376), .A2(n13377), .ZN(n13375) );
  NAND2_X1 U7412 ( .A1(n12492), .A2(n12054), .ZN(n11553) );
  NAND2_X1 U7413 ( .A1(n12684), .A2(n7534), .ZN(n12757) );
  OR2_X1 U7414 ( .A1(n14241), .A2(n14240), .ZN(n14516) );
  INV_X1 U7415 ( .A(n13871), .ZN(n7166) );
  NAND2_X1 U7416 ( .A1(n11756), .A2(n11755), .ZN(n14040) );
  NAND2_X1 U7417 ( .A1(n6910), .A2(n6909), .ZN(n13084) );
  OR2_X1 U7418 ( .A1(n13101), .A2(n7938), .ZN(n6910) );
  OR2_X1 U7419 ( .A1(n14394), .A2(n8197), .ZN(n8199) );
  AOI21_X1 U7420 ( .B1(n6949), .B2(n6571), .A(n6588), .ZN(n6948) );
  XNOR2_X1 U7421 ( .A(n8018), .B(SI_22_), .ZN(n11669) );
  NAND2_X1 U7422 ( .A1(n10545), .A2(n10544), .ZN(n10543) );
  NAND2_X1 U7423 ( .A1(n10831), .A2(n10830), .ZN(n10829) );
  OR2_X1 U7424 ( .A1(n8901), .A2(n7503), .ZN(n7502) );
  AOI21_X1 U7425 ( .B1(n8187), .B2(n6638), .A(n6582), .ZN(n10027) );
  NAND2_X1 U7426 ( .A1(n15292), .A2(n14208), .ZN(n14210) );
  INV_X2 U7427 ( .A(n14736), .ZN(n6558) );
  NAND2_X1 U7428 ( .A1(n11450), .A2(n11449), .ZN(n11590) );
  INV_X1 U7429 ( .A(n8876), .ZN(n9726) );
  NAND2_X1 U7430 ( .A1(n12849), .A2(n12664), .ZN(n9689) );
  INV_X1 U7431 ( .A(n11032), .ZN(n11968) );
  NAND3_X2 U7432 ( .A1(n6597), .A2(n7683), .A3(n7685), .ZN(n8178) );
  INV_X1 U7433 ( .A(n11884), .ZN(n6559) );
  CLKBUF_X1 U7434 ( .A(n7679), .Z(n9030) );
  NAND2_X1 U7435 ( .A1(n7967), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7692) );
  OR2_X1 U7436 ( .A1(n7691), .A2(n12851), .ZN(n7682) );
  INV_X4 U7437 ( .A(n8673), .ZN(n8711) );
  INV_X1 U7438 ( .A(n13693), .ZN(n10271) );
  OR2_X1 U7439 ( .A1(n10236), .A2(n10442), .ZN(n13467) );
  INV_X1 U7440 ( .A(n13473), .ZN(n10237) );
  INV_X4 U7441 ( .A(n11569), .ZN(n11577) );
  CLKBUF_X2 U7442 ( .A(n7691), .Z(n6564) );
  CLKBUF_X1 U7443 ( .A(n9072), .Z(n6566) );
  NAND2_X2 U7444 ( .A1(n13449), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9466) );
  INV_X1 U7445 ( .A(n8898), .ZN(n8902) );
  INV_X2 U7446 ( .A(n11671), .ZN(n11702) );
  AND2_X1 U7448 ( .A1(n12489), .A2(n12488), .ZN(n12555) );
  OR2_X1 U7449 ( .A1(n11957), .A2(n14973), .ZN(n8831) );
  NAND2_X1 U7450 ( .A1(n12258), .A2(n7442), .ZN(n8812) );
  OAI21_X1 U7451 ( .B1(n6834), .B2(n14939), .A(n6832), .ZN(n12482) );
  NOR2_X1 U7452 ( .A1(n6581), .A2(n14939), .ZN(n6822) );
  AOI21_X1 U7453 ( .B1(n7184), .B2(n7182), .A(n6681), .ZN(n6987) );
  NAND2_X1 U7454 ( .A1(n7422), .A2(n6603), .ZN(n7421) );
  AND2_X1 U7455 ( .A1(n8855), .A2(n8854), .ZN(n7541) );
  NAND2_X1 U7456 ( .A1(n11396), .A2(n11395), .ZN(n11408) );
  OR2_X1 U7457 ( .A1(n13147), .A2(n13114), .ZN(n8855) );
  AOI211_X1 U7458 ( .C1(n13148), .C2(n14731), .A(n12981), .B(n12980), .ZN(
        n12982) );
  NOR2_X1 U7459 ( .A1(n13874), .A2(n11802), .ZN(n13858) );
  NAND2_X1 U7460 ( .A1(n7095), .A2(n7099), .ZN(n12995) );
  AOI21_X1 U7461 ( .B1(n12979), .B2(n14753), .A(n12978), .ZN(n13151) );
  OR2_X1 U7462 ( .A1(n12486), .A2(n12274), .ZN(n11424) );
  OR2_X1 U7463 ( .A1(n13039), .A2(n7100), .ZN(n7095) );
  AOI21_X1 U7464 ( .B1(n13838), .B2(n14571), .A(n13837), .ZN(n14038) );
  OAI21_X1 U7465 ( .B1(n14300), .B2(n14301), .A(n6829), .ZN(n6828) );
  OR2_X1 U7466 ( .A1(n13891), .A2(n13890), .ZN(n13889) );
  NAND2_X1 U7467 ( .A1(n8666), .A2(n8665), .ZN(n12492) );
  AOI21_X1 U7468 ( .B1(n7358), .B2(n7356), .A(n7364), .ZN(n7355) );
  INV_X1 U7469 ( .A(n7358), .ZN(n7357) );
  NAND2_X1 U7470 ( .A1(n13879), .A2(n13890), .ZN(n13878) );
  NAND2_X1 U7471 ( .A1(n14294), .A2(n14292), .ZN(n14300) );
  NAND2_X1 U7472 ( .A1(n6739), .A2(n6738), .ZN(n14294) );
  NAND2_X1 U7473 ( .A1(n12081), .A2(n7174), .ZN(n12043) );
  INV_X1 U7474 ( .A(n14246), .ZN(n6739) );
  NAND2_X1 U7475 ( .A1(n7161), .A2(n7160), .ZN(n13896) );
  NOR2_X2 U7476 ( .A1(n14040), .A2(n13866), .ZN(n13851) );
  NAND2_X1 U7477 ( .A1(n6852), .A2(n6851), .ZN(n12187) );
  INV_X1 U7478 ( .A(n7163), .ZN(n7162) );
  NAND2_X1 U7479 ( .A1(n8522), .A2(n8521), .ZN(n12395) );
  XNOR2_X1 U7480 ( .A(n9017), .B(n9016), .ZN(n13258) );
  XNOR2_X1 U7481 ( .A(n12509), .B(n12360), .ZN(n12351) );
  NAND2_X1 U7482 ( .A1(n12401), .A2(n12400), .ZN(n12399) );
  XNOR2_X1 U7483 ( .A(n11670), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14150) );
  OAI21_X1 U7484 ( .B1(n11669), .B2(n8020), .A(n8001), .ZN(n6727) );
  INV_X1 U7485 ( .A(n14245), .ZN(n6738) );
  NAND2_X1 U7486 ( .A1(n8018), .A2(SI_22_), .ZN(n8001) );
  NAND2_X1 U7487 ( .A1(n11143), .A2(n8423), .ZN(n11315) );
  OAI21_X1 U7488 ( .B1(n8040), .B2(n8039), .A(n8038), .ZN(n8047) );
  NAND2_X1 U7489 ( .A1(n11145), .A2(n11144), .ZN(n11143) );
  OAI211_X1 U7490 ( .C1(n6574), .C2(n7978), .A(n6960), .B(n7266), .ZN(n8037)
         );
  NAND2_X1 U7491 ( .A1(n7090), .A2(n7089), .ZN(n11296) );
  OR2_X1 U7492 ( .A1(n10668), .A2(n10669), .ZN(n10666) );
  NAND2_X1 U7493 ( .A1(n11695), .A2(n11694), .ZN(n14094) );
  NAND2_X1 U7494 ( .A1(n7637), .A2(n7636), .ZN(n13206) );
  NAND2_X1 U7495 ( .A1(n7665), .A2(n7664), .ZN(n13228) );
  NAND2_X1 U7496 ( .A1(n10543), .A2(n7093), .ZN(n10672) );
  OR2_X1 U7497 ( .A1(n14264), .A2(n14263), .ZN(n7207) );
  OR2_X1 U7498 ( .A1(n10962), .A2(n13428), .ZN(n10960) );
  NAND2_X1 U7499 ( .A1(n7909), .A2(n7908), .ZN(n14396) );
  NAND2_X1 U7500 ( .A1(n14258), .A2(n6826), .ZN(n14264) );
  OR2_X1 U7501 ( .A1(n8892), .A2(n8895), .ZN(n8901) );
  NAND2_X1 U7502 ( .A1(n8470), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8487) );
  OR2_X1 U7503 ( .A1(n8606), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8623) );
  OR2_X1 U7504 ( .A1(n14546), .A2(n14547), .ZN(n14544) );
  NAND2_X1 U7505 ( .A1(n7852), .A2(n7851), .ZN(n10979) );
  NAND2_X1 U7506 ( .A1(n10910), .A2(n10909), .ZN(n14653) );
  NAND2_X1 U7507 ( .A1(n8469), .A2(n11062), .ZN(n7052) );
  NAND2_X1 U7508 ( .A1(n9721), .A2(n9692), .ZN(n9912) );
  NOR2_X1 U7509 ( .A1(n10016), .A2(n7350), .ZN(n7349) );
  NAND2_X1 U7510 ( .A1(n10625), .A2(n10624), .ZN(n14635) );
  INV_X1 U7511 ( .A(n11591), .ZN(n14919) );
  XNOR2_X1 U7512 ( .A(n14210), .B(n14209), .ZN(n14255) );
  NOR2_X1 U7513 ( .A1(n14528), .A2(n13701), .ZN(n13817) );
  NAND2_X1 U7514 ( .A1(n7805), .A2(n7804), .ZN(n7807) );
  NAND2_X1 U7515 ( .A1(n14566), .A2(n14565), .ZN(n14564) );
  NOR2_X1 U7516 ( .A1(n10049), .A2(n14941), .ZN(n12118) );
  AND2_X1 U7517 ( .A1(n10243), .A2(n10242), .ZN(n14603) );
  AND2_X2 U7518 ( .A1(n8177), .A2(n14751), .ZN(n14736) );
  NAND2_X1 U7519 ( .A1(n7754), .A2(n7753), .ZN(n10060) );
  OR2_X1 U7520 ( .A1(n9689), .A2(n9693), .ZN(n9691) );
  NAND2_X1 U7521 ( .A1(n10291), .A2(n14934), .ZN(n14946) );
  INV_X1 U7522 ( .A(n8178), .ZN(n7686) );
  NAND2_X1 U7523 ( .A1(n8358), .A2(n6628), .ZN(n12037) );
  INV_X1 U7524 ( .A(n12139), .ZN(n14922) );
  NAND4_X1 U7525 ( .A1(n7704), .A2(n7701), .A3(n7702), .A4(n7703), .ZN(n8876)
         );
  NAND3_X1 U7526 ( .A1(n8262), .A2(n8261), .A3(n6601), .ZN(n8278) );
  AND2_X1 U7527 ( .A1(n13466), .A2(n13613), .ZN(n6620) );
  CLKBUF_X1 U7528 ( .A(n7689), .Z(n7647) );
  INV_X2 U7529 ( .A(n6564), .ZN(n7967) );
  XNOR2_X1 U7530 ( .A(n14159), .B(n6843), .ZN(n14205) );
  NAND4_X1 U7532 ( .A1(n9744), .A2(n9743), .A3(n9742), .A4(n9741), .ZN(n13693)
         );
  INV_X2 U7533 ( .A(n6568), .ZN(n9026) );
  CLKBUF_X1 U7534 ( .A(n10236), .Z(n6824) );
  INV_X1 U7535 ( .A(n8682), .ZN(n6560) );
  XNOR2_X1 U7536 ( .A(n9155), .B(n9156), .ZN(n11952) );
  NAND2_X1 U7537 ( .A1(n7709), .A2(n7586), .ZN(n7722) );
  CLKBUF_X2 U7538 ( .A(n9072), .Z(n6567) );
  OAI211_X1 U7539 ( .C1(n9782), .C2(n6557), .A(n8257), .B(n8256), .ZN(n10050)
         );
  NAND3_X1 U7540 ( .A1(n8268), .A2(n8269), .A3(n8267), .ZN(n14932) );
  CLKBUF_X1 U7541 ( .A(n8815), .Z(n11411) );
  OAI211_X2 U7542 ( .C1(n13453), .C2(n9547), .A(n9546), .B(n9545), .ZN(n13473)
         );
  AND2_X1 U7543 ( .A1(n8240), .A2(n11627), .ZN(n8641) );
  NAND3_X1 U7544 ( .A1(n7428), .A2(n7427), .A3(n7430), .ZN(n8240) );
  CLKBUF_X2 U7545 ( .A(n8396), .Z(n8815) );
  INV_X2 U7546 ( .A(n8902), .ZN(n6561) );
  INV_X4 U7547 ( .A(n8898), .ZN(n9013) );
  NAND3_X1 U7548 ( .A1(n7426), .A2(n7425), .A3(n7430), .ZN(n8644) );
  AND2_X1 U7549 ( .A1(n9400), .A2(n14139), .ZN(n10244) );
  OR2_X1 U7550 ( .A1(n8238), .A2(n7433), .ZN(n7428) );
  NAND2_X1 U7551 ( .A1(n8238), .A2(n7432), .ZN(n7427) );
  INV_X2 U7552 ( .A(n13453), .ZN(n13444) );
  NAND2_X1 U7553 ( .A1(n13250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7564) );
  INV_X1 U7554 ( .A(n7287), .ZN(n7286) );
  AOI21_X1 U7555 ( .B1(n7262), .B2(n7735), .A(n7261), .ZN(n7260) );
  CLKBUF_X1 U7556 ( .A(n12610), .Z(n6831) );
  AND2_X1 U7557 ( .A1(n7591), .A2(n6728), .ZN(n7735) );
  XNOR2_X1 U7558 ( .A(n9436), .B(n9152), .ZN(n13636) );
  AND2_X1 U7559 ( .A1(n8213), .A2(n9130), .ZN(n8859) );
  INV_X1 U7560 ( .A(n13952), .ZN(n13965) );
  XNOR2_X1 U7561 ( .A(n7255), .B(n15162), .ZN(n14151) );
  AND2_X1 U7562 ( .A1(n11288), .A2(n9124), .ZN(n8857) );
  INV_X2 U7563 ( .A(n12602), .ZN(n12609) );
  XNOR2_X1 U7564 ( .A(n9222), .B(n9221), .ZN(n13464) );
  NAND2_X1 U7565 ( .A1(n6674), .A2(n7606), .ZN(n7288) );
  XNOR2_X1 U7566 ( .A(n7628), .B(n7561), .ZN(n8131) );
  OR2_X1 U7568 ( .A1(n8369), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8387) );
  OR2_X1 U7569 ( .A1(n7627), .A2(n8149), .ZN(n7628) );
  XNOR2_X1 U7570 ( .A(n8128), .B(n15275), .ZN(n11288) );
  XNOR2_X1 U7571 ( .A(n7949), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U7572 ( .A1(n9226), .A2(n6594), .ZN(n14142) );
  OAI21_X1 U7573 ( .B1(n8731), .B2(n7441), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8251) );
  XNOR2_X1 U7574 ( .A(n14154), .B(n7215), .ZN(n14192) );
  NAND2_X1 U7575 ( .A1(n8248), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8250) );
  NAND2_X2 U7576 ( .A1(n9020), .A2(P3_U3151), .ZN(n12606) );
  OR2_X1 U7577 ( .A1(n7468), .A2(n9479), .ZN(n9398) );
  NAND2_X1 U7578 ( .A1(n8164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8128) );
  NAND2_X2 U7579 ( .A1(n9251), .A2(P2_U3088), .ZN(n13269) );
  NAND2_X1 U7580 ( .A1(n8119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7949) );
  NAND2_X2 U7581 ( .A1(n9251), .A2(P1_U3086), .ZN(n14148) );
  OAI21_X1 U7582 ( .B1(n8119), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8121) );
  OR2_X1 U7583 ( .A1(n8335), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8355) );
  AND2_X1 U7584 ( .A1(n7439), .A2(n8237), .ZN(n7438) );
  OR2_X1 U7585 ( .A1(n9223), .A2(n7469), .ZN(n6594) );
  OR2_X1 U7586 ( .A1(n7526), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U7587 ( .A1(n9223), .A2(n6659), .ZN(n7468) );
  INV_X1 U7588 ( .A(n8393), .ZN(n7206) );
  NAND3_X1 U7589 ( .A1(n9217), .A2(n9151), .A3(n6548), .ZN(n9437) );
  NOR2_X1 U7590 ( .A1(n7353), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n7351) );
  NOR2_X1 U7591 ( .A1(n8321), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8324) );
  AND2_X1 U7592 ( .A1(n7203), .A2(n8228), .ZN(n7050) );
  AND2_X1 U7593 ( .A1(n8473), .A2(n8229), .ZN(n8230) );
  AND3_X1 U7594 ( .A1(n6757), .A2(n8232), .A3(n8231), .ZN(n8233) );
  AND2_X1 U7595 ( .A1(n7205), .A2(n8234), .ZN(n7203) );
  NAND2_X1 U7596 ( .A1(n8245), .A2(n8221), .ZN(n8301) );
  AND2_X1 U7597 ( .A1(n6733), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14196) );
  AND4_X1 U7598 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n8226)
         );
  AND2_X1 U7599 ( .A1(n8462), .A2(n8438), .ZN(n8473) );
  INV_X1 U7600 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9156) );
  NOR2_X1 U7601 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8231) );
  INV_X1 U7602 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8438) );
  NOR2_X1 U7603 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8232) );
  NOR2_X1 U7604 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n6757) );
  INV_X1 U7605 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9196) );
  NOR2_X1 U7606 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8224) );
  NOR2_X1 U7607 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8225) );
  INV_X1 U7608 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10094) );
  NOR2_X1 U7609 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9145) );
  NOR2_X1 U7610 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9146) );
  INV_X4 U7611 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7612 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8793) );
  INV_X1 U7613 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U7614 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8264) );
  INV_X1 U7615 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8228) );
  INV_X1 U7616 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8770) );
  NOR2_X2 U7617 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8245) );
  INV_X4 U7618 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7619 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7678) );
  INV_X1 U7620 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7705) );
  NOR2_X1 U7621 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7549) );
  NOR2_X1 U7622 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n7548) );
  INV_X2 U7623 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n12860) );
  NOR2_X1 U7624 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7547) );
  INV_X1 U7625 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U7626 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14195) );
  INV_X1 U7627 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7827) );
  INV_X1 U7628 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8252) );
  INV_X1 U7629 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9141) );
  INV_X4 U7630 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7631 ( .A1(n11952), .A2(n14149), .ZN(n9166) );
  NAND2_X1 U7632 ( .A1(n9709), .A2(n9708), .ZN(n9707) );
  NAND2_X1 U7633 ( .A1(n9517), .A2(n9516), .ZN(n9522) );
  NAND2_X2 U7634 ( .A1(n13306), .A2(n11881), .ZN(n13376) );
  NAND2_X2 U7635 ( .A1(n6726), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8675) );
  XNOR2_X1 U7636 ( .A(n8719), .B(n8703), .ZN(n11809) );
  INV_X1 U7637 ( .A(n11605), .ZN(n8717) );
  NOR2_X2 U7638 ( .A1(n10431), .A2(n13491), .ZN(n10388) );
  OR2_X1 U7639 ( .A1(n14578), .A2(n14596), .ZN(n10431) );
  NAND2_X2 U7640 ( .A1(n14441), .A2(n7483), .ZN(n7482) );
  NAND2_X2 U7641 ( .A1(n14443), .A2(n14442), .ZN(n14441) );
  NAND2_X2 U7642 ( .A1(n11333), .A2(n11332), .ZN(n14443) );
  OR2_X4 U7643 ( .A1(n7574), .A2(n13259), .ZN(n7690) );
  OR2_X1 U7644 ( .A1(n12969), .A2(n7123), .ZN(n7118) );
  AOI211_X2 U7645 ( .C1(n13167), .C2(n14731), .A(n13017), .B(n13016), .ZN(
        n13018) );
  NAND2_X1 U7646 ( .A1(n9162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9155) );
  OAI21_X2 U7647 ( .B1(n12395), .B2(n8546), .A(n8547), .ZN(n12381) );
  NOR2_X2 U7648 ( .A1(n13073), .A2(n13194), .ZN(n7140) );
  BUF_X8 U7649 ( .A(n11702), .Z(n6562) );
  INV_X2 U7650 ( .A(n7689), .ZN(n7679) );
  NAND2_X1 U7651 ( .A1(n8861), .A2(n9130), .ZN(n8898) );
  NAND2_X1 U7652 ( .A1(n7574), .A2(n7567), .ZN(n7691) );
  OAI21_X2 U7653 ( .B1(n8830), .B2(n11570), .A(n11567), .ZN(n11391) );
  AOI21_X2 U7654 ( .B1(n12257), .B2(n11605), .A(n11565), .ZN(n8830) );
  OAI21_X2 U7655 ( .B1(n13155), .B2(n8211), .A(n8210), .ZN(n12969) );
  NAND2_X2 U7656 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  OAI21_X2 U7657 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14201), .A(n14249), .ZN(
        n15300) );
  OAI21_X2 U7658 ( .B1(n13327), .B2(n7474), .A(n7472), .ZN(n13301) );
  NAND2_X2 U7659 ( .A1(n11845), .A2(n11844), .ZN(n13327) );
  OAI21_X2 U7660 ( .B1(n13368), .B2(n7462), .A(n7460), .ZN(n11841) );
  NAND2_X2 U7661 ( .A1(n11819), .A2(n11818), .ZN(n13368) );
  XNOR2_X2 U7662 ( .A(n9164), .B(n9163), .ZN(n9320) );
  AOI21_X2 U7663 ( .B1(n10562), .B2(n10561), .A(n6751), .ZN(n10583) );
  BUF_X2 U7664 ( .A(n7711), .Z(n6568) );
  NAND2_X2 U7665 ( .A1(n11671), .A2(n9251), .ZN(n13453) );
  NAND2_X1 U7666 ( .A1(n9557), .A2(n13636), .ZN(n14557) );
  INV_X1 U7667 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8249) );
  AOI21_X1 U7668 ( .B1(n12295), .B2(n7415), .A(n7414), .ZN(n12259) );
  NOR2_X1 U7669 ( .A1(n7418), .A2(n6579), .ZN(n7415) );
  OAI21_X1 U7670 ( .B1(n7416), .B2(n6579), .A(n6660), .ZN(n7414) );
  NAND2_X1 U7671 ( .A1(n12259), .A2(n8717), .ZN(n12258) );
  NAND2_X1 U7672 ( .A1(n6556), .A2(n9251), .ZN(n8288) );
  NAND2_X1 U7673 ( .A1(n6556), .A2(n9020), .ZN(n8396) );
  INV_X1 U7674 ( .A(n12824), .ZN(n8212) );
  AOI21_X1 U7675 ( .B1(n7114), .B2(n8194), .A(n6645), .ZN(n7113) );
  NAND2_X1 U7676 ( .A1(n7372), .A2(n6626), .ZN(n7369) );
  XNOR2_X1 U7677 ( .A(n14431), .B(n13682), .ZN(n13545) );
  NAND2_X1 U7678 ( .A1(n8058), .A2(n8057), .ZN(n8075) );
  INV_X1 U7679 ( .A(n7591), .ZN(n7261) );
  NAND2_X1 U7680 ( .A1(n7200), .A2(n11473), .ZN(n7199) );
  NAND2_X1 U7681 ( .A1(n8747), .A2(n11569), .ZN(n14943) );
  NAND2_X1 U7682 ( .A1(n7001), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8589) );
  AND2_X1 U7683 ( .A1(n6998), .A2(n6997), .ZN(n6996) );
  AND2_X1 U7684 ( .A1(n11768), .A2(n11767), .ZN(n13619) );
  INV_X1 U7685 ( .A(n13498), .ZN(n7254) );
  INV_X1 U7686 ( .A(n8910), .ZN(n8906) );
  NOR2_X1 U7687 ( .A1(n7259), .A2(n13588), .ZN(n7258) );
  NAND2_X1 U7688 ( .A1(n9835), .A2(n6758), .ZN(n9838) );
  OR2_X1 U7689 ( .A1(n9836), .A2(n15258), .ZN(n6758) );
  NAND2_X1 U7690 ( .A1(n6953), .A2(n7269), .ZN(n7940) );
  AOI21_X1 U7691 ( .B1(n7271), .B2(n7270), .A(n6667), .ZN(n7269) );
  AOI21_X1 U7692 ( .B1(n7419), .B2(n7417), .A(n6652), .ZN(n7416) );
  INV_X1 U7693 ( .A(n6603), .ZN(n7417) );
  OR2_X1 U7694 ( .A1(n12496), .A2(n12324), .ZN(n11548) );
  NOR2_X1 U7695 ( .A1(n6749), .A2(n8393), .ZN(n8773) );
  NAND2_X1 U7696 ( .A1(n8662), .A2(n8661), .ZN(n8663) );
  OR2_X1 U7697 ( .A1(n9066), .A2(n12960), .ZN(n9096) );
  NOR2_X1 U7698 ( .A1(n9060), .A2(n9050), .ZN(n9055) );
  OR2_X1 U7699 ( .A1(n13144), .A2(n8212), .ZN(n8107) );
  NAND2_X1 U7700 ( .A1(n13168), .A2(n12828), .ZN(n7106) );
  NOR2_X1 U7701 ( .A1(n6943), .A2(n6605), .ZN(n6942) );
  INV_X1 U7702 ( .A(n11154), .ZN(n7883) );
  NOR2_X1 U7703 ( .A1(n12976), .A2(n9119), .ZN(n7127) );
  NAND2_X1 U7704 ( .A1(n11778), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7446) );
  NOR2_X1 U7705 ( .A1(n7167), .A2(n6899), .ZN(n6898) );
  INV_X1 U7706 ( .A(n11801), .ZN(n6899) );
  NAND2_X1 U7707 ( .A1(n7170), .A2(n13857), .ZN(n7167) );
  INV_X1 U7708 ( .A(n11802), .ZN(n7170) );
  INV_X1 U7709 ( .A(n7155), .ZN(n7154) );
  INV_X1 U7710 ( .A(n8046), .ZN(n8044) );
  NAND2_X1 U7711 ( .A1(n7993), .A2(n7992), .ZN(n8018) );
  INV_X1 U7712 ( .A(n7638), .ZN(n7273) );
  XNOR2_X1 U7713 ( .A(n7624), .B(SI_16_), .ZN(n7638) );
  NOR2_X1 U7714 ( .A1(n6956), .A2(n6644), .ZN(n6955) );
  XNOR2_X1 U7715 ( .A(n7610), .B(SI_12_), .ZN(n7873) );
  XNOR2_X1 U7716 ( .A(n7609), .B(SI_11_), .ZN(n7860) );
  NAND2_X1 U7717 ( .A1(n7604), .A2(SI_9_), .ZN(n7606) );
  INV_X1 U7718 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U7719 ( .A1(n6730), .A2(n6729), .ZN(n6728) );
  NAND2_X1 U7720 ( .A1(n14153), .A2(n6796), .ZN(n14154) );
  NAND2_X1 U7721 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6797), .ZN(n6796) );
  INV_X1 U7722 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7723 ( .A1(n14157), .A2(n14158), .ZN(n14159) );
  AOI21_X1 U7724 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14179), .A(n14178), .ZN(
        n14230) );
  NOR2_X1 U7725 ( .A1(n14187), .A2(n14188), .ZN(n14178) );
  OAI21_X1 U7726 ( .B1(n7196), .B2(n11226), .A(n6584), .ZN(n6992) );
  AND3_X1 U7727 ( .A1(n8466), .A2(n8465), .A3(n8464), .ZN(n12459) );
  NAND2_X1 U7728 ( .A1(n10400), .A2(n7201), .ZN(n10599) );
  AND2_X1 U7729 ( .A1(n10405), .A2(n10399), .ZN(n7201) );
  NAND2_X1 U7730 ( .A1(n6985), .A2(n6984), .ZN(n12081) );
  INV_X1 U7731 ( .A(n12084), .ZN(n6984) );
  AOI21_X1 U7732 ( .B1(n10785), .B2(n10784), .A(n10783), .ZN(n10787) );
  INV_X1 U7733 ( .A(n11036), .ZN(n7198) );
  NAND2_X1 U7734 ( .A1(n12222), .A2(n6994), .ZN(n6995) );
  OR2_X1 U7735 ( .A1(n8288), .A2(n9272), .ZN(n8257) );
  OR2_X1 U7736 ( .A1(n8396), .A2(SI_2_), .ZN(n8256) );
  INV_X1 U7737 ( .A(n8641), .ZN(n8673) );
  OR2_X1 U7738 ( .A1(n8238), .A2(n6688), .ZN(n7426) );
  NAND2_X1 U7739 ( .A1(n8238), .A2(n7429), .ZN(n7425) );
  INV_X1 U7740 ( .A(n14337), .ZN(n7012) );
  OR2_X1 U7741 ( .A1(n14345), .A2(n14346), .ZN(n6852) );
  OAI21_X1 U7742 ( .B1(n12350), .B2(n7041), .A(n7039), .ZN(n12325) );
  AND2_X1 U7743 ( .A1(n7040), .A2(n11538), .ZN(n7039) );
  OR2_X1 U7744 ( .A1(n7041), .A2(n11534), .ZN(n7040) );
  NAND2_X1 U7745 ( .A1(n12222), .A2(n10202), .ZN(n11613) );
  INV_X1 U7746 ( .A(n8529), .ZN(n11409) );
  NAND2_X1 U7747 ( .A1(n8804), .A2(n11433), .ZN(n14971) );
  NOR2_X1 U7748 ( .A1(n8731), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8767) );
  OR2_X1 U7749 ( .A1(n8615), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8616) );
  AOI21_X1 U7750 ( .B1(n8506), .B2(n7059), .A(n7058), .ZN(n7057) );
  INV_X1 U7751 ( .A(n8523), .ZN(n7058) );
  INV_X1 U7752 ( .A(n8503), .ZN(n7059) );
  INV_X1 U7753 ( .A(n8506), .ZN(n7060) );
  NAND2_X1 U7754 ( .A1(n9173), .A2(n7631), .ZN(n7711) );
  NAND2_X1 U7755 ( .A1(n9173), .A2(n9251), .ZN(n9072) );
  OR2_X1 U7756 ( .A1(n13213), .A2(n12787), .ZN(n6909) );
  AOI21_X1 U7757 ( .B1(n7110), .B2(n7109), .A(n6662), .ZN(n7108) );
  INV_X1 U7758 ( .A(n7114), .ZN(n7109) );
  NAND2_X1 U7759 ( .A1(n6915), .A2(n7872), .ZN(n11155) );
  NAND2_X1 U7760 ( .A1(n11019), .A2(n11018), .ZN(n6915) );
  NAND2_X1 U7761 ( .A1(n7307), .A2(n9943), .ZN(n9948) );
  NOR2_X1 U7762 ( .A1(n14029), .A2(n14033), .ZN(n7082) );
  INV_X1 U7763 ( .A(n7373), .ZN(n7372) );
  NAND2_X1 U7764 ( .A1(n6577), .A2(n7379), .ZN(n7374) );
  INV_X1 U7765 ( .A(n13857), .ZN(n7376) );
  NAND2_X1 U7766 ( .A1(n13941), .A2(n11796), .ZN(n13926) );
  NOR2_X1 U7767 ( .A1(n7154), .A2(n6888), .ZN(n6887) );
  INV_X1 U7768 ( .A(n6602), .ZN(n7153) );
  AND2_X1 U7769 ( .A1(n7389), .A2(n13560), .ZN(n7387) );
  OAI21_X1 U7770 ( .B1(n7388), .B2(n7386), .A(n13561), .ZN(n7385) );
  INV_X1 U7771 ( .A(n13560), .ZN(n7386) );
  OAI21_X1 U7772 ( .B1(n11790), .B2(n11789), .A(n11791), .ZN(n14004) );
  NAND2_X1 U7773 ( .A1(n10906), .A2(n10905), .ZN(n10959) );
  AOI21_X1 U7774 ( .B1(n7396), .B2(n7393), .A(n6646), .ZN(n7392) );
  INV_X1 U7775 ( .A(n10631), .ZN(n7393) );
  INV_X1 U7776 ( .A(n13619), .ZN(n14029) );
  NAND2_X1 U7777 ( .A1(n9462), .A2(n13615), .ZN(n14571) );
  OR3_X1 U7778 ( .A1(n11137), .A2(n8777), .A3(n11240), .ZN(n9963) );
  NAND2_X1 U7779 ( .A1(n8716), .A2(n8715), .ZN(n12130) );
  NOR2_X1 U7780 ( .A1(n12230), .A2(n6805), .ZN(n12233) );
  NOR2_X1 U7781 ( .A1(n12226), .A2(n12519), .ZN(n6805) );
  NAND2_X1 U7782 ( .A1(n12264), .A2(n6772), .ZN(n12480) );
  NAND2_X1 U7783 ( .A1(n6773), .A2(n14924), .ZN(n6772) );
  NAND2_X1 U7784 ( .A1(n10449), .A2(n10417), .ZN(n10448) );
  INV_X1 U7785 ( .A(n6764), .ZN(n10417) );
  INV_X1 U7786 ( .A(n6927), .ZN(n13142) );
  INV_X1 U7787 ( .A(n8142), .ZN(n6937) );
  NAND2_X1 U7788 ( .A1(n6932), .A2(n14753), .ZN(n6929) );
  NOR2_X1 U7789 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  NAND2_X1 U7790 ( .A1(n6845), .A2(n6844), .ZN(n13483) );
  NAND2_X1 U7791 ( .A1(n13596), .A2(n13480), .ZN(n6844) );
  NAND2_X1 U7792 ( .A1(n13481), .A2(n6620), .ZN(n6845) );
  NOR2_X1 U7793 ( .A1(n7495), .A2(n7494), .ZN(n6874) );
  NAND2_X1 U7794 ( .A1(n7497), .A2(n6604), .ZN(n7496) );
  OR2_X1 U7795 ( .A1(n13499), .A2(n7254), .ZN(n6760) );
  NAND2_X1 U7796 ( .A1(n7254), .A2(n13499), .ZN(n6762) );
  MUX2_X1 U7797 ( .A(n13689), .B(n13506), .S(n13617), .Z(n13507) );
  AOI21_X1 U7798 ( .B1(n7501), .B2(n8907), .A(n8905), .ZN(n7500) );
  OAI21_X1 U7799 ( .B1(n8901), .B2(n7506), .A(n7505), .ZN(n8908) );
  AND2_X1 U7800 ( .A1(n13536), .A2(n7235), .ZN(n7234) );
  NAND2_X1 U7801 ( .A1(n7236), .A2(n13530), .ZN(n7235) );
  NOR2_X1 U7802 ( .A1(n7224), .A2(n7220), .ZN(n7219) );
  INV_X1 U7803 ( .A(n13557), .ZN(n7220) );
  NAND2_X1 U7804 ( .A1(n13990), .A2(n7223), .ZN(n7222) );
  INV_X1 U7805 ( .A(n13562), .ZN(n7223) );
  MUX2_X1 U7806 ( .A(n13674), .B(n13919), .S(n13617), .Z(n13589) );
  NOR2_X1 U7807 ( .A1(n8973), .A2(n8969), .ZN(n7520) );
  NAND2_X1 U7808 ( .A1(n6800), .A2(n11569), .ZN(n6799) );
  NAND2_X1 U7809 ( .A1(n11568), .A2(n11567), .ZN(n6800) );
  INV_X1 U7810 ( .A(n6863), .ZN(n6862) );
  OAI21_X1 U7811 ( .B1(n7524), .B2(n6698), .A(n6864), .ZN(n6863) );
  INV_X1 U7812 ( .A(n8998), .ZN(n6864) );
  INV_X1 U7813 ( .A(n7992), .ZN(n7268) );
  NOR2_X1 U7814 ( .A1(n6574), .A2(n7974), .ZN(n6961) );
  NAND2_X1 U7815 ( .A1(n10050), .A2(n6553), .ZN(n11439) );
  INV_X1 U7816 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7205) );
  INV_X1 U7817 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U7818 ( .A1(n6862), .A2(n6698), .ZN(n6861) );
  OR4_X1 U7819 ( .A1(n13433), .A2(n13432), .A3(n13431), .A4(n13430), .ZN(
        n13437) );
  NAND2_X1 U7820 ( .A1(n13602), .A2(n7241), .ZN(n7240) );
  INV_X1 U7821 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U7822 ( .A1(n6980), .A2(n6607), .ZN(n6978) );
  NAND2_X1 U7823 ( .A1(n12117), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U7824 ( .A1(n11965), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U7825 ( .A1(n9834), .A2(n6804), .ZN(n9873) );
  OR2_X1 U7826 ( .A1(n9836), .A2(n10329), .ZN(n6804) );
  AND3_X1 U7827 ( .A1(n7017), .A2(n7015), .A3(n6788), .ZN(n9935) );
  NAND2_X1 U7828 ( .A1(n9934), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6788) );
  AOI21_X1 U7829 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10315), .A(n10314), .ZN(
        n10482) );
  OR2_X1 U7830 ( .A1(n8726), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U7831 ( .A1(n8679), .A2(n8678), .ZN(n8694) );
  INV_X1 U7832 ( .A(n8680), .ZN(n8679) );
  INV_X1 U7833 ( .A(n7423), .ZN(n7420) );
  NAND2_X1 U7834 ( .A1(n7424), .A2(n12054), .ZN(n7423) );
  INV_X1 U7835 ( .A(n12492), .ZN(n7424) );
  INV_X1 U7836 ( .A(n12295), .ZN(n7422) );
  OR2_X1 U7837 ( .A1(n12572), .A2(n12370), .ZN(n11584) );
  NOR2_X1 U7838 ( .A1(n12373), .A2(n7037), .ZN(n7036) );
  INV_X1 U7839 ( .A(n11524), .ZN(n7037) );
  INV_X1 U7840 ( .A(n7036), .ZN(n7035) );
  INV_X1 U7841 ( .A(n11485), .ZN(n7047) );
  OR2_X1 U7842 ( .A1(n12437), .A2(n12459), .ZN(n11491) );
  NOR2_X1 U7843 ( .A1(n8444), .A2(n7049), .ZN(n7048) );
  INV_X1 U7844 ( .A(n11480), .ZN(n7049) );
  OR2_X1 U7845 ( .A1(n12136), .A2(n10855), .ZN(n11462) );
  NAND2_X1 U7846 ( .A1(n8314), .A2(n8313), .ZN(n8335) );
  INV_X1 U7847 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U7848 ( .A1(n11313), .A2(n7436), .ZN(n12451) );
  INV_X1 U7849 ( .A(n11433), .ZN(n11428) );
  AND4_X1 U7850 ( .A1(n8235), .A2(n8770), .A3(n8793), .A4(n8768), .ZN(n6616)
         );
  NOR2_X1 U7851 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8235) );
  NAND2_X1 U7852 ( .A1(n8468), .A2(n8467), .ZN(n8469) );
  NAND2_X1 U7853 ( .A1(n8363), .A2(n8365), .ZN(n7068) );
  AND2_X1 U7854 ( .A1(n12626), .A2(n7337), .ZN(n7336) );
  INV_X1 U7855 ( .A(n12625), .ZN(n7334) );
  NAND2_X1 U7856 ( .A1(n12651), .A2(n7320), .ZN(n7319) );
  INV_X1 U7857 ( .A(n12652), .ZN(n7320) );
  INV_X1 U7858 ( .A(n12723), .ZN(n7366) );
  NAND2_X1 U7859 ( .A1(n9034), .A2(n9096), .ZN(n9099) );
  OR4_X1 U7860 ( .A1(n12996), .A2(n13014), .A3(n13036), .A4(n9116), .ZN(n9117)
         );
  NAND2_X1 U7861 ( .A1(n7634), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U7862 ( .A1(n9122), .A2(n6935), .ZN(n6934) );
  INV_X1 U7863 ( .A(n8107), .ZN(n6935) );
  INV_X1 U7864 ( .A(n6934), .ZN(n6931) );
  NOR2_X1 U7865 ( .A1(n12998), .A2(n12991), .ZN(n7132) );
  NOR2_X1 U7866 ( .A1(n6550), .A2(n6605), .ZN(n6940) );
  NOR2_X2 U7867 ( .A1(n14398), .A2(n13213), .ZN(n7142) );
  NAND2_X1 U7868 ( .A1(n6661), .A2(n7842), .ZN(n7317) );
  AND2_X1 U7869 ( .A1(n7115), .A2(n6677), .ZN(n7114) );
  INV_X1 U7870 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8165) );
  INV_X1 U7871 ( .A(n11821), .ZN(n11882) );
  INV_X1 U7872 ( .A(n13464), .ZN(n9461) );
  INV_X1 U7873 ( .A(n7369), .ZN(n7368) );
  NOR2_X1 U7874 ( .A1(n13901), .A2(n14051), .ZN(n7086) );
  NOR2_X1 U7875 ( .A1(n13911), .A2(n7403), .ZN(n7402) );
  INV_X1 U7876 ( .A(n7404), .ZN(n7403) );
  OAI21_X1 U7877 ( .B1(n13930), .B2(n7164), .A(n11798), .ZN(n7163) );
  INV_X1 U7878 ( .A(n11797), .ZN(n7164) );
  NOR2_X1 U7879 ( .A1(n13930), .A2(n7405), .ZN(n7404) );
  INV_X1 U7880 ( .A(n7408), .ZN(n7405) );
  NOR2_X1 U7881 ( .A1(n14277), .A2(n14274), .ZN(n7092) );
  NAND2_X1 U7882 ( .A1(n14151), .A2(n13965), .ZN(n13463) );
  AOI21_X1 U7883 ( .B1(n7293), .B2(n7291), .A(n7290), .ZN(n7289) );
  INV_X1 U7884 ( .A(n9022), .ZN(n7290) );
  INV_X1 U7885 ( .A(n9016), .ZN(n7291) );
  INV_X1 U7886 ( .A(n7293), .ZN(n7292) );
  NAND2_X1 U7887 ( .A1(n8111), .A2(n8110), .ZN(n9017) );
  NAND2_X1 U7888 ( .A1(n7274), .A2(n6715), .ZN(n8111) );
  INV_X1 U7889 ( .A(n8108), .ZN(n7283) );
  NAND2_X1 U7890 ( .A1(n7282), .A2(SI_26_), .ZN(n7281) );
  INV_X1 U7891 ( .A(n8074), .ZN(n7282) );
  NOR2_X1 U7892 ( .A1(n7279), .A2(n8090), .ZN(n7278) );
  INV_X1 U7893 ( .A(n7280), .ZN(n7279) );
  NAND2_X1 U7894 ( .A1(n8075), .A2(n7281), .ZN(n6954) );
  NAND2_X1 U7895 ( .A1(n8074), .A2(n11238), .ZN(n7280) );
  INV_X1 U7896 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9150) );
  INV_X1 U7897 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U7898 ( .A(n8037), .B(SI_24_), .ZN(n8040) );
  INV_X1 U7899 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n15162) );
  NAND2_X1 U7900 ( .A1(n7978), .A2(n6962), .ZN(n7990) );
  INV_X1 U7901 ( .A(n7272), .ZN(n7271) );
  OAI21_X1 U7902 ( .B1(n7622), .B2(n7273), .A(n7625), .ZN(n7272) );
  NAND2_X1 U7903 ( .A1(n7655), .A2(n7619), .ZN(n7623) );
  OR2_X1 U7904 ( .A1(n10092), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U7905 ( .A1(n8276), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6841) );
  XNOR2_X1 U7906 ( .A(n14156), .B(n7213), .ZN(n14191) );
  INV_X1 U7907 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7213) );
  INV_X1 U7908 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6843) );
  AOI21_X1 U7909 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14172), .A(n14171), .ZN(
        n14173) );
  NOR2_X1 U7910 ( .A1(n14190), .A2(n14189), .ZN(n14171) );
  NOR2_X1 U7911 ( .A1(n7180), .A2(n7177), .ZN(n7176) );
  INV_X1 U7912 ( .A(n12051), .ZN(n7177) );
  INV_X1 U7913 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U7914 ( .A1(n6607), .A2(n6982), .ZN(n6979) );
  OR2_X1 U7915 ( .A1(n8540), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8556) );
  INV_X1 U7916 ( .A(n6978), .ZN(n6977) );
  AOI21_X1 U7917 ( .B1(n6978), .B2(n6979), .A(n6976), .ZN(n6975) );
  INV_X1 U7918 ( .A(n12060), .ZN(n6976) );
  INV_X1 U7919 ( .A(n11226), .ZN(n6993) );
  NOR2_X1 U7920 ( .A1(n6992), .A2(n11229), .ZN(n6990) );
  NAND2_X1 U7921 ( .A1(n8447), .A2(n11230), .ZN(n8480) );
  INV_X1 U7922 ( .A(n8448), .ZN(n8447) );
  NAND2_X1 U7923 ( .A1(n6983), .A2(n11977), .ZN(n11978) );
  OR2_X1 U7924 ( .A1(n11976), .A2(n12345), .ZN(n11977) );
  NAND2_X1 U7925 ( .A1(n12043), .A2(n12044), .ZN(n6983) );
  INV_X1 U7926 ( .A(n10786), .ZN(n7197) );
  NAND2_X1 U7927 ( .A1(n10601), .A2(n10600), .ZN(n10785) );
  NAND2_X1 U7928 ( .A1(n8513), .A2(n15103), .ZN(n8540) );
  INV_X1 U7929 ( .A(n8514), .ZN(n8513) );
  OAI21_X1 U7930 ( .B1(n9782), .B2(P3_REG2_REG_2__SCAN_IN), .A(n7014), .ZN(
        n9596) );
  NAND2_X1 U7931 ( .A1(n9782), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U7932 ( .A1(n9791), .A2(n9805), .ZN(n9793) );
  OR2_X1 U7933 ( .A1(n10317), .A2(n10316), .ZN(n6787) );
  OR2_X1 U7934 ( .A1(n14306), .A2(n12183), .ZN(n7013) );
  OR2_X1 U7935 ( .A1(n8811), .A2(n12261), .ZN(n7540) );
  OAI21_X2 U7936 ( .B1(n12276), .B2(n11557), .A(n11423), .ZN(n12257) );
  NAND2_X1 U7937 ( .A1(n7413), .A2(n7416), .ZN(n12272) );
  NAND2_X1 U7938 ( .A1(n12295), .A2(n7419), .ZN(n7413) );
  NAND2_X1 U7939 ( .A1(n12296), .A2(n12453), .ZN(n6768) );
  NAND2_X1 U7940 ( .A1(n7044), .A2(n7043), .ZN(n12348) );
  INV_X1 U7941 ( .A(n12351), .ZN(n7043) );
  NAND2_X1 U7942 ( .A1(n11516), .A2(n11523), .ZN(n12373) );
  NAND2_X1 U7943 ( .A1(n12399), .A2(n11511), .ZN(n12392) );
  AND4_X1 U7944 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n12397)
         );
  AOI21_X1 U7945 ( .B1(n7436), .B2(n11481), .A(n6621), .ZN(n7435) );
  AND2_X1 U7946 ( .A1(n11198), .A2(n8384), .ZN(n11047) );
  NAND2_X1 U7947 ( .A1(n11047), .A2(n11468), .ZN(n11046) );
  AND2_X1 U7948 ( .A1(n11470), .A2(n11469), .ZN(n11586) );
  NAND2_X1 U7949 ( .A1(n11196), .A2(n11586), .ZN(n11195) );
  NAND2_X1 U7950 ( .A1(n10288), .A2(n11590), .ZN(n10287) );
  INV_X1 U7951 ( .A(n14941), .ZN(n12456) );
  OR2_X1 U7952 ( .A1(n8288), .A2(n9260), .ZN(n8268) );
  OR2_X1 U7953 ( .A1(n10286), .A2(n10285), .ZN(n10291) );
  NAND2_X1 U7954 ( .A1(n12237), .A2(n10202), .ZN(n11580) );
  AND2_X1 U7955 ( .A1(n9963), .A2(n9319), .ZN(n9982) );
  OR2_X1 U7956 ( .A1(n8802), .A2(n8806), .ZN(n9979) );
  INV_X1 U7957 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U7958 ( .A1(n6616), .A2(n8236), .ZN(n7441) );
  NOR2_X1 U7959 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n8236) );
  XNOR2_X1 U7960 ( .A(n8775), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8778) );
  INV_X1 U7961 ( .A(n8773), .ZN(n8774) );
  NAND2_X1 U7962 ( .A1(n7069), .A2(n7070), .ZN(n8660) );
  AOI21_X1 U7963 ( .B1(n8632), .B2(n7071), .A(n6593), .ZN(n7070) );
  XNOR2_X1 U7964 ( .A(n8733), .B(n8766), .ZN(n8804) );
  AOI21_X1 U7965 ( .B1(n7057), .B2(n7060), .A(n7055), .ZN(n7054) );
  INV_X1 U7966 ( .A(n8526), .ZN(n7055) );
  AND2_X1 U7967 ( .A1(n8523), .A2(n8505), .ZN(n8506) );
  NAND2_X1 U7968 ( .A1(n8487), .A2(n7052), .ZN(n8490) );
  AND2_X1 U7969 ( .A1(n9281), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8363) );
  CLKBUF_X1 U7970 ( .A(n8364), .Z(n6750) );
  OR2_X1 U7971 ( .A1(n7955), .A2(n7954), .ZN(n7982) );
  AND2_X1 U7972 ( .A1(n7866), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7892) );
  AND2_X1 U7973 ( .A1(n10853), .A2(n10843), .ZN(n6820) );
  NAND2_X1 U7974 ( .A1(n6868), .A2(n9098), .ZN(n6866) );
  AOI21_X1 U7975 ( .B1(n9055), .B2(n7297), .A(n9092), .ZN(n7296) );
  AND2_X1 U7976 ( .A1(n9055), .A2(n9054), .ZN(n7510) );
  INV_X1 U7977 ( .A(n13259), .ZN(n7567) );
  NAND2_X1 U7978 ( .A1(n13257), .A2(n13259), .ZN(n7689) );
  OAI21_X1 U7979 ( .B1(n13454), .B2(n6568), .A(n9073), .ZN(n12956) );
  AND2_X1 U7980 ( .A1(n8107), .A2(n8105), .ZN(n9119) );
  AND2_X1 U7981 ( .A1(n8215), .A2(n8098), .ZN(n12708) );
  NAND2_X1 U7982 ( .A1(n7132), .A2(n7131), .ZN(n12970) );
  INV_X1 U7983 ( .A(n8209), .ZN(n7097) );
  NAND2_X1 U7984 ( .A1(n6948), .A2(n6952), .ZN(n6943) );
  AND2_X1 U7985 ( .A1(n6946), .A2(n13060), .ZN(n6945) );
  NAND2_X1 U7986 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  NOR2_X1 U7987 ( .A1(n13071), .A2(n6950), .ZN(n6949) );
  NOR2_X1 U7988 ( .A1(n6571), .A2(n7315), .ZN(n6950) );
  NAND2_X1 U7989 ( .A1(n13091), .A2(n12834), .ZN(n7315) );
  INV_X1 U7990 ( .A(n13084), .ZN(n7316) );
  NOR2_X1 U7991 ( .A1(n12749), .A2(n13219), .ZN(n6911) );
  NAND2_X1 U7992 ( .A1(n7919), .A2(n7545), .ZN(n7313) );
  NAND2_X1 U7993 ( .A1(n7300), .A2(n7883), .ZN(n11158) );
  OR2_X1 U7994 ( .A1(n10979), .A2(n12842), .ZN(n7115) );
  NAND2_X1 U7995 ( .A1(n10666), .A2(n6613), .ZN(n10812) );
  OAI21_X1 U7996 ( .B1(n10547), .B2(n7803), .A(n7802), .ZN(n10668) );
  NOR2_X1 U7997 ( .A1(n10675), .A2(n7094), .ZN(n7093) );
  INV_X1 U7998 ( .A(n8190), .ZN(n7094) );
  NAND2_X1 U7999 ( .A1(n7730), .A2(n9748), .ZN(n9750) );
  NAND2_X1 U8000 ( .A1(n7697), .A2(n7698), .ZN(n10067) );
  INV_X1 U8001 ( .A(n10069), .ZN(n7697) );
  INV_X1 U8002 ( .A(n10070), .ZN(n7698) );
  INV_X1 U8003 ( .A(n13002), .ZN(n13162) );
  CLKBUF_X1 U8004 ( .A(n14808), .Z(n6774) );
  NOR2_X1 U8005 ( .A1(n11387), .A2(n8163), .ZN(n9422) );
  AOI21_X1 U8006 ( .B1(n13278), .B2(n11928), .A(n11939), .ZN(n7453) );
  INV_X1 U8007 ( .A(n7453), .ZN(n7451) );
  NAND2_X1 U8008 ( .A1(n13359), .A2(n13358), .ZN(n7467) );
  AOI21_X1 U8009 ( .B1(n7458), .B2(n7459), .A(n7456), .ZN(n7455) );
  INV_X1 U8010 ( .A(n13349), .ZN(n7456) );
  MUX2_X1 U8011 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14152), .S(n11671), .Z(n9658)
         );
  NOR2_X1 U8012 ( .A1(n14455), .A2(n7484), .ZN(n7483) );
  INV_X1 U8013 ( .A(n11341), .ZN(n7484) );
  OAI22_X1 U8014 ( .A1(n9656), .A2(n7412), .B1(n10237), .B2(n11884), .ZN(n9737) );
  AOI22_X1 U8015 ( .A1(n11821), .A2(n13473), .B1(n9654), .B2(n13696), .ZN(
        n9655) );
  NOR2_X1 U8016 ( .A1(n7476), .A2(n13386), .ZN(n7475) );
  INV_X1 U8017 ( .A(n7535), .ZN(n7476) );
  INV_X1 U8018 ( .A(n7463), .ZN(n7462) );
  AOI21_X1 U8019 ( .B1(n7463), .B2(n7461), .A(n6650), .ZN(n7460) );
  OR2_X1 U8020 ( .A1(n11085), .A2(n11084), .ZN(n11178) );
  AND2_X1 U8021 ( .A1(n13641), .A2(n13642), .ZN(n6846) );
  AND2_X1 U8022 ( .A1(n11678), .A2(n11677), .ZN(n15203) );
  OR2_X1 U8023 ( .A1(n11769), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9743) );
  NAND4_X1 U8024 ( .A1(n9402), .A2(n9401), .A3(n7446), .A4(n7445), .ZN(n10236)
         );
  NAND2_X1 U8025 ( .A1(n10245), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7445) );
  AOI21_X1 U8026 ( .B1(n14472), .B2(n10877), .A(n10876), .ZN(n10878) );
  NAND2_X1 U8027 ( .A1(n13447), .A2(n13446), .ZN(n13646) );
  NAND2_X1 U8028 ( .A1(n13457), .A2(n13456), .ZN(n13824) );
  OR2_X1 U8029 ( .A1(n13454), .A2(n13453), .ZN(n13457) );
  AOI21_X1 U8030 ( .B1(n7169), .B2(n7166), .A(n6655), .ZN(n7165) );
  NAND2_X1 U8031 ( .A1(n13889), .A2(n6898), .ZN(n6897) );
  NAND2_X1 U8032 ( .A1(n13872), .A2(n13871), .ZN(n7168) );
  INV_X1 U8033 ( .A(n7167), .ZN(n7169) );
  INV_X1 U8034 ( .A(n7380), .ZN(n7377) );
  XNOR2_X1 U8035 ( .A(n14040), .B(n6969), .ZN(n13857) );
  INV_X1 U8036 ( .A(n7168), .ZN(n13874) );
  NAND2_X1 U8037 ( .A1(n7086), .A2(n7085), .ZN(n13866) );
  AOI21_X1 U8038 ( .B1(n7087), .B2(n13673), .A(n13897), .ZN(n13879) );
  NAND2_X1 U8039 ( .A1(n14072), .A2(n15203), .ZN(n7406) );
  NAND2_X1 U8040 ( .A1(n13945), .A2(n7404), .ZN(n7407) );
  NOR2_X1 U8041 ( .A1(n13964), .A2(n13954), .ZN(n13944) );
  NAND2_X1 U8042 ( .A1(n13926), .A2(n13930), .ZN(n13925) );
  NOR2_X1 U8043 ( .A1(n6886), .A2(n13946), .ZN(n6884) );
  INV_X1 U8044 ( .A(n11794), .ZN(n7157) );
  NAND2_X1 U8045 ( .A1(n7159), .A2(n13568), .ZN(n7158) );
  AND2_X1 U8046 ( .A1(n13958), .A2(n7158), .ZN(n7155) );
  AND2_X1 U8047 ( .A1(n13989), .A2(n7382), .ZN(n13972) );
  NOR2_X1 U8048 ( .A1(n13974), .A2(n7383), .ZN(n7382) );
  INV_X1 U8049 ( .A(n13563), .ZN(n7383) );
  OR2_X1 U8050 ( .A1(n6891), .A2(n6888), .ZN(n11795) );
  NOR2_X1 U8051 ( .A1(n14004), .A2(n11793), .ZN(n6891) );
  AOI21_X1 U8052 ( .B1(n7389), .B2(n13433), .A(n6664), .ZN(n7388) );
  NAND2_X1 U8053 ( .A1(n6902), .A2(n6901), .ZN(n11790) );
  AOI21_X1 U8054 ( .B1(n6903), .B2(n13545), .A(n6649), .ZN(n6901) );
  AND2_X1 U8055 ( .A1(n13549), .A2(n7390), .ZN(n7389) );
  INV_X1 U8056 ( .A(n13432), .ZN(n7390) );
  OR2_X1 U8057 ( .A1(n11837), .A2(n11838), .ZN(n13549) );
  NOR2_X1 U8058 ( .A1(n11258), .A2(n6904), .ZN(n6903) );
  INV_X1 U8059 ( .A(n11255), .ZN(n6904) );
  NAND2_X1 U8060 ( .A1(n11170), .A2(n11169), .ZN(n11242) );
  NAND2_X1 U8061 ( .A1(n7092), .A2(n7091), .ZN(n11175) );
  AOI21_X1 U8062 ( .B1(n6878), .B2(n6880), .A(n6648), .ZN(n6876) );
  NAND2_X1 U8063 ( .A1(n10632), .A2(n10631), .ZN(n10694) );
  NOR2_X1 U8064 ( .A1(n7395), .A2(n7394), .ZN(n10695) );
  INV_X1 U8065 ( .A(n10693), .ZN(n7394) );
  INV_X1 U8066 ( .A(n10694), .ZN(n7395) );
  NAND2_X1 U8067 ( .A1(n10692), .A2(n10691), .ZN(n13514) );
  XNOR2_X1 U8068 ( .A(n13514), .B(n13687), .ZN(n13426) );
  NAND2_X1 U8069 ( .A1(n7151), .A2(n10621), .ZN(n10687) );
  OAI21_X1 U8070 ( .B1(n10522), .B2(n6669), .A(n10525), .ZN(n14546) );
  AND4_X1 U8071 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n13490) );
  AND2_X1 U8072 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10251) );
  AND2_X1 U8073 ( .A1(n7410), .A2(n7409), .ZN(n14565) );
  NAND2_X1 U8074 ( .A1(n10237), .A2(n13696), .ZN(n7409) );
  NAND2_X1 U8075 ( .A1(n13467), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U8076 ( .A1(n7412), .A2(n13473), .ZN(n7411) );
  XNOR2_X1 U8077 ( .A(n13696), .B(n13473), .ZN(n13417) );
  AND2_X1 U8078 ( .A1(n9672), .A2(n9669), .ZN(n11784) );
  AND2_X1 U8079 ( .A1(n9455), .A2(n9454), .ZN(n10390) );
  AND2_X1 U8080 ( .A1(n14628), .A2(n14642), .ZN(n14639) );
  AND2_X1 U8081 ( .A1(n9557), .A2(n9556), .ZN(n14636) );
  AND2_X1 U8082 ( .A1(n10364), .A2(n9325), .ZN(n10231) );
  AND2_X1 U8083 ( .A1(n7294), .A2(n9019), .ZN(n7293) );
  INV_X1 U8084 ( .A(n9068), .ZN(n7294) );
  NAND2_X1 U8085 ( .A1(n9017), .A2(n9016), .ZN(n7295) );
  XNOR2_X1 U8086 ( .A(n8075), .B(n8059), .ZN(n13267) );
  OR2_X1 U8087 ( .A1(n9629), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n10103) );
  OAI21_X1 U8088 ( .B1(n7822), .B2(n7288), .A(n7286), .ZN(n7861) );
  INV_X1 U8089 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U8090 ( .A1(n7260), .A2(n6925), .ZN(n7746) );
  NAND2_X1 U8091 ( .A1(n7722), .A2(n6919), .ZN(n6925) );
  INV_X1 U8092 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6733) );
  XNOR2_X1 U8093 ( .A(n6830), .B(n14196), .ZN(n14198) );
  INV_X1 U8094 ( .A(n14195), .ZN(n6830) );
  INV_X1 U8095 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7215) );
  XNOR2_X1 U8096 ( .A(n14191), .B(n6734), .ZN(n14203) );
  OAI22_X1 U8097 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14879), .B1(n14230), 
        .B2(n14180), .ZN(n14236) );
  OAI21_X1 U8098 ( .B1(n14239), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n14509), .ZN(
        n14241) );
  OR2_X1 U8099 ( .A1(n11411), .A2(n15059), .ZN(n8704) );
  NAND2_X1 U8100 ( .A1(n11809), .A2(n11409), .ZN(n8705) );
  NAND2_X1 U8101 ( .A1(n7191), .A2(n12454), .ZN(n7190) );
  INV_X1 U8102 ( .A(n11963), .ZN(n7191) );
  XNOR2_X1 U8103 ( .A(n11983), .B(n11985), .ZN(n12006) );
  NAND2_X1 U8104 ( .A1(n11033), .A2(n7199), .ZN(n11035) );
  AND2_X1 U8105 ( .A1(n11033), .A2(n6575), .ZN(n11100) );
  AND2_X1 U8106 ( .A1(n10162), .A2(n10161), .ZN(n10164) );
  NAND2_X1 U8107 ( .A1(n10164), .A2(n10163), .ZN(n10400) );
  NAND2_X1 U8108 ( .A1(n8620), .A2(n8619), .ZN(n12338) );
  NAND2_X1 U8109 ( .A1(n11989), .A2(n11988), .ZN(n12050) );
  NAND2_X1 U8110 ( .A1(n12074), .A2(n12075), .ZN(n11989) );
  OR2_X1 U8111 ( .A1(n11973), .A2(n12370), .ZN(n11974) );
  NAND2_X2 U8112 ( .A1(n8605), .A2(n8604), .ZN(n12509) );
  AND3_X1 U8113 ( .A1(n8655), .A2(n8654), .A3(n8653), .ZN(n12324) );
  NAND2_X1 U8114 ( .A1(n8638), .A2(n8637), .ZN(n12327) );
  NOR2_X1 U8115 ( .A1(n7075), .A2(n11609), .ZN(n11610) );
  INV_X1 U8116 ( .A(n12274), .ZN(n12296) );
  INV_X1 U8117 ( .A(n12359), .ZN(n12385) );
  NOR2_X1 U8118 ( .A1(n14912), .A2(n7005), .ZN(n7003) );
  AND2_X1 U8119 ( .A1(n7007), .A2(n7008), .ZN(n7005) );
  NAND2_X1 U8120 ( .A1(n7008), .A2(n7011), .ZN(n7006) );
  OR2_X1 U8121 ( .A1(n12186), .A2(n12210), .ZN(n6851) );
  AND2_X1 U8122 ( .A1(n8750), .A2(n8749), .ZN(n12248) );
  INV_X1 U8123 ( .A(n14934), .ZN(n12468) );
  OR2_X1 U8124 ( .A1(n14979), .A2(n12549), .ZN(n6837) );
  NOR2_X1 U8125 ( .A1(n12480), .A2(n6656), .ZN(n12548) );
  XNOR2_X1 U8126 ( .A(n8771), .B(n8770), .ZN(n11137) );
  OAI21_X1 U8127 ( .B1(n8769), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8771) );
  OAI211_X1 U8128 ( .C1(n8767), .C2(n7189), .A(n7187), .B(n7185), .ZN(n8777)
         );
  INV_X1 U8129 ( .A(n7188), .ZN(n7187) );
  OAI22_X1 U8130 ( .A1(n6576), .A2(n7189), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_24__SCAN_IN), .ZN(n7188) );
  INV_X1 U8131 ( .A(n12222), .ZN(n12237) );
  NAND2_X1 U8132 ( .A1(n8531), .A2(n6998), .ZN(n8588) );
  NAND2_X1 U8133 ( .A1(n7878), .A2(n7877), .ZN(n14689) );
  NAND2_X1 U8134 ( .A1(n9909), .A2(n9914), .ZN(n10010) );
  NAND2_X1 U8135 ( .A1(n10190), .A2(n10189), .ZN(n10449) );
  AOI21_X1 U8136 ( .B1(n7349), .B2(n7347), .A(n7346), .ZN(n7345) );
  AND2_X1 U8137 ( .A1(n7331), .A2(n10423), .ZN(n7330) );
  OAI21_X1 U8138 ( .B1(n10690), .B2(n6568), .A(n7831), .ZN(n10895) );
  NAND2_X1 U8139 ( .A1(n9429), .A2(n14751), .ZN(n14690) );
  OR2_X1 U8140 ( .A1(n9428), .A2(n9414), .ZN(n12792) );
  NAND2_X1 U8141 ( .A1(n7891), .A2(n7890), .ZN(n14410) );
  AND2_X1 U8142 ( .A1(n6558), .A2(n14748), .ZN(n14731) );
  AND2_X1 U8143 ( .A1(n7134), .A2(n13140), .ZN(n6936) );
  NOR2_X1 U8144 ( .A1(n14427), .A2(n7464), .ZN(n7463) );
  INV_X1 U8145 ( .A(n11827), .ZN(n7464) );
  NAND2_X1 U8146 ( .A1(n13366), .A2(n11827), .ZN(n14428) );
  NAND2_X1 U8147 ( .A1(n11293), .A2(n11292), .ZN(n14106) );
  NAND2_X1 U8148 ( .A1(n11692), .A2(n11691), .ZN(n13435) );
  NAND2_X1 U8149 ( .A1(n13368), .A2(n13367), .ZN(n13366) );
  AND2_X1 U8150 ( .A1(n11784), .A2(n10390), .ZN(n14433) );
  NOR2_X1 U8151 ( .A1(n10558), .A2(n6752), .ZN(n6751) );
  AOI21_X1 U8152 ( .B1(n9485), .B2(n9636), .A(n9627), .ZN(n9632) );
  INV_X1 U8153 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U8154 ( .A1(n13818), .A2(n13819), .ZN(n6780) );
  NOR2_X1 U8155 ( .A1(n13816), .A2(n6778), .ZN(n6777) );
  NAND2_X1 U8156 ( .A1(n6779), .A2(n13952), .ZN(n6778) );
  NAND2_X1 U8157 ( .A1(n13820), .A2(n13965), .ZN(n6781) );
  AND2_X1 U8158 ( .A1(n13669), .A2(n13662), .ZN(n11776) );
  NAND2_X1 U8159 ( .A1(n6894), .A2(n6900), .ZN(n6893) );
  AND2_X1 U8160 ( .A1(n7084), .A2(n7083), .ZN(n14027) );
  OR2_X1 U8161 ( .A1(n14575), .A2(n10275), .ZN(n14012) );
  INV_X1 U8162 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U8163 ( .A1(n6912), .A2(n7823), .ZN(n10690) );
  OR2_X1 U8164 ( .A1(n7822), .A2(n7821), .ZN(n6912) );
  XNOR2_X1 U8165 ( .A(n14198), .B(n14199), .ZN(n15304) );
  OAI21_X1 U8166 ( .B1(n14260), .B2(n14259), .A(n6827), .ZN(n6826) );
  INV_X1 U8167 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14305) );
  INV_X1 U8168 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U8169 ( .A1(n8888), .A2(n8887), .ZN(n7533) );
  NAND2_X1 U8170 ( .A1(n7504), .A2(n8907), .ZN(n7503) );
  INV_X1 U8171 ( .A(n7506), .ZN(n7504) );
  INV_X1 U8172 ( .A(n7505), .ZN(n7501) );
  NOR2_X1 U8173 ( .A1(n6609), .A2(n8900), .ZN(n7506) );
  NAND2_X1 U8174 ( .A1(n6609), .A2(n8900), .ZN(n7505) );
  NOR2_X1 U8175 ( .A1(n13510), .A2(n13509), .ZN(n7252) );
  NAND2_X1 U8176 ( .A1(n7253), .A2(n13513), .ZN(n7251) );
  NAND2_X1 U8177 ( .A1(n7230), .A2(n13521), .ZN(n7228) );
  INV_X1 U8178 ( .A(n13521), .ZN(n7226) );
  AOI21_X1 U8179 ( .B1(n6640), .B2(n8919), .A(n8918), .ZN(n7518) );
  NAND2_X1 U8180 ( .A1(n6632), .A2(n8919), .ZN(n7519) );
  NOR2_X1 U8181 ( .A1(n6640), .A2(n8919), .ZN(n6859) );
  NAND2_X1 U8182 ( .A1(n8910), .A2(n6632), .ZN(n6858) );
  OAI21_X1 U8183 ( .B1(n7229), .B2(n7227), .A(n7225), .ZN(n13524) );
  NAND2_X1 U8184 ( .A1(n7226), .A2(n13520), .ZN(n7225) );
  AND2_X1 U8185 ( .A1(n13516), .A2(n13515), .ZN(n7229) );
  NAND2_X1 U8186 ( .A1(n13519), .A2(n7228), .ZN(n7227) );
  AND2_X1 U8187 ( .A1(n13532), .A2(n7238), .ZN(n7237) );
  INV_X1 U8188 ( .A(n13530), .ZN(n7238) );
  AND2_X1 U8189 ( .A1(n13547), .A2(n13546), .ZN(n13548) );
  AND2_X1 U8190 ( .A1(n8948), .A2(n7499), .ZN(n7498) );
  AND2_X1 U8191 ( .A1(n7222), .A2(n13565), .ZN(n7221) );
  NAND2_X1 U8192 ( .A1(n7249), .A2(n13581), .ZN(n7247) );
  OAI21_X1 U8193 ( .B1(n7256), .B2(n13587), .A(n7257), .ZN(n13593) );
  NAND2_X1 U8194 ( .A1(n13588), .A2(n7259), .ZN(n7257) );
  NAND2_X1 U8195 ( .A1(n8982), .A2(n6702), .ZN(n7513) );
  OAI21_X1 U8196 ( .B1(n8978), .B2(n8977), .A(n6706), .ZN(n6870) );
  NAND2_X1 U8197 ( .A1(n7525), .A2(n8994), .ZN(n7524) );
  NAND2_X1 U8198 ( .A1(n8995), .A2(n7523), .ZN(n7522) );
  INV_X1 U8199 ( .A(n8994), .ZN(n7523) );
  INV_X1 U8200 ( .A(n7922), .ZN(n7626) );
  AND2_X1 U8201 ( .A1(n6617), .A2(n7273), .ZN(n7270) );
  AOI21_X1 U8202 ( .B1(n7286), .B2(n7288), .A(n7285), .ZN(n7284) );
  INV_X1 U8203 ( .A(n7860), .ZN(n7285) );
  INV_X1 U8204 ( .A(n9933), .ZN(n7018) );
  OR2_X1 U8205 ( .A1(n13465), .A2(n13636), .ZN(n13466) );
  INV_X1 U8206 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9148) );
  AND2_X1 U8207 ( .A1(n8025), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U8208 ( .A1(n8017), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U8209 ( .A1(n7944), .A2(n9717), .ZN(n7962) );
  NOR2_X1 U8210 ( .A1(n6959), .A2(n6958), .ZN(n6957) );
  INV_X1 U8211 ( .A(n7603), .ZN(n6958) );
  NOR2_X1 U8212 ( .A1(n6959), .A2(n7286), .ZN(n6956) );
  NAND2_X1 U8213 ( .A1(n7214), .A2(n14155), .ZN(n14156) );
  NAND2_X1 U8214 ( .A1(n12037), .A2(n10838), .ZN(n11463) );
  INV_X1 U8215 ( .A(n14932), .ZN(n14931) );
  NOR2_X1 U8216 ( .A1(n8803), .A2(n11428), .ZN(n6994) );
  OR2_X1 U8217 ( .A1(n7432), .A2(n15270), .ZN(n7429) );
  NAND2_X1 U8218 ( .A1(n7019), .A2(n9874), .ZN(n7016) );
  INV_X1 U8219 ( .A(n9838), .ZN(n7019) );
  NAND2_X1 U8220 ( .A1(n9838), .A2(n9837), .ZN(n9869) );
  NAND2_X1 U8221 ( .A1(n9927), .A2(n9928), .ZN(n10117) );
  NAND2_X1 U8222 ( .A1(n12195), .A2(n12196), .ZN(n12198) );
  OR2_X1 U8223 ( .A1(n11959), .A2(n12026), .ZN(n11574) );
  OR2_X1 U8224 ( .A1(n8694), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U8225 ( .A1(n8668), .A2(n8667), .ZN(n8680) );
  INV_X1 U8226 ( .A(n8669), .ZN(n8668) );
  OR2_X1 U8227 ( .A1(n8651), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8669) );
  OR2_X1 U8228 ( .A1(n12327), .A2(n12335), .ZN(n11542) );
  NAND2_X1 U8229 ( .A1(n8622), .A2(n8621), .ZN(n8639) );
  INV_X1 U8230 ( .A(n8623), .ZN(n8622) );
  NAND2_X1 U8231 ( .A1(n11473), .A2(n14967), .ZN(n7029) );
  NOR2_X1 U8232 ( .A1(n11473), .A2(n14967), .ZN(n7028) );
  INV_X1 U8233 ( .A(n7028), .ZN(n7027) );
  OR2_X1 U8234 ( .A1(n12037), .A2(n10838), .ZN(n11464) );
  NAND2_X1 U8235 ( .A1(n12138), .A2(n10298), .ZN(n11445) );
  NAND2_X1 U8236 ( .A1(n11437), .A2(n11436), .ZN(n10081) );
  AND2_X1 U8237 ( .A1(n15270), .A2(P3_IR_REG_30__SCAN_IN), .ZN(n7432) );
  OAI22_X1 U8238 ( .A1(n8533), .A2(n7431), .B1(P3_IR_REG_31__SCAN_IN), .B2(
        P3_IR_REG_30__SCAN_IN), .ZN(n7430) );
  NOR2_X1 U8239 ( .A1(n15270), .A2(P3_IR_REG_30__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U8240 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7434), .ZN(n7433) );
  INV_X1 U8241 ( .A(n8634), .ZN(n7072) );
  INV_X1 U8242 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8234) );
  AND2_X1 U8243 ( .A1(n8233), .A2(n7205), .ZN(n7204) );
  INV_X1 U8244 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6997) );
  AND2_X1 U8245 ( .A1(n8530), .A2(n8534), .ZN(n7000) );
  AND2_X1 U8246 ( .A1(n8230), .A2(n8228), .ZN(n7437) );
  NAND2_X1 U8247 ( .A1(n8227), .A2(n8226), .ZN(n8393) );
  INV_X1 U8248 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U8249 ( .A1(n8252), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8275) );
  AND2_X1 U8250 ( .A1(n7366), .A2(n12756), .ZN(n7362) );
  NAND2_X1 U8251 ( .A1(n6663), .A2(n9004), .ZN(n7531) );
  NOR2_X1 U8252 ( .A1(n9056), .A2(n9057), .ZN(n7297) );
  OR2_X1 U8253 ( .A1(n9091), .A2(n9046), .ZN(n9060) );
  INV_X1 U8254 ( .A(n7100), .ZN(n7098) );
  NAND2_X1 U8255 ( .A1(n8005), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8028) );
  INV_X1 U8256 ( .A(n6949), .ZN(n6947) );
  INV_X1 U8257 ( .A(n6917), .ZN(n6916) );
  OAI21_X1 U8258 ( .B1(n11018), .B2(n6918), .A(n7884), .ZN(n6917) );
  INV_X1 U8259 ( .A(n7872), .ZN(n6918) );
  NOR2_X1 U8260 ( .A1(n6569), .A2(n10680), .ZN(n7149) );
  NAND2_X1 U8261 ( .A1(n9952), .A2(n9956), .ZN(n9953) );
  NAND2_X1 U8262 ( .A1(n7125), .A2(n7124), .ZN(n7123) );
  NAND2_X1 U8263 ( .A1(n7527), .A2(n7629), .ZN(n7526) );
  INV_X1 U8264 ( .A(n7528), .ZN(n7527) );
  NAND2_X1 U8265 ( .A1(n7640), .A2(n7351), .ZN(n8119) );
  OR2_X1 U8266 ( .A1(n7770), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7788) );
  AOI21_X1 U8267 ( .B1(n13286), .B2(n11889), .A(n13348), .ZN(n7458) );
  INV_X1 U8268 ( .A(n13286), .ZN(n7459) );
  INV_X1 U8269 ( .A(n13367), .ZN(n7461) );
  OR4_X1 U8270 ( .A1(n13439), .A2(n13974), .A3(n13958), .A4(n13438), .ZN(
        n13440) );
  INV_X1 U8271 ( .A(n13610), .ZN(n7245) );
  AND2_X1 U8272 ( .A1(n13621), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U8273 ( .A1(n7244), .A2(n13610), .ZN(n7243) );
  INV_X1 U8274 ( .A(n13622), .ZN(n7244) );
  OAI22_X1 U8275 ( .A1(n11380), .A2(n11379), .B1(n11378), .B2(n11377), .ZN(
        n13807) );
  NAND2_X1 U8276 ( .A1(n14045), .A2(n11745), .ZN(n7380) );
  NOR2_X1 U8277 ( .A1(n13913), .A2(n13919), .ZN(n7088) );
  NAND2_X1 U8278 ( .A1(n6889), .A2(n11793), .ZN(n6883) );
  NOR2_X2 U8279 ( .A1(n11175), .A2(n14431), .ZN(n7090) );
  INV_X1 U8280 ( .A(n6879), .ZN(n6878) );
  OAI21_X1 U8281 ( .B1(n13428), .B2(n6880), .A(n13429), .ZN(n6879) );
  INV_X1 U8282 ( .A(n10912), .ZN(n6880) );
  NOR2_X1 U8283 ( .A1(n14559), .A2(n13506), .ZN(n7081) );
  NAND2_X1 U8284 ( .A1(n10436), .A2(n14573), .ZN(n13479) );
  NAND2_X1 U8285 ( .A1(n10268), .A2(n10267), .ZN(n14567) );
  OR2_X1 U8286 ( .A1(n13417), .A2(n10266), .ZN(n10268) );
  NAND2_X1 U8287 ( .A1(n9160), .A2(n7470), .ZN(n7469) );
  INV_X1 U8288 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U8289 ( .A1(n7940), .A2(SI_18_), .ZN(n7941) );
  XNOR2_X1 U8290 ( .A(n7613), .B(n9328), .ZN(n7885) );
  NOR2_X2 U8291 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9476) );
  NOR2_X1 U8292 ( .A1(n6924), .A2(n7593), .ZN(n6923) );
  NAND2_X1 U8293 ( .A1(n6666), .A2(n7590), .ZN(n6907) );
  INV_X1 U8294 ( .A(n12107), .ZN(n7181) );
  NAND2_X1 U8295 ( .A1(n7194), .A2(n6608), .ZN(n6991) );
  NAND2_X1 U8296 ( .A1(n10787), .A2(n10786), .ZN(n11033) );
  NAND2_X1 U8297 ( .A1(n8479), .A2(n8478), .ZN(n8495) );
  INV_X1 U8298 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8478) );
  OR2_X1 U8299 ( .A1(n8404), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8424) );
  OR2_X1 U8300 ( .A1(n8424), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U8301 ( .A(n10050), .B(n11032), .ZN(n10160) );
  XNOR2_X1 U8302 ( .A(n12588), .B(n11032), .ZN(n11966) );
  NAND2_X1 U8303 ( .A1(n11998), .A2(n12409), .ZN(n6982) );
  OR2_X1 U8304 ( .A1(n8495), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U8305 ( .A1(n8311), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U8306 ( .A1(n6560), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U8307 ( .A1(n9856), .A2(n9594), .ZN(n9595) );
  NAND2_X1 U8308 ( .A1(n9596), .A2(n9595), .ZN(n9790) );
  NAND2_X1 U8309 ( .A1(n9586), .A2(n9585), .ZN(n9787) );
  INV_X1 U8310 ( .A(n7026), .ZN(n7025) );
  XNOR2_X1 U8311 ( .A(n9873), .B(n9837), .ZN(n9876) );
  NOR2_X1 U8312 ( .A1(n9839), .A2(n9840), .ZN(n9871) );
  OR2_X1 U8313 ( .A1(n8361), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8378) );
  OR2_X1 U8314 ( .A1(n7020), .A2(n10115), .ZN(n9937) );
  XNOR2_X1 U8315 ( .A(n10486), .B(n10483), .ZN(n10310) );
  NAND2_X1 U8316 ( .A1(n10310), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U8317 ( .A1(n6787), .A2(n6635), .ZN(n7024) );
  NAND2_X1 U8318 ( .A1(n10490), .A2(n10491), .ZN(n12195) );
  AOI21_X1 U8319 ( .B1(n7024), .B2(n7023), .A(n7021), .ZN(n12176) );
  NOR2_X1 U8320 ( .A1(n12144), .A2(n7022), .ZN(n7021) );
  INV_X1 U8321 ( .A(n12174), .ZN(n7023) );
  OR2_X1 U8322 ( .A1(n14881), .A2(n14880), .ZN(n14884) );
  OR2_X1 U8323 ( .A1(n14901), .A2(n14900), .ZN(n14904) );
  OR2_X1 U8324 ( .A1(n14330), .A2(n14329), .ZN(n14332) );
  AND2_X1 U8325 ( .A1(n8531), .A2(n8530), .ZN(n8535) );
  NAND2_X1 U8326 ( .A1(n8531), .A2(n7000), .ZN(n8568) );
  AOI21_X1 U8327 ( .B1(n14347), .B2(n12213), .A(n12212), .ZN(n12230) );
  OR2_X1 U8328 ( .A1(n12224), .A2(n12220), .ZN(n7011) );
  INV_X1 U8329 ( .A(n7009), .ZN(n7008) );
  OAI21_X1 U8330 ( .B1(n12188), .B2(n7011), .A(n7010), .ZN(n7009) );
  NAND2_X1 U8331 ( .A1(n12224), .A2(n12220), .ZN(n7010) );
  AND2_X1 U8332 ( .A1(n14336), .A2(n12185), .ZN(n12186) );
  NAND2_X1 U8333 ( .A1(n11413), .A2(n11412), .ZN(n11415) );
  NAND2_X1 U8334 ( .A1(n11574), .A2(n11572), .ZN(n11582) );
  AND2_X1 U8335 ( .A1(n8718), .A2(n11563), .ZN(n7442) );
  INV_X1 U8336 ( .A(n8756), .ZN(n12316) );
  INV_X1 U8337 ( .A(n12345), .ZN(n12323) );
  AND2_X1 U8338 ( .A1(n11542), .A2(n11543), .ZN(n12326) );
  NAND2_X1 U8339 ( .A1(n8595), .A2(n8594), .ZN(n8606) );
  INV_X1 U8340 ( .A(n8596), .ZN(n8595) );
  AND2_X1 U8341 ( .A1(n11585), .A2(n11584), .ZN(n12361) );
  AOI21_X1 U8342 ( .B1(n7036), .B2(n7034), .A(n11520), .ZN(n7033) );
  NOR2_X1 U8343 ( .A1(n7035), .A2(n7032), .ZN(n7031) );
  NAND2_X1 U8344 ( .A1(n8555), .A2(n8554), .ZN(n8572) );
  INV_X1 U8345 ( .A(n8556), .ZN(n8555) );
  OR2_X1 U8346 ( .A1(n8572), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8596) );
  AND2_X1 U8347 ( .A1(n11502), .A2(n11508), .ZN(n12412) );
  INV_X1 U8348 ( .A(n7046), .ZN(n7045) );
  OAI21_X1 U8349 ( .B1(n7048), .B2(n7047), .A(n12449), .ZN(n7046) );
  INV_X1 U8350 ( .A(n11315), .ZN(n8445) );
  NAND2_X1 U8351 ( .A1(n11141), .A2(n7048), .ZN(n11319) );
  NAND2_X1 U8352 ( .A1(n11046), .A2(n8403), .ZN(n11145) );
  NAND2_X1 U8353 ( .A1(n8386), .A2(n8385), .ZN(n8404) );
  INV_X1 U8354 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8385) );
  INV_X1 U8355 ( .A(n8387), .ZN(n8386) );
  INV_X1 U8356 ( .A(n11586), .ZN(n8383) );
  NAND2_X1 U8357 ( .A1(n10829), .A2(n8368), .ZN(n11199) );
  NAND2_X1 U8358 ( .A1(n8354), .A2(n8353), .ZN(n8369) );
  INV_X1 U8359 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8353) );
  INV_X1 U8360 ( .A(n11594), .ZN(n8350) );
  AND2_X1 U8361 ( .A1(n11462), .A2(n11460), .ZN(n11594) );
  INV_X1 U8362 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n8294) );
  AOI21_X1 U8363 ( .B1(n11591), .B2(n14918), .A(n8282), .ZN(n10174) );
  NAND2_X1 U8364 ( .A1(n10042), .A2(n11437), .ZN(n14915) );
  CLKBUF_X1 U8365 ( .A(n10081), .Z(n14937) );
  INV_X1 U8366 ( .A(n14971), .ZN(n14966) );
  OR2_X1 U8367 ( .A1(n8780), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8368 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7189) );
  AND2_X1 U8369 ( .A1(n6576), .A2(n8768), .ZN(n7186) );
  NAND2_X1 U8370 ( .A1(n8675), .A2(n8664), .ZN(n8674) );
  XNOR2_X1 U8371 ( .A(n8794), .B(n8793), .ZN(n9962) );
  AND2_X1 U8372 ( .A1(n8602), .A2(n8584), .ZN(n8585) );
  AND2_X1 U8373 ( .A1(n7000), .A2(n6999), .ZN(n6998) );
  INV_X1 U8374 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8375 ( .A1(n8509), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U8376 ( .A1(n7437), .A2(n8410), .ZN(n8509) );
  AND2_X1 U8377 ( .A1(n9543), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8454) );
  CLKBUF_X1 U8378 ( .A(n8393), .Z(n8394) );
  AOI21_X1 U8379 ( .B1(n7066), .B2(n7065), .A(n6668), .ZN(n7064) );
  INV_X1 U8380 ( .A(n8365), .ZN(n7065) );
  XNOR2_X1 U8381 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8397) );
  XNOR2_X1 U8382 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8341) );
  XNOR2_X1 U8383 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8327) );
  XNOR2_X1 U8384 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8303) );
  INV_X1 U8385 ( .A(n8245), .ZN(n6759) );
  CLKBUF_X1 U8386 ( .A(n8275), .Z(n6789) );
  OR2_X1 U8387 ( .A1(n7795), .A2(n7794), .ZN(n7813) );
  INV_X1 U8388 ( .A(n12846), .ZN(n10193) );
  OR2_X1 U8389 ( .A1(n8081), .A2(n12680), .ZN(n8097) );
  INV_X1 U8390 ( .A(n7362), .ZN(n7356) );
  AND2_X1 U8391 ( .A1(n12672), .A2(n12671), .ZN(n7364) );
  XNOR2_X1 U8392 ( .A(n10060), .B(n6554), .ZN(n10006) );
  NAND2_X1 U8393 ( .A1(n7570), .A2(n7569), .ZN(n7931) );
  NAND2_X1 U8394 ( .A1(n7336), .A2(n7334), .ZN(n7333) );
  INV_X1 U8395 ( .A(n7336), .ZN(n7335) );
  INV_X1 U8396 ( .A(n9683), .ZN(n7324) );
  AND2_X1 U8397 ( .A1(n9688), .A2(n9521), .ZN(n7325) );
  XNOR2_X1 U8398 ( .A(n14794), .B(n12663), .ZN(n9913) );
  INV_X1 U8399 ( .A(n9914), .ZN(n7347) );
  INV_X1 U8400 ( .A(n10187), .ZN(n7346) );
  NAND2_X1 U8401 ( .A1(n10457), .A2(n10416), .ZN(n6764) );
  NAND2_X1 U8402 ( .A1(n7984), .A2(n7983), .ZN(n7996) );
  INV_X1 U8403 ( .A(n7982), .ZN(n7984) );
  NAND2_X1 U8404 ( .A1(n7571), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7955) );
  INV_X1 U8405 ( .A(n7933), .ZN(n7571) );
  NOR2_X1 U8406 ( .A1(n7365), .A2(n7359), .ZN(n7358) );
  INV_X1 U8407 ( .A(n7361), .ZN(n7359) );
  OR2_X1 U8408 ( .A1(n12799), .A2(n12670), .ZN(n7365) );
  NAND2_X1 U8409 ( .A1(n7366), .A2(n12662), .ZN(n7361) );
  NAND2_X1 U8410 ( .A1(n12757), .A2(n7362), .ZN(n7360) );
  NAND2_X1 U8411 ( .A1(n14384), .A2(n12625), .ZN(n12732) );
  NAND2_X1 U8412 ( .A1(n7640), .A2(n7352), .ZN(n7947) );
  INV_X1 U8413 ( .A(n7353), .ZN(n7352) );
  INV_X1 U8414 ( .A(n7120), .ZN(n7119) );
  OAI21_X1 U8415 ( .B1(n7123), .B2(n7127), .A(n7121), .ZN(n7120) );
  NAND2_X1 U8416 ( .A1(n7126), .A2(n9122), .ZN(n7121) );
  NAND2_X1 U8417 ( .A1(n6934), .A2(n7124), .ZN(n6932) );
  NOR2_X1 U8418 ( .A1(n6930), .A2(n13189), .ZN(n6928) );
  NOR2_X1 U8419 ( .A1(n6933), .A2(n6931), .ZN(n6930) );
  NOR2_X1 U8420 ( .A1(n9122), .A2(n6935), .ZN(n6933) );
  INV_X1 U8421 ( .A(n7132), .ZN(n12986) );
  OR2_X1 U8422 ( .A1(n7103), .A2(n7101), .ZN(n7100) );
  INV_X1 U8423 ( .A(n7106), .ZN(n7101) );
  NAND2_X1 U8424 ( .A1(n6675), .A2(n7106), .ZN(n7099) );
  OR2_X1 U8425 ( .A1(n7104), .A2(n7105), .ZN(n7103) );
  INV_X1 U8426 ( .A(n9102), .ZN(n7104) );
  NAND2_X1 U8427 ( .A1(n7139), .A2(n7138), .ZN(n13021) );
  AND2_X1 U8428 ( .A1(n13179), .A2(n12830), .ZN(n7105) );
  INV_X1 U8429 ( .A(n6782), .ZN(n13039) );
  NOR2_X1 U8430 ( .A1(n6940), .A2(n6951), .ZN(n6939) );
  NAND2_X1 U8431 ( .A1(n13084), .A2(n6942), .ZN(n6941) );
  NOR2_X1 U8432 ( .A1(n12777), .A2(n13053), .ZN(n6951) );
  NAND2_X1 U8433 ( .A1(n7140), .A2(n13185), .ZN(n13047) );
  NOR2_X1 U8434 ( .A1(n7145), .A2(n13206), .ZN(n7141) );
  INV_X1 U8435 ( .A(n14398), .ZN(n7143) );
  NAND2_X1 U8436 ( .A1(n7309), .A2(n6572), .ZN(n7308) );
  INV_X1 U8437 ( .A(n7311), .ZN(n7309) );
  NOR2_X1 U8438 ( .A1(n13116), .A2(n13119), .ZN(n13115) );
  NOR2_X1 U8439 ( .A1(n11364), .A2(n7312), .ZN(n7311) );
  INV_X1 U8440 ( .A(n7920), .ZN(n7312) );
  NAND2_X1 U8441 ( .A1(n7892), .A2(n7568), .ZN(n7912) );
  OR2_X1 U8442 ( .A1(n7912), .A2(n15161), .ZN(n7914) );
  INV_X1 U8443 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15161) );
  OR2_X1 U8444 ( .A1(n6613), .A2(n7317), .ZN(n6905) );
  OR2_X1 U8445 ( .A1(n7813), .A2(n7812), .ZN(n7834) );
  NOR2_X1 U8446 ( .A1(n7834), .A2(n7833), .ZN(n7854) );
  NAND2_X1 U8447 ( .A1(n10676), .A2(n7149), .ZN(n10978) );
  NAND2_X1 U8448 ( .A1(n10676), .A2(n14803), .ZN(n10818) );
  INV_X1 U8449 ( .A(n14378), .ZN(n12800) );
  AND2_X1 U8450 ( .A1(n11220), .A2(n11288), .ZN(n14745) );
  AND2_X1 U8451 ( .A1(n7127), .A2(n9122), .ZN(n7122) );
  NAND2_X1 U8452 ( .A1(n8027), .A2(n8026), .ZN(n13168) );
  NAND2_X1 U8453 ( .A1(n7112), .A2(n7113), .ZN(n11153) );
  NAND2_X1 U8454 ( .A1(n10973), .A2(n7114), .ZN(n7112) );
  INV_X1 U8455 ( .A(n14795), .ZN(n14819) );
  NAND2_X1 U8456 ( .A1(n7560), .A2(n7529), .ZN(n7528) );
  INV_X1 U8457 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7560) );
  INV_X1 U8458 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7529) );
  XNOR2_X1 U8459 ( .A(n8151), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8173) );
  NOR2_X1 U8460 ( .A1(n8153), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8150) );
  CLKBUF_X1 U8461 ( .A(n8152), .Z(n8153) );
  AND2_X1 U8462 ( .A1(n7633), .A2(n6872), .ZN(n6871) );
  AND2_X1 U8463 ( .A1(n7632), .A2(n6873), .ZN(n6872) );
  INV_X1 U8464 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6873) );
  INV_X1 U8465 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n15275) );
  OR2_X1 U8466 ( .A1(n7875), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7887) );
  OR2_X1 U8467 ( .A1(n7725), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U8468 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  NAND2_X1 U8469 ( .A1(n11680), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11730) );
  NOR2_X1 U8470 ( .A1(n11853), .A2(n7479), .ZN(n7478) );
  INV_X1 U8471 ( .A(n7480), .ZN(n7479) );
  NAND2_X1 U8472 ( .A1(n7493), .A2(n7492), .ZN(n7491) );
  INV_X1 U8473 ( .A(n10800), .ZN(n7492) );
  INV_X1 U8474 ( .A(n10799), .ZN(n7493) );
  AND2_X1 U8475 ( .A1(n11920), .A2(n11918), .ZN(n13319) );
  NAND2_X1 U8476 ( .A1(n11843), .A2(n11842), .ZN(n7480) );
  NAND2_X1 U8477 ( .A1(n13375), .A2(n11890), .ZN(n13285) );
  AND2_X1 U8478 ( .A1(n13321), .A2(n11907), .ZN(n13349) );
  INV_X1 U8479 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10950) );
  AND2_X1 U8480 ( .A1(n9660), .A2(n9659), .ZN(n9709) );
  AOI21_X1 U8481 ( .B1(n9654), .B2(n9658), .A(n7546), .ZN(n9659) );
  AND2_X1 U8482 ( .A1(n9657), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n7546) );
  OAI211_X1 U8483 ( .C1(n10442), .C2(n11882), .A(n7444), .B(n7443), .ZN(n9708)
         );
  NAND2_X1 U8484 ( .A1(n9654), .A2(n6824), .ZN(n7444) );
  OR2_X1 U8485 ( .A1(n10364), .A2(n9661), .ZN(n7443) );
  NAND2_X1 U8486 ( .A1(n10925), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11069) );
  OR2_X1 U8487 ( .A1(n11069), .A2(n11068), .ZN(n11085) );
  NOR2_X1 U8488 ( .A1(n13308), .A2(n7466), .ZN(n7465) );
  INV_X1 U8489 ( .A(n11874), .ZN(n7466) );
  AND2_X1 U8490 ( .A1(n10917), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10925) );
  NOR2_X1 U8491 ( .A1(n11697), .A2(n11696), .ZN(n11705) );
  OR2_X1 U8492 ( .A1(n11300), .A2(n11299), .ZN(n11697) );
  OR2_X1 U8493 ( .A1(n11852), .A2(n11851), .ZN(n7535) );
  NAND2_X1 U8494 ( .A1(n13327), .A2(n7478), .ZN(n7477) );
  NOR2_X1 U8495 ( .A1(n11178), .A2(n11177), .ZN(n11248) );
  AOI21_X1 U8496 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13733) );
  NAND2_X1 U8497 ( .A1(n7471), .A2(n9200), .ZN(n9194) );
  OAI21_X1 U8498 ( .B1(n13787), .B2(n13785), .A(n13786), .ZN(n13784) );
  AOI21_X1 U8499 ( .B1(n14290), .B2(n10152), .A(n10151), .ZN(n10155) );
  AOI21_X1 U8500 ( .B1(n7368), .B2(n7375), .A(n6658), .ZN(n7367) );
  INV_X1 U8501 ( .A(n6895), .ZN(n6894) );
  INV_X1 U8502 ( .A(n11804), .ZN(n6900) );
  NAND2_X1 U8503 ( .A1(n13851), .A2(n13841), .ZN(n13840) );
  NOR2_X1 U8504 ( .A1(n6896), .A2(n13845), .ZN(n6895) );
  INV_X1 U8505 ( .A(n7165), .ZN(n6896) );
  INV_X1 U8506 ( .A(n7086), .ZN(n13880) );
  NAND2_X1 U8507 ( .A1(n7401), .A2(n7399), .ZN(n13898) );
  OAI22_X1 U8508 ( .A1(n13911), .A2(n7406), .B1(n13674), .B2(n14065), .ZN(
        n7400) );
  NAND2_X1 U8509 ( .A1(n7088), .A2(n7087), .ZN(n13901) );
  AOI21_X1 U8510 ( .B1(n7162), .B2(n7164), .A(n6647), .ZN(n7160) );
  INV_X1 U8511 ( .A(n7088), .ZN(n13914) );
  AND2_X1 U8512 ( .A1(n11705), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11715) );
  AND2_X1 U8513 ( .A1(n11715), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11717) );
  OR2_X1 U8514 ( .A1(n13958), .A2(n11711), .ZN(n7381) );
  AND2_X1 U8515 ( .A1(n11714), .A2(n11713), .ZN(n13962) );
  INV_X1 U8516 ( .A(n7090), .ZN(n11260) );
  INV_X1 U8517 ( .A(n7092), .ZN(n14278) );
  OR2_X1 U8518 ( .A1(n10634), .A2(n10950), .ZN(n10697) );
  AND2_X1 U8519 ( .A1(n10693), .A2(n10627), .ZN(n13425) );
  NAND2_X1 U8520 ( .A1(n7081), .A2(n14554), .ZN(n10645) );
  NOR2_X1 U8521 ( .A1(n10516), .A2(n10515), .ZN(n10528) );
  NAND2_X1 U8522 ( .A1(n10510), .A2(n10509), .ZN(n10620) );
  NAND2_X1 U8523 ( .A1(n14554), .A2(n10538), .ZN(n14555) );
  NAND2_X1 U8524 ( .A1(n10384), .A2(n10383), .ZN(n10522) );
  NAND2_X1 U8525 ( .A1(n7150), .A2(n10272), .ZN(n10379) );
  XNOR2_X1 U8526 ( .A(n14603), .B(n13490), .ZN(n13419) );
  OR2_X1 U8527 ( .A1(n11910), .A2(n9459), .ZN(n10273) );
  NAND2_X1 U8528 ( .A1(n9463), .A2(n10265), .ZN(n13468) );
  OR2_X1 U8529 ( .A1(n13931), .A2(n14550), .ZN(n14074) );
  NAND2_X1 U8530 ( .A1(n13945), .A2(n7408), .ZN(n13929) );
  XNOR2_X1 U8531 ( .A(n9168), .B(n9153), .ZN(n10361) );
  XNOR2_X1 U8532 ( .A(n9025), .B(n9024), .ZN(n13445) );
  OAI21_X1 U8533 ( .B1(n9017), .B2(n7292), .A(n7289), .ZN(n9025) );
  AOI21_X1 U8534 ( .B1(n7278), .B2(n7276), .A(n6718), .ZN(n7275) );
  INV_X1 U8535 ( .A(n7281), .ZN(n7276) );
  OR2_X1 U8536 ( .A1(n8075), .A2(n7277), .ZN(n7274) );
  INV_X1 U8537 ( .A(n7278), .ZN(n7277) );
  XNOR2_X1 U8538 ( .A(n8078), .B(n8077), .ZN(n13265) );
  NAND2_X1 U8539 ( .A1(n6954), .A2(n7280), .ZN(n8078) );
  INV_X1 U8540 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9152) );
  INV_X1 U8541 ( .A(n9435), .ZN(n9439) );
  OAI21_X1 U8542 ( .B1(n7623), .B2(n7273), .A(n7271), .ZN(n7924) );
  NAND2_X1 U8543 ( .A1(n7623), .A2(n7622), .ZN(n7639) );
  NAND2_X1 U8544 ( .A1(n7823), .A2(n7606), .ZN(n7845) );
  NAND2_X1 U8545 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U8546 ( .A1(n7735), .A2(n7736), .ZN(n7738) );
  NAND2_X1 U8547 ( .A1(n7724), .A2(n7589), .ZN(n7736) );
  NAND2_X1 U8548 ( .A1(n7722), .A2(n7721), .ZN(n7724) );
  OAI21_X1 U8549 ( .B1(n7631), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6850), .ZN(
        n7581) );
  NAND2_X1 U8550 ( .A1(n7631), .A2(n8252), .ZN(n6850) );
  NAND2_X1 U8551 ( .A1(n6737), .A2(n6735), .ZN(n14194) );
  NAND2_X1 U8552 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6736), .ZN(n6735) );
  XNOR2_X1 U8553 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14193) );
  NOR2_X1 U8554 ( .A1(n15289), .A2(n14204), .ZN(n14206) );
  NAND2_X1 U8555 ( .A1(n14162), .A2(n14161), .ZN(n14212) );
  NOR2_X1 U8556 ( .A1(n14253), .A2(n14213), .ZN(n14215) );
  OAI21_X1 U8557 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14170), .A(n14169), .ZN(
        n14189) );
  NAND2_X1 U8558 ( .A1(n7208), .A2(n7207), .ZN(n14227) );
  NAND2_X1 U8559 ( .A1(n7209), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7208) );
  OAI21_X1 U8560 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14177), .A(n14176), .ZN(
        n14188) );
  XNOR2_X1 U8561 ( .A(n10830), .B(n11032), .ZN(n12030) );
  AOI22_X1 U8562 ( .A1(n12099), .A2(n11972), .B1(n12359), .B2(n11971), .ZN(
        n12014) );
  AOI21_X1 U8563 ( .B1(n7179), .B2(n7183), .A(n6657), .ZN(n7178) );
  NAND2_X1 U8564 ( .A1(n10085), .A2(n10043), .ZN(n10084) );
  OR2_X1 U8565 ( .A1(n11975), .A2(n12131), .ZN(n7174) );
  NAND2_X1 U8566 ( .A1(n6991), .A2(n6989), .ZN(n11228) );
  INV_X1 U8567 ( .A(n6992), .ZN(n6989) );
  AND4_X1 U8568 ( .A1(n8519), .A2(n8518), .A3(n8517), .A4(n8516), .ZN(n12398)
         );
  INV_X1 U8569 ( .A(n6973), .ZN(n12061) );
  AOI21_X1 U8570 ( .B1(n12000), .B2(n6974), .A(n6977), .ZN(n6973) );
  INV_X1 U8571 ( .A(n6979), .ZN(n6974) );
  OAI21_X1 U8572 ( .B1(n12000), .B2(n6977), .A(n6975), .ZN(n12059) );
  OAI21_X1 U8573 ( .B1(n6970), .B2(n6972), .A(n6971), .ZN(n12068) );
  AOI21_X1 U8574 ( .B1(n6975), .B2(n6977), .A(n6671), .ZN(n6971) );
  NAND2_X1 U8575 ( .A1(n11984), .A2(n6744), .ZN(n12074) );
  NAND2_X1 U8576 ( .A1(n11983), .A2(n6745), .ZN(n6744) );
  INV_X1 U8577 ( .A(n11985), .ZN(n6745) );
  AND2_X1 U8578 ( .A1(n10400), .A2(n10399), .ZN(n10406) );
  NAND2_X1 U8579 ( .A1(n6608), .A2(n7193), .ZN(n6988) );
  NAND2_X1 U8580 ( .A1(n11281), .A2(n11280), .ZN(n11962) );
  AOI21_X1 U8581 ( .B1(n7194), .B2(n6575), .A(n7195), .ZN(n11227) );
  AND3_X1 U8582 ( .A1(n8443), .A2(n8442), .A3(n8441), .ZN(n11105) );
  AND4_X1 U8583 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n12370)
         );
  INV_X1 U8584 ( .A(n12118), .ZN(n12112) );
  OR2_X1 U8585 ( .A1(n11411), .A2(n11238), .ZN(n8692) );
  NAND2_X1 U8586 ( .A1(n9980), .A2(n12453), .ZN(n12120) );
  OAI21_X1 U8587 ( .B1(n12000), .B2(n11965), .A(n6982), .ZN(n12116) );
  NAND2_X1 U8588 ( .A1(n9971), .A2(n9970), .ZN(n12124) );
  NAND2_X1 U8589 ( .A1(n9975), .A2(n9982), .ZN(n12126) );
  INV_X1 U8590 ( .A(n11622), .ZN(n6795) );
  AOI21_X1 U8591 ( .B1(n12249), .B2(n8312), .A(n8730), .ZN(n12261) );
  INV_X1 U8592 ( .A(n12360), .ZN(n12131) );
  INV_X1 U8593 ( .A(n12370), .ZN(n12346) );
  INV_X1 U8594 ( .A(n12397), .ZN(n12132) );
  INV_X1 U8595 ( .A(n12398), .ZN(n12423) );
  AND2_X1 U8596 ( .A1(n9817), .A2(n9793), .ZN(n9794) );
  NAND2_X1 U8597 ( .A1(n7025), .A2(n9817), .ZN(n9818) );
  INV_X1 U8598 ( .A(n6787), .ZN(n10484) );
  INV_X1 U8599 ( .A(n7024), .ZN(n12175) );
  INV_X1 U8600 ( .A(n7013), .ZN(n14338) );
  XNOR2_X1 U8601 ( .A(n12186), .B(n12210), .ZN(n14345) );
  INV_X1 U8602 ( .A(n6852), .ZN(n14344) );
  INV_X1 U8603 ( .A(n11415), .ZN(n14364) );
  XNOR2_X1 U8604 ( .A(n11391), .B(n11582), .ZN(n11957) );
  INV_X1 U8605 ( .A(n6833), .ZN(n6832) );
  XNOR2_X1 U8606 ( .A(n12275), .B(n12272), .ZN(n6834) );
  OAI22_X1 U8607 ( .A1(n12273), .A2(n14943), .B1(n14941), .B2(n12274), .ZN(
        n6833) );
  AOI21_X1 U8608 ( .B1(n12284), .B2(n6822), .A(n6821), .ZN(n12489) );
  INV_X1 U8609 ( .A(n12286), .ZN(n6821) );
  AOI21_X1 U8610 ( .B1(n6769), .B2(n12450), .A(n6766), .ZN(n12494) );
  NAND2_X1 U8611 ( .A1(n6768), .A2(n6767), .ZN(n6766) );
  NAND2_X1 U8612 ( .A1(n12297), .A2(n12456), .ZN(n6767) );
  NAND2_X1 U8613 ( .A1(n8650), .A2(n8649), .ZN(n12496) );
  NAND2_X1 U8614 ( .A1(n12348), .A2(n11534), .ZN(n12336) );
  NAND2_X1 U8615 ( .A1(n7038), .A2(n11524), .ZN(n12375) );
  NAND2_X1 U8616 ( .A1(n12392), .A2(n12391), .ZN(n7038) );
  AND2_X1 U8617 ( .A1(n12387), .A2(n12386), .ZN(n12523) );
  NAND2_X1 U8618 ( .A1(n11195), .A2(n11470), .ZN(n11045) );
  INV_X1 U8619 ( .A(n12470), .ZN(n12428) );
  NAND2_X1 U8620 ( .A1(n10287), .A2(n8309), .ZN(n10743) );
  INV_X1 U8621 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U8622 ( .A1(n9982), .A2(n9981), .ZN(n14934) );
  INV_X1 U8623 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U8624 ( .A1(n8593), .A2(n8592), .ZN(n12572) );
  NAND2_X1 U8625 ( .A1(n8553), .A2(n8552), .ZN(n12579) );
  INV_X1 U8626 ( .A(n11961), .ZN(n12584) );
  AND2_X1 U8627 ( .A1(n8494), .A2(n8493), .ZN(n12592) );
  NAND2_X1 U8628 ( .A1(n8477), .A2(n8476), .ZN(n12596) );
  AND3_X1 U8629 ( .A1(n8349), .A2(n8348), .A3(n8347), .ZN(n10855) );
  NAND2_X1 U8630 ( .A1(n8782), .A2(n8781), .ZN(n10283) );
  INV_X1 U8631 ( .A(n7441), .ZN(n7439) );
  NAND2_X1 U8632 ( .A1(n7073), .A2(n8634), .ZN(n8648) );
  NAND2_X1 U8633 ( .A1(n7074), .A2(n8631), .ZN(n7073) );
  INV_X1 U8634 ( .A(n8633), .ZN(n7074) );
  XNOR2_X1 U8635 ( .A(n8735), .B(n8734), .ZN(n11433) );
  INV_X1 U8636 ( .A(SI_19_), .ZN(n9717) );
  OAI21_X1 U8637 ( .B1(n8504), .B2(n7060), .A(n7057), .ZN(n8527) );
  NAND2_X1 U8638 ( .A1(n8507), .A2(n8506), .ZN(n8524) );
  NAND2_X1 U8639 ( .A1(n8504), .A2(n8503), .ZN(n8507) );
  INV_X1 U8640 ( .A(SI_13_), .ZN(n9328) );
  INV_X1 U8641 ( .A(SI_11_), .ZN(n9290) );
  INV_X1 U8642 ( .A(SI_10_), .ZN(n9285) );
  INV_X1 U8643 ( .A(n10309), .ZN(n10315) );
  OAI21_X1 U8644 ( .B1(n6750), .B2(n8363), .A(n8365), .ZN(n8377) );
  INV_X1 U8645 ( .A(n9926), .ZN(n9934) );
  XNOR2_X1 U8646 ( .A(n8302), .B(P3_IR_REG_4__SCAN_IN), .ZN(n9836) );
  XNOR2_X1 U8647 ( .A(n8266), .B(n8265), .ZN(n9601) );
  OR2_X1 U8648 ( .A1(n14382), .A2(n14381), .ZN(n14384) );
  NAND2_X1 U8649 ( .A1(n10763), .A2(n10762), .ZN(n10844) );
  NAND2_X1 U8650 ( .A1(n12757), .A2(n12756), .ZN(n12755) );
  AOI21_X1 U8651 ( .B1(n12786), .B2(n7341), .A(n7339), .ZN(n12648) );
  INV_X1 U8652 ( .A(n7340), .ZN(n7339) );
  AOI21_X1 U8653 ( .B1(n7341), .B2(n12785), .A(n12692), .ZN(n7340) );
  AND2_X1 U8654 ( .A1(n7343), .A2(n7341), .ZN(n12767) );
  OR2_X1 U8655 ( .A1(n12653), .A2(n10011), .ZN(n7318) );
  NAND2_X1 U8656 ( .A1(n10010), .A2(n7349), .ZN(n10188) );
  NAND2_X1 U8657 ( .A1(n10010), .A2(n10009), .ZN(n10017) );
  AND2_X1 U8658 ( .A1(n7360), .A2(n7358), .ZN(n12808) );
  NAND2_X1 U8659 ( .A1(n7360), .A2(n7361), .ZN(n12798) );
  INV_X1 U8660 ( .A(n11288), .ZN(n9136) );
  AND2_X1 U8661 ( .A1(n7510), .A2(n9098), .ZN(n6867) );
  NAND2_X1 U8662 ( .A1(n6866), .A2(n9097), .ZN(n6865) );
  NAND2_X1 U8663 ( .A1(n8072), .A2(n8071), .ZN(n12826) );
  NAND2_X1 U8664 ( .A1(n7681), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7683) );
  OR2_X1 U8665 ( .A1(n7689), .A2(n7688), .ZN(n7694) );
  OR2_X1 U8666 ( .A1(n7690), .A2(n9181), .ZN(n7693) );
  INV_X1 U8667 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n11652) );
  INV_X1 U8668 ( .A(n9066), .ZN(n13134) );
  INV_X1 U8669 ( .A(n12956), .ZN(n13137) );
  NAND2_X1 U8670 ( .A1(n8061), .A2(n8060), .ZN(n12991) );
  NAND2_X1 U8671 ( .A1(n8050), .A2(n8049), .ZN(n13002) );
  NAND2_X1 U8672 ( .A1(n6938), .A2(n6550), .ZN(n13044) );
  OR2_X1 U8673 ( .A1(n7316), .A2(n6943), .ZN(n6938) );
  NAND2_X1 U8674 ( .A1(n6944), .A2(n6948), .ZN(n13061) );
  NAND2_X1 U8675 ( .A1(n7316), .A2(n6949), .ZN(n6944) );
  AOI21_X1 U8676 ( .B1(n7316), .B2(n7315), .A(n6571), .ZN(n13072) );
  NAND2_X1 U8677 ( .A1(n7313), .A2(n7920), .ZN(n11365) );
  NAND2_X1 U8678 ( .A1(n7107), .A2(n7108), .ZN(n11207) );
  NAND2_X1 U8679 ( .A1(n11158), .A2(n7884), .ZN(n11217) );
  OAI21_X1 U8680 ( .B1(n10973), .B2(n8194), .A(n7115), .ZN(n11017) );
  NAND2_X1 U8681 ( .A1(n10812), .A2(n7842), .ZN(n10974) );
  AND2_X1 U8682 ( .A1(n10666), .A2(n7820), .ZN(n10814) );
  NAND2_X1 U8683 ( .A1(n10543), .A2(n8190), .ZN(n10674) );
  NAND2_X1 U8684 ( .A1(n8187), .A2(n8186), .ZN(n10055) );
  INV_X1 U8685 ( .A(n14731), .ZN(n13129) );
  NAND2_X1 U8686 ( .A1(n9948), .A2(n7744), .ZN(n10054) );
  NAND2_X1 U8687 ( .A1(n6558), .A2(n9426), .ZN(n14739) );
  OR2_X1 U8688 ( .A1(n9173), .A2(n12857), .ZN(n7137) );
  NAND2_X1 U8689 ( .A1(n9173), .A2(n7136), .ZN(n7135) );
  INV_X1 U8690 ( .A(n14739), .ZN(n14393) );
  OR2_X1 U8691 ( .A1(n9422), .A2(n8167), .ZN(n14764) );
  INV_X1 U8692 ( .A(n9130), .ZN(n11220) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11043) );
  INV_X1 U8694 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10228) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15273) );
  INV_X1 U8696 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10415) );
  INV_X1 U8697 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10101) );
  INV_X1 U8698 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9623) );
  INV_X1 U8699 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9331) );
  AND2_X1 U8700 ( .A1(n7830), .A2(n7846), .ZN(n14702) );
  INV_X1 U8701 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9281) );
  INV_X1 U8702 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9277) );
  INV_X1 U8703 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9261) );
  INV_X1 U8704 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9256) );
  INV_X1 U8705 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9253) );
  INV_X1 U8706 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9255) );
  AOI21_X1 U8707 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(n10587) );
  AOI22_X1 U8708 ( .A1(n10344), .A2(n10343), .B1(n10342), .B2(n10341), .ZN(
        n13294) );
  INV_X1 U8709 ( .A(n7475), .ZN(n7474) );
  AOI21_X1 U8710 ( .B1(n7475), .B2(n7473), .A(n6654), .ZN(n7472) );
  INV_X1 U8711 ( .A(n7478), .ZN(n7473) );
  NOR2_X1 U8712 ( .A1(n11945), .A2(n7451), .ZN(n7448) );
  OAI22_X1 U8713 ( .A1(n7451), .A2(n7450), .B1(n11945), .B2(n7453), .ZN(n7449)
         );
  NOR2_X1 U8714 ( .A1(n13278), .A2(n11945), .ZN(n7450) );
  INV_X1 U8715 ( .A(n11945), .ZN(n7452) );
  INV_X1 U8716 ( .A(n6824), .ZN(n9671) );
  NAND2_X1 U8717 ( .A1(n7467), .A2(n11874), .ZN(n13309) );
  AND2_X1 U8718 ( .A1(n11350), .A2(n7485), .ZN(n7481) );
  NAND2_X1 U8719 ( .A1(n11655), .A2(n11654), .ZN(n14051) );
  NAND2_X1 U8720 ( .A1(n13327), .A2(n7480), .ZN(n13340) );
  NAND2_X1 U8721 ( .A1(n13285), .A2(n13286), .ZN(n13284) );
  INV_X1 U8722 ( .A(n14603), .ZN(n13491) );
  AND2_X1 U8723 ( .A1(n10947), .A2(n7490), .ZN(n7486) );
  AND2_X1 U8724 ( .A1(n7487), .A2(n7490), .ZN(n10948) );
  NAND2_X1 U8725 ( .A1(n14441), .A2(n11341), .ZN(n14454) );
  INV_X1 U8726 ( .A(n7482), .ZN(n14453) );
  NAND2_X1 U8727 ( .A1(n7477), .A2(n7535), .ZN(n13385) );
  INV_X1 U8728 ( .A(n13387), .ZN(n13662) );
  AOI21_X1 U8729 ( .B1(n13659), .B2(n13660), .A(n6786), .ZN(n6785) );
  NAND4_X1 U8730 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n13691) );
  NOR2_X1 U8731 ( .A1(n9229), .A2(n9228), .ZN(n13773) );
  OR2_X1 U8732 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  AOI21_X1 U8733 ( .B1(n10879), .B2(n14537), .A(n14529), .ZN(n10881) );
  INV_X1 U8734 ( .A(n13646), .ZN(n14022) );
  INV_X1 U8735 ( .A(n13824), .ZN(n14025) );
  NAND2_X1 U8736 ( .A1(n6897), .A2(n7165), .ZN(n13844) );
  OAI21_X1 U8737 ( .B1(n13878), .B2(n7375), .A(n7372), .ZN(n13836) );
  NAND2_X1 U8738 ( .A1(n7168), .A2(n7169), .ZN(n13856) );
  OR2_X1 U8739 ( .A1(n13874), .A2(n13873), .ZN(n14048) );
  NAND2_X1 U8740 ( .A1(n13925), .A2(n11797), .ZN(n13912) );
  AND2_X1 U8741 ( .A1(n7406), .A2(n7407), .ZN(n13910) );
  INV_X1 U8742 ( .A(n13944), .ZN(n13933) );
  NAND2_X1 U8743 ( .A1(n11687), .A2(n11686), .ZN(n13954) );
  NAND2_X1 U8744 ( .A1(n6885), .A2(n7152), .ZN(n13943) );
  OAI21_X1 U8745 ( .B1(n14004), .B2(n11793), .A(n6887), .ZN(n6885) );
  INV_X1 U8746 ( .A(n13962), .ZN(n14083) );
  NAND2_X1 U8747 ( .A1(n7156), .A2(n7155), .ZN(n13957) );
  NAND2_X1 U8748 ( .A1(n11795), .A2(n6602), .ZN(n7156) );
  NAND2_X1 U8749 ( .A1(n13989), .A2(n13563), .ZN(n13973) );
  NAND2_X1 U8750 ( .A1(n11795), .A2(n11794), .ZN(n13971) );
  NAND2_X1 U8751 ( .A1(n6890), .A2(n11792), .ZN(n13988) );
  INV_X1 U8752 ( .A(n6891), .ZN(n6890) );
  NAND2_X1 U8753 ( .A1(n7384), .A2(n7388), .ZN(n14005) );
  NAND2_X1 U8754 ( .A1(n11294), .A2(n7389), .ZN(n7384) );
  NAND2_X1 U8755 ( .A1(n7391), .A2(n13549), .ZN(n11295) );
  OR2_X1 U8756 ( .A1(n11294), .A2(n13433), .ZN(n7391) );
  NAND2_X1 U8757 ( .A1(n11256), .A2(n6903), .ZN(n11310) );
  NAND2_X1 U8758 ( .A1(n11256), .A2(n11255), .ZN(n11257) );
  NAND2_X1 U8759 ( .A1(n11058), .A2(n11057), .ZN(n14274) );
  NAND2_X1 U8760 ( .A1(n6877), .A2(n10912), .ZN(n11054) );
  NAND2_X1 U8761 ( .A1(n10959), .A2(n13428), .ZN(n6877) );
  NAND2_X1 U8762 ( .A1(n10916), .A2(n10915), .ZN(n14450) );
  NAND2_X1 U8763 ( .A1(n10694), .A2(n7396), .ZN(n10923) );
  INV_X1 U8764 ( .A(n14581), .ZN(n14016) );
  NAND2_X1 U8765 ( .A1(n11671), .A2(n7398), .ZN(n9546) );
  NOR2_X1 U8766 ( .A1(n9251), .A2(n7263), .ZN(n7398) );
  NAND2_X1 U8767 ( .A1(n10231), .A2(n10230), .ZN(n14010) );
  AND2_X2 U8768 ( .A1(n9564), .A2(n9563), .ZN(n14679) );
  NAND2_X1 U8769 ( .A1(n6811), .A2(n6809), .ZN(n14117) );
  INV_X1 U8770 ( .A(n6810), .ZN(n6809) );
  NAND2_X1 U8771 ( .A1(n14021), .A2(n14577), .ZN(n6811) );
  OAI21_X1 U8772 ( .B1(n14022), .B2(n14655), .A(n14023), .ZN(n6810) );
  NOR3_X1 U8773 ( .A1(n14027), .A2(n14028), .A3(n6631), .ZN(n14030) );
  OR2_X1 U8774 ( .A1(n14026), .A2(n14639), .ZN(n14031) );
  AND3_X2 U8775 ( .A1(n9563), .A2(n11783), .A3(n9672), .ZN(n14663) );
  INV_X1 U8776 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8777 ( .A1(n9071), .A2(n9070), .ZN(n13454) );
  NAND2_X1 U8778 ( .A1(n7295), .A2(n7293), .ZN(n9071) );
  INV_X1 U8779 ( .A(n9399), .ZN(n14139) );
  XNOR2_X1 U8780 ( .A(n8109), .B(n8108), .ZN(n13261) );
  NAND2_X1 U8781 ( .A1(n7274), .A2(n7275), .ZN(n8109) );
  XNOR2_X1 U8782 ( .A(n9161), .B(n9160), .ZN(n14149) );
  OR2_X1 U8783 ( .A1(n11669), .A2(n9020), .ZN(n11670) );
  CLKBUF_X1 U8784 ( .A(n14151), .Z(n6847) );
  INV_X1 U8785 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10772) );
  INV_X1 U8786 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10096) );
  INV_X1 U8787 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10338) );
  INV_X1 U8788 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10106) );
  INV_X1 U8789 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9644) );
  INV_X1 U8790 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9543) );
  OR2_X1 U8791 ( .A1(n9484), .A2(n9483), .ZN(n9636) );
  INV_X1 U8792 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9389) );
  INV_X1 U8793 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n15110) );
  INV_X1 U8794 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9315) );
  INV_X1 U8795 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9298) );
  INV_X1 U8796 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9282) );
  OR2_X1 U8797 ( .A1(n9218), .A2(n9217), .ZN(n10504) );
  NAND2_X1 U8798 ( .A1(n7745), .A2(n7746), .ZN(n7748) );
  AOI21_X1 U8799 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14202), .A(n15299), .ZN(
        n15291) );
  NOR2_X1 U8800 ( .A1(n14255), .A2(n14254), .ZN(n14253) );
  INV_X1 U8801 ( .A(n14221), .ZN(n7212) );
  NOR2_X1 U8802 ( .A1(n14227), .A2(n14228), .ZN(n14494) );
  NAND2_X1 U8803 ( .A1(n14493), .A2(n14495), .ZN(n14499) );
  INV_X1 U8804 ( .A(n14233), .ZN(n7211) );
  INV_X1 U8805 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6840) );
  NOR2_X2 U8806 ( .A1(n9963), .A2(n9169), .ZN(P3_U3897) );
  OR2_X1 U8807 ( .A1(n11621), .A2(n11620), .ZN(n6793) );
  AND2_X1 U8808 ( .A1(n12218), .A2(n6791), .ZN(n6790) );
  OR2_X1 U8809 ( .A1(n12219), .A2(n14882), .ZN(n6791) );
  NAND2_X1 U8810 ( .A1(n14843), .A2(n7006), .ZN(n7004) );
  AOI211_X1 U8811 ( .C1(n12240), .C2(n14903), .A(n12239), .B(n12238), .ZN(
        n12241) );
  OAI21_X1 U8812 ( .B1(n11960), .B2(n14949), .A(n6770), .ZN(P3_U3204) );
  INV_X1 U8813 ( .A(n6771), .ZN(n6770) );
  OAI21_X1 U8814 ( .B1(n11957), .B2(n12431), .A(n7051), .ZN(n6771) );
  AOI21_X1 U8815 ( .B1(n11959), .B2(n12470), .A(n11958), .ZN(n7051) );
  OAI21_X1 U8816 ( .B1(n8839), .B2(n12544), .A(n8838), .ZN(n8840) );
  NOR2_X1 U8817 ( .A1(n6630), .A2(n6814), .ZN(n6813) );
  OAI21_X1 U8818 ( .B1(n12548), .B2(n14986), .A(n6801), .ZN(P3_U3486) );
  INV_X1 U8819 ( .A(n6802), .ZN(n6801) );
  OAI21_X1 U8820 ( .B1(n12550), .B2(n12544), .A(n6803), .ZN(n6802) );
  OR2_X1 U8821 ( .A1(n14989), .A2(n12481), .ZN(n6803) );
  AOI21_X1 U8822 ( .B1(n11959), .B2(n8834), .A(n8833), .ZN(n8835) );
  NOR2_X1 U8823 ( .A1(n6629), .A2(n6818), .ZN(n6817) );
  NOR2_X1 U8824 ( .A1(n14979), .A2(n15211), .ZN(n6818) );
  INV_X1 U8825 ( .A(n6836), .ZN(n6835) );
  OAI21_X1 U8826 ( .B1(n12550), .B2(n12597), .A(n6837), .ZN(n6836) );
  OAI21_X1 U8827 ( .B1(n10449), .B2(n7332), .A(n7330), .ZN(n10755) );
  NAND2_X1 U8828 ( .A1(n8856), .A2(n7541), .ZN(P2_U3237) );
  AOI21_X1 U8829 ( .B1(n13146), .B2(n8847), .A(n14736), .ZN(n8848) );
  NAND2_X1 U8830 ( .A1(n7133), .A2(n6721), .ZN(P2_U3496) );
  NAND2_X1 U8831 ( .A1(n13235), .A2(n14814), .ZN(n7133) );
  NAND2_X1 U8832 ( .A1(n13366), .A2(n7463), .ZN(n14430) );
  NAND2_X1 U8833 ( .A1(n6781), .A2(n6776), .ZN(n13823) );
  NAND2_X1 U8834 ( .A1(n6780), .A2(n6777), .ZN(n6776) );
  INV_X1 U8835 ( .A(n11806), .ZN(n7173) );
  INV_X1 U8836 ( .A(n7207), .ZN(n14262) );
  INV_X1 U8837 ( .A(n14294), .ZN(n14293) );
  INV_X1 U8838 ( .A(n14301), .ZN(n6742) );
  XNOR2_X1 U8839 ( .A(n14304), .B(n7217), .ZN(n7216) );
  XNOR2_X1 U8840 ( .A(n14303), .B(n14305), .ZN(n7217) );
  OAI21_X1 U8841 ( .B1(n11418), .B2(n12243), .A(n11414), .ZN(n11608) );
  INV_X1 U8842 ( .A(n11608), .ZN(n7079) );
  AND2_X1 U8843 ( .A1(n13206), .A2(n12750), .ZN(n6571) );
  OR2_X1 U8844 ( .A1(n14380), .A2(n13228), .ZN(n6572) );
  NOR2_X1 U8845 ( .A1(n11415), .A2(n11417), .ZN(n11607) );
  OR2_X1 U8846 ( .A1(n6634), .A2(n7028), .ZN(n6573) );
  OR2_X1 U8847 ( .A1(n8016), .A2(n7988), .ZN(n6574) );
  INV_X1 U8848 ( .A(n13228), .ZN(n7146) );
  INV_X2 U8849 ( .A(n8902), .ZN(n8999) );
  AND2_X1 U8850 ( .A1(n7198), .A2(n7199), .ZN(n6575) );
  INV_X1 U8851 ( .A(n12436), .ZN(n12409) );
  INV_X1 U8852 ( .A(n10560), .ZN(n6752) );
  AND2_X1 U8853 ( .A1(n8766), .A2(n8793), .ZN(n6576) );
  OR2_X1 U8854 ( .A1(n7166), .A2(n7377), .ZN(n6577) );
  NAND2_X1 U8855 ( .A1(n11279), .A2(n11318), .ZN(n7193) );
  AND3_X1 U8856 ( .A1(n8230), .A2(n8233), .A3(n7050), .ZN(n6578) );
  NAND2_X1 U8857 ( .A1(n7921), .A2(n7146), .ZN(n7145) );
  NOR2_X1 U8858 ( .A1(n12277), .A2(n12285), .ZN(n6579) );
  NAND4_X1 U8859 ( .A1(n9554), .A2(n9553), .A3(n9552), .A4(n9551), .ZN(n13694)
         );
  AND2_X1 U8860 ( .A1(n7421), .A2(n7419), .ZN(n6581) );
  AND2_X1 U8861 ( .A1(n10060), .A2(n12847), .ZN(n6582) );
  AND2_X1 U8862 ( .A1(n11517), .A2(n11524), .ZN(n12391) );
  INV_X1 U8863 ( .A(n12391), .ZN(n7034) );
  OR2_X1 U8864 ( .A1(n8884), .A2(n8883), .ZN(n6583) );
  AND2_X1 U8865 ( .A1(n7342), .A2(n12646), .ZN(n7341) );
  INV_X1 U8866 ( .A(n7183), .ZN(n7182) );
  NAND2_X1 U8867 ( .A1(n6595), .A2(n11992), .ZN(n7183) );
  OR2_X1 U8868 ( .A1(n11225), .A2(n11231), .ZN(n6584) );
  XNOR2_X1 U8869 ( .A(n8717), .B(n12257), .ZN(n12479) );
  INV_X1 U8870 ( .A(n12479), .ZN(n6773) );
  OR2_X1 U8871 ( .A1(n9010), .A2(n9009), .ZN(n6585) );
  OR2_X1 U8872 ( .A1(n13600), .A2(n13599), .ZN(n6586) );
  OAI21_X1 U8873 ( .B1(n7099), .B2(n7097), .A(n6670), .ZN(n7096) );
  AND2_X1 U8874 ( .A1(n7149), .A2(n7148), .ZN(n6587) );
  NOR2_X1 U8875 ( .A1(n13200), .A2(n12833), .ZN(n6588) );
  INV_X1 U8876 ( .A(n11582), .ZN(n7076) );
  AND2_X1 U8877 ( .A1(n7119), .A2(n7116), .ZN(n6589) );
  INV_X1 U8878 ( .A(n12384), .ZN(n12410) );
  AND2_X1 U8879 ( .A1(n8383), .A2(n8368), .ZN(n6590) );
  AND2_X1 U8880 ( .A1(n7018), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8881 ( .A1(n11586), .A2(n7027), .ZN(n6592) );
  INV_X1 U8882 ( .A(n11144), .ZN(n6754) );
  INV_X2 U8883 ( .A(n9654), .ZN(n11884) );
  INV_X1 U8884 ( .A(n7988), .ZN(n7989) );
  AND2_X1 U8885 ( .A1(n15202), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6593) );
  AND2_X1 U8886 ( .A1(n9593), .A2(n9592), .ZN(n14843) );
  INV_X2 U8887 ( .A(n6620), .ZN(n13596) );
  AND2_X1 U8888 ( .A1(n8410), .A2(n8228), .ZN(n8413) );
  OR2_X1 U8889 ( .A1(n11993), .A2(n12285), .ZN(n6595) );
  OR2_X1 U8890 ( .A1(n14007), .A2(n14094), .ZN(n6596) );
  NAND2_X1 U8891 ( .A1(n7929), .A2(n7928), .ZN(n13213) );
  AND2_X1 U8892 ( .A1(n7682), .A2(n7684), .ZN(n6597) );
  INV_X1 U8893 ( .A(n13670), .ZN(n6969) );
  NAND2_X1 U8894 ( .A1(n7137), .A2(n7135), .ZN(n8869) );
  XNOR2_X1 U8895 ( .A(n13139), .B(n8118), .ZN(n9122) );
  INV_X1 U8896 ( .A(n9122), .ZN(n7124) );
  NAND2_X1 U8897 ( .A1(n9141), .A2(n9200), .ZN(n9202) );
  OR2_X1 U8898 ( .A1(n10355), .A2(n10354), .ZN(n6598) );
  AND2_X1 U8899 ( .A1(n7477), .A2(n7475), .ZN(n6599) );
  AND2_X1 U8900 ( .A1(n6799), .A2(n6798), .ZN(n6600) );
  AND2_X1 U8901 ( .A1(n8263), .A2(n8260), .ZN(n6601) );
  NOR2_X1 U8902 ( .A1(n13047), .A2(n13179), .ZN(n7139) );
  INV_X1 U8903 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8768) );
  NOR2_X1 U8904 ( .A1(n13566), .A2(n7157), .ZN(n6602) );
  NAND2_X1 U8905 ( .A1(n12492), .A2(n12309), .ZN(n6603) );
  OR2_X1 U8906 ( .A1(n8326), .A2(n8325), .ZN(n9837) );
  OR2_X1 U8907 ( .A1(n8873), .A2(n8872), .ZN(n6604) );
  AND2_X1 U8908 ( .A1(n13053), .A2(n12777), .ZN(n6605) );
  NAND2_X1 U8909 ( .A1(n6897), .A2(n6895), .ZN(n6606) );
  NAND2_X1 U8910 ( .A1(n11966), .A2(n12398), .ZN(n6607) );
  AND2_X1 U8911 ( .A1(n6993), .A2(n6575), .ZN(n6608) );
  AND2_X1 U8912 ( .A1(n8897), .A2(n8896), .ZN(n6609) );
  AND2_X1 U8913 ( .A1(n8912), .A2(n8911), .ZN(n6610) );
  AND2_X1 U8914 ( .A1(n7631), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6611) );
  INV_X1 U8915 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9395) );
  AND2_X1 U8916 ( .A1(n10813), .A2(n7820), .ZN(n6613) );
  INV_X1 U8917 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15116) );
  OR2_X1 U8918 ( .A1(n9579), .A2(n9805), .ZN(n6614) );
  INV_X1 U8919 ( .A(n13696), .ZN(n7412) );
  OR2_X1 U8920 ( .A1(n13886), .A2(n13672), .ZN(n6615) );
  INV_X1 U8921 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n15270) );
  OR2_X1 U8922 ( .A1(n7626), .A2(SI_17_), .ZN(n6617) );
  INV_X1 U8923 ( .A(n11511), .ZN(n7032) );
  NOR2_X1 U8924 ( .A1(n13039), .A2(n7105), .ZN(n6618) );
  INV_X1 U8925 ( .A(n10979), .ZN(n7148) );
  INV_X1 U8926 ( .A(n13278), .ZN(n7454) );
  NAND2_X1 U8927 ( .A1(n7646), .A2(n7645), .ZN(n13219) );
  NAND2_X1 U8928 ( .A1(n7980), .A2(n7979), .ZN(n13053) );
  OR2_X1 U8929 ( .A1(n9173), .A2(n9254), .ZN(n6619) );
  INV_X1 U8930 ( .A(n13025), .ZN(n7138) );
  AND2_X1 U8931 ( .A1(n12437), .A2(n11233), .ZN(n6621) );
  OR2_X1 U8932 ( .A1(n14094), .A2(n13678), .ZN(n6622) );
  AND4_X1 U8933 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n6623)
         );
  NOR2_X1 U8934 ( .A1(n8394), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8410) );
  OR2_X1 U8935 ( .A1(n10060), .A2(n12847), .ZN(n6624) );
  OR2_X1 U8936 ( .A1(n7148), .A2(n12842), .ZN(n6625) );
  OR2_X1 U8937 ( .A1(n13841), .A2(n13669), .ZN(n6626) );
  INV_X1 U8938 ( .A(n12303), .ZN(n6747) );
  INV_X1 U8939 ( .A(n13603), .ZN(n7241) );
  INV_X1 U8940 ( .A(n12785), .ZN(n7344) );
  XNOR2_X1 U8941 ( .A(n13149), .B(n12825), .ZN(n12976) );
  OR2_X1 U8942 ( .A1(n14410), .A2(n12839), .ZN(n6627) );
  INV_X1 U8943 ( .A(n8803), .ZN(n10202) );
  NAND2_X1 U8944 ( .A1(n11566), .A2(n11567), .ZN(n11563) );
  AND3_X1 U8945 ( .A1(n8359), .A2(n8357), .A3(n8360), .ZN(n6628) );
  NOR2_X1 U8946 ( .A1(n8811), .A2(n12597), .ZN(n6629) );
  NOR2_X1 U8947 ( .A1(n8811), .A2(n12544), .ZN(n6630) );
  INV_X1 U8948 ( .A(n7419), .ZN(n7418) );
  NOR2_X1 U8949 ( .A1(n12291), .A2(n7420), .ZN(n7419) );
  AND2_X1 U8950 ( .A1(n14029), .A2(n14636), .ZN(n6631) );
  OR2_X1 U8951 ( .A1(n6610), .A2(n8914), .ZN(n6632) );
  AND2_X1 U8952 ( .A1(n11101), .A2(n12133), .ZN(n6633) );
  AND2_X1 U8953 ( .A1(n11470), .A2(n7029), .ZN(n6634) );
  OR2_X1 U8954 ( .A1(n10483), .A2(n10482), .ZN(n6635) );
  OR2_X1 U8955 ( .A1(n12259), .A2(n8717), .ZN(n6636) );
  AND2_X1 U8956 ( .A1(n7098), .A2(n8209), .ZN(n6637) );
  INV_X1 U8957 ( .A(n14033), .ZN(n13841) );
  NAND2_X1 U8958 ( .A1(n11758), .A2(n11757), .ZN(n14033) );
  AND2_X1 U8959 ( .A1(n6624), .A2(n8186), .ZN(n6638) );
  AND2_X1 U8960 ( .A1(n8779), .A2(n10039), .ZN(n6639) );
  AND2_X1 U8961 ( .A1(n6610), .A2(n8914), .ZN(n6640) );
  NAND2_X1 U8962 ( .A1(n14689), .A2(n12840), .ZN(n6641) );
  AND2_X1 U8963 ( .A1(n13605), .A2(n13604), .ZN(n6642) );
  INV_X1 U8964 ( .A(n7130), .ZN(n8850) );
  NOR2_X1 U8965 ( .A1(n13144), .A2(n12970), .ZN(n7130) );
  OR2_X1 U8966 ( .A1(n8988), .A2(n8987), .ZN(n6643) );
  AND2_X1 U8967 ( .A1(n7609), .A2(n9290), .ZN(n6644) );
  AND2_X1 U8968 ( .A1(n11027), .A2(n12841), .ZN(n6645) );
  AND2_X1 U8969 ( .A1(n13514), .A2(n10945), .ZN(n6646) );
  INV_X1 U8970 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7629) );
  INV_X1 U8971 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8533) );
  NOR2_X1 U8972 ( .A1(n13919), .A2(n13674), .ZN(n6647) );
  NOR2_X1 U8973 ( .A1(n14450), .A2(n13685), .ZN(n6648) );
  NOR2_X1 U8974 ( .A1(n11837), .A2(n13681), .ZN(n6649) );
  NOR2_X1 U8975 ( .A1(n11833), .A2(n11832), .ZN(n6650) );
  NOR2_X1 U8976 ( .A1(n13962), .A2(n13573), .ZN(n6651) );
  AND2_X1 U8977 ( .A1(n12486), .A2(n12296), .ZN(n6652) );
  AND2_X1 U8978 ( .A1(n7524), .A2(n6698), .ZN(n6653) );
  INV_X1 U8979 ( .A(n7379), .ZN(n7378) );
  NAND2_X1 U8980 ( .A1(n7380), .A2(n6615), .ZN(n7379) );
  OR2_X1 U8981 ( .A1(n13299), .A2(n13300), .ZN(n6654) );
  INV_X1 U8982 ( .A(n7129), .ZN(n7128) );
  NAND2_X1 U8983 ( .A1(n13149), .A2(n12825), .ZN(n7129) );
  AND2_X1 U8984 ( .A1(n13855), .A2(n6969), .ZN(n6655) );
  INV_X1 U8985 ( .A(n7180), .ZN(n7179) );
  OR2_X1 U8986 ( .A1(n12020), .A2(n6681), .ZN(n7180) );
  AND2_X1 U8987 ( .A1(n6773), .A2(n14958), .ZN(n6656) );
  OAI21_X1 U8988 ( .B1(n7883), .B2(n7299), .A(n7901), .ZN(n7298) );
  INV_X1 U8989 ( .A(n7884), .ZN(n7299) );
  NOR2_X1 U8990 ( .A1(n12019), .A2(n12130), .ZN(n6657) );
  NOR2_X1 U8991 ( .A1(n14033), .A2(n11803), .ZN(n6658) );
  OR2_X1 U8992 ( .A1(n7469), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8993 ( .A1(n12277), .A2(n12285), .ZN(n6660) );
  OR2_X1 U8994 ( .A1(n10979), .A2(n9104), .ZN(n6661) );
  INV_X1 U8995 ( .A(n13439), .ZN(n13946) );
  NOR2_X1 U8996 ( .A1(n14689), .A2(n12840), .ZN(n6662) );
  INV_X1 U8997 ( .A(n7196), .ZN(n7195) );
  AOI21_X1 U8998 ( .B1(n6575), .B2(n7197), .A(n6633), .ZN(n7196) );
  AND2_X1 U8999 ( .A1(n9001), .A2(n9000), .ZN(n6663) );
  INV_X1 U9000 ( .A(n7314), .ZN(n6952) );
  AND2_X1 U9001 ( .A1(n13194), .A2(n8993), .ZN(n7314) );
  INV_X1 U9002 ( .A(n7126), .ZN(n7125) );
  OAI22_X1 U9003 ( .A1(n9119), .A2(n7129), .B1(n8212), .B2(n8852), .ZN(n7126)
         );
  NOR2_X1 U9004 ( .A1(n11688), .A2(n13680), .ZN(n6664) );
  INV_X1 U9005 ( .A(n7397), .ZN(n7396) );
  NAND2_X1 U9006 ( .A1(n13426), .A2(n10693), .ZN(n7397) );
  AND2_X1 U9007 ( .A1(n6905), .A2(n6625), .ZN(n6665) );
  AND2_X1 U9008 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n6666) );
  AND2_X1 U9009 ( .A1(n7626), .A2(SI_17_), .ZN(n6667) );
  AND2_X1 U9010 ( .A1(n9298), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6668) );
  NAND2_X1 U9011 ( .A1(n7376), .A2(n6577), .ZN(n7375) );
  INV_X1 U9012 ( .A(n7067), .ZN(n7066) );
  NAND2_X1 U9013 ( .A1(n8376), .A2(n7068), .ZN(n7067) );
  AND2_X1 U9014 ( .A1(n13497), .A2(n10523), .ZN(n6669) );
  NAND2_X1 U9015 ( .A1(n13162), .A2(n12795), .ZN(n6670) );
  AND2_X1 U9016 ( .A1(n11967), .A2(n12384), .ZN(n6671) );
  OR2_X1 U9017 ( .A1(n9004), .A2(n6663), .ZN(n6672) );
  AND2_X1 U9018 ( .A1(n7202), .A2(n6639), .ZN(n6673) );
  INV_X1 U9019 ( .A(n6889), .ZN(n6888) );
  AND2_X1 U9020 ( .A1(n6622), .A2(n11792), .ZN(n6889) );
  OR2_X1 U9021 ( .A1(n7607), .A2(n9285), .ZN(n6674) );
  NAND2_X1 U9022 ( .A1(n11982), .A2(n11981), .ZN(n11983) );
  NAND2_X1 U9023 ( .A1(n9103), .A2(n13014), .ZN(n6675) );
  OR2_X1 U9024 ( .A1(n13855), .A2(n13670), .ZN(n6676) );
  OR2_X1 U9025 ( .A1(n11027), .A2(n12841), .ZN(n6677) );
  OR2_X1 U9026 ( .A1(n12101), .A2(n12359), .ZN(n11516) );
  OR2_X1 U9027 ( .A1(n8887), .A2(n8888), .ZN(n6678) );
  AND2_X1 U9028 ( .A1(n13563), .A2(n13564), .ZN(n13990) );
  INV_X1 U9029 ( .A(n13990), .ZN(n7224) );
  AND2_X1 U9030 ( .A1(n7108), .A2(n6627), .ZN(n6679) );
  AND2_X1 U9031 ( .A1(n6898), .A2(n6900), .ZN(n6680) );
  AND2_X1 U9032 ( .A1(n7181), .A2(n6595), .ZN(n6681) );
  AND2_X1 U9033 ( .A1(n10754), .A2(n10753), .ZN(n6682) );
  AND2_X1 U9034 ( .A1(n12021), .A2(n7078), .ZN(n6683) );
  AND2_X1 U9035 ( .A1(n7271), .A2(n6617), .ZN(n6684) );
  INV_X1 U9036 ( .A(n13532), .ZN(n7236) );
  AND2_X1 U9037 ( .A1(n6572), .A2(n7545), .ZN(n6685) );
  AND2_X1 U9038 ( .A1(n12650), .A2(n12649), .ZN(n6686) );
  OR2_X1 U9039 ( .A1(n8922), .A2(n8923), .ZN(n6687) );
  AND2_X1 U9040 ( .A1(n7433), .A2(n15270), .ZN(n6688) );
  OR2_X1 U9041 ( .A1(n13602), .A2(n7241), .ZN(n6689) );
  OR2_X1 U9042 ( .A1(n7516), .A2(n7515), .ZN(n6690) );
  AND2_X1 U9043 ( .A1(n11969), .A2(n12132), .ZN(n6691) );
  NAND2_X1 U9044 ( .A1(n7245), .A2(n13622), .ZN(n6692) );
  NAND2_X1 U9045 ( .A1(n7864), .A2(n7863), .ZN(n11027) );
  AND2_X1 U9046 ( .A1(n12452), .A2(n8446), .ZN(n7436) );
  AND2_X1 U9047 ( .A1(n6672), .A2(n6861), .ZN(n6693) );
  OR2_X1 U9048 ( .A1(n7154), .A2(n6883), .ZN(n6694) );
  INV_X1 U9049 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U9050 ( .A1(n7113), .A2(n6641), .ZN(n7111) );
  AND2_X1 U9051 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n6695) );
  AND2_X1 U9052 ( .A1(n6908), .A2(n6907), .ZN(n7583) );
  INV_X1 U9053 ( .A(n7193), .ZN(n7192) );
  OR2_X1 U9054 ( .A1(n6862), .A2(n6653), .ZN(n6696) );
  INV_X1 U9055 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7354) );
  OR2_X1 U9056 ( .A1(n7454), .A2(n7452), .ZN(n6697) );
  INV_X2 U9057 ( .A(n11750), .ZN(n13449) );
  NAND2_X1 U9058 ( .A1(n11246), .A2(n11245), .ZN(n11837) );
  INV_X1 U9059 ( .A(n11837), .ZN(n7089) );
  NAND2_X1 U9060 ( .A1(n11663), .A2(n11662), .ZN(n13900) );
  INV_X1 U9061 ( .A(n13900), .ZN(n7087) );
  INV_X1 U9062 ( .A(n12764), .ZN(n7342) );
  NAND2_X1 U9063 ( .A1(n8080), .A2(n8079), .ZN(n13149) );
  INV_X1 U9064 ( .A(n13149), .ZN(n7131) );
  AND2_X1 U9065 ( .A1(n8997), .A2(n8996), .ZN(n6698) );
  NAND2_X1 U9066 ( .A1(n7313), .A2(n7311), .ZN(n6699) );
  OR2_X1 U9067 ( .A1(n11190), .A2(n13545), .ZN(n11256) );
  OR2_X1 U9068 ( .A1(n14398), .A2(n13228), .ZN(n6700) );
  INV_X1 U9069 ( .A(SI_1_), .ZN(n7265) );
  INV_X1 U9070 ( .A(n14045), .ZN(n7085) );
  OR2_X1 U9071 ( .A1(n12558), .A2(n12544), .ZN(n6701) );
  NAND2_X1 U9072 ( .A1(n7640), .A2(n7634), .ZN(n7925) );
  AND2_X1 U9073 ( .A1(n8980), .A2(n8979), .ZN(n6702) );
  INV_X1 U9074 ( .A(n7140), .ZN(n13062) );
  INV_X1 U9075 ( .A(n7152), .ZN(n6886) );
  AOI21_X1 U9076 ( .B1(n7155), .B2(n7153), .A(n6651), .ZN(n7152) );
  INV_X1 U9077 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6734) );
  INV_X1 U9078 ( .A(n7147), .ZN(n13103) );
  NAND2_X1 U9079 ( .A1(n7144), .A2(n7142), .ZN(n7147) );
  AND2_X1 U9080 ( .A1(n7156), .A2(n7158), .ZN(n6703) );
  OR2_X1 U9081 ( .A1(n13972), .A2(n11711), .ZN(n6704) );
  AND2_X1 U9082 ( .A1(n7391), .A2(n7389), .ZN(n6705) );
  NAND2_X1 U9083 ( .A1(n8445), .A2(n8444), .ZN(n11313) );
  INV_X1 U9084 ( .A(n8995), .ZN(n7525) );
  OR2_X1 U9085 ( .A1(n8982), .A2(n6702), .ZN(n6706) );
  AND2_X1 U9086 ( .A1(n7144), .A2(n7143), .ZN(n6707) );
  INV_X1 U9087 ( .A(n7145), .ZN(n7144) );
  AND2_X1 U9088 ( .A1(n7482), .A2(n7485), .ZN(n6708) );
  AND2_X1 U9089 ( .A1(n11313), .A2(n8446), .ZN(n6709) );
  OR2_X1 U9090 ( .A1(n9014), .A2(n9015), .ZN(n6710) );
  OR2_X1 U9091 ( .A1(n7512), .A2(n7511), .ZN(n6711) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U9093 ( .A1(n7202), .A2(n8779), .ZN(n10040) );
  NAND2_X1 U9094 ( .A1(n10527), .A2(n13423), .ZN(n10632) );
  INV_X2 U9095 ( .A(n14986), .ZN(n14989) );
  AND2_X1 U9096 ( .A1(n6587), .A2(n10676), .ZN(n6712) );
  NAND2_X1 U9097 ( .A1(n11319), .A2(n11485), .ZN(n12448) );
  AND2_X1 U9098 ( .A1(n14856), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U9099 ( .A1(n11704), .A2(n11703), .ZN(n14089) );
  INV_X1 U9100 ( .A(n14089), .ZN(n7159) );
  XOR2_X1 U9101 ( .A(n8021), .B(SI_23_), .Z(n6714) );
  AND2_X1 U9102 ( .A1(n7275), .A2(n7283), .ZN(n6715) );
  NOR2_X1 U9103 ( .A1(n8647), .A2(n7072), .ZN(n7071) );
  AND2_X1 U9104 ( .A1(n11141), .A2(n11480), .ZN(n6716) );
  AND2_X1 U9105 ( .A1(n6991), .A2(n6990), .ZN(n6717) );
  AND2_X1 U9106 ( .A1(n8089), .A2(SI_27_), .ZN(n6718) );
  NAND2_X1 U9107 ( .A1(n8767), .A2(n8766), .ZN(n6719) );
  INV_X2 U9108 ( .A(n12619), .ZN(n10011) );
  NOR2_X1 U9109 ( .A1(n9409), .A2(n14748), .ZN(n6720) );
  INV_X1 U9110 ( .A(n13817), .ZN(n6779) );
  INV_X1 U9111 ( .A(n14458), .ZN(n14440) );
  NAND2_X1 U9112 ( .A1(n8130), .A2(n8129), .ZN(n14753) );
  AND2_X1 U9113 ( .A1(n6774), .A2(n14809), .ZN(n14799) );
  INV_X1 U9114 ( .A(n14799), .ZN(n7116) );
  OR2_X1 U9115 ( .A1(n14814), .A2(n15256), .ZN(n6721) );
  NOR2_X1 U9116 ( .A1(n9871), .A2(n9870), .ZN(n6722) );
  INV_X1 U9117 ( .A(n14635), .ZN(n7080) );
  NAND2_X1 U9118 ( .A1(n11067), .A2(n11066), .ZN(n14476) );
  INV_X1 U9119 ( .A(n14476), .ZN(n7091) );
  NAND2_X1 U9120 ( .A1(n8739), .A2(n10039), .ZN(n12450) );
  OR2_X1 U9121 ( .A1(n13266), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6723) );
  AND2_X1 U9122 ( .A1(n8764), .A2(n8798), .ZN(n14920) );
  NAND2_X1 U9123 ( .A1(n12188), .A2(n12224), .ZN(n7007) );
  NAND2_X1 U9124 ( .A1(n15228), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6724) );
  INV_X1 U9125 ( .A(SI_4_), .ZN(n6729) );
  INV_X1 U9126 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7263) );
  INV_X1 U9127 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6827) );
  INV_X1 U9128 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6736) );
  INV_X1 U9129 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n7022) );
  INV_X1 U9130 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6842) );
  INV_X1 U9131 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6965) );
  INV_X1 U9132 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9133 ( .A1(n8721), .A2(n8720), .ZN(n8814) );
  OAI22_X1 U9134 ( .A1(n11408), .A2(n11407), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n11807), .ZN(n11398) );
  INV_X2 U9135 ( .A(n11418), .ZN(n12547) );
  OR2_X2 U9136 ( .A1(n11609), .A2(n7544), .ZN(n11419) );
  NAND2_X1 U9137 ( .A1(n8549), .A2(n8548), .ZN(n8564) );
  NAND2_X1 U9138 ( .A1(n8306), .A2(n8305), .ZN(n8328) );
  NAND2_X1 U9139 ( .A1(n6725), .A2(n8291), .ZN(n8304) );
  NAND2_X1 U9140 ( .A1(n8344), .A2(n8343), .ZN(n8364) );
  AND2_X2 U9141 ( .A1(n6753), .A2(n6598), .ZN(n10562) );
  NAND2_X1 U9142 ( .A1(n11919), .A2(n13319), .ZN(n13323) );
  NAND2_X1 U9143 ( .A1(n6824), .A2(n11940), .ZN(n9660) );
  NAND2_X1 U9144 ( .A1(n8290), .A2(n8289), .ZN(n6725) );
  NAND2_X1 U9145 ( .A1(n8420), .A2(n8419), .ZN(n8432) );
  NAND2_X1 U9146 ( .A1(n7482), .A2(n7481), .ZN(n11819) );
  INV_X1 U9147 ( .A(n9151), .ZN(n10091) );
  NAND4_X2 U9148 ( .A1(n9217), .A2(n6623), .A3(n9151), .A4(n6548), .ZN(n9223)
         );
  AND4_X2 U9149 ( .A1(n9476), .A2(n9146), .A3(n9145), .A4(n9147), .ZN(n9151)
         );
  NAND2_X1 U9150 ( .A1(n13294), .A2(n13293), .ZN(n13292) );
  INV_X1 U9151 ( .A(n8663), .ZN(n6726) );
  NAND2_X1 U9152 ( .A1(n7061), .A2(n6724), .ZN(n7063) );
  OAI22_X2 U9153 ( .A1(n8814), .A2(n8813), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(
        n13264), .ZN(n11394) );
  OAI21_X2 U9154 ( .B1(n8364), .B2(n7067), .A(n7064), .ZN(n8398) );
  NAND2_X1 U9155 ( .A1(n10355), .A2(n10354), .ZN(n10612) );
  NAND2_X1 U9156 ( .A1(n13292), .A2(n10353), .ZN(n10355) );
  NAND2_X1 U9157 ( .A1(n11400), .A2(n11399), .ZN(n11418) );
  NAND2_X1 U9158 ( .A1(n8586), .A2(n8585), .ZN(n8603) );
  NOR2_X1 U9159 ( .A1(n12277), .A2(n12260), .ZN(n11557) );
  NAND2_X1 U9160 ( .A1(n11237), .A2(n11409), .ZN(n8693) );
  NAND2_X1 U9161 ( .A1(n8583), .A2(n8582), .ZN(n8586) );
  NAND2_X1 U9162 ( .A1(n8566), .A2(n8565), .ZN(n8581) );
  NAND2_X1 U9163 ( .A1(n8400), .A2(n8399), .ZN(n8418) );
  AND2_X1 U9164 ( .A1(n11606), .A2(n11605), .ZN(n7078) );
  NAND4_X1 U9165 ( .A1(n6683), .A2(n7079), .A3(n7076), .A4(n7077), .ZN(n7075)
         );
  OAI22_X1 U9166 ( .A1(n8971), .A2(n7520), .B1(n8970), .B2(n8972), .ZN(n8978)
         );
  INV_X1 U9167 ( .A(n8877), .ZN(n7495) );
  NAND2_X1 U9168 ( .A1(n7502), .A2(n7500), .ZN(n8910) );
  OAI21_X1 U9169 ( .B1(n6870), .B2(n6869), .A(n7513), .ZN(n8988) );
  OAI21_X1 U9170 ( .B1(n9129), .B2(n11044), .A(n9133), .ZN(n9135) );
  NAND2_X1 U9171 ( .A1(n7616), .A2(n7615), .ZN(n7655) );
  OAI21_X1 U9172 ( .B1(n8276), .B2(n6842), .A(n6841), .ZN(n7587) );
  NAND2_X1 U9173 ( .A1(n6806), .A2(n6955), .ZN(n7874) );
  NAND2_X1 U9174 ( .A1(n7767), .A2(n7766), .ZN(n7769) );
  NAND2_X1 U9175 ( .A1(n7735), .A2(n7721), .ZN(n6924) );
  INV_X1 U9176 ( .A(n6963), .ZN(n6730) );
  NAND2_X1 U9177 ( .A1(n7056), .A2(n7054), .ZN(n8549) );
  NAND2_X1 U9178 ( .A1(n8564), .A2(n8563), .ZN(n8566) );
  NAND2_X1 U9179 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U9180 ( .A1(n8045), .A2(n8044), .ZN(n8058) );
  NAND2_X1 U9181 ( .A1(n7042), .A2(n11539), .ZN(n7041) );
  NAND2_X1 U9182 ( .A1(n12301), .A2(n11553), .ZN(n12292) );
  NAND2_X1 U9183 ( .A1(n7676), .A2(n7583), .ZN(n6906) );
  OAI21_X1 U9184 ( .B1(n13857), .B2(n7374), .A(n6676), .ZN(n7373) );
  AOI21_X1 U9185 ( .B1(n14027), .B2(n14581), .A(n7172), .ZN(n7171) );
  NAND2_X1 U9186 ( .A1(n6775), .A2(n6731), .ZN(n6853) );
  INV_X1 U9187 ( .A(n6732), .ZN(n6731) );
  OAI21_X1 U9188 ( .B1(n11578), .B2(n11569), .A(n7077), .ZN(n6732) );
  OAI22_X2 U9189 ( .A1(n7248), .A2(n7246), .B1(n13581), .B2(n7249), .ZN(n13585) );
  NAND2_X1 U9190 ( .A1(n13505), .A2(n13504), .ZN(n13510) );
  OR2_X1 U9191 ( .A1(n13517), .A2(n13518), .ZN(n13519) );
  NAND2_X1 U9192 ( .A1(n13572), .A2(n13571), .ZN(n13577) );
  NAND2_X1 U9193 ( .A1(n13595), .A2(n13594), .ZN(n13600) );
  NAND2_X1 U9194 ( .A1(n6761), .A2(n6760), .ZN(n13503) );
  NAND2_X1 U9195 ( .A1(n6763), .A2(n13665), .ZN(P1_U3242) );
  NAND2_X1 U9196 ( .A1(n14194), .A2(n14193), .ZN(n14153) );
  OAI21_X1 U9197 ( .B1(n14507), .B2(n14506), .A(n6840), .ZN(n6839) );
  XNOR2_X1 U9198 ( .A(n14220), .B(n7212), .ZN(n14257) );
  NOR2_X1 U9199 ( .A1(n15297), .A2(n15298), .ZN(n15296) );
  XNOR2_X1 U9200 ( .A(n14232), .B(n7211), .ZN(n14504) );
  NAND2_X1 U9201 ( .A1(n14196), .A2(n14195), .ZN(n6737) );
  NAND2_X1 U9202 ( .A1(n14502), .A2(n14234), .ZN(n14507) );
  NAND2_X1 U9203 ( .A1(n14256), .A2(n14222), .ZN(n14260) );
  NAND2_X1 U9204 ( .A1(n14505), .A2(n6839), .ZN(n14511) );
  INV_X1 U9205 ( .A(n9723), .ZN(n7327) );
  NAND2_X1 U9206 ( .A1(n8214), .A2(n14748), .ZN(n14808) );
  OAI211_X2 U9207 ( .C1(n14382), .C2(n7335), .A(n12635), .B(n7333), .ZN(n12746) );
  NAND2_X1 U9208 ( .A1(n8124), .A2(n7640), .ZN(n8126) );
  AOI211_X2 U9209 ( .C1(n12764), .C2(n12765), .A(n12648), .B(n12771), .ZN(
        n12763) );
  OAI211_X2 U9210 ( .C1(n6568), .C2(n10239), .A(n7728), .B(n7727), .ZN(n9757)
         );
  NAND2_X1 U9211 ( .A1(n14257), .A2(n15241), .ZN(n14256) );
  NAND2_X1 U9212 ( .A1(n14504), .A2(n14503), .ZN(n14502) );
  NAND2_X1 U9213 ( .A1(n12745), .A2(n12641), .ZN(n12786) );
  XNOR2_X1 U9214 ( .A(n14215), .B(n14216), .ZN(n15297) );
  NAND2_X1 U9215 ( .A1(n14497), .A2(n14496), .ZN(n14493) );
  XNOR2_X1 U9216 ( .A(n6740), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9217 ( .A1(n14302), .A2(n6741), .ZN(n6740) );
  NAND2_X1 U9218 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  INV_X1 U9219 ( .A(n14300), .ZN(n6743) );
  NAND2_X1 U9220 ( .A1(n14516), .A2(n15017), .ZN(n14513) );
  NAND2_X1 U9221 ( .A1(n14192), .A2(n15112), .ZN(n7214) );
  NOR2_X2 U9222 ( .A1(n8155), .A2(n6580), .ZN(n7627) );
  NAND2_X1 U9223 ( .A1(n6748), .A2(n6747), .ZN(n12301) );
  NAND2_X1 U9224 ( .A1(n14915), .A2(n14919), .ZN(n14914) );
  NAND2_X1 U9225 ( .A1(n10828), .A2(n11589), .ZN(n10827) );
  NAND2_X1 U9226 ( .A1(n10279), .A2(n11447), .ZN(n10278) );
  OAI21_X1 U9227 ( .B1(n11141), .B2(n7047), .A(n7045), .ZN(n8752) );
  OAI21_X2 U9228 ( .B1(n12419), .B2(n12421), .A(n11507), .ZN(n12413) );
  OAI21_X2 U9229 ( .B1(n12362), .B2(n11521), .A(n11522), .ZN(n12350) );
  AOI21_X1 U9230 ( .B1(n11421), .B2(n11420), .A(n11419), .ZN(n11422) );
  INV_X1 U9231 ( .A(n12304), .ZN(n6748) );
  OAI21_X2 U9232 ( .B1(n12445), .B2(n8753), .A(n11496), .ZN(n12419) );
  XNOR2_X1 U9233 ( .A(n8849), .B(n9119), .ZN(n13147) );
  OAI22_X2 U9234 ( .A1(n13059), .A2(n8207), .B1(n13194), .B2(n12832), .ZN(
        n13046) );
  NAND2_X1 U9235 ( .A1(n8193), .A2(n8192), .ZN(n10973) );
  AOI21_X2 U9236 ( .B1(n6782), .B2(n6637), .A(n7096), .ZN(n12983) );
  NAND2_X1 U9237 ( .A1(n13092), .A2(n8204), .ZN(n13070) );
  NAND2_X1 U9238 ( .A1(n13100), .A2(n13102), .ZN(n13099) );
  NAND2_X1 U9239 ( .A1(n13037), .A2(n13036), .ZN(n6782) );
  NAND2_X2 U9240 ( .A1(n7206), .A2(n6578), .ZN(n8731) );
  OAI21_X1 U9241 ( .B1(n6986), .B2(n12126), .A(n11997), .ZN(P3_U3154) );
  INV_X1 U9242 ( .A(n8278), .ZN(n6746) );
  OAI21_X2 U9243 ( .B1(n12357), .B2(n11583), .A(n11584), .ZN(n12344) );
  NOR2_X1 U9244 ( .A1(n12380), .A2(n7539), .ZN(n12369) );
  NAND2_X2 U9245 ( .A1(n6746), .A2(n14932), .ZN(n11437) );
  NAND2_X1 U9246 ( .A1(n10719), .A2(n8352), .ZN(n10831) );
  OR2_X1 U9247 ( .A1(n12137), .A2(n10401), .ZN(n11450) );
  INV_X1 U9248 ( .A(n11590), .ZN(n11447) );
  INV_X1 U9249 ( .A(n11196), .ZN(n6755) );
  NAND4_X1 U9250 ( .A1(n6616), .A2(n8230), .A3(n8233), .A4(n7050), .ZN(n6749)
         );
  NAND2_X1 U9251 ( .A1(n10827), .A2(n11464), .ZN(n11196) );
  OAI21_X1 U9252 ( .B1(n6755), .B2(n6592), .A(n6573), .ZN(n11140) );
  NAND2_X1 U9253 ( .A1(n11142), .A2(n6754), .ZN(n11141) );
  OAI21_X2 U9254 ( .B1(n12292), .B2(n11426), .A(n11424), .ZN(n12276) );
  NAND2_X1 U9255 ( .A1(n6765), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U9256 ( .A1(n7063), .A2(n8702), .ZN(n8719) );
  NAND2_X1 U9257 ( .A1(n10587), .A2(n10586), .ZN(n10798) );
  NAND2_X1 U9258 ( .A1(n10612), .A2(n10613), .ZN(n6753) );
  NAND2_X1 U9259 ( .A1(n13407), .A2(n13406), .ZN(n13405) );
  NAND2_X1 U9260 ( .A1(n13323), .A2(n11920), .ZN(n13395) );
  NAND2_X1 U9261 ( .A1(n12420), .A2(n8502), .ZN(n12407) );
  NAND2_X1 U9262 ( .A1(n12422), .A2(n12421), .ZN(n12420) );
  NAND2_X1 U9263 ( .A1(n12411), .A2(n11508), .ZN(n12401) );
  NAND2_X1 U9264 ( .A1(n10278), .A2(n11450), .ZN(n10740) );
  NAND2_X1 U9265 ( .A1(n10715), .A2(n11462), .ZN(n10828) );
  NAND2_X1 U9266 ( .A1(n10171), .A2(n11446), .ZN(n10279) );
  NAND2_X1 U9267 ( .A1(n11627), .A2(n11812), .ZN(n8682) );
  NOR2_X2 U9268 ( .A1(n12381), .A2(n12391), .ZN(n12380) );
  NAND2_X1 U9269 ( .A1(n10172), .A2(n8293), .ZN(n10288) );
  CLKBUF_X1 U9270 ( .A(n14931), .Z(n6756) );
  NAND2_X1 U9271 ( .A1(n11960), .A2(n8831), .ZN(n8837) );
  NAND2_X1 U9272 ( .A1(n6856), .A2(n7435), .ZN(n12435) );
  NAND2_X1 U9273 ( .A1(n10169), .A2(n11595), .ZN(n10171) );
  NAND2_X1 U9274 ( .A1(n8280), .A2(n8279), .ZN(n14918) );
  NAND2_X4 U9275 ( .A1(n8705), .A2(n8704), .ZN(n12477) );
  NOR2_X1 U9276 ( .A1(n10114), .A2(n10115), .ZN(n10313) );
  INV_X1 U9277 ( .A(n8469), .ZN(n6765) );
  NOR2_X1 U9278 ( .A1(n12180), .A2(n14870), .ZN(n14892) );
  NOR2_X1 U9279 ( .A1(n12177), .A2(n14845), .ZN(n14852) );
  NOR2_X1 U9280 ( .A1(n14850), .A2(n6713), .ZN(n12179) );
  XNOR2_X1 U9281 ( .A(n12179), .B(n14875), .ZN(n14871) );
  NAND3_X1 U9282 ( .A1(n13496), .A2(n13495), .A3(n6762), .ZN(n6761) );
  OR2_X1 U9283 ( .A1(n13586), .A2(n7258), .ZN(n7256) );
  OAI22_X1 U9284 ( .A1(n7250), .A2(n7252), .B1(n13513), .B2(n7253), .ZN(n13517) );
  OAI21_X1 U9285 ( .B1(n13658), .B2(n6784), .A(n11368), .ZN(n6763) );
  XNOR2_X2 U9286 ( .A(n9224), .B(n9395), .ZN(n9233) );
  NAND3_X1 U9287 ( .A1(n6586), .A2(n13601), .A3(n6689), .ZN(n7239) );
  OAI21_X1 U9288 ( .B1(n13556), .B2(n13555), .A(n13554), .ZN(n13559) );
  AOI21_X1 U9289 ( .B1(n7330), .B2(n7332), .A(n6682), .ZN(n7328) );
  NAND2_X1 U9290 ( .A1(n7457), .A2(n7455), .ZN(n13318) );
  NAND2_X1 U9291 ( .A1(n7806), .A2(n7807), .ZN(n10622) );
  INV_X1 U9292 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6968) );
  NAND2_X1 U9293 ( .A1(n6906), .A2(n7585), .ZN(n7709) );
  INV_X1 U9294 ( .A(n10420), .ZN(n7332) );
  NAND2_X1 U9295 ( .A1(n6764), .A2(n10420), .ZN(n7331) );
  NAND2_X1 U9296 ( .A1(n8434), .A2(n8433), .ZN(n8455) );
  NAND2_X1 U9297 ( .A1(n8330), .A2(n8329), .ZN(n8342) );
  OR2_X1 U9298 ( .A1(n11579), .A2(n11577), .ZN(n6775) );
  NAND2_X1 U9299 ( .A1(n8418), .A2(n8417), .ZN(n8420) );
  NAND2_X1 U9300 ( .A1(n8432), .A2(n8431), .ZN(n8434) );
  NAND2_X1 U9301 ( .A1(n8398), .A2(n8397), .ZN(n8400) );
  NAND2_X2 U9302 ( .A1(n8617), .A2(n8616), .ZN(n8633) );
  OAI21_X1 U9303 ( .B1(n8689), .B2(n8688), .A(n8690), .ZN(n8701) );
  XNOR2_X1 U9304 ( .A(n12295), .B(n6747), .ZN(n6769) );
  NAND2_X1 U9305 ( .A1(n12258), .A2(n6636), .ZN(n12263) );
  NAND2_X1 U9306 ( .A1(n8752), .A2(n11491), .ZN(n12445) );
  NAND2_X1 U9307 ( .A1(n7440), .A2(n7438), .ZN(n12598) );
  INV_X2 U9308 ( .A(n7590), .ZN(n7631) );
  NAND2_X1 U9309 ( .A1(n6963), .A2(SI_4_), .ZN(n7591) );
  NAND2_X1 U9310 ( .A1(n13651), .A2(n6785), .ZN(n6784) );
  AND2_X2 U9311 ( .A1(n7321), .A2(n7322), .ZN(n9721) );
  NAND2_X1 U9312 ( .A1(n7343), .A2(n12646), .ZN(n12765) );
  NAND2_X1 U9313 ( .A1(n10844), .A2(n6820), .ZN(n11115) );
  NOR2_X1 U9314 ( .A1(n12763), .A2(n6686), .ZN(n12716) );
  OAI21_X1 U9315 ( .B1(n12757), .B2(n7357), .A(n7355), .ZN(n7363) );
  INV_X1 U9316 ( .A(n10009), .ZN(n7350) );
  NAND2_X1 U9317 ( .A1(n7329), .A2(n7328), .ZN(n10760) );
  INV_X1 U9318 ( .A(n7349), .ZN(n7348) );
  NAND2_X1 U9319 ( .A1(n8614), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8617) );
  OR2_X1 U9320 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  INV_X1 U9321 ( .A(n6975), .ZN(n6972) );
  INV_X1 U9322 ( .A(n12083), .ZN(n6985) );
  XNOR2_X1 U9323 ( .A(n6987), .B(n12020), .ZN(n6986) );
  AOI21_X1 U9324 ( .B1(n12068), .B2(n11970), .A(n6691), .ZN(n12099) );
  OAI22_X1 U9325 ( .A1(n12997), .A2(n12996), .B1(n13162), .B2(n12827), .ZN(
        n12984) );
  NAND2_X1 U9326 ( .A1(n10067), .A2(n9770), .ZN(n7715) );
  NAND2_X1 U9327 ( .A1(n7310), .A2(n7308), .ZN(n13116) );
  NOR2_X1 U9328 ( .A1(n13115), .A2(n6911), .ZN(n13101) );
  OAI22_X1 U9329 ( .A1(n13019), .A2(n8015), .B1(n7138), .B2(n12829), .ZN(
        n13007) );
  NOR2_X2 U9330 ( .A1(n9204), .A2(n9203), .ZN(n13712) );
  NAND2_X2 U9331 ( .A1(n7686), .A2(n8869), .ZN(n9770) );
  NAND2_X1 U9332 ( .A1(n13142), .A2(n6936), .ZN(n13235) );
  NAND2_X1 U9333 ( .A1(n13221), .A2(n8201), .ZN(n13100) );
  NAND2_X1 U9334 ( .A1(n6783), .A2(n9082), .ZN(n9089) );
  OAI22_X1 U9335 ( .A1(n9093), .A2(n9094), .B1(n9081), .B2(n9080), .ZN(n6783)
         );
  NAND2_X1 U9336 ( .A1(n7295), .A2(n9019), .ZN(n9069) );
  INV_X1 U9337 ( .A(n8047), .ZN(n8045) );
  OAI21_X1 U9338 ( .B1(n7821), .B2(n7288), .A(n7608), .ZN(n7287) );
  INV_X2 U9339 ( .A(n7590), .ZN(n8276) );
  INV_X1 U9340 ( .A(n7400), .ZN(n7399) );
  OAI21_X1 U9341 ( .B1(n7370), .B2(n7369), .A(n7367), .ZN(n11775) );
  NAND2_X1 U9342 ( .A1(n7807), .A2(n6957), .ZN(n6806) );
  AOI21_X2 U9343 ( .B1(n13850), .B2(n14571), .A(n13849), .ZN(n14042) );
  OAI21_X1 U9344 ( .B1(n14032), .B2(n14276), .A(n7173), .ZN(n7172) );
  NAND2_X1 U9345 ( .A1(n7371), .A2(n6577), .ZN(n13848) );
  OAI21_X1 U9346 ( .B1(n14026), .B2(n14020), .A(n7171), .ZN(P1_U3356) );
  NAND3_X1 U9347 ( .A1(n13649), .A2(n13648), .A3(n13650), .ZN(n6786) );
  NAND2_X1 U9348 ( .A1(n7623), .A2(n6684), .ZN(n6953) );
  OR2_X1 U9349 ( .A1(n13593), .A2(n13592), .ZN(n13594) );
  OAI21_X1 U9350 ( .B1(n7631), .B2(n6965), .A(n6964), .ZN(n6963) );
  NOR2_X1 U9351 ( .A1(n14872), .A2(n14871), .ZN(n14870) );
  NAND2_X1 U9352 ( .A1(n9790), .A2(n9789), .ZN(n9792) );
  NOR2_X1 U9353 ( .A1(n14307), .A2(n14308), .ZN(n14306) );
  NOR2_X1 U9354 ( .A1(n14852), .A2(n14851), .ZN(n14850) );
  NOR2_X1 U9355 ( .A1(n14892), .A2(n14891), .ZN(n14890) );
  NOR2_X1 U9356 ( .A1(n11322), .A2(n14844), .ZN(n14845) );
  NAND2_X1 U9357 ( .A1(n7013), .A2(n7012), .ZN(n14336) );
  NAND2_X1 U9358 ( .A1(n6792), .A2(n6790), .ZN(P3_U3200) );
  NAND2_X1 U9359 ( .A1(n12189), .A2(n14843), .ZN(n6792) );
  NAND2_X1 U9360 ( .A1(n7063), .A2(n7062), .ZN(n8721) );
  NOR2_X2 U9361 ( .A1(n12547), .A2(n12128), .ZN(n11609) );
  NAND2_X1 U9362 ( .A1(n6794), .A2(n6793), .ZN(P3_U3296) );
  OAI21_X1 U9363 ( .B1(n6854), .B2(n11615), .A(n6795), .ZN(n6794) );
  NOR2_X1 U9364 ( .A1(n15290), .A2(n15291), .ZN(n15289) );
  XNOR2_X1 U9365 ( .A(n14203), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15290) );
  INV_X1 U9366 ( .A(n8731), .ZN(n7440) );
  OR2_X1 U9367 ( .A1(n8955), .A2(n8954), .ZN(n8961) );
  NAND2_X1 U9368 ( .A1(n11570), .A2(n11577), .ZN(n6798) );
  AOI21_X1 U9369 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n6869) );
  AOI21_X1 U9370 ( .B1(n7507), .B2(n6867), .A(n6865), .ZN(n9133) );
  AOI21_X1 U9371 ( .B1(n8988), .B2(n8987), .A(n8985), .ZN(n8986) );
  AOI21_X1 U9372 ( .B1(n8884), .B2(n8883), .A(n8881), .ZN(n8882) );
  INV_X1 U9373 ( .A(n8240), .ZN(n11812) );
  AOI21_X1 U9374 ( .B1(n12263), .B2(n12450), .A(n12262), .ZN(n12264) );
  NAND2_X1 U9375 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U9376 ( .A1(n9879), .A2(n9878), .ZN(n9927) );
  NAND2_X1 U9377 ( .A1(n7631), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U9378 ( .A1(n13578), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U9379 ( .A1(n7234), .A2(n7237), .ZN(n7233) );
  NAND2_X1 U9380 ( .A1(n6807), .A2(n13283), .ZN(P1_U3214) );
  NAND2_X1 U9381 ( .A1(n6808), .A2(n14440), .ZN(n6807) );
  OAI21_X1 U9382 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n6808) );
  NAND2_X1 U9383 ( .A1(n13980), .A2(n13962), .ZN(n13964) );
  NOR2_X2 U9384 ( .A1(n14653), .A2(n10964), .ZN(n10963) );
  NAND2_X1 U9385 ( .A1(n13462), .A2(n13463), .ZN(n13465) );
  AND2_X4 U9386 ( .A1(n9399), .A2(n11808), .ZN(n10245) );
  NAND2_X1 U9387 ( .A1(n7468), .A2(n6881), .ZN(n14134) );
  NAND3_X1 U9388 ( .A1(n6812), .A2(n8812), .A3(n12450), .ZN(n8750) );
  NAND2_X1 U9389 ( .A1(n8740), .A2(n12021), .ZN(n6812) );
  NAND2_X1 U9390 ( .A1(n6816), .A2(n6813), .ZN(P3_U3487) );
  NOR2_X1 U9391 ( .A1(n14989), .A2(n6815), .ZN(n6814) );
  NAND2_X1 U9392 ( .A1(n8810), .A2(n14989), .ZN(n6816) );
  NAND2_X1 U9393 ( .A1(n6819), .A2(n6817), .ZN(P3_U3455) );
  NAND2_X1 U9394 ( .A1(n8810), .A2(n14979), .ZN(n6819) );
  INV_X1 U9395 ( .A(n7363), .ZN(n12677) );
  NAND2_X1 U9396 ( .A1(n12491), .A2(n6701), .ZN(P3_U3484) );
  NAND2_X1 U9397 ( .A1(n7421), .A2(n7423), .ZN(n12283) );
  NAND2_X1 U9398 ( .A1(n13468), .A2(n13639), .ZN(n13469) );
  OAI21_X1 U9399 ( .B1(n6642), .B2(n6823), .A(n7242), .ZN(n13635) );
  NAND2_X1 U9400 ( .A1(n6848), .A2(n6692), .ZN(n6823) );
  INV_X1 U9401 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9144) );
  INV_X1 U9402 ( .A(n14151), .ZN(n9433) );
  NAND2_X1 U9403 ( .A1(n7976), .A2(n7975), .ZN(n6962) );
  NAND2_X1 U9404 ( .A1(n7787), .A2(n7600), .ZN(n7805) );
  NAND2_X1 U9405 ( .A1(n13489), .A2(n13488), .ZN(n13494) );
  OAI21_X1 U9406 ( .B1(n9223), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9225) );
  OAI21_X2 U9407 ( .B1(n10239), .B2(n13453), .A(n10238), .ZN(n14596) );
  OAI21_X1 U9408 ( .B1(n13494), .B2(n13493), .A(n13492), .ZN(n13496) );
  NAND2_X1 U9409 ( .A1(n13600), .A2(n13599), .ZN(n13598) );
  NAND2_X1 U9410 ( .A1(n13552), .A2(n13551), .ZN(n13556) );
  OAI21_X1 U9411 ( .B1(n13577), .B2(n13576), .A(n13575), .ZN(n13579) );
  NAND2_X1 U9412 ( .A1(n7107), .A2(n6679), .ZN(n8196) );
  NAND2_X1 U9413 ( .A1(n13120), .A2(n13119), .ZN(n13221) );
  NAND2_X1 U9414 ( .A1(n8185), .A2(n8184), .ZN(n9944) );
  AOI21_X2 U9415 ( .B1(n12969), .B2(n12968), .A(n7128), .ZN(n8849) );
  NAND2_X1 U9416 ( .A1(n8203), .A2(n13083), .ZN(n13092) );
  AOI21_X1 U9417 ( .B1(n11357), .B2(n11364), .A(n8200), .ZN(n13120) );
  AOI21_X1 U9418 ( .B1(n13046), .B2(n13045), .A(n8208), .ZN(n13037) );
  NAND2_X1 U9419 ( .A1(n10026), .A2(n10027), .ZN(n10025) );
  XNOR2_X1 U9420 ( .A(n14206), .B(n7210), .ZN(n15294) );
  NOR2_X1 U9421 ( .A1(n14499), .A2(n14500), .ZN(n14498) );
  NAND2_X1 U9422 ( .A1(n6828), .A2(n14302), .ZN(n7218) );
  NAND2_X1 U9423 ( .A1(n7785), .A2(n7784), .ZN(n7787) );
  NAND2_X1 U9424 ( .A1(n7990), .A2(n7989), .ZN(n7993) );
  NAND2_X1 U9425 ( .A1(n13277), .A2(n13278), .ZN(n13276) );
  INV_X1 U9426 ( .A(n6921), .ZN(n6920) );
  NAND2_X1 U9427 ( .A1(n7722), .A2(n6923), .ZN(n6922) );
  INV_X1 U9428 ( .A(n13589), .ZN(n7259) );
  NAND2_X1 U9429 ( .A1(n12413), .A2(n12412), .ZN(n12411) );
  NAND2_X1 U9430 ( .A1(n12433), .A2(n8486), .ZN(n12422) );
  NAND2_X1 U9431 ( .A1(n12435), .A2(n12434), .ZN(n12433) );
  NAND2_X1 U9432 ( .A1(n6838), .A2(n6835), .ZN(P3_U3454) );
  OR2_X1 U9433 ( .A1(n12548), .A2(n14977), .ZN(n6838) );
  NAND2_X1 U9434 ( .A1(n11315), .A2(n7436), .ZN(n6856) );
  INV_X1 U9435 ( .A(n14207), .ZN(n7210) );
  NAND2_X1 U9436 ( .A1(n14300), .A2(n14301), .ZN(n14302) );
  NAND2_X1 U9437 ( .A1(n15294), .A2(n15293), .ZN(n15292) );
  XNOR2_X1 U9438 ( .A(n12660), .B(n12658), .ZN(n12685) );
  NAND2_X1 U9439 ( .A1(n14264), .A2(n14263), .ZN(n7209) );
  INV_X1 U9440 ( .A(n7589), .ZN(n7262) );
  NAND2_X1 U9441 ( .A1(n7769), .A2(n7597), .ZN(n7785) );
  NAND2_X1 U9442 ( .A1(n6922), .A2(n6920), .ZN(n7767) );
  NAND2_X1 U9443 ( .A1(n7338), .A2(n7344), .ZN(n7343) );
  XNOR2_X1 U9444 ( .A(n7218), .B(n7216), .ZN(SUB_1596_U4) );
  NAND2_X1 U9445 ( .A1(n11617), .A2(n11616), .ZN(n6855) );
  OAI21_X1 U9446 ( .B1(n11581), .B2(n11580), .A(n6855), .ZN(n6854) );
  NAND2_X1 U9447 ( .A1(n13654), .A2(n6846), .ZN(n13651) );
  NAND2_X1 U9448 ( .A1(n13635), .A2(n13634), .ZN(n13654) );
  NAND2_X1 U9449 ( .A1(n13609), .A2(n13608), .ZN(n6848) );
  NAND2_X1 U9450 ( .A1(n6849), .A2(n7221), .ZN(n13567) );
  NAND3_X1 U9451 ( .A1(n13559), .A2(n13558), .A3(n7219), .ZN(n6849) );
  NAND2_X1 U9452 ( .A1(n7239), .A2(n7240), .ZN(n13606) );
  INV_X1 U9453 ( .A(n13579), .ZN(n7248) );
  NAND2_X1 U9454 ( .A1(n7582), .A2(n7672), .ZN(n7676) );
  NAND2_X1 U9455 ( .A1(n9793), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7026) );
  INV_X1 U9456 ( .A(n9792), .ZN(n9791) );
  NAND2_X1 U9457 ( .A1(n9819), .A2(n9820), .ZN(n9835) );
  XNOR2_X1 U9458 ( .A(n12182), .B(n14323), .ZN(n14307) );
  AOI21_X2 U9459 ( .B1(n6853), .B2(n7079), .A(n11609), .ZN(n11614) );
  AOI21_X2 U9460 ( .B1(n11571), .B2(n6600), .A(n11582), .ZN(n11576) );
  NAND2_X1 U9461 ( .A1(n8660), .A2(n8659), .ZN(n8662) );
  NAND2_X2 U9462 ( .A1(n8658), .A2(n8657), .ZN(n12295) );
  AND2_X2 U9463 ( .A1(n8857), .A2(n11044), .ZN(n8861) );
  OAI21_X1 U9464 ( .B1(n8909), .B2(n6858), .A(n6859), .ZN(n6857) );
  OR2_X1 U9465 ( .A1(n8909), .A2(n8906), .ZN(n8915) );
  NAND2_X1 U9466 ( .A1(n6860), .A2(n6693), .ZN(n7530) );
  NAND2_X1 U9467 ( .A1(n7521), .A2(n6696), .ZN(n6860) );
  NAND2_X1 U9468 ( .A1(n9061), .A2(n7296), .ZN(n6868) );
  NAND2_X1 U9469 ( .A1(n6871), .A2(n8124), .ZN(n8164) );
  AND2_X2 U9470 ( .A1(n7633), .A2(n7632), .ZN(n7640) );
  OAI22_X1 U9471 ( .A1(n7496), .A2(n6874), .B1(n8878), .B2(n8877), .ZN(n8884)
         );
  NAND2_X1 U9472 ( .A1(n10959), .A2(n6878), .ZN(n6875) );
  NAND2_X1 U9473 ( .A1(n6875), .A2(n6876), .ZN(n14267) );
  NAND3_X1 U9474 ( .A1(n6884), .A2(n6882), .A3(n6694), .ZN(n13941) );
  NAND2_X1 U9475 ( .A1(n14004), .A2(n6887), .ZN(n6882) );
  NAND2_X1 U9476 ( .A1(n13889), .A2(n6680), .ZN(n6892) );
  NAND2_X1 U9477 ( .A1(n6892), .A2(n6893), .ZN(n11805) );
  NAND2_X1 U9478 ( .A1(n13889), .A2(n11801), .ZN(n13872) );
  NAND2_X1 U9479 ( .A1(n11190), .A2(n6903), .ZN(n6902) );
  INV_X1 U9480 ( .A(n6906), .ZN(n7708) );
  NAND2_X1 U9481 ( .A1(n7631), .A2(n6695), .ZN(n6908) );
  NAND2_X1 U9482 ( .A1(n11019), .A2(n6916), .ZN(n6913) );
  NAND2_X1 U9483 ( .A1(n6913), .A2(n6914), .ZN(n7903) );
  AOI21_X1 U9484 ( .B1(n6916), .B2(n6918), .A(n7298), .ZN(n6914) );
  INV_X1 U9485 ( .A(n6924), .ZN(n6919) );
  OAI21_X1 U9486 ( .B1(n7260), .B2(n7593), .A(n7594), .ZN(n6921) );
  NAND2_X1 U9487 ( .A1(n8844), .A2(n6928), .ZN(n6926) );
  OAI211_X1 U9488 ( .C1(n8844), .C2(n6929), .A(n6937), .B(n6926), .ZN(n6927)
         );
  XNOR2_X2 U9489 ( .A(n7940), .B(SI_18_), .ZN(n7943) );
  NAND2_X1 U9490 ( .A1(n7807), .A2(n7603), .ZN(n7822) );
  INV_X1 U9491 ( .A(n7284), .ZN(n6959) );
  NAND2_X1 U9492 ( .A1(n7976), .A2(n6961), .ZN(n6960) );
  NAND4_X1 U9493 ( .A1(n14305), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n15028), 
        .A4(P2_ADDR_REG_19__SCAN_IN), .ZN(n6966) );
  NAND4_X1 U9494 ( .A1(n7580), .A2(n11652), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6968), .ZN(n6967) );
  INV_X1 U9495 ( .A(n12000), .ZN(n6970) );
  OAI22_X1 U9496 ( .A1(n10787), .A2(n6988), .B1(n7192), .B2(n6990), .ZN(n11281) );
  NAND2_X4 U9497 ( .A1(n6995), .A2(n6673), .ZN(n11032) );
  NAND2_X1 U9498 ( .A1(n8531), .A2(n6996), .ZN(n7001) );
  NAND2_X1 U9499 ( .A1(n12187), .A2(n7003), .ZN(n7002) );
  OAI211_X1 U9500 ( .C1(n12187), .C2(n7004), .A(n7002), .B(n12241), .ZN(
        P3_U3201) );
  NAND2_X1 U9501 ( .A1(n12187), .A2(n12188), .ZN(n12221) );
  NAND2_X1 U9502 ( .A1(n9870), .A2(n7018), .ZN(n7017) );
  NAND2_X1 U9503 ( .A1(n7016), .A2(n9869), .ZN(n9839) );
  NAND3_X1 U9504 ( .A1(n7016), .A2(n9869), .A3(n6591), .ZN(n7015) );
  NOR2_X1 U9505 ( .A1(n9937), .A2(n9936), .ZN(n10114) );
  NOR2_X1 U9506 ( .A1(n9935), .A2(n10110), .ZN(n10115) );
  AND2_X1 U9507 ( .A1(n9935), .A2(n10110), .ZN(n7020) );
  NAND2_X1 U9508 ( .A1(n7026), .A2(n9817), .ZN(n9819) );
  NAND2_X1 U9509 ( .A1(n12399), .A2(n7031), .ZN(n7030) );
  NAND2_X1 U9510 ( .A1(n7030), .A2(n7033), .ZN(n12362) );
  NAND2_X1 U9511 ( .A1(n12351), .A2(n11534), .ZN(n7042) );
  INV_X1 U9512 ( .A(n12350), .ZN(n7044) );
  AND2_X2 U9513 ( .A1(n7053), .A2(n7052), .ZN(n8470) );
  NAND2_X1 U9514 ( .A1(n8504), .A2(n7057), .ZN(n7056) );
  INV_X1 U9515 ( .A(n8701), .ZN(n7061) );
  AND2_X1 U9516 ( .A1(n6723), .A2(n8702), .ZN(n7062) );
  OAI21_X2 U9517 ( .B1(n8674), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8675), .ZN(
        n8689) );
  NAND2_X1 U9518 ( .A1(n8633), .A2(n7071), .ZN(n7069) );
  INV_X1 U9519 ( .A(n11607), .ZN(n7077) );
  NAND2_X1 U9520 ( .A1(n14646), .A2(n7543), .ZN(n10964) );
  AND3_X2 U9521 ( .A1(n7080), .A2(n7081), .A3(n14554), .ZN(n7543) );
  NAND2_X1 U9522 ( .A1(n13851), .A2(n7082), .ZN(n7083) );
  INV_X1 U9523 ( .A(n7083), .ZN(n13832) );
  AOI21_X1 U9524 ( .B1(n13840), .B2(n14029), .A(n6570), .ZN(n7084) );
  NOR2_X2 U9525 ( .A1(n6596), .A2(n14089), .ZN(n13980) );
  OR2_X2 U9526 ( .A1(n10973), .A2(n7111), .ZN(n7107) );
  NAND2_X1 U9527 ( .A1(n12969), .A2(n7122), .ZN(n7117) );
  NAND3_X1 U9528 ( .A1(n7118), .A2(n7117), .A3(n7119), .ZN(n13141) );
  NAND3_X1 U9529 ( .A1(n7118), .A2(n7117), .A3(n6589), .ZN(n7134) );
  INV_X2 U9530 ( .A(n6566), .ZN(n7951) );
  XNOR2_X2 U9531 ( .A(n7630), .B(n7629), .ZN(n8140) );
  NOR2_X2 U9532 ( .A1(n8850), .A2(n13139), .ZN(n12964) );
  NOR2_X2 U9533 ( .A1(n10057), .A2(n10219), .ZN(n10550) );
  NOR2_X2 U9534 ( .A1(n9766), .A2(n9757), .ZN(n9952) );
  OAI22_X1 U9535 ( .A1(n9547), .A2(n9251), .B1(n7631), .B2(n9255), .ZN(n7136)
         );
  NAND3_X1 U9536 ( .A1(n6587), .A2(n14820), .A3(n10676), .ZN(n11160) );
  NAND2_X1 U9537 ( .A1(n10379), .A2(n10378), .ZN(n10381) );
  NAND2_X1 U9538 ( .A1(n10430), .A2(n13482), .ZN(n7150) );
  NAND2_X1 U9539 ( .A1(n10270), .A2(n10269), .ZN(n10430) );
  NAND2_X1 U9540 ( .A1(n10687), .A2(n10686), .ZN(n10689) );
  NAND2_X1 U9541 ( .A1(n10620), .A2(n10619), .ZN(n7151) );
  NAND2_X1 U9542 ( .A1(n13926), .A2(n7162), .ZN(n7161) );
  XNOR2_X1 U9543 ( .A(n11805), .B(n13459), .ZN(n14026) );
  NAND2_X1 U9544 ( .A1(n12050), .A2(n12051), .ZN(n7184) );
  NAND2_X1 U9545 ( .A1(n7175), .A2(n7178), .ZN(n12023) );
  NAND2_X1 U9546 ( .A1(n12050), .A2(n7176), .ZN(n7175) );
  NAND2_X1 U9547 ( .A1(n7184), .A2(n11992), .ZN(n12106) );
  NAND2_X1 U9548 ( .A1(n8767), .A2(n6576), .ZN(n8769) );
  NAND2_X1 U9549 ( .A1(n8767), .A2(n7186), .ZN(n7185) );
  NAND2_X2 U9550 ( .A1(n11962), .A2(n7190), .ZN(n12000) );
  INV_X1 U9551 ( .A(n10787), .ZN(n7194) );
  INV_X1 U9552 ( .A(n11034), .ZN(n7200) );
  NAND2_X1 U9553 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  NAND3_X1 U9554 ( .A1(n7206), .A2(n7204), .A3(n7437), .ZN(n8736) );
  MUX2_X1 U9555 ( .A(n11437), .B(n10041), .S(n11032), .Z(n10085) );
  OAI211_X2 U9556 ( .C1(n13453), .C2(n9733), .A(n9732), .B(n9731), .ZN(n14573)
         );
  XNOR2_X1 U9557 ( .A(n12848), .B(n14794), .ZN(n9943) );
  NAND2_X1 U9558 ( .A1(n12012), .A2(n11974), .ZN(n12083) );
  NAND2_X1 U9559 ( .A1(n10046), .A2(n10047), .ZN(n10162) );
  INV_X1 U9560 ( .A(n9757), .ZN(n14789) );
  INV_X1 U9561 ( .A(n10173), .ZN(n11595) );
  NAND2_X1 U9562 ( .A1(n11446), .A2(n11445), .ZN(n10173) );
  AND2_X2 U9563 ( .A1(n14513), .A2(n14515), .ZN(n14246) );
  NOR2_X2 U9564 ( .A1(n15296), .A2(n14217), .ZN(n14220) );
  INV_X1 U9565 ( .A(n13520), .ZN(n7230) );
  NAND2_X1 U9566 ( .A1(n7231), .A2(n7232), .ZN(n13552) );
  NAND2_X1 U9567 ( .A1(n13531), .A2(n7234), .ZN(n7231) );
  AND2_X1 U9568 ( .A1(n13548), .A2(n7233), .ZN(n7232) );
  INV_X1 U9569 ( .A(n13580), .ZN(n7249) );
  NAND2_X1 U9570 ( .A1(n13511), .A2(n7251), .ZN(n7250) );
  INV_X1 U9571 ( .A(n13512), .ZN(n7253) );
  NOR2_X2 U9572 ( .A1(n9437), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U9573 ( .A1(n13503), .A2(n13502), .ZN(n13501) );
  NOR2_X1 U9574 ( .A1(n9219), .A2(n9479), .ZN(n7255) );
  NOR2_X2 U9575 ( .A1(n9220), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n9219) );
  OAI21_X1 U9576 ( .B1(n8276), .B2(n7263), .A(n7265), .ZN(n7264) );
  OAI21_X1 U9577 ( .B1(n7264), .B2(n6611), .A(n7583), .ZN(n7674) );
  INV_X1 U9578 ( .A(n11155), .ZN(n7300) );
  NAND2_X1 U9579 ( .A1(n9750), .A2(n9945), .ZN(n7307) );
  NAND2_X1 U9580 ( .A1(n7303), .A2(n7301), .ZN(n7765) );
  AND2_X1 U9581 ( .A1(n7302), .A2(n7762), .ZN(n7301) );
  OR2_X1 U9582 ( .A1(n7306), .A2(n9943), .ZN(n7302) );
  NAND2_X1 U9583 ( .A1(n9750), .A2(n7304), .ZN(n7303) );
  NOR2_X1 U9584 ( .A1(n7306), .A2(n7305), .ZN(n7304) );
  INV_X1 U9585 ( .A(n9945), .ZN(n7305) );
  INV_X1 U9586 ( .A(n7744), .ZN(n7306) );
  NAND2_X1 U9587 ( .A1(n7919), .A2(n6685), .ZN(n7310) );
  OAI21_X2 U9588 ( .B1(n10666), .B2(n7317), .A(n6665), .ZN(n11019) );
  INV_X1 U9589 ( .A(n9765), .ZN(n14780) );
  NAND2_X1 U9590 ( .A1(n7714), .A2(n9752), .ZN(n8181) );
  NAND2_X1 U9591 ( .A1(n9726), .A2(n9765), .ZN(n9752) );
  OAI21_X2 U9592 ( .B1(n8152), .B2(n7528), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7630) );
  NOR2_X2 U9593 ( .A1(n12775), .A2(n7318), .ZN(n12784) );
  NAND3_X1 U9594 ( .A1(n7324), .A2(n7327), .A3(n9688), .ZN(n7321) );
  NAND3_X1 U9595 ( .A1(n7325), .A2(n9522), .A3(n7327), .ZN(n7322) );
  OAI211_X1 U9596 ( .C1(n7324), .C2(n9522), .A(n9688), .B(n7323), .ZN(n9724)
         );
  NAND2_X1 U9597 ( .A1(n9683), .A2(n7326), .ZN(n7323) );
  NAND2_X1 U9598 ( .A1(n9522), .A2(n9521), .ZN(n9684) );
  INV_X1 U9599 ( .A(n9521), .ZN(n7326) );
  NAND2_X1 U9600 ( .A1(n10449), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U9601 ( .A1(n14381), .A2(n12625), .ZN(n7337) );
  INV_X1 U9602 ( .A(n12786), .ZN(n7338) );
  OAI21_X1 U9603 ( .B1(n9909), .B2(n7348), .A(n7345), .ZN(n10190) );
  INV_X1 U9604 ( .A(n13878), .ZN(n7370) );
  NAND2_X1 U9605 ( .A1(n13878), .A2(n6615), .ZN(n13863) );
  NAND2_X1 U9606 ( .A1(n13878), .A2(n7378), .ZN(n7371) );
  OR2_X2 U9607 ( .A1(n13972), .A2(n7381), .ZN(n13960) );
  AOI21_X1 U9608 ( .B1(n11294), .B2(n7387), .A(n7385), .ZN(n13991) );
  OAI21_X2 U9609 ( .B1(n10632), .B2(n7397), .A(n7392), .ZN(n10962) );
  NAND2_X1 U9610 ( .A1(n13945), .A2(n7402), .ZN(n7401) );
  INV_X1 U9611 ( .A(n7407), .ZN(n13928) );
  OR2_X1 U9612 ( .A1(n13954), .A2(n11725), .ZN(n7408) );
  INV_X2 U9613 ( .A(n14573), .ZN(n14590) );
  AND2_X2 U9614 ( .A1(n13478), .A2(n13479), .ZN(n14566) );
  XNOR2_X1 U9615 ( .A(n8238), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U9616 ( .A1(n10829), .A2(n6590), .ZN(n11198) );
  NAND3_X1 U9617 ( .A1(n10287), .A2(n8333), .A3(n8309), .ZN(n10741) );
  NAND2_X1 U9618 ( .A1(n12258), .A2(n8718), .ZN(n8740) );
  NAND2_X1 U9619 ( .A1(n8812), .A2(n7540), .ZN(n8818) );
  NAND2_X1 U9620 ( .A1(n13394), .A2(n7448), .ZN(n7447) );
  OAI211_X1 U9621 ( .C1(n13394), .C2(n6697), .A(n7449), .B(n7447), .ZN(n11951)
         );
  NAND2_X1 U9622 ( .A1(n13394), .A2(n11929), .ZN(n13277) );
  NAND2_X1 U9623 ( .A1(n13375), .A2(n7458), .ZN(n7457) );
  NOR2_X4 U9624 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9200) );
  NAND2_X1 U9625 ( .A1(n11343), .A2(n11344), .ZN(n7485) );
  NAND2_X1 U9626 ( .A1(n10798), .A2(n7491), .ZN(n10801) );
  INV_X1 U9627 ( .A(n7487), .ZN(n10939) );
  NOR2_X1 U9628 ( .A1(n10802), .A2(n7489), .ZN(n7488) );
  INV_X1 U9629 ( .A(n7491), .ZN(n7489) );
  NAND2_X1 U9630 ( .A1(n10940), .A2(n10941), .ZN(n7490) );
  INV_X1 U9631 ( .A(n8878), .ZN(n7494) );
  INV_X1 U9632 ( .A(n8871), .ZN(n7497) );
  NOR2_X1 U9633 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  INV_X1 U9634 ( .A(n8946), .ZN(n7499) );
  NAND2_X1 U9635 ( .A1(n7508), .A2(n6710), .ZN(n7507) );
  NAND3_X1 U9636 ( .A1(n7509), .A2(n6585), .A3(n6711), .ZN(n7508) );
  INV_X1 U9637 ( .A(n9008), .ZN(n7509) );
  INV_X1 U9638 ( .A(n9015), .ZN(n7511) );
  INV_X1 U9639 ( .A(n9014), .ZN(n7512) );
  NAND3_X1 U9640 ( .A1(n7517), .A2(n6857), .A3(n6690), .ZN(n7514) );
  NAND2_X1 U9641 ( .A1(n7514), .A2(n6687), .ZN(n8930) );
  INV_X1 U9642 ( .A(n8923), .ZN(n7515) );
  INV_X1 U9643 ( .A(n8922), .ZN(n7516) );
  OAI21_X1 U9644 ( .B1(n8915), .B2(n7519), .A(n7518), .ZN(n7517) );
  NAND3_X1 U9645 ( .A1(n8989), .A2(n6643), .A3(n7522), .ZN(n7521) );
  NAND2_X1 U9646 ( .A1(n7559), .A2(n7558), .ZN(n8152) );
  NAND2_X1 U9647 ( .A1(n7530), .A2(n7531), .ZN(n9010) );
  NAND3_X1 U9648 ( .A1(n8885), .A2(n6583), .A3(n6678), .ZN(n7532) );
  NAND2_X1 U9649 ( .A1(n7532), .A2(n7533), .ZN(n8894) );
  INV_X1 U9650 ( .A(n8848), .ZN(n8856) );
  NOR2_X2 U9651 ( .A1(n11296), .A2(n14106), .ZN(n14008) );
  CLKBUF_X1 U9652 ( .A(n8682), .Z(n8823) );
  OR2_X1 U9653 ( .A1(n8682), .A2(n8258), .ZN(n8262) );
  BUF_X1 U9654 ( .A(n9434), .Z(n9435) );
  NOR2_X2 U9655 ( .A1(n13021), .A2(n13168), .ZN(n13010) );
  INV_X1 U9656 ( .A(n8859), .ZN(n9409) );
  NAND2_X1 U9657 ( .A1(n12685), .A2(n12657), .ZN(n12684) );
  NAND4_X2 U9658 ( .A1(n8273), .A2(n8272), .A3(n8271), .A4(n8270), .ZN(n8751)
         );
  AOI21_X1 U9659 ( .B1(n13138), .B2(n14731), .A(n8219), .ZN(n8220) );
  NAND4_X2 U9660 ( .A1(n8286), .A2(n8285), .A3(n8284), .A4(n8283), .ZN(n12138)
         );
  INV_X1 U9661 ( .A(n8746), .ZN(n12223) );
  INV_X1 U9662 ( .A(n8301), .ZN(n8227) );
  INV_X1 U9663 ( .A(n8930), .ZN(n8933) );
  XNOR2_X1 U9664 ( .A(n8818), .B(n7076), .ZN(n8829) );
  NAND2_X1 U9665 ( .A1(n11391), .A2(n11574), .ZN(n11421) );
  NAND2_X2 U9666 ( .A1(n9166), .A2(n9165), .ZN(n9653) );
  INV_X1 U9667 ( .A(n12380), .ZN(n12383) );
  CLKBUF_X2 U9668 ( .A(n8278), .Z(n12139) );
  OR2_X1 U9669 ( .A1(n10144), .A2(n10143), .ZN(n14824) );
  OR2_X1 U9670 ( .A1(n10144), .A2(n10134), .ZN(n14834) );
  NAND2_X1 U9671 ( .A1(n14979), .A2(n14966), .ZN(n12597) );
  INV_X1 U9672 ( .A(n12597), .ZN(n8834) );
  AND2_X2 U9673 ( .A1(n8809), .A2(n9982), .ZN(n14979) );
  INV_X1 U9674 ( .A(n14575), .ZN(n14002) );
  OR2_X1 U9675 ( .A1(n12660), .A2(n12659), .ZN(n7534) );
  OR2_X1 U9676 ( .A1(n11841), .A2(n11840), .ZN(n7536) );
  AND2_X1 U9677 ( .A1(n11178), .A2(n11177), .ZN(n7537) );
  OR2_X1 U9678 ( .A1(n13141), .A2(n13114), .ZN(n7538) );
  AND2_X1 U9679 ( .A1(n12579), .A2(n12132), .ZN(n7539) );
  AND2_X1 U9680 ( .A1(n14747), .A2(n8863), .ZN(n7542) );
  AND2_X1 U9681 ( .A1(n11607), .A2(n11418), .ZN(n7544) );
  OR2_X1 U9682 ( .A1(n14396), .A2(n11359), .ZN(n7545) );
  INV_X1 U9683 ( .A(n11481), .ZN(n8444) );
  AOI21_X1 U9684 ( .B1(n13475), .B2(n13472), .A(n13471), .ZN(n13477) );
  INV_X1 U9685 ( .A(n8931), .ZN(n8932) );
  NAND2_X1 U9686 ( .A1(n13529), .A2(n13528), .ZN(n13531) );
  AND2_X1 U9687 ( .A1(n13545), .A2(n13535), .ZN(n13536) );
  OAI21_X1 U9688 ( .B1(n9013), .B2(n12750), .A(n8981), .ZN(n8982) );
  INV_X1 U9689 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8229) );
  INV_X1 U9690 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7553) );
  AND4_X1 U9691 ( .A1(n7632), .A2(n7552), .A3(n7551), .A4(n8165), .ZN(n7556)
         );
  INV_X1 U9692 ( .A(n11330), .ZN(n11331) );
  INV_X1 U9693 ( .A(n11979), .ZN(n11980) );
  OR2_X1 U9694 ( .A1(n14863), .A2(n14862), .ZN(n12154) );
  INV_X1 U9695 ( .A(n12592), .ZN(n8501) );
  INV_X1 U9696 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8221) );
  INV_X1 U9697 ( .A(n8007), .ZN(n8005) );
  INV_X1 U9698 ( .A(n7914), .ZN(n7570) );
  INV_X1 U9699 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7833) );
  INV_X1 U9700 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9701 ( .A1(n11329), .A2(n11331), .ZN(n11332) );
  AND2_X1 U9702 ( .A1(n14045), .A2(n13671), .ZN(n11802) );
  INV_X1 U9703 ( .A(n7843), .ZN(n7607) );
  NAND2_X1 U9704 ( .A1(n11978), .A2(n11980), .ZN(n11981) );
  INV_X1 U9705 ( .A(n8480), .ZN(n8479) );
  INV_X1 U9706 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U9707 ( .A1(n8707), .A2(n8706), .ZN(n8726) );
  NAND2_X1 U9708 ( .A1(n8776), .A2(n8778), .ZN(n8780) );
  INV_X1 U9709 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8766) );
  AND2_X1 U9710 ( .A1(n8503), .A2(n8488), .ZN(n8489) );
  XNOR2_X1 U9711 ( .A(n8869), .B(n6554), .ZN(n9518) );
  OR2_X1 U9712 ( .A1(n8028), .A2(n12758), .ZN(n8063) );
  OR2_X1 U9713 ( .A1(n7996), .A2(n12779), .ZN(n8007) );
  OR2_X1 U9714 ( .A1(n7931), .A2(n15272), .ZN(n7933) );
  INV_X1 U9715 ( .A(n13078), .ZN(n13200) );
  OR2_X1 U9716 ( .A1(n9708), .A2(n11910), .ZN(n9662) );
  INV_X1 U9717 ( .A(n13330), .ZN(n11844) );
  INV_X1 U9718 ( .A(n13433), .ZN(n11258) );
  INV_X1 U9719 ( .A(n11952), .ZN(n9322) );
  OR2_X1 U9720 ( .A1(n7977), .A2(n10201), .ZN(n7978) );
  NOR2_X1 U9721 ( .A1(n9478), .A2(n9477), .ZN(n9482) );
  INV_X1 U9722 ( .A(n12285), .ZN(n12260) );
  INV_X1 U9723 ( .A(n10487), .ZN(n10483) );
  AND2_X1 U9724 ( .A1(n9589), .A2(n9587), .ZN(n9593) );
  AND4_X1 U9725 ( .A1(n8577), .A2(n8576), .A3(n8575), .A4(n8574), .ZN(n12359)
         );
  AND2_X1 U9726 ( .A1(n11513), .A2(n11511), .ZN(n12400) );
  OR2_X1 U9727 ( .A1(n12135), .A2(n14959), .ZN(n11470) );
  NAND2_X1 U9728 ( .A1(n14986), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8838) );
  AND2_X1 U9729 ( .A1(n9961), .A2(n10281), .ZN(n10282) );
  NAND2_X1 U9730 ( .A1(n11550), .A2(n11553), .ZN(n12303) );
  INV_X1 U9731 ( .A(n8815), .ZN(n8591) );
  AND3_X1 U9732 ( .A1(n8382), .A2(n8381), .A3(n8380), .ZN(n14959) );
  INV_X1 U9733 ( .A(n12450), .ZN(n14939) );
  AND2_X1 U9734 ( .A1(n8548), .A2(n8525), .ZN(n8526) );
  INV_X1 U9735 ( .A(n14754), .ZN(n12801) );
  AND2_X1 U9736 ( .A1(n7854), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7866) );
  AND2_X1 U9737 ( .A1(n9136), .A2(n9130), .ZN(n9413) );
  INV_X1 U9738 ( .A(n12838), .ZN(n11359) );
  OR2_X1 U9739 ( .A1(n7690), .A2(n7699), .ZN(n7703) );
  AND2_X1 U9740 ( .A1(n9412), .A2(n14745), .ZN(n14795) );
  NOR2_X1 U9741 ( .A1(n11730), .A2(n15150), .ZN(n11729) );
  OR2_X1 U9742 ( .A1(n9648), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9455) );
  INV_X1 U9743 ( .A(n14433), .ZN(n14456) );
  AND2_X1 U9744 ( .A1(n11717), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11680) );
  OR2_X1 U9745 ( .A1(n13638), .A2(n13701), .ZN(n13388) );
  INV_X1 U9746 ( .A(n13388), .ZN(n13398) );
  OR2_X1 U9747 ( .A1(n13462), .A2(n10274), .ZN(n14642) );
  AOI22_X1 U9748 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14164), .B1(n14212), .B2(
        n14163), .ZN(n14166) );
  INV_X1 U9749 ( .A(n11474), .ZN(n14967) );
  INV_X1 U9750 ( .A(n12126), .ZN(n12058) );
  AND2_X1 U9751 ( .A1(n11406), .A2(n11405), .ZN(n12243) );
  AND2_X1 U9752 ( .A1(n8687), .A2(n8686), .ZN(n12274) );
  AND4_X1 U9753 ( .A1(n8611), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(n12360)
         );
  INV_X1 U9754 ( .A(n12197), .ZN(n14836) );
  INV_X1 U9755 ( .A(n14313), .ZN(n14895) );
  INV_X1 U9756 ( .A(n14357), .ZN(n14906) );
  INV_X1 U9757 ( .A(n14943), .ZN(n12453) );
  INV_X1 U9758 ( .A(n12431), .ZN(n12471) );
  AND2_X1 U9759 ( .A1(n12461), .A2(n14966), .ZN(n12470) );
  OR2_X1 U9760 ( .A1(n12243), .A2(n12242), .ZN(n14363) );
  AND2_X1 U9761 ( .A1(n14920), .A2(n12478), .ZN(n14973) );
  AND2_X1 U9762 ( .A1(n12541), .A2(n12540), .ZN(n12593) );
  INV_X1 U9763 ( .A(n14973), .ZN(n14963) );
  INV_X1 U9764 ( .A(n8804), .ZN(n11619) );
  NOR2_X1 U9765 ( .A1(n8537), .A2(n8536), .ZN(n14326) );
  INV_X1 U9766 ( .A(n12792), .ZN(n14688) );
  OR2_X1 U9767 ( .A1(n8097), .A2(n8096), .ZN(n8215) );
  OR2_X1 U9768 ( .A1(n12802), .A2(n6563), .ZN(n8072) );
  INV_X1 U9769 ( .A(n11644), .ZN(n14725) );
  INV_X1 U9770 ( .A(n12976), .ZN(n12968) );
  NAND2_X1 U9771 ( .A1(n14767), .A2(n8176), .ZN(n14751) );
  AND2_X1 U9772 ( .A1(n6558), .A2(n14753), .ZN(n13131) );
  INV_X1 U9773 ( .A(n9751), .ZN(n9748) );
  INV_X1 U9774 ( .A(n14753), .ZN(n13189) );
  OR2_X1 U9775 ( .A1(n10133), .A2(n10132), .ZN(n10144) );
  NAND2_X1 U9776 ( .A1(n8173), .A2(n8160), .ZN(n14759) );
  OR2_X1 U9777 ( .A1(n7887), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7906) );
  NOR2_X1 U9778 ( .A1(n10697), .A2(n10696), .ZN(n10917) );
  AND2_X1 U9779 ( .A1(n10365), .A2(n10231), .ZN(n14451) );
  AND2_X1 U9780 ( .A1(n14451), .A2(n14636), .ZN(n14447) );
  OR2_X1 U9781 ( .A1(n11769), .A2(n13839), .ZN(n11765) );
  INV_X1 U9782 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14164) );
  INV_X1 U9783 ( .A(n14534), .ZN(n13813) );
  INV_X1 U9784 ( .A(n6570), .ZN(n14577) );
  INV_X1 U9785 ( .A(n13566), .ZN(n13974) );
  AND2_X1 U9786 ( .A1(n11784), .A2(n10391), .ZN(n14581) );
  INV_X1 U9787 ( .A(n14012), .ZN(n14572) );
  AND2_X1 U9788 ( .A1(n9672), .A2(n10390), .ZN(n9564) );
  INV_X1 U9789 ( .A(n14636), .ZN(n14655) );
  INV_X1 U9790 ( .A(n14571), .ZN(n14550) );
  INV_X1 U9791 ( .A(n14639), .ZN(n14660) );
  AND2_X1 U9792 ( .A1(n10231), .A2(n10362), .ZN(n9672) );
  INV_X1 U9793 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9160) );
  AND2_X1 U9794 ( .A1(n9630), .A2(n10103), .ZN(n11056) );
  INV_X1 U9795 ( .A(n9319), .ZN(n9169) );
  INV_X1 U9796 ( .A(n6545), .ZN(n12121) );
  INV_X1 U9797 ( .A(n12124), .ZN(n11042) );
  AND2_X1 U9798 ( .A1(n11406), .A2(n8745), .ZN(n12026) );
  INV_X1 U9799 ( .A(n12324), .ZN(n12297) );
  INV_X2 U9800 ( .A(P3_U3897), .ZN(n12140) );
  INV_X1 U9801 ( .A(n14903), .ZN(n14882) );
  NAND2_X1 U9802 ( .A1(n14946), .A2(n14945), .ZN(n12431) );
  NAND2_X1 U9803 ( .A1(n14989), .A2(n14966), .ZN(n12544) );
  OR3_X1 U9804 ( .A1(n10285), .A2(n8800), .A3(n8799), .ZN(n14986) );
  INV_X1 U9805 ( .A(n14979), .ZN(n14977) );
  NAND2_X1 U9806 ( .A1(n8780), .A2(n9319), .ZN(n9329) );
  AND2_X1 U9807 ( .A1(n9962), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9319) );
  INV_X1 U9808 ( .A(n8778), .ZN(n11240) );
  INV_X1 U9809 ( .A(SI_16_), .ZN(n9531) );
  INV_X1 U9810 ( .A(SI_12_), .ZN(n9280) );
  OR2_X1 U9811 ( .A1(n9428), .A2(n9412), .ZN(n12806) );
  NAND2_X1 U9812 ( .A1(n9698), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14694) );
  INV_X1 U9813 ( .A(n13213), .ZN(n13110) );
  INV_X1 U9814 ( .A(n14690), .ZN(n12821) );
  NAND2_X1 U9815 ( .A1(n8088), .A2(n8087), .ZN(n12825) );
  INV_X1 U9816 ( .A(n14718), .ZN(n14706) );
  INV_X1 U9817 ( .A(n14760), .ZN(n14761) );
  INV_X1 U9818 ( .A(n14764), .ZN(n14767) );
  INV_X1 U9819 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13273) );
  INV_X1 U9820 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10770) );
  INV_X1 U9821 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9541) );
  AND2_X1 U9822 ( .A1(n9232), .A2(n9231), .ZN(n14525) );
  NAND2_X1 U9823 ( .A1(n10366), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14463) );
  INV_X1 U9824 ( .A(n14447), .ZN(n13414) );
  INV_X1 U9825 ( .A(n13819), .ZN(n14536) );
  INV_X1 U9826 ( .A(n14002), .ZN(n14276) );
  AND2_X1 U9827 ( .A1(n10263), .A2(n14010), .ZN(n14575) );
  OR2_X1 U9828 ( .A1(n14575), .A2(n10273), .ZN(n14020) );
  INV_X1 U9829 ( .A(n14679), .ZN(n14676) );
  OR3_X1 U9830 ( .A1(n14115), .A2(n14114), .A3(n14113), .ZN(n14133) );
  INV_X1 U9831 ( .A(n14663), .ZN(n14661) );
  AND2_X1 U9832 ( .A1(n10361), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9325) );
  INV_X1 U9833 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10198) );
  AND2_X1 U9834 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9175), .ZN(P2_U3947) );
  OAI211_X1 U9835 ( .C1(n13142), .C2(n14736), .A(n7538), .B(n8220), .ZN(
        P2_U3236) );
  INV_X1 U9836 ( .A(n13695), .ZN(P1_U4016) );
  AND3_X2 U9837 ( .A1(n7549), .A2(n7548), .A3(n7547), .ZN(n7634) );
  NOR2_X1 U9838 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7550) );
  NAND2_X1 U9839 ( .A1(n7634), .A2(n7550), .ZN(n8123) );
  INV_X1 U9840 ( .A(n8123), .ZN(n7557) );
  AND3_X2 U9841 ( .A1(n7827), .A2(n7705), .A3(n7847), .ZN(n7632) );
  NAND2_X1 U9842 ( .A1(n7948), .A2(n7354), .ZN(n8122) );
  INV_X1 U9843 ( .A(n8122), .ZN(n7552) );
  NOR2_X1 U9844 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7551) );
  NOR2_X1 U9845 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7555) );
  NOR2_X2 U9846 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7554) );
  INV_X2 U9847 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n15098) );
  NAND4_X1 U9848 ( .A1(n7555), .A2(n7554), .A3(n15098), .A4(n7553), .ZN(n7824)
         );
  NOR2_X2 U9849 ( .A1(n7824), .A2(n7725), .ZN(n7633) );
  NAND3_X1 U9850 ( .A1(n7557), .A2(n7556), .A3(n7633), .ZN(n8155) );
  INV_X1 U9851 ( .A(n8155), .ZN(n7559) );
  INV_X1 U9852 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7561) );
  NAND2_X1 U9853 ( .A1(n7627), .A2(n7561), .ZN(n7565) );
  INV_X1 U9854 ( .A(n7565), .ZN(n7563) );
  INV_X1 U9855 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9856 ( .A1(n7563), .A2(n7562), .ZN(n13250) );
  XNOR2_X2 U9857 ( .A(n7564), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7574) );
  INV_X1 U9858 ( .A(n7574), .ZN(n13257) );
  NAND2_X1 U9859 ( .A1(n7565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9860 ( .A1(n7679), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9861 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7756) );
  INV_X1 U9862 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7755) );
  NOR2_X1 U9863 ( .A1(n7756), .A2(n7755), .ZN(n7775) );
  NAND2_X1 U9864 ( .A1(n7775), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7795) );
  INV_X1 U9865 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7794) );
  INV_X1 U9866 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7812) );
  AND2_X1 U9867 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7568) );
  AND2_X1 U9868 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n7569) );
  INV_X1 U9869 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15272) );
  INV_X1 U9870 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U9871 ( .A1(n7933), .A2(n15268), .ZN(n7572) );
  NAND2_X1 U9872 ( .A1(n7955), .A2(n7572), .ZN(n13088) );
  OR2_X1 U9873 ( .A1(n6563), .A2(n13088), .ZN(n7578) );
  INV_X1 U9874 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7573) );
  OR2_X1 U9875 ( .A1(n7690), .A2(n7573), .ZN(n7577) );
  INV_X1 U9876 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7575) );
  OR2_X1 U9877 ( .A1(n8101), .A2(n7575), .ZN(n7576) );
  NAND4_X1 U9878 ( .A1(n7579), .A2(n7578), .A3(n7577), .A4(n7576), .ZN(n12834)
         );
  INV_X1 U9879 ( .A(n12834), .ZN(n12750) );
  INV_X1 U9880 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9457) );
  INV_X1 U9881 ( .A(SI_0_), .ZN(n9456) );
  NOR2_X1 U9882 ( .A1(n7581), .A2(n9456), .ZN(n7672) );
  INV_X1 U9883 ( .A(n7674), .ZN(n7582) );
  MUX2_X1 U9884 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7631), .Z(n7584) );
  NAND2_X1 U9885 ( .A1(n7584), .A2(SI_2_), .ZN(n7586) );
  OAI21_X1 U9886 ( .B1(n7584), .B2(SI_2_), .A(n7586), .ZN(n7707) );
  INV_X1 U9887 ( .A(n7707), .ZN(n7585) );
  NAND2_X1 U9888 ( .A1(n7587), .A2(SI_3_), .ZN(n7589) );
  OAI21_X1 U9889 ( .B1(SI_3_), .B2(n7587), .A(n7589), .ZN(n7588) );
  INV_X1 U9890 ( .A(n7588), .ZN(n7721) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8276), .Z(n7592) );
  NAND2_X1 U9892 ( .A1(n7592), .A2(SI_5_), .ZN(n7594) );
  OAI21_X1 U9893 ( .B1(n7592), .B2(SI_5_), .A(n7594), .ZN(n7593) );
  INV_X1 U9894 ( .A(n7593), .ZN(n7745) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8276), .Z(n7595) );
  NAND2_X1 U9896 ( .A1(n7595), .A2(SI_6_), .ZN(n7597) );
  OAI21_X1 U9897 ( .B1(SI_6_), .B2(n7595), .A(n7597), .ZN(n7596) );
  INV_X1 U9898 ( .A(n7596), .ZN(n7766) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8276), .Z(n7598) );
  NAND2_X1 U9900 ( .A1(n7598), .A2(SI_7_), .ZN(n7600) );
  OAI21_X1 U9901 ( .B1(SI_7_), .B2(n7598), .A(n7600), .ZN(n7599) );
  INV_X1 U9902 ( .A(n7599), .ZN(n7784) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7631), .Z(n7601) );
  NAND2_X1 U9904 ( .A1(n7601), .A2(SI_8_), .ZN(n7603) );
  OAI21_X1 U9905 ( .B1(SI_8_), .B2(n7601), .A(n7603), .ZN(n7602) );
  INV_X1 U9906 ( .A(n7602), .ZN(n7804) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n8276), .Z(n7604) );
  OAI21_X1 U9908 ( .B1(n7604), .B2(SI_9_), .A(n7606), .ZN(n7605) );
  INV_X1 U9909 ( .A(n7605), .ZN(n7821) );
  MUX2_X1 U9910 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n8276), .Z(n7843) );
  NAND2_X1 U9911 ( .A1(n7607), .A2(n9285), .ZN(n7608) );
  MUX2_X1 U9912 ( .A(n9543), .B(n9541), .S(n8276), .Z(n7609) );
  MUX2_X1 U9913 ( .A(n9644), .B(n9623), .S(n8276), .Z(n7610) );
  NAND2_X1 U9914 ( .A1(n7874), .A2(n7873), .ZN(n7612) );
  NAND2_X1 U9915 ( .A1(n7610), .A2(n9280), .ZN(n7611) );
  NAND2_X1 U9916 ( .A1(n7612), .A2(n7611), .ZN(n7886) );
  MUX2_X1 U9917 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n7631), .Z(n7613) );
  NAND2_X1 U9918 ( .A1(n7886), .A2(n7885), .ZN(n7616) );
  INV_X1 U9919 ( .A(n7613), .ZN(n7614) );
  NAND2_X1 U9920 ( .A1(n7614), .A2(n9328), .ZN(n7615) );
  INV_X1 U9921 ( .A(SI_14_), .ZN(n9392) );
  MUX2_X1 U9922 ( .A(n10106), .B(n10101), .S(n7631), .Z(n7904) );
  MUX2_X1 U9923 ( .A(n10338), .B(n10415), .S(n9020), .Z(n7659) );
  INV_X1 U9924 ( .A(n7659), .ZN(n7617) );
  NAND2_X1 U9925 ( .A1(n7617), .A2(SI_15_), .ZN(n7620) );
  OAI21_X1 U9926 ( .B1(n9392), .B2(n7904), .A(n7620), .ZN(n7618) );
  INV_X1 U9927 ( .A(n7618), .ZN(n7619) );
  INV_X1 U9928 ( .A(n7904), .ZN(n7657) );
  NOR2_X1 U9929 ( .A1(n7657), .A2(SI_14_), .ZN(n7621) );
  INV_X1 U9930 ( .A(SI_15_), .ZN(n9474) );
  AOI22_X1 U9931 ( .A1(n7621), .A2(n7620), .B1(n9474), .B2(n7659), .ZN(n7622)
         );
  MUX2_X1 U9932 ( .A(n10096), .B(n15273), .S(n9020), .Z(n7624) );
  NAND2_X1 U9933 ( .A1(n7624), .A2(n9531), .ZN(n7625) );
  MUX2_X1 U9934 ( .A(n10198), .B(n10228), .S(n9020), .Z(n7922) );
  MUX2_X1 U9935 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9020), .Z(n7939) );
  XNOR2_X1 U9936 ( .A(n7943), .B(n7939), .ZN(n11693) );
  NAND2_X1 U9937 ( .A1(n11693), .A2(n9026), .ZN(n7637) );
  INV_X2 U9938 ( .A(n9173), .ZN(n7950) );
  NAND2_X1 U9939 ( .A1(n7947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7635) );
  XNOR2_X1 U9940 ( .A(n7635), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U9941 ( .A1(n7951), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7950), .B2(
        n12949), .ZN(n7636) );
  INV_X1 U9942 ( .A(n13206), .ZN(n13091) );
  XNOR2_X1 U9943 ( .A(n7639), .B(n7638), .ZN(n11290) );
  NAND2_X1 U9944 ( .A1(n11290), .A2(n9026), .ZN(n7646) );
  INV_X1 U9945 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9946 ( .A1(n7640), .A2(n7641), .ZN(n7875) );
  INV_X1 U9947 ( .A(n7906), .ZN(n7643) );
  INV_X1 U9948 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7642) );
  NAND2_X1 U9949 ( .A1(n7643), .A2(n7642), .ZN(n7662) );
  OAI21_X1 U9950 ( .B1(n7662), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7644) );
  XNOR2_X1 U9951 ( .A(n7644), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U9952 ( .A1(n7951), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7950), .B2(
        n11133), .ZN(n7645) );
  INV_X1 U9953 ( .A(n13219), .ZN(n7921) );
  NAND2_X1 U9954 ( .A1(n9029), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7654) );
  INV_X1 U9955 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7648) );
  OR2_X1 U9956 ( .A1(n7647), .A2(n7648), .ZN(n7653) );
  INV_X1 U9957 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7667) );
  INV_X1 U9958 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7649) );
  OAI21_X1 U9959 ( .B1(n7914), .B2(n7667), .A(n7649), .ZN(n7650) );
  NAND2_X1 U9960 ( .A1(n7650), .A2(n7931), .ZN(n13121) );
  OR2_X1 U9961 ( .A1(n6564), .A2(n13121), .ZN(n7652) );
  INV_X1 U9962 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13125) );
  OR2_X1 U9963 ( .A1(n8101), .A2(n13125), .ZN(n7651) );
  NAND4_X1 U9964 ( .A1(n7654), .A2(n7653), .A3(n7652), .A4(n7651), .ZN(n12836)
         );
  XNOR2_X1 U9965 ( .A(n7655), .B(SI_14_), .ZN(n7905) );
  INV_X1 U9966 ( .A(n7905), .ZN(n7658) );
  INV_X1 U9967 ( .A(n7655), .ZN(n7656) );
  OAI22_X1 U9968 ( .A1(n7658), .A2(n7657), .B1(n7656), .B2(SI_14_), .ZN(n7661)
         );
  XNOR2_X1 U9969 ( .A(n7659), .B(SI_15_), .ZN(n7660) );
  XNOR2_X1 U9970 ( .A(n7661), .B(n7660), .ZN(n11243) );
  NAND2_X1 U9971 ( .A1(n11243), .A2(n9026), .ZN(n7665) );
  NAND2_X1 U9972 ( .A1(n7662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7663) );
  XNOR2_X1 U9973 ( .A(n7663), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14719) );
  AOI22_X1 U9974 ( .A1(n7951), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7950), .B2(
        n14719), .ZN(n7664) );
  NAND2_X1 U9975 ( .A1(n9029), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7671) );
  INV_X1 U9976 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7666) );
  OR2_X1 U9977 ( .A1(n7647), .A2(n7666), .ZN(n7670) );
  XNOR2_X1 U9978 ( .A(n7914), .B(n7667), .ZN(n12817) );
  OR2_X1 U9979 ( .A1(n6563), .A2(n12817), .ZN(n7669) );
  INV_X1 U9980 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11360) );
  OR2_X1 U9981 ( .A1(n8101), .A2(n11360), .ZN(n7668) );
  NAND4_X1 U9982 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n12837)
         );
  INV_X1 U9983 ( .A(n7672), .ZN(n7673) );
  NAND2_X1 U9984 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  NAND2_X1 U9985 ( .A1(n7676), .A2(n7675), .ZN(n9547) );
  NAND2_X1 U9986 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7677) );
  XNOR2_X1 U9987 ( .A(n7678), .B(n7677), .ZN(n12857) );
  NAND2_X1 U9988 ( .A1(n7679), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7685) );
  INV_X1 U9989 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7680) );
  OR2_X1 U9990 ( .A1(n7690), .A2(n7680), .ZN(n7684) );
  INV_X1 U9991 ( .A(n8135), .ZN(n7681) );
  INV_X1 U9992 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n12851) );
  INV_X1 U9993 ( .A(n8869), .ZN(n14772) );
  NAND2_X1 U9994 ( .A1(n8178), .A2(n14772), .ZN(n7687) );
  NAND2_X2 U9995 ( .A1(n9770), .A2(n7687), .ZN(n10070) );
  NAND2_X1 U9996 ( .A1(n7681), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7695) );
  INV_X1 U9997 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7688) );
  INV_X1 U9998 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9181) );
  NAND4_X2 U9999 ( .A1(n7695), .A2(n7694), .A3(n7693), .A4(n7692), .ZN(n8862)
         );
  NAND2_X1 U10000 ( .A1(n8276), .A2(SI_0_), .ZN(n7696) );
  XNOR2_X1 U10001 ( .A(n7696), .B(n8252), .ZN(n13274) );
  MUX2_X1 U10002 ( .A(n12860), .B(n13274), .S(n9173), .Z(n14747) );
  OR2_X1 U10003 ( .A1(n8862), .A2(n14747), .ZN(n10069) );
  NAND2_X1 U10004 ( .A1(n7679), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7704) );
  INV_X1 U10005 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7699) );
  INV_X1 U10006 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7700) );
  OR2_X1 U10007 ( .A1(n8135), .A2(n7700), .ZN(n7702) );
  INV_X1 U10008 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9525) );
  OR2_X1 U10009 ( .A1(n6563), .A2(n9525), .ZN(n7701) );
  NAND2_X1 U10010 ( .A1(n7725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7706) );
  XNOR2_X1 U10011 ( .A(n7706), .B(n7705), .ZN(n9254) );
  NAND2_X1 U10012 ( .A1(n7708), .A2(n7707), .ZN(n7710) );
  NAND2_X1 U10013 ( .A1(n7710), .A2(n7709), .ZN(n9733) );
  OR2_X1 U10014 ( .A1(n7711), .A2(n9733), .ZN(n7713) );
  OR2_X1 U10015 ( .A1(n6566), .A2(n9253), .ZN(n7712) );
  NAND2_X1 U10016 ( .A1(n8876), .A2(n14780), .ZN(n7714) );
  INV_X1 U10017 ( .A(n8181), .ZN(n9763) );
  NAND2_X1 U10018 ( .A1(n7715), .A2(n9763), .ZN(n9772) );
  NAND2_X1 U10019 ( .A1(n9772), .A2(n9752), .ZN(n7730) );
  NAND2_X1 U10020 ( .A1(n7679), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7720) );
  INV_X1 U10021 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7716) );
  OR2_X1 U10022 ( .A1(n7690), .A2(n7716), .ZN(n7719) );
  INV_X1 U10023 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9756) );
  OR2_X1 U10024 ( .A1(n8101), .A2(n9756), .ZN(n7718) );
  OR2_X1 U10025 ( .A1(n6563), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7717) );
  NAND4_X2 U10026 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n12849) );
  OR2_X1 U10027 ( .A1(n7722), .A2(n7721), .ZN(n7723) );
  NAND2_X1 U10028 ( .A1(n7724), .A2(n7723), .ZN(n10239) );
  NAND2_X1 U10029 ( .A1(n7739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7726) );
  INV_X1 U10030 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U10031 ( .A(n7726), .B(n7740), .ZN(n9333) );
  OR2_X1 U10032 ( .A1(n9173), .A2(n9333), .ZN(n7728) );
  OR2_X1 U10033 ( .A1(n6567), .A2(n9256), .ZN(n7727) );
  OR2_X1 U10034 ( .A1(n12849), .A2(n14789), .ZN(n9945) );
  NAND2_X1 U10035 ( .A1(n12849), .A2(n14789), .ZN(n7729) );
  NAND2_X1 U10036 ( .A1(n9945), .A2(n7729), .ZN(n9751) );
  NAND2_X1 U10037 ( .A1(n7679), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7734) );
  INV_X1 U10038 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9335) );
  OR2_X1 U10039 ( .A1(n7690), .A2(n9335), .ZN(n7733) );
  OAI21_X1 U10040 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7756), .ZN(n9955) );
  OR2_X1 U10041 ( .A1(n6563), .A2(n9955), .ZN(n7732) );
  INV_X1 U10042 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9951) );
  OR2_X1 U10043 ( .A1(n8135), .A2(n9951), .ZN(n7731) );
  NAND4_X1 U10044 ( .A1(n7734), .A2(n7733), .A3(n7732), .A4(n7731), .ZN(n12848) );
  OR2_X1 U10045 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  AND2_X1 U10046 ( .A1(n7738), .A2(n7737), .ZN(n10241) );
  NAND2_X1 U10047 ( .A1(n10241), .A2(n9026), .ZN(n7743) );
  INV_X1 U10048 ( .A(n7739), .ZN(n7826) );
  NAND2_X1 U10049 ( .A1(n7826), .A2(n7740), .ZN(n7749) );
  NAND2_X1 U10050 ( .A1(n7749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7741) );
  XNOR2_X1 U10051 ( .A(n7741), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9379) );
  AOI22_X1 U10052 ( .A1(n7951), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7950), .B2(
        n9379), .ZN(n7742) );
  NAND2_X1 U10053 ( .A1(n7743), .A2(n7742), .ZN(n14794) );
  INV_X1 U10054 ( .A(n14794), .ZN(n9956) );
  OR2_X1 U10055 ( .A1(n12848), .A2(n9956), .ZN(n7744) );
  OR2_X1 U10056 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  NAND2_X1 U10057 ( .A1(n7748), .A2(n7747), .ZN(n10356) );
  OR2_X1 U10058 ( .A1(n10356), .A2(n6568), .ZN(n7754) );
  INV_X1 U10059 ( .A(n7749), .ZN(n7751) );
  INV_X1 U10060 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10061 ( .A1(n7751), .A2(n7750), .ZN(n7770) );
  NAND2_X1 U10062 ( .A1(n7770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U10063 ( .A(n7752), .B(P2_IR_REG_5__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U10064 ( .A1(n7951), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7950), .B2(
        n12870), .ZN(n7753) );
  INV_X1 U10065 ( .A(n10060), .ZN(n10137) );
  NAND2_X1 U10066 ( .A1(n7679), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7761) );
  INV_X1 U10067 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10061) );
  OR2_X1 U10068 ( .A1(n8101), .A2(n10061), .ZN(n7760) );
  AND2_X1 U10069 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  OR2_X1 U10070 ( .A1(n7757), .A2(n7775), .ZN(n9910) );
  OR2_X1 U10071 ( .A1(n6563), .A2(n9910), .ZN(n7759) );
  INV_X1 U10072 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9336) );
  OR2_X1 U10073 ( .A1(n7690), .A2(n9336), .ZN(n7758) );
  NAND4_X1 U10074 ( .A1(n7761), .A2(n7760), .A3(n7759), .A4(n7758), .ZN(n12847) );
  NAND2_X1 U10075 ( .A1(n10137), .A2(n12847), .ZN(n7762) );
  INV_X1 U10076 ( .A(n12847), .ZN(n7763) );
  NAND2_X1 U10077 ( .A1(n7763), .A2(n10060), .ZN(n7764) );
  NAND2_X1 U10078 ( .A1(n7765), .A2(n7764), .ZN(n10024) );
  OR2_X1 U10079 ( .A1(n7767), .A2(n7766), .ZN(n7768) );
  NAND2_X1 U10080 ( .A1(n7769), .A2(n7768), .ZN(n10503) );
  OR2_X1 U10081 ( .A1(n10503), .A2(n6568), .ZN(n7773) );
  NAND2_X1 U10082 ( .A1(n7788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7771) );
  XNOR2_X1 U10083 ( .A(n7771), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9347) );
  AOI22_X1 U10084 ( .A1(n7951), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7950), .B2(
        n9347), .ZN(n7772) );
  NAND2_X1 U10085 ( .A1(n7773), .A2(n7772), .ZN(n10219) );
  NAND2_X1 U10086 ( .A1(n9029), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7781) );
  INV_X1 U10087 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7774) );
  OR2_X1 U10088 ( .A1(n7647), .A2(n7774), .ZN(n7780) );
  OR2_X1 U10089 ( .A1(n7775), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U10090 ( .A1(n7795), .A2(n7776), .ZN(n10030) );
  OR2_X1 U10091 ( .A1(n6564), .A2(n10030), .ZN(n7779) );
  INV_X1 U10092 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7777) );
  OR2_X1 U10093 ( .A1(n8135), .A2(n7777), .ZN(n7778) );
  NAND4_X1 U10094 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n12846) );
  XNOR2_X1 U10095 ( .A(n10219), .B(n10193), .ZN(n10026) );
  INV_X1 U10096 ( .A(n10026), .ZN(n8188) );
  NAND2_X1 U10097 ( .A1(n10024), .A2(n8188), .ZN(n7783) );
  NAND2_X1 U10098 ( .A1(n10219), .A2(n10193), .ZN(n7782) );
  NAND2_X1 U10099 ( .A1(n7783), .A2(n7782), .ZN(n10547) );
  OR2_X1 U10100 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U10101 ( .A1(n7787), .A2(n7786), .ZN(n10511) );
  OR2_X1 U10102 ( .A1(n10511), .A2(n6568), .ZN(n7792) );
  INV_X1 U10103 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U10104 ( .A1(n7789), .A2(n15098), .ZN(n7808) );
  NAND2_X1 U10105 ( .A1(n7808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7790) );
  XNOR2_X1 U10106 ( .A(n7790), .B(P2_IR_REG_7__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U10107 ( .A1(n7951), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7950), .B2(
        n12898), .ZN(n7791) );
  NAND2_X1 U10108 ( .A1(n7792), .A2(n7791), .ZN(n10552) );
  NAND2_X1 U10109 ( .A1(n9029), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7800) );
  INV_X1 U10110 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7793) );
  OR2_X1 U10111 ( .A1(n7647), .A2(n7793), .ZN(n7799) );
  NAND2_X1 U10112 ( .A1(n7795), .A2(n7794), .ZN(n7796) );
  NAND2_X1 U10113 ( .A1(n7813), .A2(n7796), .ZN(n14733) );
  OR2_X1 U10114 ( .A1(n6564), .A2(n14733), .ZN(n7798) );
  INV_X1 U10115 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9348) );
  OR2_X1 U10116 ( .A1(n8101), .A2(n9348), .ZN(n7797) );
  NAND4_X1 U10117 ( .A1(n7800), .A2(n7799), .A3(n7798), .A4(n7797), .ZN(n12845) );
  INV_X1 U10118 ( .A(n12845), .ZN(n7801) );
  AND2_X1 U10119 ( .A1(n10552), .A2(n7801), .ZN(n7803) );
  OR2_X1 U10120 ( .A1(n10552), .A2(n7801), .ZN(n7802) );
  OR2_X1 U10121 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  OR2_X1 U10122 ( .A1(n10622), .A2(n6568), .ZN(n7811) );
  OAI21_X1 U10123 ( .B1(n7808), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7809) );
  XNOR2_X1 U10124 ( .A(n7809), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9570) );
  AOI22_X1 U10125 ( .A1(n7951), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7950), .B2(
        n9570), .ZN(n7810) );
  NAND2_X2 U10126 ( .A1(n7811), .A2(n7810), .ZN(n10680) );
  NAND2_X1 U10127 ( .A1(n9030), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7819) );
  INV_X1 U10128 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10678) );
  OR2_X1 U10129 ( .A1(n8101), .A2(n10678), .ZN(n7818) );
  NAND2_X1 U10130 ( .A1(n7813), .A2(n7812), .ZN(n7814) );
  NAND2_X1 U10131 ( .A1(n7834), .A2(n7814), .ZN(n10677) );
  OR2_X1 U10132 ( .A1(n6564), .A2(n10677), .ZN(n7817) );
  INV_X1 U10133 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7815) );
  OR2_X1 U10134 ( .A1(n7690), .A2(n7815), .ZN(n7816) );
  NAND4_X1 U10135 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n12844) );
  XNOR2_X1 U10136 ( .A(n10680), .B(n12844), .ZN(n10675) );
  INV_X1 U10137 ( .A(n10675), .ZN(n10669) );
  INV_X1 U10138 ( .A(n12844), .ZN(n10424) );
  NAND2_X1 U10139 ( .A1(n10680), .A2(n10424), .ZN(n7820) );
  INV_X1 U10140 ( .A(n7824), .ZN(n7825) );
  NAND2_X1 U10141 ( .A1(n7826), .A2(n7825), .ZN(n7829) );
  NAND2_X1 U10142 ( .A1(n7829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7828) );
  MUX2_X1 U10143 ( .A(n7828), .B(P2_IR_REG_31__SCAN_IN), .S(n7827), .Z(n7830)
         );
  OR2_X1 U10144 ( .A1(n7829), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7846) );
  AOI22_X1 U10145 ( .A1(n7951), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7950), .B2(
        n14702), .ZN(n7831) );
  NAND2_X1 U10146 ( .A1(n7679), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7840) );
  INV_X1 U10147 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7832) );
  OR2_X1 U10148 ( .A1(n7690), .A2(n7832), .ZN(n7839) );
  INV_X1 U10149 ( .A(n7854), .ZN(n7836) );
  NAND2_X1 U10150 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  NAND2_X1 U10151 ( .A1(n7836), .A2(n7835), .ZN(n10820) );
  OR2_X1 U10152 ( .A1(n6564), .A2(n10820), .ZN(n7838) );
  INV_X1 U10153 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10821) );
  OR2_X1 U10154 ( .A1(n8101), .A2(n10821), .ZN(n7837) );
  NAND4_X1 U10155 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n12843) );
  XNOR2_X1 U10156 ( .A(n6569), .B(n12843), .ZN(n10813) );
  INV_X1 U10157 ( .A(n12843), .ZN(n7841) );
  OR2_X1 U10158 ( .A1(n6569), .A2(n7841), .ZN(n7842) );
  XNOR2_X1 U10159 ( .A(n7843), .B(SI_10_), .ZN(n7844) );
  XNOR2_X1 U10160 ( .A(n7845), .B(n7844), .ZN(n10907) );
  NAND2_X1 U10161 ( .A1(n10907), .A2(n9026), .ZN(n7852) );
  NAND2_X1 U10162 ( .A1(n7846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7848) );
  MUX2_X1 U10163 ( .A(n7848), .B(P2_IR_REG_31__SCAN_IN), .S(n7847), .Z(n7850)
         );
  INV_X1 U10164 ( .A(n7640), .ZN(n7849) );
  NAND2_X1 U10165 ( .A1(n7850), .A2(n7849), .ZN(n9888) );
  INV_X1 U10166 ( .A(n9888), .ZN(n9896) );
  AOI22_X1 U10167 ( .A1(n7951), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7950), 
        .B2(n9896), .ZN(n7851) );
  NAND2_X1 U10168 ( .A1(n9029), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7859) );
  INV_X1 U10169 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7853) );
  OR2_X1 U10170 ( .A1(n7647), .A2(n7853), .ZN(n7858) );
  NOR2_X1 U10171 ( .A1(n7854), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10172 ( .A1(n7866), .A2(n7855), .ZN(n10980) );
  OR2_X1 U10173 ( .A1(n6564), .A2(n10980), .ZN(n7857) );
  INV_X1 U10174 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10981) );
  OR2_X1 U10175 ( .A1(n8135), .A2(n10981), .ZN(n7856) );
  NAND4_X1 U10176 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n12842) );
  INV_X1 U10177 ( .A(n12842), .ZN(n9104) );
  XNOR2_X1 U10178 ( .A(n7861), .B(n7860), .ZN(n10913) );
  NAND2_X1 U10179 ( .A1(n10913), .A2(n9026), .ZN(n7864) );
  INV_X1 U10180 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8149) );
  OR2_X1 U10181 ( .A1(n7640), .A2(n8149), .ZN(n7862) );
  XNOR2_X1 U10182 ( .A(n7862), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U10183 ( .A1(n7951), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7950), 
        .B2(n12917), .ZN(n7863) );
  NAND2_X1 U10184 ( .A1(n9029), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7871) );
  INV_X1 U10185 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7865) );
  OR2_X1 U10186 ( .A1(n7647), .A2(n7865), .ZN(n7870) );
  NOR2_X1 U10187 ( .A1(n7866), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7867) );
  OR2_X1 U10188 ( .A1(n7892), .A2(n7867), .ZN(n11023) );
  OR2_X1 U10189 ( .A1(n6563), .A2(n11023), .ZN(n7869) );
  INV_X1 U10190 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11024) );
  OR2_X1 U10191 ( .A1(n8101), .A2(n11024), .ZN(n7868) );
  NAND4_X1 U10192 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n12841) );
  INV_X1 U10193 ( .A(n12841), .ZN(n8927) );
  XNOR2_X1 U10194 ( .A(n11027), .B(n8927), .ZN(n11016) );
  INV_X1 U10195 ( .A(n11016), .ZN(n11018) );
  NAND2_X1 U10196 ( .A1(n11027), .A2(n8927), .ZN(n7872) );
  XNOR2_X1 U10197 ( .A(n7874), .B(n7873), .ZN(n11055) );
  NAND2_X1 U10198 ( .A1(n11055), .A2(n9026), .ZN(n7878) );
  NAND2_X1 U10199 ( .A1(n7875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U10200 ( .A(n7876), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10201 ( .A1(n7951), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7950), 
        .B2(n9897), .ZN(n7877) );
  NAND2_X1 U10202 ( .A1(n9030), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10203 ( .A1(n8135), .A2(n15207), .ZN(n7881) );
  INV_X1 U10204 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9891) );
  OR2_X1 U10205 ( .A1(n7690), .A2(n9891), .ZN(n7880) );
  XNOR2_X1 U10206 ( .A(n7892), .B(P2_REG3_REG_12__SCAN_IN), .ZN(n14693) );
  OR2_X1 U10207 ( .A1(n6564), .A2(n14693), .ZN(n7879) );
  NAND4_X1 U10208 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n12840) );
  INV_X1 U10209 ( .A(n12840), .ZN(n11120) );
  XNOR2_X1 U10210 ( .A(n14689), .B(n11120), .ZN(n11154) );
  OR2_X1 U10211 ( .A1(n14689), .A2(n11120), .ZN(n7884) );
  XNOR2_X1 U10212 ( .A(n7886), .B(n7885), .ZN(n11061) );
  NAND2_X1 U10213 ( .A1(n11061), .A2(n9026), .ZN(n7891) );
  NAND2_X1 U10214 ( .A1(n7887), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7888) );
  MUX2_X1 U10215 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7888), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n7889) );
  NAND2_X1 U10216 ( .A1(n7889), .A2(n7906), .ZN(n10999) );
  INV_X1 U10217 ( .A(n10999), .ZN(n14710) );
  AOI22_X1 U10218 ( .A1(n7951), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7950), 
        .B2(n14710), .ZN(n7890) );
  NAND2_X1 U10219 ( .A1(n7679), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U10220 ( .A1(n7892), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7894) );
  INV_X1 U10221 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10222 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  NAND2_X1 U10223 ( .A1(n7895), .A2(n7912), .ZN(n11208) );
  OR2_X1 U10224 ( .A1(n6564), .A2(n11208), .ZN(n7899) );
  INV_X1 U10225 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7896) );
  OR2_X1 U10226 ( .A1(n8101), .A2(n7896), .ZN(n7898) );
  INV_X1 U10227 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10987) );
  OR2_X1 U10228 ( .A1(n7690), .A2(n10987), .ZN(n7897) );
  NAND4_X1 U10229 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n12839) );
  INV_X1 U10230 ( .A(n12839), .ZN(n14379) );
  NAND2_X1 U10231 ( .A1(n14410), .A2(n14379), .ZN(n7901) );
  OR2_X1 U10232 ( .A1(n14410), .A2(n14379), .ZN(n7902) );
  NAND2_X1 U10233 ( .A1(n7903), .A2(n7902), .ZN(n14388) );
  INV_X1 U10234 ( .A(n14388), .ZN(n7919) );
  XNOR2_X1 U10235 ( .A(n7905), .B(n7904), .ZN(n11171) );
  NAND2_X1 U10236 ( .A1(n11171), .A2(n9026), .ZN(n7909) );
  NAND2_X1 U10237 ( .A1(n7906), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7907) );
  XNOR2_X1 U10238 ( .A(n7907), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U10239 ( .A1(n7951), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7950), 
        .B2(n12938), .ZN(n7908) );
  NAND2_X1 U10240 ( .A1(n9030), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7918) );
  INV_X1 U10241 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7910) );
  OR2_X1 U10242 ( .A1(n7690), .A2(n7910), .ZN(n7917) );
  INV_X1 U10243 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7911) );
  OR2_X1 U10244 ( .A1(n8101), .A2(n7911), .ZN(n7916) );
  NAND2_X1 U10245 ( .A1(n7912), .A2(n15161), .ZN(n7913) );
  NAND2_X1 U10246 ( .A1(n7914), .A2(n7913), .ZN(n14391) );
  OR2_X1 U10247 ( .A1(n6563), .A2(n14391), .ZN(n7915) );
  NAND4_X1 U10248 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n12838) );
  NAND2_X1 U10249 ( .A1(n14396), .A2(n11359), .ZN(n7920) );
  INV_X1 U10250 ( .A(n12837), .ZN(n14380) );
  XNOR2_X1 U10251 ( .A(n13228), .B(n14380), .ZN(n11364) );
  INV_X1 U10252 ( .A(n12836), .ZN(n12749) );
  XNOR2_X1 U10253 ( .A(n13219), .B(n12749), .ZN(n13119) );
  XNOR2_X1 U10254 ( .A(n7922), .B(SI_17_), .ZN(n7923) );
  XNOR2_X1 U10255 ( .A(n7924), .B(n7923), .ZN(n11689) );
  NAND2_X1 U10256 ( .A1(n11689), .A2(n9026), .ZN(n7929) );
  NAND2_X1 U10257 ( .A1(n7925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7926) );
  MUX2_X1 U10258 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7926), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7927) );
  AND2_X1 U10259 ( .A1(n7927), .A2(n7947), .ZN(n11636) );
  AOI22_X1 U10260 ( .A1(n7951), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7950), 
        .B2(n11636), .ZN(n7928) );
  NAND2_X1 U10261 ( .A1(n9029), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7937) );
  INV_X1 U10262 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7930) );
  OR2_X1 U10263 ( .A1(n7647), .A2(n7930), .ZN(n7936) );
  NAND2_X1 U10264 ( .A1(n7931), .A2(n15272), .ZN(n7932) );
  NAND2_X1 U10265 ( .A1(n7933), .A2(n7932), .ZN(n13106) );
  OR2_X1 U10266 ( .A1(n6564), .A2(n13106), .ZN(n7935) );
  INV_X1 U10267 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13107) );
  OR2_X1 U10268 ( .A1(n8135), .A2(n13107), .ZN(n7934) );
  NAND4_X1 U10269 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n12835) );
  NOR2_X1 U10270 ( .A1(n13110), .A2(n12835), .ZN(n7938) );
  INV_X1 U10271 ( .A(n12835), .ZN(n12787) );
  INV_X1 U10272 ( .A(n7939), .ZN(n7942) );
  OAI21_X2 U10273 ( .B1(n7943), .B2(n7942), .A(n7941), .ZN(n7964) );
  MUX2_X1 U10274 ( .A(n10772), .B(n10770), .S(n9020), .Z(n7944) );
  INV_X1 U10275 ( .A(n7944), .ZN(n7945) );
  NAND2_X1 U10276 ( .A1(n7945), .A2(SI_19_), .ZN(n7946) );
  NAND2_X1 U10277 ( .A1(n7962), .A2(n7946), .ZN(n7963) );
  XNOR2_X1 U10278 ( .A(n7964), .B(n7963), .ZN(n11701) );
  NAND2_X1 U10279 ( .A1(n11701), .A2(n9026), .ZN(n7953) );
  INV_X1 U10280 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7948) );
  AOI22_X1 U10281 ( .A1(n7951), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9124), 
        .B2(n7950), .ZN(n7952) );
  INV_X1 U10282 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10283 ( .A1(n7955), .A2(n7954), .ZN(n7956) );
  NAND2_X1 U10284 ( .A1(n7982), .A2(n7956), .ZN(n13074) );
  INV_X1 U10285 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n11642) );
  OR2_X1 U10286 ( .A1(n7690), .A2(n11642), .ZN(n7959) );
  INV_X1 U10287 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7957) );
  OR2_X1 U10288 ( .A1(n7647), .A2(n7957), .ZN(n7958) );
  AND2_X1 U10289 ( .A1(n7959), .A2(n7958), .ZN(n7961) );
  NAND2_X1 U10290 ( .A1(n7681), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7960) );
  OAI211_X1 U10291 ( .C1(n13074), .C2(n6563), .A(n7961), .B(n7960), .ZN(n12833) );
  INV_X1 U10292 ( .A(n12833), .ZN(n12788) );
  OAI21_X2 U10293 ( .B1(n7964), .B2(n7963), .A(n7962), .ZN(n7977) );
  INV_X1 U10294 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11110) );
  MUX2_X1 U10295 ( .A(n11110), .B(n11043), .S(n9020), .Z(n7974) );
  XNOR2_X1 U10296 ( .A(n7976), .B(n7974), .ZN(n11712) );
  NAND2_X1 U10297 ( .A1(n11712), .A2(n9026), .ZN(n7966) );
  OR2_X1 U10298 ( .A1(n6567), .A2(n11043), .ZN(n7965) );
  NAND2_X2 U10299 ( .A1(n7966), .A2(n7965), .ZN(n13194) );
  XNOR2_X1 U10300 ( .A(n7982), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U10301 ( .A1(n13063), .A2(n7967), .ZN(n7973) );
  INV_X1 U10302 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10303 ( .A1(n9030), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10304 ( .A1(n9029), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7968) );
  OAI211_X1 U10305 ( .C1(n8101), .C2(n7970), .A(n7969), .B(n7968), .ZN(n7971)
         );
  INV_X1 U10306 ( .A(n7971), .ZN(n7972) );
  NAND2_X1 U10307 ( .A1(n7973), .A2(n7972), .ZN(n12832) );
  XNOR2_X1 U10308 ( .A(n13194), .B(n12832), .ZN(n13060) );
  INV_X1 U10309 ( .A(n12832), .ZN(n8993) );
  INV_X1 U10310 ( .A(n7974), .ZN(n7975) );
  INV_X1 U10311 ( .A(SI_20_), .ZN(n10201) );
  MUX2_X1 U10312 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9020), .Z(n7991) );
  XNOR2_X1 U10313 ( .A(n7991), .B(SI_21_), .ZN(n7988) );
  XNOR2_X1 U10314 ( .A(n7990), .B(n7988), .ZN(n11685) );
  NAND2_X1 U10315 ( .A1(n11685), .A2(n9026), .ZN(n7980) );
  INV_X1 U10316 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11221) );
  OR2_X1 U10317 ( .A1(n6567), .A2(n11221), .ZN(n7979) );
  INV_X1 U10318 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13050) );
  INV_X1 U10319 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7981) );
  INV_X1 U10320 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12719) );
  OAI21_X1 U10321 ( .B1(n7982), .B2(n7981), .A(n12719), .ZN(n7985) );
  AND2_X1 U10322 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n7983) );
  NAND2_X1 U10323 ( .A1(n7985), .A2(n7996), .ZN(n13049) );
  OR2_X1 U10324 ( .A1(n13049), .A2(n6564), .ZN(n7987) );
  AOI22_X1 U10325 ( .A1(n9030), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n9029), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n7986) );
  OAI211_X1 U10326 ( .C1(n8135), .C2(n13050), .A(n7987), .B(n7986), .ZN(n12831) );
  INV_X1 U10327 ( .A(n12831), .ZN(n12777) );
  INV_X1 U10328 ( .A(n13053), .ZN(n13185) );
  NAND2_X1 U10329 ( .A1(n7991), .A2(SI_21_), .ZN(n7992) );
  MUX2_X1 U10330 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9020), .Z(n8019) );
  XNOR2_X1 U10331 ( .A(n11669), .B(n8019), .ZN(n11287) );
  NAND2_X1 U10332 ( .A1(n11287), .A2(n9026), .ZN(n7995) );
  INV_X1 U10333 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15202) );
  OR2_X1 U10334 ( .A1(n6567), .A2(n15202), .ZN(n7994) );
  NAND2_X2 U10335 ( .A1(n7995), .A2(n7994), .ZN(n13179) );
  INV_X1 U10336 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8000) );
  INV_X1 U10337 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U10338 ( .A1(n7996), .A2(n12779), .ZN(n7997) );
  NAND2_X1 U10339 ( .A1(n8007), .A2(n7997), .ZN(n13032) );
  OR2_X1 U10340 ( .A1(n13032), .A2(n6563), .ZN(n7999) );
  AOI22_X1 U10341 ( .A1(n9030), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n9029), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n7998) );
  OAI211_X1 U10342 ( .C1(n8101), .C2(n8000), .A(n7999), .B(n7998), .ZN(n12830)
         );
  INV_X1 U10343 ( .A(n12830), .ZN(n12653) );
  XNOR2_X1 U10344 ( .A(n13179), .B(n12653), .ZN(n13036) );
  OAI22_X1 U10345 ( .A1(n13029), .A2(n13036), .B1(n12653), .B2(n13179), .ZN(
        n13019) );
  INV_X1 U10346 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8002) );
  INV_X1 U10347 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11373) );
  MUX2_X1 U10348 ( .A(n8002), .B(n11373), .S(n9020), .Z(n8021) );
  NAND2_X1 U10349 ( .A1(n11726), .A2(n9026), .ZN(n8004) );
  OR2_X1 U10350 ( .A1(n6567), .A2(n11373), .ZN(n8003) );
  NAND2_X2 U10351 ( .A1(n8004), .A2(n8003), .ZN(n13025) );
  INV_X1 U10352 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10353 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  NAND2_X1 U10354 ( .A1(n8028), .A2(n8008), .ZN(n12686) );
  OR2_X1 U10355 ( .A1(n12686), .A2(n6564), .ZN(n8014) );
  INV_X1 U10356 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10357 ( .A1(n9030), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8010) );
  INV_X1 U10358 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15226) );
  OR2_X1 U10359 ( .A1(n7690), .A2(n15226), .ZN(n8009) );
  OAI211_X1 U10360 ( .C1(n8011), .C2(n8101), .A(n8010), .B(n8009), .ZN(n8012)
         );
  INV_X1 U10361 ( .A(n8012), .ZN(n8013) );
  NAND2_X1 U10362 ( .A1(n8014), .A2(n8013), .ZN(n12829) );
  INV_X1 U10363 ( .A(n12829), .ZN(n12778) );
  NOR2_X1 U10364 ( .A1(n13025), .A2(n12778), .ZN(n8015) );
  INV_X1 U10365 ( .A(SI_23_), .ZN(n10714) );
  NAND2_X1 U10366 ( .A1(n8021), .A2(n10714), .ZN(n8023) );
  OAI21_X1 U10367 ( .B1(SI_22_), .B2(n8019), .A(n8023), .ZN(n8016) );
  INV_X1 U10368 ( .A(n8016), .ZN(n8017) );
  INV_X1 U10369 ( .A(n8019), .ZN(n8020) );
  INV_X1 U10370 ( .A(SI_22_), .ZN(n8636) );
  NOR2_X1 U10371 ( .A1(n8020), .A2(n8636), .ZN(n8024) );
  INV_X1 U10372 ( .A(n8021), .ZN(n8022) );
  AOI22_X1 U10373 ( .A1(n8024), .A2(n8023), .B1(n8022), .B2(SI_23_), .ZN(n8025) );
  MUX2_X1 U10374 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8276), .Z(n8036) );
  XNOR2_X1 U10375 ( .A(n8040), .B(n8036), .ZN(n11661) );
  NAND2_X1 U10376 ( .A1(n11661), .A2(n9026), .ZN(n8027) );
  INV_X1 U10377 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11388) );
  OR2_X1 U10378 ( .A1(n6567), .A2(n11388), .ZN(n8026) );
  INV_X1 U10379 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12758) );
  NAND2_X1 U10380 ( .A1(n8028), .A2(n12758), .ZN(n8029) );
  AND2_X1 U10381 ( .A1(n8063), .A2(n8029), .ZN(n13011) );
  NAND2_X1 U10382 ( .A1(n13011), .A2(n7967), .ZN(n8035) );
  INV_X1 U10383 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10384 ( .A1(n9029), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10385 ( .A1(n7679), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8030) );
  OAI211_X1 U10386 ( .C1(n8032), .C2(n8101), .A(n8031), .B(n8030), .ZN(n8033)
         );
  INV_X1 U10387 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10388 ( .A1(n8035), .A2(n8034), .ZN(n12828) );
  INV_X1 U10389 ( .A(n12828), .ZN(n12724) );
  XNOR2_X1 U10390 ( .A(n13168), .B(n12724), .ZN(n13014) );
  INV_X1 U10391 ( .A(n13014), .ZN(n13006) );
  INV_X1 U10392 ( .A(n8036), .ZN(n8039) );
  NAND2_X1 U10393 ( .A1(n8037), .A2(SI_24_), .ZN(n8038) );
  INV_X1 U10394 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11624) );
  MUX2_X1 U10395 ( .A(n11624), .B(n13273), .S(n9020), .Z(n8041) );
  NAND2_X1 U10396 ( .A1(n8041), .A2(n11138), .ZN(n8057) );
  INV_X1 U10397 ( .A(n8041), .ZN(n8042) );
  NAND2_X1 U10398 ( .A1(n8042), .A2(SI_25_), .ZN(n8043) );
  NAND2_X1 U10399 ( .A1(n8057), .A2(n8043), .ZN(n8046) );
  NAND2_X1 U10400 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U10401 ( .A1(n8058), .A2(n8048), .ZN(n11653) );
  NAND2_X1 U10402 ( .A1(n11653), .A2(n9026), .ZN(n8050) );
  OR2_X1 U10403 ( .A1(n6567), .A2(n13273), .ZN(n8049) );
  XNOR2_X1 U10404 ( .A(n8063), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U10405 ( .A1(n12999), .A2(n7967), .ZN(n8056) );
  INV_X1 U10406 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8053) );
  NAND2_X1 U10407 ( .A1(n7679), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U10408 ( .A1(n9029), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8051) );
  OAI211_X1 U10409 ( .C1(n8053), .C2(n8101), .A(n8052), .B(n8051), .ZN(n8054)
         );
  INV_X1 U10410 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U10411 ( .A1(n8056), .A2(n8055), .ZN(n12827) );
  INV_X1 U10412 ( .A(n12827), .ZN(n12795) );
  XNOR2_X1 U10413 ( .A(n13002), .B(n12795), .ZN(n12996) );
  INV_X1 U10414 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14146) );
  INV_X1 U10415 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15228) );
  MUX2_X1 U10416 ( .A(n14146), .B(n15228), .S(n9020), .Z(n8074) );
  XNOR2_X1 U10417 ( .A(n8074), .B(SI_26_), .ZN(n8059) );
  NAND2_X1 U10418 ( .A1(n13267), .A2(n9026), .ZN(n8061) );
  OR2_X1 U10419 ( .A1(n6567), .A2(n15228), .ZN(n8060) );
  INV_X1 U10420 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n15026) );
  INV_X1 U10421 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8062) );
  OAI21_X1 U10422 ( .B1(n8063), .B2(n15026), .A(n8062), .ZN(n8066) );
  INV_X1 U10423 ( .A(n8063), .ZN(n8065) );
  AND2_X1 U10424 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n8064) );
  NAND2_X1 U10425 ( .A1(n8065), .A2(n8064), .ZN(n8081) );
  NAND2_X1 U10426 ( .A1(n8066), .A2(n8081), .ZN(n12802) );
  INV_X1 U10427 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10428 ( .A1(n7679), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10429 ( .A1(n9029), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8067) );
  OAI211_X1 U10430 ( .C1(n8069), .C2(n8101), .A(n8068), .B(n8067), .ZN(n8070)
         );
  INV_X1 U10431 ( .A(n8070), .ZN(n8071) );
  INV_X1 U10432 ( .A(n12826), .ZN(n8211) );
  OR2_X1 U10433 ( .A1(n12991), .A2(n8211), .ZN(n9101) );
  NAND2_X1 U10434 ( .A1(n12984), .A2(n9101), .ZN(n8073) );
  NAND2_X1 U10435 ( .A1(n12991), .A2(n8211), .ZN(n9100) );
  NAND2_X1 U10436 ( .A1(n8073), .A2(n9100), .ZN(n12977) );
  INV_X1 U10437 ( .A(SI_26_), .ZN(n11238) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9020), .Z(n8089) );
  INV_X1 U10439 ( .A(n8089), .ZN(n8076) );
  XNOR2_X1 U10440 ( .A(n8076), .B(SI_27_), .ZN(n8077) );
  NAND2_X1 U10441 ( .A1(n13265), .A2(n9026), .ZN(n8080) );
  INV_X1 U10442 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13266) );
  OR2_X1 U10443 ( .A1(n6567), .A2(n13266), .ZN(n8079) );
  INV_X1 U10444 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U10445 ( .A1(n8081), .A2(n12680), .ZN(n8082) );
  NAND2_X1 U10446 ( .A1(n8097), .A2(n8082), .ZN(n12972) );
  OR2_X1 U10447 ( .A1(n12972), .A2(n6563), .ZN(n8088) );
  INV_X1 U10448 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U10449 ( .A1(n7679), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U10450 ( .A1(n9029), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8083) );
  OAI211_X1 U10451 ( .C1(n8101), .C2(n8085), .A(n8084), .B(n8083), .ZN(n8086)
         );
  INV_X1 U10452 ( .A(n8086), .ZN(n8087) );
  NAND2_X1 U10453 ( .A1(n12977), .A2(n12976), .ZN(n12975) );
  NOR2_X1 U10454 ( .A1(n8089), .A2(SI_27_), .ZN(n8090) );
  INV_X1 U10455 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11390) );
  INV_X1 U10456 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13264) );
  MUX2_X1 U10457 ( .A(n11390), .B(n13264), .S(n9020), .Z(n8091) );
  INV_X1 U10458 ( .A(SI_28_), .ZN(n12607) );
  NAND2_X1 U10459 ( .A1(n8091), .A2(n12607), .ZN(n8110) );
  INV_X1 U10460 ( .A(n8091), .ZN(n8092) );
  NAND2_X1 U10461 ( .A1(n8092), .A2(SI_28_), .ZN(n8093) );
  NAND2_X1 U10462 ( .A1(n8110), .A2(n8093), .ZN(n8108) );
  NAND2_X1 U10463 ( .A1(n13261), .A2(n9026), .ZN(n8095) );
  OR2_X1 U10464 ( .A1(n6567), .A2(n13264), .ZN(n8094) );
  INV_X1 U10465 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10466 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U10467 ( .A1(n12708), .A2(n7967), .ZN(n8104) );
  INV_X1 U10468 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U10469 ( .A1(n9029), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10470 ( .A1(n9030), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8099) );
  OAI211_X1 U10471 ( .C1(n8851), .C2(n8101), .A(n8100), .B(n8099), .ZN(n8102)
         );
  INV_X1 U10472 ( .A(n8102), .ZN(n8103) );
  NAND2_X1 U10473 ( .A1(n8104), .A2(n8103), .ZN(n12824) );
  NAND2_X1 U10474 ( .A1(n13144), .A2(n8212), .ZN(n8105) );
  INV_X1 U10475 ( .A(n12825), .ZN(n8106) );
  NAND2_X1 U10476 ( .A1(n13149), .A2(n8106), .ZN(n8843) );
  NAND3_X1 U10477 ( .A1(n12975), .A2(n9119), .A3(n8843), .ZN(n8844) );
  INV_X1 U10478 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14141) );
  INV_X1 U10479 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15002) );
  MUX2_X1 U10480 ( .A(n14141), .B(n15002), .S(n9020), .Z(n9018) );
  XNOR2_X1 U10481 ( .A(n9018), .B(SI_29_), .ZN(n9016) );
  NAND2_X1 U10482 ( .A1(n13258), .A2(n9026), .ZN(n8113) );
  OR2_X1 U10483 ( .A1(n6567), .A2(n15002), .ZN(n8112) );
  NAND2_X2 U10484 ( .A1(n8113), .A2(n8112), .ZN(n13139) );
  INV_X1 U10485 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U10486 ( .A1(n7681), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8115) );
  INV_X1 U10487 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n15097) );
  OR2_X1 U10488 ( .A1(n7690), .A2(n15097), .ZN(n8114) );
  OAI211_X1 U10489 ( .C1(n7647), .C2(n15256), .A(n8115), .B(n8114), .ZN(n8116)
         );
  INV_X1 U10490 ( .A(n8116), .ZN(n8117) );
  OAI21_X1 U10491 ( .B1(n8215), .B2(n6564), .A(n8117), .ZN(n12823) );
  INV_X1 U10492 ( .A(n12823), .ZN(n8118) );
  INV_X1 U10493 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8120) );
  XNOR2_X1 U10494 ( .A(n8121), .B(n8120), .ZN(n8213) );
  NOR2_X1 U10495 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U10496 ( .A1(n8126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8125) );
  MUX2_X1 U10497 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8125), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8127) );
  AND2_X2 U10498 ( .A1(n8127), .A2(n8164), .ZN(n9130) );
  OR2_X1 U10499 ( .A1(n11044), .A2(n11220), .ZN(n8130) );
  NAND2_X1 U10500 ( .A1(n9124), .A2(n9136), .ZN(n8129) );
  INV_X1 U10501 ( .A(n8131), .ZN(n8132) );
  NAND2_X1 U10502 ( .A1(n8132), .A2(n9413), .ZN(n14378) );
  INV_X1 U10503 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8133) );
  OR2_X1 U10504 ( .A1(n7690), .A2(n8133), .ZN(n8139) );
  INV_X1 U10505 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8134) );
  OR2_X1 U10506 ( .A1(n8135), .A2(n8134), .ZN(n8138) );
  INV_X1 U10507 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8136) );
  OR2_X1 U10508 ( .A1(n7647), .A2(n8136), .ZN(n8137) );
  AND3_X1 U10509 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n9077) );
  NAND2_X1 U10510 ( .A1(n8131), .A2(n9413), .ZN(n14754) );
  INV_X1 U10511 ( .A(P2_B_REG_SCAN_IN), .ZN(n8158) );
  NOR2_X1 U10512 ( .A1(n8140), .A2(n8158), .ZN(n8141) );
  OR2_X1 U10513 ( .A1(n14754), .A2(n8141), .ZN(n12958) );
  OAI22_X1 U10514 ( .A1(n8212), .A2(n14378), .B1(n9077), .B2(n12958), .ZN(
        n8142) );
  INV_X1 U10515 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15048) );
  INV_X1 U10516 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15065) );
  NAND2_X1 U10517 ( .A1(n15048), .A2(n15065), .ZN(n15221) );
  OR4_X1 U10518 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8143) );
  NOR4_X1 U10519 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n15221), .A4(n8143), .ZN(n8162) );
  INV_X1 U10520 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14992) );
  INV_X1 U10521 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15045) );
  INV_X1 U10522 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15084) );
  INV_X1 U10523 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15109) );
  NAND4_X1 U10524 ( .A1(n14992), .A2(n15045), .A3(n15084), .A4(n15109), .ZN(
        n15222) );
  NOR4_X1 U10525 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8147) );
  NOR4_X1 U10526 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8146) );
  NOR4_X1 U10527 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8145) );
  NOR4_X1 U10528 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8144) );
  NAND4_X1 U10529 ( .A1(n8147), .A2(n8146), .A3(n8145), .A4(n8144), .ZN(n8148)
         );
  NOR4_X1 U10530 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        n15222), .A4(n8148), .ZN(n8161) );
  OR2_X1 U10531 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U10532 ( .A1(n8153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8154) );
  XNOR2_X1 U10533 ( .A(n8154), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10534 ( .A1(n8155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8156) );
  MUX2_X1 U10535 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8156), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8157) );
  NAND2_X1 U10536 ( .A1(n8157), .A2(n8153), .ZN(n11387) );
  XNOR2_X1 U10537 ( .A(n11387), .B(n8158), .ZN(n8159) );
  OR2_X1 U10538 ( .A1(n8169), .A2(n8159), .ZN(n8160) );
  AOI21_X1 U10539 ( .B1(n8162), .B2(n8161), .A(n14759), .ZN(n9416) );
  INV_X1 U10540 ( .A(n9416), .ZN(n9408) );
  NAND2_X1 U10541 ( .A1(n8169), .A2(n8173), .ZN(n8163) );
  OAI21_X1 U10542 ( .B1(n8164), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8166) );
  XNOR2_X1 U10543 ( .A(n8166), .B(n8165), .ZN(n9419) );
  NAND2_X1 U10544 ( .A1(n9419), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10545 ( .A1(n11044), .A2(n14748), .ZN(n9412) );
  AND2_X1 U10546 ( .A1(n9412), .A2(n9413), .ZN(n9421) );
  NOR2_X1 U10547 ( .A1(n14764), .A2(n9421), .ZN(n8168) );
  NAND2_X1 U10548 ( .A1(n9408), .A2(n8168), .ZN(n10133) );
  OR2_X1 U10549 ( .A1(n14759), .A2(P2_D_REG_1__SCAN_IN), .ZN(n8171) );
  INV_X1 U10550 ( .A(n8173), .ZN(n13268) );
  INV_X1 U10551 ( .A(n8169), .ZN(n13270) );
  NAND2_X1 U10552 ( .A1(n13268), .A2(n13270), .ZN(n8170) );
  NAND2_X1 U10553 ( .A1(n8171), .A2(n8170), .ZN(n14766) );
  INV_X1 U10554 ( .A(n14766), .ZN(n9406) );
  OR2_X1 U10555 ( .A1(n14759), .A2(P2_D_REG_0__SCAN_IN), .ZN(n8174) );
  INV_X1 U10556 ( .A(n11387), .ZN(n8172) );
  OR2_X1 U10557 ( .A1(n8173), .A2(n8172), .ZN(n14762) );
  NAND2_X1 U10558 ( .A1(n8174), .A2(n14762), .ZN(n10134) );
  NAND2_X1 U10559 ( .A1(n9406), .A2(n10134), .ZN(n8175) );
  OR2_X1 U10560 ( .A1(n10133), .A2(n8175), .ZN(n8177) );
  NAND2_X1 U10561 ( .A1(n8861), .A2(n11220), .ZN(n10131) );
  INV_X1 U10562 ( .A(n10131), .ZN(n8176) );
  INV_X1 U10563 ( .A(n12991), .ZN(n13155) );
  INV_X1 U10564 ( .A(n14747), .ZN(n9676) );
  NAND2_X1 U10565 ( .A1(n8862), .A2(n9676), .ZN(n10066) );
  NAND2_X1 U10566 ( .A1(n10070), .A2(n10066), .ZN(n8180) );
  OR2_X1 U10567 ( .A1(n8178), .A2(n8869), .ZN(n8179) );
  NAND2_X1 U10568 ( .A1(n8180), .A2(n8179), .ZN(n9764) );
  NAND2_X1 U10569 ( .A1(n9764), .A2(n8181), .ZN(n8183) );
  OR2_X1 U10570 ( .A1(n8876), .A2(n9765), .ZN(n8182) );
  NAND2_X1 U10571 ( .A1(n8183), .A2(n8182), .ZN(n9749) );
  NAND2_X1 U10572 ( .A1(n9749), .A2(n9751), .ZN(n8185) );
  OR2_X1 U10573 ( .A1(n12849), .A2(n9757), .ZN(n8184) );
  INV_X1 U10574 ( .A(n9943), .ZN(n9946) );
  NAND2_X1 U10575 ( .A1(n9944), .A2(n9946), .ZN(n8187) );
  OR2_X1 U10576 ( .A1(n12848), .A2(n14794), .ZN(n8186) );
  OR2_X1 U10577 ( .A1(n10219), .A2(n12846), .ZN(n8189) );
  NAND2_X1 U10578 ( .A1(n10025), .A2(n8189), .ZN(n10545) );
  XNOR2_X1 U10579 ( .A(n10552), .B(n12845), .ZN(n10546) );
  INV_X1 U10580 ( .A(n10546), .ZN(n10544) );
  OR2_X1 U10581 ( .A1(n10552), .A2(n12845), .ZN(n8190) );
  NAND2_X1 U10582 ( .A1(n10680), .A2(n12844), .ZN(n8191) );
  NAND2_X1 U10583 ( .A1(n10672), .A2(n8191), .ZN(n10811) );
  INV_X1 U10584 ( .A(n10813), .ZN(n10810) );
  NAND2_X1 U10585 ( .A1(n10811), .A2(n10810), .ZN(n8193) );
  NAND2_X1 U10586 ( .A1(n6569), .A2(n12843), .ZN(n8192) );
  AND2_X1 U10587 ( .A1(n10979), .A2(n12842), .ZN(n8194) );
  NAND2_X1 U10588 ( .A1(n14410), .A2(n12839), .ZN(n8195) );
  NAND2_X1 U10589 ( .A1(n8196), .A2(n8195), .ZN(n14394) );
  AND2_X1 U10590 ( .A1(n14396), .A2(n12838), .ZN(n8197) );
  OR2_X1 U10591 ( .A1(n14396), .A2(n12838), .ZN(n8198) );
  NOR2_X1 U10592 ( .A1(n13228), .A2(n12837), .ZN(n8200) );
  NAND2_X1 U10593 ( .A1(n13219), .A2(n12836), .ZN(n8201) );
  XNOR2_X1 U10594 ( .A(n13213), .B(n12787), .ZN(n13102) );
  NAND2_X1 U10595 ( .A1(n13213), .A2(n12835), .ZN(n8202) );
  NAND2_X1 U10596 ( .A1(n13099), .A2(n8202), .ZN(n13094) );
  INV_X1 U10597 ( .A(n13094), .ZN(n8203) );
  XNOR2_X1 U10598 ( .A(n13206), .B(n12750), .ZN(n13083) );
  INV_X1 U10599 ( .A(n13083), .ZN(n13095) );
  OR2_X1 U10600 ( .A1(n13206), .A2(n12834), .ZN(n8204) );
  NOR2_X1 U10601 ( .A1(n13078), .A2(n12833), .ZN(n8205) );
  NAND2_X1 U10602 ( .A1(n13078), .A2(n12833), .ZN(n8206) );
  AND2_X1 U10603 ( .A1(n13194), .A2(n12832), .ZN(n8207) );
  XNOR2_X1 U10604 ( .A(n13053), .B(n12831), .ZN(n13043) );
  INV_X1 U10605 ( .A(n13043), .ZN(n13045) );
  NOR2_X1 U10606 ( .A1(n13053), .A2(n12831), .ZN(n8208) );
  NAND2_X1 U10607 ( .A1(n13025), .A2(n12829), .ZN(n9102) );
  OR2_X1 U10608 ( .A1(n13025), .A2(n12829), .ZN(n9103) );
  NAND2_X1 U10609 ( .A1(n13002), .A2(n12827), .ZN(n8209) );
  INV_X1 U10610 ( .A(n13144), .ZN(n8852) );
  XNOR2_X1 U10611 ( .A(n8859), .B(n11288), .ZN(n8214) );
  INV_X1 U10612 ( .A(n6774), .ZN(n14816) );
  OAI21_X2 U10613 ( .B1(n6720), .B2(n14816), .A(n6558), .ZN(n13114) );
  INV_X1 U10614 ( .A(n11027), .ZN(n14820) );
  NAND2_X1 U10615 ( .A1(n14772), .A2(n14747), .ZN(n10074) );
  OR2_X1 U10616 ( .A1(n10074), .A2(n9765), .ZN(n9766) );
  INV_X1 U10617 ( .A(n10552), .ZN(n14740) );
  AND2_X2 U10618 ( .A1(n10550), .A2(n14740), .ZN(n10676) );
  INV_X1 U10619 ( .A(n10680), .ZN(n14803) );
  OR2_X2 U10620 ( .A1(n11160), .A2(n14689), .ZN(n11212) );
  OR2_X2 U10621 ( .A1(n14410), .A2(n11212), .ZN(n14397) );
  OR2_X2 U10622 ( .A1(n14396), .A2(n14397), .ZN(n14398) );
  NAND2_X1 U10623 ( .A1(n13087), .A2(n13200), .ZN(n13073) );
  NAND2_X1 U10624 ( .A1(n13010), .A2(n13162), .ZN(n12998) );
  NAND2_X2 U10625 ( .A1(n11044), .A2(n14745), .ZN(n12619) );
  AOI211_X1 U10626 ( .C1(n13139), .C2(n8850), .A(n12664), .B(n12964), .ZN(
        n13138) );
  INV_X1 U10627 ( .A(n13139), .ZN(n8218) );
  INV_X1 U10628 ( .A(n11044), .ZN(n14749) );
  AND2_X1 U10629 ( .A1(n14749), .A2(n14745), .ZN(n9426) );
  INV_X1 U10630 ( .A(n8215), .ZN(n8216) );
  INV_X1 U10631 ( .A(n14751), .ZN(n14734) );
  AOI22_X1 U10632 ( .A1(n8216), .A2(n14734), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14736), .ZN(n8217) );
  OAI21_X1 U10633 ( .B1(n8218), .B2(n14739), .A(n8217), .ZN(n8219) );
  NAND2_X2 U10634 ( .A1(n12598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8238) );
  INV_X1 U10635 ( .A(n8239), .ZN(n11627) );
  NAND2_X1 U10636 ( .A1(n6560), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8244) );
  INV_X1 U10637 ( .A(n8644), .ZN(n8310) );
  NAND2_X1 U10638 ( .A1(n8310), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10639 ( .A1(n8641), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10640 ( .A1(n8312), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8241) );
  INV_X1 U10641 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10642 ( .A1(n8773), .A2(n8247), .ZN(n8248) );
  INV_X1 U10643 ( .A(n8275), .ZN(n8253) );
  NAND2_X1 U10644 ( .A1(n8253), .A2(n8264), .ZN(n8255) );
  NAND2_X1 U10645 ( .A1(n9255), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10646 ( .A1(n8255), .A2(n8254), .ZN(n8290) );
  XNOR2_X1 U10647 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8289) );
  XNOR2_X1 U10648 ( .A(n8290), .B(n8289), .ZN(n9272) );
  NAND2_X2 U10649 ( .A1(n11438), .A2(n11439), .ZN(n11591) );
  NAND2_X1 U10650 ( .A1(n8312), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8263) );
  INV_X1 U10651 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10652 ( .A1(n8641), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8261) );
  INV_X1 U10653 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8259) );
  OR2_X1 U10654 ( .A1(n8644), .A2(n8259), .ZN(n8260) );
  OR2_X1 U10655 ( .A1(n8396), .A2(n7265), .ZN(n8269) );
  XNOR2_X1 U10656 ( .A(n8264), .B(n6789), .ZN(n9260) );
  INV_X1 U10657 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10658 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8265) );
  OR2_X1 U10659 ( .A1(n6556), .A2(n9601), .ZN(n8267) );
  NAND2_X1 U10660 ( .A1(n8278), .A2(n14931), .ZN(n11436) );
  NAND2_X1 U10661 ( .A1(n8312), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10662 ( .A1(n8641), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10663 ( .A1(n8310), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10664 ( .A1(n9457), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10665 ( .A1(n6789), .A2(n8274), .ZN(n8277) );
  MUX2_X1 U10666 ( .A(n8277), .B(SI_0_), .S(n8276), .Z(n12611) );
  MUX2_X1 U10667 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12611), .S(n6557), .Z(n10474)
         );
  NAND2_X1 U10668 ( .A1(n8751), .A2(n10474), .ZN(n10086) );
  NAND2_X1 U10669 ( .A1(n10081), .A2(n10086), .ZN(n8280) );
  NAND2_X1 U10670 ( .A1(n14922), .A2(n6756), .ZN(n8279) );
  INV_X1 U10671 ( .A(n10050), .ZN(n14916) );
  NOR2_X1 U10672 ( .A1(n6553), .A2(n14916), .ZN(n8282) );
  NAND2_X1 U10673 ( .A1(n8710), .A2(n8295), .ZN(n8286) );
  NAND2_X1 U10674 ( .A1(n8311), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10675 ( .A1(n8641), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10676 ( .A1(n8310), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10677 ( .A1(n8301), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8287) );
  XNOR2_X1 U10678 ( .A(n8287), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U10679 ( .A1(n9253), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U10680 ( .A(n8304), .B(n8303), .ZN(n9264) );
  OR2_X1 U10681 ( .A1(n8815), .A2(SI_3_), .ZN(n8292) );
  INV_X1 U10682 ( .A(n10298), .ZN(n12469) );
  NAND2_X1 U10683 ( .A1(n12138), .A2(n12469), .ZN(n8293) );
  NAND2_X1 U10684 ( .A1(n8310), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10685 ( .A1(n8311), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10686 ( .A1(n8295), .A2(n8294), .ZN(n8315) );
  NAND2_X1 U10687 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8296) );
  NAND2_X1 U10688 ( .A1(n8315), .A2(n8296), .ZN(n10396) );
  NAND2_X1 U10689 ( .A1(n8710), .A2(n10396), .ZN(n8298) );
  NAND2_X1 U10690 ( .A1(n8641), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8297) );
  NAND4_X1 U10691 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n12137) );
  OR2_X1 U10692 ( .A1(n8301), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10693 ( .A1(n8321), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10694 ( .A1(n8304), .A2(n8303), .ZN(n8306) );
  NAND2_X1 U10695 ( .A1(n9256), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8305) );
  XNOR2_X1 U10696 ( .A(n8328), .B(n8327), .ZN(n9266) );
  OR2_X1 U10697 ( .A1(n8529), .A2(n9266), .ZN(n8308) );
  OR2_X1 U10698 ( .A1(n8815), .A2(SI_4_), .ZN(n8307) );
  OAI211_X1 U10699 ( .C1(n9836), .C2(n9579), .A(n8308), .B(n8307), .ZN(n10401)
         );
  NAND2_X1 U10700 ( .A1(n12137), .A2(n10401), .ZN(n11449) );
  INV_X1 U10701 ( .A(n10401), .ZN(n10410) );
  NAND2_X1 U10702 ( .A1(n12137), .A2(n10410), .ZN(n8309) );
  NAND2_X1 U10703 ( .A1(n8310), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10704 ( .A1(n8311), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8319) );
  INV_X1 U10705 ( .A(n8315), .ZN(n8314) );
  NAND2_X1 U10706 ( .A1(n8315), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10707 ( .A1(n8335), .A2(n8316), .ZN(n10595) );
  NAND2_X1 U10708 ( .A1(n8710), .A2(n10595), .ZN(n8318) );
  NAND2_X1 U10709 ( .A1(n8711), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8317) );
  NAND4_X1 U10710 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n10720) );
  NOR2_X1 U10711 ( .A1(n8324), .A2(n8533), .ZN(n8322) );
  MUX2_X1 U10712 ( .A(n8533), .B(n8322), .S(P3_IR_REG_5__SCAN_IN), .Z(n8326)
         );
  INV_X1 U10713 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10714 ( .A1(n8324), .A2(n8323), .ZN(n8361) );
  INV_X1 U10715 ( .A(n8361), .ZN(n8325) );
  INV_X1 U10716 ( .A(n9837), .ZN(n9874) );
  NAND2_X1 U10717 ( .A1(n8328), .A2(n8327), .ZN(n8330) );
  NAND2_X1 U10718 ( .A1(n9261), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8329) );
  XNOR2_X1 U10719 ( .A(n8342), .B(n8341), .ZN(n9269) );
  OR2_X1 U10720 ( .A1(n8529), .A2(n9269), .ZN(n8332) );
  OR2_X1 U10721 ( .A1(n8815), .A2(SI_5_), .ZN(n8331) );
  OAI211_X1 U10722 ( .C1(n9874), .C2(n9579), .A(n8332), .B(n8331), .ZN(n10862)
         );
  OR2_X1 U10723 ( .A1(n10720), .A2(n10862), .ZN(n11454) );
  NAND2_X1 U10724 ( .A1(n10720), .A2(n10862), .ZN(n11458) );
  NAND2_X1 U10725 ( .A1(n11454), .A2(n11458), .ZN(n8333) );
  INV_X1 U10726 ( .A(n8333), .ZN(n11588) );
  INV_X1 U10727 ( .A(n10720), .ZN(n10660) );
  NAND2_X1 U10728 ( .A1(n10660), .A2(n10862), .ZN(n8334) );
  NAND2_X1 U10729 ( .A1(n10741), .A2(n8334), .ZN(n10717) );
  INV_X1 U10730 ( .A(n10717), .ZN(n8351) );
  INV_X2 U10731 ( .A(n8644), .ZN(n8819) );
  NAND2_X1 U10732 ( .A1(n8819), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10733 ( .A1(n8311), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10734 ( .A1(n8335), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10735 ( .A1(n8355), .A2(n8336), .ZN(n10654) );
  NAND2_X1 U10736 ( .A1(n8710), .A2(n10654), .ZN(n8338) );
  NAND2_X1 U10737 ( .A1(n8711), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8337) );
  NAND4_X1 U10738 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n12136) );
  INV_X1 U10739 ( .A(SI_6_), .ZN(n9275) );
  OR2_X1 U10740 ( .A1(n8815), .A2(n9275), .ZN(n8349) );
  NAND2_X1 U10741 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  NAND2_X1 U10742 ( .A1(n9277), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8343) );
  XNOR2_X1 U10743 ( .A(n9281), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8345) );
  XNOR2_X1 U10744 ( .A(n6750), .B(n8345), .ZN(n9276) );
  OR2_X1 U10745 ( .A1(n8529), .A2(n9276), .ZN(n8348) );
  NAND2_X1 U10746 ( .A1(n8361), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8346) );
  OR2_X1 U10747 ( .A1(n9579), .A2(n9934), .ZN(n8347) );
  NAND2_X1 U10748 ( .A1(n12136), .A2(n10855), .ZN(n11460) );
  NAND2_X1 U10749 ( .A1(n8351), .A2(n8350), .ZN(n10719) );
  INV_X1 U10750 ( .A(n10855), .ZN(n10663) );
  NAND2_X1 U10751 ( .A1(n12136), .A2(n10663), .ZN(n8352) );
  NAND2_X1 U10752 ( .A1(n8819), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8360) );
  INV_X1 U10753 ( .A(n8355), .ZN(n8354) );
  NAND2_X1 U10754 ( .A1(n8355), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U10755 ( .A1(n8369), .A2(n8356), .ZN(n10871) );
  NAND2_X1 U10756 ( .A1(n8710), .A2(n10871), .ZN(n8358) );
  NAND2_X1 U10757 ( .A1(n8711), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8357) );
  NAND2_X1 U10758 ( .A1(n8378), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10759 ( .A(n8362), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U10760 ( .A1(n9282), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8365) );
  XNOR2_X1 U10761 ( .A(n9298), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8375) );
  XNOR2_X1 U10762 ( .A(n8377), .B(n8375), .ZN(n9286) );
  OR2_X1 U10763 ( .A1(n8529), .A2(n9286), .ZN(n8367) );
  OR2_X1 U10764 ( .A1(n8815), .A2(SI_7_), .ZN(n8366) );
  OAI211_X1 U10765 ( .C1(n10110), .C2(n9579), .A(n8367), .B(n8366), .ZN(n10838) );
  NAND2_X1 U10766 ( .A1(n11464), .A2(n11463), .ZN(n10830) );
  INV_X1 U10767 ( .A(n10838), .ZN(n10872) );
  NAND2_X1 U10768 ( .A1(n12037), .A2(n10872), .ZN(n8368) );
  NAND2_X1 U10769 ( .A1(n8819), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10770 ( .A1(n8311), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U10771 ( .A1(n8369), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10772 ( .A1(n8387), .A2(n8370), .ZN(n12038) );
  NAND2_X1 U10773 ( .A1(n8710), .A2(n12038), .ZN(n8372) );
  NAND2_X1 U10774 ( .A1(n8711), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8371) );
  NAND4_X1 U10775 ( .A1(n8374), .A2(n8373), .A3(n8372), .A4(n8371), .ZN(n12135) );
  INV_X1 U10776 ( .A(SI_8_), .ZN(n9294) );
  OR2_X1 U10777 ( .A1(n8815), .A2(n9294), .ZN(n8382) );
  INV_X1 U10778 ( .A(n8375), .ZN(n8376) );
  XNOR2_X1 U10779 ( .A(n8398), .B(n8397), .ZN(n9295) );
  OR2_X1 U10780 ( .A1(n8529), .A2(n9295), .ZN(n8381) );
  OAI21_X1 U10781 ( .B1(n8378), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U10782 ( .A(n8379), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10309) );
  OR2_X1 U10783 ( .A1(n9579), .A2(n10315), .ZN(n8380) );
  NAND2_X1 U10784 ( .A1(n12135), .A2(n14959), .ZN(n11469) );
  INV_X1 U10785 ( .A(n12135), .ZN(n10789) );
  NAND2_X1 U10786 ( .A1(n10789), .A2(n14959), .ZN(n8384) );
  NAND2_X1 U10787 ( .A1(n8819), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10788 ( .A1(n8311), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10789 ( .A1(n8387), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10790 ( .A1(n8404), .A2(n8388), .ZN(n11050) );
  NAND2_X1 U10791 ( .A1(n8710), .A2(n11050), .ZN(n8390) );
  NAND2_X1 U10792 ( .A1(n8711), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8389) );
  NAND4_X1 U10793 ( .A1(n8392), .A2(n8391), .A3(n8390), .A4(n8389), .ZN(n12134) );
  NAND2_X1 U10794 ( .A1(n8394), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8395) );
  INV_X1 U10795 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n15004) );
  XNOR2_X1 U10796 ( .A(n8395), .B(n15004), .ZN(n10487) );
  OR2_X1 U10797 ( .A1(n8815), .A2(SI_9_), .ZN(n8402) );
  NAND2_X1 U10798 ( .A1(n9315), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8399) );
  XNOR2_X1 U10799 ( .A(n9331), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n8416) );
  XNOR2_X1 U10800 ( .A(n8418), .B(n8416), .ZN(n9291) );
  OR2_X1 U10801 ( .A1(n8529), .A2(n9291), .ZN(n8401) );
  OAI211_X1 U10802 ( .C1(n10483), .C2(n9579), .A(n8402), .B(n8401), .ZN(n11474) );
  XNOR2_X1 U10803 ( .A(n12134), .B(n11474), .ZN(n11468) );
  NAND2_X1 U10804 ( .A1(n12134), .A2(n14967), .ZN(n8403) );
  NAND2_X1 U10805 ( .A1(n8311), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10806 ( .A1(n8819), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10807 ( .A1(n8404), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10808 ( .A1(n8424), .A2(n8405), .ZN(n11031) );
  NAND2_X1 U10809 ( .A1(n8710), .A2(n11031), .ZN(n8407) );
  NAND2_X1 U10810 ( .A1(n8711), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8406) );
  NAND4_X1 U10811 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n12133) );
  NOR2_X1 U10812 ( .A1(n8410), .A2(n8533), .ZN(n8411) );
  MUX2_X1 U10813 ( .A(n8533), .B(n8411), .S(P3_IR_REG_10__SCAN_IN), .Z(n8412)
         );
  INV_X1 U10814 ( .A(n8412), .ZN(n8415) );
  INV_X1 U10815 ( .A(n8413), .ZN(n8414) );
  NAND2_X1 U10816 ( .A1(n8415), .A2(n8414), .ZN(n12194) );
  INV_X1 U10817 ( .A(n12194), .ZN(n12144) );
  OR2_X1 U10818 ( .A1(n8815), .A2(SI_10_), .ZN(n8422) );
  INV_X1 U10819 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U10820 ( .A1(n15110), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8419) );
  XNOR2_X1 U10821 ( .A(n9389), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8430) );
  XNOR2_X1 U10822 ( .A(n8432), .B(n8430), .ZN(n9283) );
  OR2_X1 U10823 ( .A1(n8529), .A2(n9283), .ZN(n8421) );
  OAI211_X1 U10824 ( .C1(n12144), .C2(n9579), .A(n8422), .B(n8421), .ZN(n14972) );
  OR2_X1 U10825 ( .A1(n12133), .A2(n14972), .ZN(n11479) );
  NAND2_X1 U10826 ( .A1(n12133), .A2(n14972), .ZN(n11480) );
  NAND2_X1 U10827 ( .A1(n11479), .A2(n11480), .ZN(n11144) );
  INV_X1 U10828 ( .A(n14972), .ZN(n11150) );
  NAND2_X1 U10829 ( .A1(n12133), .A2(n11150), .ZN(n8423) );
  NAND2_X1 U10830 ( .A1(n8819), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U10831 ( .A1(n11401), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10832 ( .A1(n8424), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10833 ( .A1(n8448), .A2(n8425), .ZN(n11320) );
  NAND2_X1 U10834 ( .A1(n8710), .A2(n11320), .ZN(n8427) );
  NAND2_X1 U10835 ( .A1(n8711), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8426) );
  NAND4_X1 U10836 ( .A1(n8429), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(n12455) );
  INV_X1 U10837 ( .A(n8430), .ZN(n8431) );
  NAND2_X1 U10838 ( .A1(n9389), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8433) );
  XNOR2_X1 U10839 ( .A(n9541), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8435) );
  XNOR2_X1 U10840 ( .A(n8455), .B(n8435), .ZN(n9288) );
  OR2_X1 U10841 ( .A1(n8529), .A2(n9288), .ZN(n8443) );
  OR2_X1 U10842 ( .A1(n11411), .A2(SI_11_), .ZN(n8442) );
  NOR2_X1 U10843 ( .A1(n8413), .A2(n8533), .ZN(n8436) );
  MUX2_X1 U10844 ( .A(n8533), .B(n8436), .S(P3_IR_REG_11__SCAN_IN), .Z(n8437)
         );
  INV_X1 U10845 ( .A(n8437), .ZN(n8440) );
  AND2_X1 U10846 ( .A1(n8413), .A2(n8438), .ZN(n8461) );
  INV_X1 U10847 ( .A(n8461), .ZN(n8439) );
  NAND2_X1 U10848 ( .A1(n8440), .A2(n8439), .ZN(n12197) );
  OR2_X1 U10849 ( .A1(n9579), .A2(n14836), .ZN(n8441) );
  XNOR2_X1 U10850 ( .A(n12455), .B(n11105), .ZN(n11481) );
  INV_X1 U10851 ( .A(n12455), .ZN(n11231) );
  INV_X1 U10852 ( .A(n11105), .ZN(n11486) );
  NAND2_X1 U10853 ( .A1(n11231), .A2(n11486), .ZN(n8446) );
  NAND2_X1 U10854 ( .A1(n11401), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10855 ( .A1(n8711), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10856 ( .A1(n8448), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U10857 ( .A1(n8480), .A2(n8449), .ZN(n12460) );
  NAND2_X1 U10858 ( .A1(n8710), .A2(n12460), .ZN(n8451) );
  NAND2_X1 U10859 ( .A1(n8819), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8450) );
  NAND4_X1 U10860 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n12437) );
  NAND2_X1 U10861 ( .A1(n9541), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10862 ( .A1(n9644), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10863 ( .A1(n9623), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10864 ( .A1(n8467), .A2(n8457), .ZN(n8458) );
  NAND2_X1 U10865 ( .A1(n8459), .A2(n8458), .ZN(n8460) );
  NAND2_X1 U10866 ( .A1(n8468), .A2(n8460), .ZN(n9279) );
  OR2_X1 U10867 ( .A1(n8529), .A2(n9279), .ZN(n8466) );
  OR2_X1 U10868 ( .A1(n11411), .A2(n9280), .ZN(n8465) );
  OR2_X1 U10869 ( .A1(n8461), .A2(n8533), .ZN(n8463) );
  XNOR2_X1 U10870 ( .A(n8463), .B(n8462), .ZN(n14856) );
  OR2_X1 U10871 ( .A1(n9579), .A2(n14856), .ZN(n8464) );
  NAND2_X1 U10872 ( .A1(n12437), .A2(n12459), .ZN(n11490) );
  NAND2_X1 U10873 ( .A1(n11491), .A2(n11490), .ZN(n12452) );
  INV_X1 U10874 ( .A(n12459), .ZN(n11233) );
  INV_X1 U10875 ( .A(n8470), .ZN(n8471) );
  INV_X1 U10876 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U10877 ( .A1(n8471), .A2(n9720), .ZN(n8472) );
  NAND2_X1 U10878 ( .A1(n8487), .A2(n8472), .ZN(n9327) );
  NAND2_X1 U10879 ( .A1(n9327), .A2(n11409), .ZN(n8477) );
  INV_X1 U10880 ( .A(n9579), .ZN(n8590) );
  NAND2_X1 U10881 ( .A1(n8413), .A2(n8473), .ZN(n8474) );
  NAND2_X1 U10882 ( .A1(n8474), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8475) );
  XNOR2_X1 U10883 ( .A(n8475), .B(n8229), .ZN(n12201) );
  AOI22_X1 U10884 ( .A1(n8591), .A2(n9328), .B1(n8590), .B2(n12201), .ZN(n8476) );
  NAND2_X1 U10885 ( .A1(n8819), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U10886 ( .A1(n11401), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10887 ( .A1(n8480), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U10888 ( .A1(n8495), .A2(n8481), .ZN(n12440) );
  NAND2_X1 U10889 ( .A1(n8710), .A2(n12440), .ZN(n8483) );
  NAND2_X1 U10890 ( .A1(n8711), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8482) );
  NAND4_X1 U10891 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n12454) );
  OR2_X1 U10892 ( .A1(n12596), .A2(n12454), .ZN(n11497) );
  NAND2_X1 U10893 ( .A1(n12596), .A2(n12454), .ZN(n11496) );
  NAND2_X1 U10894 ( .A1(n11497), .A2(n11496), .ZN(n12434) );
  INV_X1 U10895 ( .A(n12454), .ZN(n11964) );
  OR2_X1 U10896 ( .A1(n12596), .A2(n11964), .ZN(n8486) );
  NAND2_X1 U10897 ( .A1(n10106), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10898 ( .A1(n10101), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8488) );
  OR2_X1 U10899 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  NAND2_X2 U10900 ( .A1(n8490), .A2(n8489), .ZN(n8504) );
  AND2_X1 U10901 ( .A1(n8504), .A2(n8491), .ZN(n9390) );
  NAND2_X1 U10902 ( .A1(n9390), .A2(n11409), .ZN(n8494) );
  NAND2_X1 U10903 ( .A1(n8509), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8492) );
  XNOR2_X1 U10904 ( .A(n8492), .B(P3_IR_REG_14__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U10905 ( .A1(n8591), .A2(SI_14_), .B1(n8590), .B2(n14905), .ZN(
        n8493) );
  NAND2_X1 U10906 ( .A1(n8819), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U10907 ( .A1(n11401), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10908 ( .A1(n8495), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10909 ( .A1(n8514), .A2(n8496), .ZN(n12426) );
  NAND2_X1 U10910 ( .A1(n8710), .A2(n12426), .ZN(n8498) );
  NAND2_X1 U10911 ( .A1(n8711), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8497) );
  NAND4_X1 U10912 ( .A1(n8500), .A2(n8499), .A3(n8498), .A4(n8497), .ZN(n12436) );
  NAND2_X1 U10913 ( .A1(n12592), .A2(n12436), .ZN(n11500) );
  NAND2_X1 U10914 ( .A1(n8501), .A2(n12409), .ZN(n11507) );
  NAND2_X1 U10915 ( .A1(n11500), .A2(n11507), .ZN(n12421) );
  NAND2_X1 U10916 ( .A1(n8501), .A2(n12436), .ZN(n8502) );
  NAND2_X1 U10917 ( .A1(n10338), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10918 ( .A1(n10415), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8505) );
  AND2_X1 U10919 ( .A1(n8524), .A2(n8508), .ZN(n9472) );
  NAND2_X1 U10920 ( .A1(n9472), .A2(n11409), .ZN(n8512) );
  OR2_X1 U10921 ( .A1(n8531), .A2(n8533), .ZN(n8510) );
  XNOR2_X1 U10922 ( .A(n8510), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14323) );
  AOI22_X1 U10923 ( .A1(n8591), .A2(SI_15_), .B1(n8590), .B2(n14323), .ZN(
        n8511) );
  AND2_X2 U10924 ( .A1(n8512), .A2(n8511), .ZN(n12588) );
  NAND2_X1 U10925 ( .A1(n8819), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10926 ( .A1(n11401), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10927 ( .A1(n8514), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10928 ( .A1(n8540), .A2(n8515), .ZN(n12414) );
  NAND2_X1 U10929 ( .A1(n8710), .A2(n12414), .ZN(n8517) );
  NAND2_X1 U10930 ( .A1(n8711), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8516) );
  NAND2_X1 U10931 ( .A1(n12588), .A2(n12398), .ZN(n8520) );
  NAND2_X1 U10932 ( .A1(n12407), .A2(n8520), .ZN(n8522) );
  INV_X1 U10933 ( .A(n12588), .ZN(n8754) );
  NAND2_X1 U10934 ( .A1(n8754), .A2(n12423), .ZN(n8521) );
  NAND2_X1 U10935 ( .A1(n10096), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10936 ( .A1(n15273), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8525) );
  OR2_X1 U10937 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  NAND2_X1 U10938 ( .A1(n8549), .A2(n8528), .ZN(n9530) );
  OR2_X1 U10939 ( .A1(n9530), .A2(n8529), .ZN(n8539) );
  INV_X1 U10940 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8530) );
  NOR2_X1 U10941 ( .A1(n8535), .A2(n8533), .ZN(n8532) );
  MUX2_X1 U10942 ( .A(n8533), .B(n8532), .S(P3_IR_REG_16__SCAN_IN), .Z(n8537)
         );
  INV_X1 U10943 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8534) );
  INV_X1 U10944 ( .A(n8568), .ZN(n8536) );
  AOI22_X1 U10945 ( .A1(n8591), .A2(SI_16_), .B1(n8590), .B2(n14326), .ZN(
        n8538) );
  NAND2_X1 U10946 ( .A1(n8539), .A2(n8538), .ZN(n11961) );
  NAND2_X1 U10947 ( .A1(n8819), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10948 ( .A1(n11401), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10949 ( .A1(n8540), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10950 ( .A1(n8556), .A2(n8541), .ZN(n12402) );
  NAND2_X1 U10951 ( .A1(n8710), .A2(n12402), .ZN(n8543) );
  NAND2_X1 U10952 ( .A1(n8711), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8542) );
  NAND4_X1 U10953 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n12384) );
  AND2_X1 U10954 ( .A1(n11961), .A2(n12384), .ZN(n8546) );
  NAND2_X1 U10955 ( .A1(n12584), .A2(n12410), .ZN(n8547) );
  NAND2_X1 U10956 ( .A1(n10198), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10957 ( .A1(n10228), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10958 ( .A1(n8565), .A2(n8550), .ZN(n8562) );
  XNOR2_X1 U10959 ( .A(n8564), .B(n8562), .ZN(n9624) );
  NAND2_X1 U10960 ( .A1(n9624), .A2(n11409), .ZN(n8553) );
  NAND2_X1 U10961 ( .A1(n8568), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U10962 ( .A(n8551), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U10963 ( .A1(n8591), .A2(SI_17_), .B1(n8590), .B2(n12210), .ZN(
        n8552) );
  NAND2_X1 U10964 ( .A1(n8819), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10965 ( .A1(n11401), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8560) );
  INV_X1 U10966 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10967 ( .A1(n8556), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10968 ( .A1(n8572), .A2(n8557), .ZN(n12388) );
  NAND2_X1 U10969 ( .A1(n8710), .A2(n12388), .ZN(n8559) );
  NAND2_X1 U10970 ( .A1(n8711), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8558) );
  OR2_X1 U10971 ( .A1(n12579), .A2(n12397), .ZN(n11517) );
  NAND2_X1 U10972 ( .A1(n12579), .A2(n12397), .ZN(n11524) );
  INV_X1 U10973 ( .A(n8562), .ZN(n8563) );
  INV_X1 U10974 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U10975 ( .A1(n10651), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8582) );
  INV_X1 U10976 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10653) );
  NAND2_X1 U10977 ( .A1(n10653), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10978 ( .A1(n8582), .A2(n8567), .ZN(n8579) );
  XNOR2_X1 U10979 ( .A(n8581), .B(n8579), .ZN(n9713) );
  NAND2_X1 U10980 ( .A1(n9713), .A2(n11409), .ZN(n8571) );
  NAND2_X1 U10981 ( .A1(n8588), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U10982 ( .A(n8569), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U10983 ( .A1(n8591), .A2(SI_18_), .B1(n8590), .B2(n12226), .ZN(
        n8570) );
  NAND2_X1 U10984 ( .A1(n8571), .A2(n8570), .ZN(n12101) );
  NAND2_X1 U10985 ( .A1(n8819), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U10986 ( .A1(n11401), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U10987 ( .A1(n8572), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U10988 ( .A1(n8596), .A2(n8573), .ZN(n12376) );
  NAND2_X1 U10989 ( .A1(n8710), .A2(n12376), .ZN(n8575) );
  NAND2_X1 U10990 ( .A1(n8711), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U10991 ( .A1(n12101), .A2(n12359), .ZN(n11523) );
  NAND2_X1 U10992 ( .A1(n12369), .A2(n12373), .ZN(n12368) );
  OR2_X1 U10993 ( .A1(n12101), .A2(n12385), .ZN(n8578) );
  NAND2_X1 U10994 ( .A1(n12368), .A2(n8578), .ZN(n12357) );
  INV_X1 U10995 ( .A(n8579), .ZN(n8580) );
  NAND2_X1 U10996 ( .A1(n10772), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10997 ( .A1(n10770), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8584) );
  OR2_X1 U10998 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U10999 ( .A1(n8603), .A2(n8587), .ZN(n9718) );
  NAND2_X1 U11000 ( .A1(n9718), .A2(n11409), .ZN(n8593) );
  AOI22_X1 U11001 ( .A1(n8591), .A2(n9717), .B1(n8590), .B2(n12237), .ZN(n8592) );
  NAND2_X1 U11002 ( .A1(n11401), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11003 ( .A1(n8819), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8600) );
  INV_X1 U11004 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U11005 ( .A1(n8596), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11006 ( .A1(n8606), .A2(n8597), .ZN(n12363) );
  NAND2_X1 U11007 ( .A1(n8710), .A2(n12363), .ZN(n8599) );
  NAND2_X1 U11008 ( .A1(n8711), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8598) );
  AND2_X1 U11009 ( .A1(n12572), .A2(n12370), .ZN(n11583) );
  XNOR2_X2 U11010 ( .A(n8615), .B(n11043), .ZN(n8614) );
  XNOR2_X1 U11011 ( .A(n8614), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U11012 ( .A1(n10199), .A2(n11409), .ZN(n8605) );
  OR2_X1 U11013 ( .A1(n11411), .A2(n10201), .ZN(n8604) );
  NAND2_X1 U11014 ( .A1(n11401), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8611) );
  NAND2_X1 U11015 ( .A1(n8711), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U11016 ( .A1(n8606), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U11017 ( .A1(n8623), .A2(n8607), .ZN(n12352) );
  NAND2_X1 U11018 ( .A1(n8710), .A2(n12352), .ZN(n8609) );
  NAND2_X1 U11019 ( .A1(n8819), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U11020 ( .A1(n12344), .A2(n12351), .ZN(n8613) );
  NAND2_X1 U11021 ( .A1(n12509), .A2(n12131), .ZN(n8612) );
  INV_X1 U11022 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U11023 ( .A1(n11223), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U11024 ( .A1(n11221), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8618) );
  AND2_X1 U11025 ( .A1(n8634), .A2(n8618), .ZN(n8631) );
  XNOR2_X1 U11026 ( .A(n8633), .B(n8631), .ZN(n10294) );
  NAND2_X1 U11027 ( .A1(n10294), .A2(n11409), .ZN(n8620) );
  INV_X1 U11028 ( .A(SI_21_), .ZN(n10295) );
  OR2_X1 U11029 ( .A1(n11411), .A2(n10295), .ZN(n8619) );
  INV_X1 U11030 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11031 ( .A1(n8623), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11032 ( .A1(n8639), .A2(n8624), .ZN(n12339) );
  NAND2_X1 U11033 ( .A1(n12339), .A2(n8710), .ZN(n8628) );
  NAND2_X1 U11034 ( .A1(n8819), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11035 ( .A1(n11401), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11036 ( .A1(n8711), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8625) );
  NAND4_X1 U11037 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n12345) );
  AND2_X1 U11038 ( .A1(n12338), .A2(n12345), .ZN(n8629) );
  OR2_X1 U11039 ( .A1(n12338), .A2(n12345), .ZN(n8630) );
  INV_X1 U11040 ( .A(n8631), .ZN(n8632) );
  INV_X1 U11041 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8635) );
  XNOR2_X1 U11042 ( .A(n8635), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8647) );
  XNOR2_X1 U11043 ( .A(n8648), .B(n8647), .ZN(n10468) );
  NAND2_X1 U11044 ( .A1(n10468), .A2(n11409), .ZN(n8638) );
  OR2_X1 U11045 ( .A1(n11411), .A2(n8636), .ZN(n8637) );
  INV_X1 U11046 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12503) );
  NAND2_X1 U11047 ( .A1(n8639), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U11048 ( .A1(n8651), .A2(n8640), .ZN(n12328) );
  NAND2_X1 U11049 ( .A1(n12328), .A2(n8710), .ZN(n8643) );
  AOI22_X1 U11050 ( .A1(n11401), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n8711), 
        .B2(P3_REG2_REG_22__SCAN_IN), .ZN(n8642) );
  OAI211_X1 U11051 ( .C1(n8644), .C2(n12503), .A(n8643), .B(n8642), .ZN(n12310) );
  NOR2_X1 U11052 ( .A1(n12327), .A2(n12310), .ZN(n8645) );
  NAND2_X1 U11053 ( .A1(n12327), .A2(n12310), .ZN(n8646) );
  XNOR2_X1 U11054 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8659) );
  XNOR2_X1 U11055 ( .A(n8660), .B(n8659), .ZN(n10712) );
  NAND2_X1 U11056 ( .A1(n10712), .A2(n11409), .ZN(n8650) );
  OR2_X1 U11057 ( .A1(n11411), .A2(n10714), .ZN(n8649) );
  NAND2_X1 U11058 ( .A1(n8651), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11059 ( .A1(n8669), .A2(n8652), .ZN(n12312) );
  NAND2_X1 U11060 ( .A1(n12312), .A2(n8710), .ZN(n8655) );
  AOI22_X1 U11061 ( .A1(n11401), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n8711), 
        .B2(P3_REG2_REG_23__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U11062 ( .A1(n8819), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11063 ( .A1(n12496), .A2(n12324), .ZN(n8656) );
  NAND2_X1 U11064 ( .A1(n11548), .A2(n8656), .ZN(n8756) );
  NAND2_X1 U11065 ( .A1(n12308), .A2(n8756), .ZN(n8658) );
  NAND2_X1 U11066 ( .A1(n12496), .A2(n12297), .ZN(n8657) );
  NAND2_X1 U11067 ( .A1(n11373), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11068 ( .A1(n8663), .A2(n11388), .ZN(n8664) );
  INV_X1 U11069 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11954) );
  XNOR2_X1 U11070 ( .A(n8674), .B(n11954), .ZN(n10956) );
  NAND2_X1 U11071 ( .A1(n10956), .A2(n11409), .ZN(n8666) );
  INV_X1 U11072 ( .A(SI_24_), .ZN(n10957) );
  OR2_X1 U11073 ( .A1(n11411), .A2(n10957), .ZN(n8665) );
  INV_X1 U11074 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12299) );
  INV_X1 U11075 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11076 ( .A1(n8669), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11077 ( .A1(n8680), .A2(n8670), .ZN(n12298) );
  NAND2_X1 U11078 ( .A1(n12298), .A2(n8710), .ZN(n8672) );
  AOI22_X1 U11079 ( .A1(n11401), .A2(P3_REG0_REG_24__SCAN_IN), .B1(n8819), 
        .B2(P3_REG1_REG_24__SCAN_IN), .ZN(n8671) );
  OAI211_X1 U11080 ( .C1(n8673), .C2(n12299), .A(n8672), .B(n8671), .ZN(n12309) );
  XNOR2_X1 U11081 ( .A(n13273), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8688) );
  XNOR2_X1 U11082 ( .A(n8689), .B(n8688), .ZN(n11136) );
  NAND2_X1 U11083 ( .A1(n11136), .A2(n11409), .ZN(n8677) );
  OR2_X1 U11084 ( .A1(n11411), .A2(n11138), .ZN(n8676) );
  NAND2_X2 U11085 ( .A1(n8677), .A2(n8676), .ZN(n12486) );
  INV_X1 U11086 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11087 ( .A1(n8680), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11088 ( .A1(n8694), .A2(n8681), .ZN(n12287) );
  NAND2_X1 U11089 ( .A1(n12287), .A2(n8710), .ZN(n8687) );
  INV_X1 U11090 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12556) );
  NAND2_X1 U11091 ( .A1(n8819), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U11092 ( .A1(n8711), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8683) );
  OAI211_X1 U11093 ( .C1(n8823), .C2(n12556), .A(n8684), .B(n8683), .ZN(n8685)
         );
  INV_X1 U11094 ( .A(n8685), .ZN(n8686) );
  NAND2_X1 U11095 ( .A1(n12486), .A2(n12274), .ZN(n8757) );
  AND2_X2 U11096 ( .A1(n11424), .A2(n8757), .ZN(n12291) );
  NAND2_X1 U11097 ( .A1(n13273), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8690) );
  XNOR2_X1 U11098 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8691) );
  XNOR2_X1 U11099 ( .A(n8701), .B(n8691), .ZN(n11237) );
  NAND2_X2 U11100 ( .A1(n8693), .A2(n8692), .ZN(n12277) );
  NAND2_X1 U11101 ( .A1(n8694), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U11102 ( .A1(n8708), .A2(n8695), .ZN(n12278) );
  NAND2_X1 U11103 ( .A1(n12278), .A2(n8710), .ZN(n8700) );
  INV_X1 U11104 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U11105 ( .A1(n8819), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11106 ( .A1(n8711), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8696) );
  OAI211_X1 U11107 ( .C1(n8823), .C2(n12552), .A(n8697), .B(n8696), .ZN(n8698)
         );
  INV_X1 U11108 ( .A(n8698), .ZN(n8699) );
  NAND2_X2 U11109 ( .A1(n8700), .A2(n8699), .ZN(n12285) );
  NAND2_X1 U11110 ( .A1(n14146), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8702) );
  INV_X1 U11111 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U11112 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13266), .B2(n14144), .ZN(n8703) );
  INV_X1 U11113 ( .A(SI_27_), .ZN(n15059) );
  INV_X1 U11114 ( .A(n8708), .ZN(n8707) );
  INV_X1 U11115 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11116 ( .A1(n8708), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11117 ( .A1(n8726), .A2(n8709), .ZN(n12266) );
  NAND2_X1 U11118 ( .A1(n12266), .A2(n8312), .ZN(n8716) );
  INV_X1 U11119 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U11120 ( .A1(n8819), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11121 ( .A1(n8711), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8712) );
  OAI211_X1 U11122 ( .C1(n8823), .C2(n12549), .A(n8713), .B(n8712), .ZN(n8714)
         );
  INV_X1 U11123 ( .A(n8714), .ZN(n8715) );
  XNOR2_X2 U11124 ( .A(n12477), .B(n12130), .ZN(n11605) );
  OR2_X1 U11125 ( .A1(n12477), .A2(n12130), .ZN(n8718) );
  NAND2_X1 U11126 ( .A1(n13266), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8720) );
  AOI22_X1 U11127 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13264), .B2(n11390), .ZN(n8722) );
  INV_X1 U11128 ( .A(n8722), .ZN(n8723) );
  XNOR2_X1 U11129 ( .A(n8814), .B(n8723), .ZN(n12605) );
  NAND2_X1 U11130 ( .A1(n12605), .A2(n11409), .ZN(n8725) );
  OR2_X1 U11131 ( .A1(n11411), .A2(n12607), .ZN(n8724) );
  NAND2_X1 U11132 ( .A1(n8726), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U11133 ( .A1(n8741), .A2(n8727), .ZN(n12249) );
  INV_X1 U11134 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n15211) );
  NAND2_X1 U11135 ( .A1(n8819), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11136 ( .A1(n8711), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8728) );
  OAI211_X1 U11137 ( .C1(n8823), .C2(n15211), .A(n8729), .B(n8728), .ZN(n8730)
         );
  NAND2_X1 U11138 ( .A1(n12253), .A2(n12261), .ZN(n11567) );
  INV_X1 U11139 ( .A(n8767), .ZN(n8732) );
  NAND2_X1 U11140 ( .A1(n8732), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11141 ( .A1(n12222), .A2(n11619), .ZN(n8739) );
  NAND2_X1 U11142 ( .A1(n8731), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8735) );
  INV_X1 U11143 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U11144 ( .A1(n8736), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U11145 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8737), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8738) );
  AND2_X1 U11146 ( .A1(n8738), .A2(n8731), .ZN(n8803) );
  NAND2_X1 U11147 ( .A1(n11428), .A2(n8803), .ZN(n10039) );
  INV_X1 U11148 ( .A(n8741), .ZN(n11955) );
  NAND2_X1 U11149 ( .A1(n11955), .A2(n8710), .ZN(n11406) );
  INV_X1 U11150 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11151 ( .A1(n8819), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11152 ( .A1(n8711), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8742) );
  OAI211_X1 U11153 ( .C1(n8823), .C2(n8832), .A(n8743), .B(n8742), .ZN(n8744)
         );
  INV_X1 U11154 ( .A(n8744), .ZN(n8745) );
  INV_X1 U11155 ( .A(n6831), .ZN(n8826) );
  NAND2_X1 U11156 ( .A1(n8826), .A2(n12223), .ZN(n9591) );
  NAND2_X1 U11157 ( .A1(n9579), .A2(n9591), .ZN(n8747) );
  AND2_X2 U11158 ( .A1(n11619), .A2(n11428), .ZN(n11569) );
  INV_X1 U11159 ( .A(n12130), .ZN(n12273) );
  NAND3_X1 U11160 ( .A1(n9579), .A2(n9591), .A3(n11569), .ZN(n14941) );
  OAI22_X1 U11161 ( .A1(n12026), .A2(n14943), .B1(n12273), .B2(n14941), .ZN(
        n8748) );
  INV_X1 U11162 ( .A(n8748), .ZN(n8749) );
  INV_X1 U11163 ( .A(n10474), .ZN(n10100) );
  NAND2_X1 U11164 ( .A1(n14930), .A2(n11436), .ZN(n10042) );
  NAND2_X1 U11165 ( .A1(n14914), .A2(n11438), .ZN(n10169) );
  NAND2_X1 U11166 ( .A1(n10740), .A2(n11588), .ZN(n10739) );
  NAND2_X1 U11167 ( .A1(n10739), .A2(n11454), .ZN(n10716) );
  NAND2_X1 U11168 ( .A1(n10716), .A2(n11594), .ZN(n10715) );
  INV_X1 U11169 ( .A(n10830), .ZN(n11589) );
  INV_X1 U11170 ( .A(n12134), .ZN(n11473) );
  OR2_X1 U11171 ( .A1(n12455), .A2(n11486), .ZN(n11485) );
  INV_X1 U11172 ( .A(n12452), .ZN(n12449) );
  INV_X1 U11173 ( .A(n11497), .ZN(n8753) );
  NAND2_X1 U11174 ( .A1(n12588), .A2(n12423), .ZN(n11502) );
  NAND2_X1 U11175 ( .A1(n8754), .A2(n12398), .ZN(n11508) );
  NAND2_X1 U11176 ( .A1(n12584), .A2(n12384), .ZN(n11513) );
  NAND2_X1 U11177 ( .A1(n11961), .A2(n12410), .ZN(n11511) );
  AND2_X1 U11178 ( .A1(n12572), .A2(n12346), .ZN(n11521) );
  OR2_X1 U11179 ( .A1(n12572), .A2(n12346), .ZN(n11522) );
  OR2_X1 U11180 ( .A1(n12509), .A2(n12360), .ZN(n11534) );
  NAND2_X1 U11181 ( .A1(n12338), .A2(n12323), .ZN(n11539) );
  OR2_X1 U11182 ( .A1(n12338), .A2(n12323), .ZN(n11538) );
  INV_X1 U11183 ( .A(n12310), .ZN(n12335) );
  NAND2_X1 U11184 ( .A1(n12327), .A2(n12335), .ZN(n11543) );
  NAND2_X1 U11185 ( .A1(n12325), .A2(n11543), .ZN(n8755) );
  NAND2_X1 U11186 ( .A1(n8755), .A2(n11542), .ZN(n12317) );
  NAND2_X1 U11187 ( .A1(n12318), .A2(n11548), .ZN(n12304) );
  OR2_X1 U11188 ( .A1(n12492), .A2(n12054), .ZN(n11550) );
  INV_X1 U11189 ( .A(n8757), .ZN(n11426) );
  AND2_X1 U11190 ( .A1(n12477), .A2(n12273), .ZN(n11565) );
  XNOR2_X1 U11191 ( .A(n8830), .B(n11563), .ZN(n12254) );
  NAND2_X1 U11192 ( .A1(n11619), .A2(n10202), .ZN(n8758) );
  AOI21_X1 U11193 ( .B1(n12222), .B2(n8758), .A(n11428), .ZN(n8761) );
  NAND2_X1 U11194 ( .A1(n11433), .A2(n10202), .ZN(n8759) );
  AND2_X1 U11195 ( .A1(n8804), .A2(n8759), .ZN(n8760) );
  OR2_X1 U11196 ( .A1(n8761), .A2(n8760), .ZN(n9972) );
  NOR2_X1 U11197 ( .A1(n11580), .A2(n14966), .ZN(n8762) );
  NAND2_X1 U11198 ( .A1(n9972), .A2(n8762), .ZN(n8764) );
  AND2_X1 U11199 ( .A1(n11619), .A2(n8803), .ZN(n8763) );
  NAND2_X1 U11200 ( .A1(n12237), .A2(n8763), .ZN(n8798) );
  OR2_X1 U11201 ( .A1(n11613), .A2(n11619), .ZN(n12478) );
  NAND2_X1 U11202 ( .A1(n12254), .A2(n14963), .ZN(n8765) );
  NAND2_X1 U11203 ( .A1(n12248), .A2(n8765), .ZN(n8810) );
  XNOR2_X1 U11204 ( .A(n8777), .B(P3_B_REG_SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11205 ( .A1(n8772), .A2(n11137), .ZN(n8776) );
  NAND2_X1 U11206 ( .A1(n8774), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11207 ( .A1(n8777), .A2(n11240), .ZN(n8779) );
  OR2_X1 U11208 ( .A1(n8780), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U11209 ( .A1(n11137), .A2(n11240), .ZN(n8781) );
  NAND2_X1 U11210 ( .A1(n10040), .A2(n10283), .ZN(n8802) );
  NOR2_X1 U11211 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .ZN(
        n15218) );
  NOR4_X1 U11212 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8785) );
  NOR4_X1 U11213 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8784) );
  NOR4_X1 U11214 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8783) );
  NAND4_X1 U11215 ( .A1(n15218), .A2(n8785), .A3(n8784), .A4(n8783), .ZN(n8791) );
  NOR4_X1 U11216 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8789) );
  NOR4_X1 U11217 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8788) );
  NOR4_X1 U11218 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8787) );
  NOR4_X1 U11219 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8786) );
  NAND4_X1 U11220 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8790)
         );
  NOR2_X1 U11221 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  OR2_X1 U11222 ( .A1(n8780), .A2(n8792), .ZN(n8801) );
  NAND2_X1 U11223 ( .A1(n6719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8794) );
  AND2_X1 U11224 ( .A1(n8801), .A2(n9982), .ZN(n8795) );
  NAND2_X1 U11225 ( .A1(n8802), .A2(n8795), .ZN(n10285) );
  OAI22_X1 U11226 ( .A1(n12222), .A2(n8804), .B1(n8803), .B2(n14971), .ZN(
        n8796) );
  AOI21_X1 U11227 ( .B1(n8796), .B2(n11580), .A(n11569), .ZN(n8797) );
  NOR2_X1 U11228 ( .A1(n10040), .A2(n8797), .ZN(n8800) );
  NAND2_X1 U11229 ( .A1(n11580), .A2(n11569), .ZN(n9961) );
  NAND2_X1 U11230 ( .A1(n8798), .A2(n11577), .ZN(n10281) );
  NOR2_X1 U11231 ( .A1(n10283), .A2(n10282), .ZN(n8799) );
  INV_X1 U11232 ( .A(n12253), .ZN(n8811) );
  INV_X1 U11233 ( .A(n8801), .ZN(n8806) );
  INV_X1 U11234 ( .A(n9972), .ZN(n8808) );
  OR2_X1 U11235 ( .A1(n11580), .A2(n11577), .ZN(n9988) );
  NAND2_X1 U11236 ( .A1(n11433), .A2(n8803), .ZN(n11611) );
  NOR2_X1 U11237 ( .A1(n8804), .A2(n11611), .ZN(n8805) );
  NAND2_X1 U11238 ( .A1(n12222), .A2(n8805), .ZN(n9974) );
  AND2_X1 U11239 ( .A1(n9988), .A2(n9974), .ZN(n8807) );
  OR3_X1 U11240 ( .A1(n10040), .A2(n10283), .A3(n8806), .ZN(n9984) );
  OAI22_X1 U11241 ( .A1(n9979), .A2(n8808), .B1(n8807), .B2(n9984), .ZN(n8809)
         );
  NOR2_X1 U11242 ( .A1(n11390), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U11243 ( .A(n14141), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n11392) );
  XNOR2_X1 U11244 ( .A(n11394), .B(n11392), .ZN(n11625) );
  NAND2_X1 U11245 ( .A1(n11625), .A2(n11409), .ZN(n8817) );
  INV_X1 U11246 ( .A(SI_29_), .ZN(n11626) );
  OR2_X1 U11247 ( .A1(n11411), .A2(n11626), .ZN(n8816) );
  NAND2_X1 U11248 ( .A1(n11959), .A2(n12026), .ZN(n11572) );
  INV_X1 U11249 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11250 ( .A1(n8819), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11251 ( .A1(n8711), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U11252 ( .C1(n8823), .C2(n8822), .A(n8821), .B(n8820), .ZN(n8824)
         );
  INV_X1 U11253 ( .A(n8824), .ZN(n8825) );
  AND2_X1 U11254 ( .A1(n11406), .A2(n8825), .ZN(n11417) );
  AND2_X1 U11255 ( .A1(n8826), .A2(P3_B_REG_SCAN_IN), .ZN(n8827) );
  OR2_X1 U11256 ( .A1(n14943), .A2(n8827), .ZN(n12242) );
  OAI22_X1 U11257 ( .A1(n12261), .A2(n14941), .B1(n11417), .B2(n12242), .ZN(
        n8828) );
  AOI21_X2 U11258 ( .B1(n8829), .B2(n12450), .A(n8828), .ZN(n11960) );
  INV_X1 U11259 ( .A(n11566), .ZN(n11570) );
  NAND2_X1 U11260 ( .A1(n8837), .A2(n14979), .ZN(n8836) );
  INV_X1 U11261 ( .A(n11959), .ZN(n8839) );
  NOR2_X1 U11262 ( .A1(n14979), .A2(n8832), .ZN(n8833) );
  NAND2_X1 U11263 ( .A1(n8836), .A2(n8835), .ZN(P3_U3456) );
  INV_X1 U11264 ( .A(n8837), .ZN(n8842) );
  INV_X1 U11265 ( .A(n8840), .ZN(n8841) );
  OAI21_X1 U11266 ( .B1(n8842), .B2(n14986), .A(n8841), .ZN(P3_U3488) );
  AND2_X1 U11267 ( .A1(n12975), .A2(n8843), .ZN(n8845) );
  OAI211_X1 U11268 ( .C1(n8845), .C2(n9119), .A(n8844), .B(n14753), .ZN(n8846)
         );
  AOI22_X1 U11269 ( .A1(n12823), .A2(n12801), .B1(n12825), .B2(n12800), .ZN(
        n12710) );
  NAND2_X1 U11270 ( .A1(n12708), .A2(n14734), .ZN(n8847) );
  AOI211_X1 U11271 ( .C1(n13144), .C2(n12970), .A(n13104), .B(n7130), .ZN(
        n13143) );
  OAI22_X1 U11272 ( .A1(n8852), .A2(n14739), .B1(n6558), .B2(n8851), .ZN(n8853) );
  AOI21_X1 U11273 ( .B1(n13143), .B2(n14731), .A(n8853), .ZN(n8854) );
  INV_X1 U11274 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U11275 ( .A1(n8859), .A2(n8858), .ZN(n8863) );
  INV_X1 U11276 ( .A(n8862), .ZN(n8860) );
  NAND2_X1 U11277 ( .A1(n7542), .A2(n8860), .ZN(n8866) );
  OAI211_X1 U11278 ( .C1(n8863), .C2(n14747), .A(n8862), .B(n8898), .ZN(n8865)
         );
  NAND2_X1 U11279 ( .A1(n9676), .A2(n8902), .ZN(n8864) );
  NAND3_X1 U11280 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8873) );
  NAND2_X1 U11281 ( .A1(n8178), .A2(n8898), .ZN(n8868) );
  NAND2_X1 U11282 ( .A1(n8869), .A2(n8902), .ZN(n8867) );
  NAND2_X1 U11283 ( .A1(n8868), .A2(n8867), .ZN(n8872) );
  AOI22_X1 U11284 ( .A1(n8178), .A2(n8902), .B1(n8898), .B2(n8869), .ZN(n8870)
         );
  AOI21_X1 U11285 ( .B1(n8873), .B2(n8872), .A(n8870), .ZN(n8871) );
  NAND2_X1 U11286 ( .A1(n8876), .A2(n8902), .ZN(n8875) );
  NAND2_X1 U11287 ( .A1(n9765), .A2(n8898), .ZN(n8874) );
  NAND2_X1 U11288 ( .A1(n8875), .A2(n8874), .ZN(n8878) );
  AOI22_X1 U11289 ( .A1(n8876), .A2(n8898), .B1(n8902), .B2(n9765), .ZN(n8877)
         );
  NAND2_X1 U11290 ( .A1(n12849), .A2(n8999), .ZN(n8880) );
  NAND2_X1 U11291 ( .A1(n9757), .A2(n9013), .ZN(n8879) );
  NAND2_X1 U11292 ( .A1(n8880), .A2(n8879), .ZN(n8883) );
  AOI22_X1 U11293 ( .A1(n12849), .A2(n9013), .B1(n8999), .B2(n9757), .ZN(n8881) );
  INV_X1 U11294 ( .A(n8882), .ZN(n8885) );
  AOI22_X1 U11295 ( .A1(n12848), .A2(n9013), .B1(n6561), .B2(n14794), .ZN(
        n8888) );
  NAND2_X1 U11296 ( .A1(n12848), .A2(n6561), .ZN(n8886) );
  OAI21_X1 U11297 ( .B1(n9956), .B2(n8999), .A(n8886), .ZN(n8887) );
  NAND2_X1 U11298 ( .A1(n10060), .A2(n9013), .ZN(n8890) );
  NAND2_X1 U11299 ( .A1(n12847), .A2(n8999), .ZN(n8889) );
  NAND2_X1 U11300 ( .A1(n8890), .A2(n8889), .ZN(n8893) );
  AOI22_X1 U11301 ( .A1(n8999), .A2(n10060), .B1(n12847), .B2(n9013), .ZN(
        n8891) );
  AOI21_X1 U11302 ( .B1(n8894), .B2(n8893), .A(n8891), .ZN(n8892) );
  NOR2_X1 U11303 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  NAND2_X1 U11304 ( .A1(n10219), .A2(n8999), .ZN(n8897) );
  NAND2_X1 U11305 ( .A1(n12846), .A2(n9013), .ZN(n8896) );
  NAND2_X1 U11306 ( .A1(n10219), .A2(n9013), .ZN(n8899) );
  OAI21_X1 U11307 ( .B1(n9013), .B2(n10193), .A(n8899), .ZN(n8900) );
  NAND2_X1 U11308 ( .A1(n10552), .A2(n9013), .ZN(n8904) );
  NAND2_X1 U11309 ( .A1(n12845), .A2(n8999), .ZN(n8903) );
  NAND2_X1 U11310 ( .A1(n8904), .A2(n8903), .ZN(n8907) );
  AOI22_X1 U11311 ( .A1(n10552), .A2(n8999), .B1(n9013), .B2(n12845), .ZN(
        n8905) );
  NOR2_X1 U11312 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  NAND2_X1 U11313 ( .A1(n10680), .A2(n8999), .ZN(n8912) );
  NAND2_X1 U11314 ( .A1(n12844), .A2(n9013), .ZN(n8911) );
  NAND2_X1 U11315 ( .A1(n10680), .A2(n9013), .ZN(n8913) );
  OAI21_X1 U11316 ( .B1(n9013), .B2(n10424), .A(n8913), .ZN(n8914) );
  NAND2_X1 U11317 ( .A1(n6569), .A2(n9013), .ZN(n8917) );
  NAND2_X1 U11318 ( .A1(n12843), .A2(n8999), .ZN(n8916) );
  NAND2_X1 U11319 ( .A1(n8917), .A2(n8916), .ZN(n8919) );
  AOI22_X1 U11320 ( .A1(n6569), .A2(n6561), .B1(n9013), .B2(n12843), .ZN(n8918) );
  NAND2_X1 U11321 ( .A1(n10979), .A2(n8999), .ZN(n8921) );
  NAND2_X1 U11322 ( .A1(n12842), .A2(n9013), .ZN(n8920) );
  NAND2_X1 U11323 ( .A1(n8921), .A2(n8920), .ZN(n8923) );
  AOI22_X1 U11324 ( .A1(n10979), .A2(n9013), .B1(n8999), .B2(n12842), .ZN(
        n8922) );
  NAND2_X1 U11325 ( .A1(n11027), .A2(n9013), .ZN(n8925) );
  NAND2_X1 U11326 ( .A1(n12841), .A2(n8999), .ZN(n8924) );
  NAND2_X1 U11327 ( .A1(n8925), .A2(n8924), .ZN(n8931) );
  NAND2_X1 U11328 ( .A1(n8930), .A2(n8931), .ZN(n8929) );
  NAND2_X1 U11329 ( .A1(n11027), .A2(n8999), .ZN(n8926) );
  OAI21_X1 U11330 ( .B1(n8927), .B2(n6561), .A(n8926), .ZN(n8928) );
  NAND2_X1 U11331 ( .A1(n8929), .A2(n8928), .ZN(n8935) );
  NAND2_X1 U11332 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U11333 ( .A1(n8935), .A2(n8934), .ZN(n8940) );
  NAND2_X1 U11334 ( .A1(n14689), .A2(n6561), .ZN(n8937) );
  NAND2_X1 U11335 ( .A1(n12840), .A2(n9013), .ZN(n8936) );
  NAND2_X1 U11336 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  AOI22_X1 U11337 ( .A1(n14689), .A2(n9013), .B1(n6561), .B2(n12840), .ZN(
        n8938) );
  AOI21_X1 U11338 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n8942) );
  NOR2_X1 U11339 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  OR2_X1 U11340 ( .A1(n8942), .A2(n8941), .ZN(n8947) );
  NAND2_X1 U11341 ( .A1(n14410), .A2(n9013), .ZN(n8944) );
  NAND2_X1 U11342 ( .A1(n12839), .A2(n8999), .ZN(n8943) );
  NAND2_X1 U11343 ( .A1(n8944), .A2(n8943), .ZN(n8948) );
  NAND2_X1 U11344 ( .A1(n14410), .A2(n8999), .ZN(n8945) );
  OAI21_X1 U11345 ( .B1(n14379), .B2(n8999), .A(n8945), .ZN(n8946) );
  NAND2_X1 U11346 ( .A1(n14396), .A2(n8999), .ZN(n8950) );
  NAND2_X1 U11347 ( .A1(n12838), .A2(n9013), .ZN(n8949) );
  NAND2_X1 U11348 ( .A1(n8950), .A2(n8949), .ZN(n8952) );
  AOI22_X1 U11349 ( .A1(n14396), .A2(n9013), .B1(n8999), .B2(n12838), .ZN(
        n8951) );
  AOI21_X1 U11350 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8955) );
  NAND2_X1 U11351 ( .A1(n13228), .A2(n9013), .ZN(n8957) );
  NAND2_X1 U11352 ( .A1(n12837), .A2(n8999), .ZN(n8956) );
  NAND2_X1 U11353 ( .A1(n8957), .A2(n8956), .ZN(n8962) );
  NAND2_X1 U11354 ( .A1(n8961), .A2(n8962), .ZN(n8960) );
  NAND2_X1 U11355 ( .A1(n13228), .A2(n6561), .ZN(n8958) );
  OAI21_X1 U11356 ( .B1(n14380), .B2(n6561), .A(n8958), .ZN(n8959) );
  NAND2_X1 U11357 ( .A1(n8960), .A2(n8959), .ZN(n8966) );
  INV_X1 U11358 ( .A(n8961), .ZN(n8964) );
  INV_X1 U11359 ( .A(n8962), .ZN(n8963) );
  NAND2_X1 U11360 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  NAND2_X1 U11361 ( .A1(n8966), .A2(n8965), .ZN(n8971) );
  NAND2_X1 U11362 ( .A1(n13219), .A2(n6561), .ZN(n8968) );
  NAND2_X1 U11363 ( .A1(n12836), .A2(n9013), .ZN(n8967) );
  NAND2_X1 U11364 ( .A1(n8968), .A2(n8967), .ZN(n8970) );
  INV_X1 U11365 ( .A(n8970), .ZN(n8969) );
  AOI22_X1 U11366 ( .A1(n13219), .A2(n9013), .B1(n6561), .B2(n12836), .ZN(
        n8972) );
  INV_X1 U11367 ( .A(n8972), .ZN(n8973) );
  NAND2_X1 U11368 ( .A1(n13213), .A2(n9013), .ZN(n8975) );
  NAND2_X1 U11369 ( .A1(n12835), .A2(n6561), .ZN(n8974) );
  NAND2_X1 U11370 ( .A1(n8975), .A2(n8974), .ZN(n8977) );
  AOI22_X1 U11371 ( .A1(n13213), .A2(n6561), .B1(n9013), .B2(n12835), .ZN(
        n8976) );
  NAND2_X1 U11372 ( .A1(n13206), .A2(n8999), .ZN(n8980) );
  NAND2_X1 U11373 ( .A1(n12834), .A2(n9013), .ZN(n8979) );
  NAND2_X1 U11374 ( .A1(n13206), .A2(n9013), .ZN(n8981) );
  NAND2_X1 U11375 ( .A1(n13078), .A2(n9013), .ZN(n8984) );
  NAND2_X1 U11376 ( .A1(n12833), .A2(n6561), .ZN(n8983) );
  NAND2_X1 U11377 ( .A1(n8984), .A2(n8983), .ZN(n8987) );
  AOI22_X1 U11378 ( .A1(n13078), .A2(n8999), .B1(n9013), .B2(n12833), .ZN(
        n8985) );
  INV_X1 U11379 ( .A(n8986), .ZN(n8989) );
  NAND2_X1 U11380 ( .A1(n13194), .A2(n8999), .ZN(n8991) );
  NAND2_X1 U11381 ( .A1(n12832), .A2(n9013), .ZN(n8990) );
  NAND2_X1 U11382 ( .A1(n8991), .A2(n8990), .ZN(n8995) );
  NAND2_X1 U11383 ( .A1(n13194), .A2(n9013), .ZN(n8992) );
  OAI21_X1 U11384 ( .B1(n9013), .B2(n8993), .A(n8992), .ZN(n8994) );
  NAND2_X1 U11385 ( .A1(n13053), .A2(n9013), .ZN(n8997) );
  NAND2_X1 U11386 ( .A1(n12831), .A2(n6561), .ZN(n8996) );
  AOI22_X1 U11387 ( .A1(n13053), .A2(n6561), .B1(n9013), .B2(n12831), .ZN(
        n8998) );
  NAND2_X1 U11388 ( .A1(n13179), .A2(n6561), .ZN(n9001) );
  NAND2_X1 U11389 ( .A1(n12830), .A2(n9013), .ZN(n9000) );
  NAND2_X1 U11390 ( .A1(n13179), .A2(n9013), .ZN(n9003) );
  NAND2_X1 U11391 ( .A1(n12830), .A2(n6561), .ZN(n9002) );
  NAND2_X1 U11392 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  NAND2_X1 U11393 ( .A1(n13025), .A2(n9013), .ZN(n9006) );
  NAND2_X1 U11394 ( .A1(n12829), .A2(n8999), .ZN(n9005) );
  NAND2_X1 U11395 ( .A1(n9006), .A2(n9005), .ZN(n9009) );
  AOI22_X1 U11396 ( .A1(n13025), .A2(n8999), .B1(n9013), .B2(n12829), .ZN(
        n9007) );
  AOI21_X1 U11397 ( .B1(n9010), .B2(n9009), .A(n9007), .ZN(n9008) );
  NAND2_X1 U11398 ( .A1(n13168), .A2(n6561), .ZN(n9012) );
  NAND2_X1 U11399 ( .A1(n12828), .A2(n9013), .ZN(n9011) );
  NAND2_X1 U11400 ( .A1(n9012), .A2(n9011), .ZN(n9015) );
  AOI22_X1 U11401 ( .A1(n13168), .A2(n9013), .B1(n6561), .B2(n12828), .ZN(
        n9014) );
  NAND2_X1 U11402 ( .A1(n9018), .A2(n11626), .ZN(n9019) );
  MUX2_X1 U11403 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9020), .Z(n9021) );
  NAND2_X1 U11404 ( .A1(n9021), .A2(SI_30_), .ZN(n9022) );
  OAI21_X1 U11405 ( .B1(n9021), .B2(SI_30_), .A(n9022), .ZN(n9068) );
  MUX2_X1 U11406 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9020), .Z(n9023) );
  XNOR2_X1 U11407 ( .A(n9023), .B(SI_31_), .ZN(n9024) );
  NAND2_X1 U11408 ( .A1(n13445), .A2(n9026), .ZN(n9028) );
  INV_X1 U11409 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13252) );
  OR2_X1 U11410 ( .A1(n6567), .A2(n13252), .ZN(n9027) );
  NAND2_X1 U11411 ( .A1(n9028), .A2(n9027), .ZN(n9066) );
  INV_X1 U11412 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11413 ( .A1(n9029), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11414 ( .A1(n9030), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9031) );
  OAI211_X1 U11415 ( .C1(n8101), .C2(n9033), .A(n9032), .B(n9031), .ZN(n12960)
         );
  NAND2_X1 U11416 ( .A1(n9066), .A2(n12960), .ZN(n9034) );
  AND2_X1 U11417 ( .A1(n12823), .A2(n8999), .ZN(n9035) );
  AOI21_X1 U11418 ( .B1(n13139), .B2(n9013), .A(n9035), .ZN(n9081) );
  NAND2_X1 U11419 ( .A1(n13139), .A2(n6561), .ZN(n9037) );
  NAND2_X1 U11420 ( .A1(n12823), .A2(n9013), .ZN(n9036) );
  NAND2_X1 U11421 ( .A1(n9037), .A2(n9036), .ZN(n9080) );
  NAND2_X1 U11422 ( .A1(n9081), .A2(n9080), .ZN(n9086) );
  AND2_X1 U11423 ( .A1(n12824), .A2(n6561), .ZN(n9038) );
  AOI21_X1 U11424 ( .B1(n13144), .B2(n9013), .A(n9038), .ZN(n9084) );
  NAND2_X1 U11425 ( .A1(n13144), .A2(n8999), .ZN(n9040) );
  NAND2_X1 U11426 ( .A1(n12824), .A2(n9013), .ZN(n9039) );
  NAND2_X1 U11427 ( .A1(n9040), .A2(n9039), .ZN(n9083) );
  NAND2_X1 U11428 ( .A1(n9084), .A2(n9083), .ZN(n9041) );
  AND2_X1 U11429 ( .A1(n9086), .A2(n9041), .ZN(n9042) );
  NAND2_X1 U11430 ( .A1(n9099), .A2(n9042), .ZN(n9091) );
  AND2_X1 U11431 ( .A1(n12825), .A2(n8999), .ZN(n9043) );
  AOI21_X1 U11432 ( .B1(n13149), .B2(n9013), .A(n9043), .ZN(n9063) );
  NAND2_X1 U11433 ( .A1(n13149), .A2(n6561), .ZN(n9045) );
  NAND2_X1 U11434 ( .A1(n12825), .A2(n9013), .ZN(n9044) );
  NAND2_X1 U11435 ( .A1(n9045), .A2(n9044), .ZN(n9062) );
  AND2_X1 U11436 ( .A1(n9063), .A2(n9062), .ZN(n9046) );
  AND2_X1 U11437 ( .A1(n12826), .A2(n8999), .ZN(n9047) );
  AOI21_X1 U11438 ( .B1(n12991), .B2(n9013), .A(n9047), .ZN(n9059) );
  NAND2_X1 U11439 ( .A1(n12991), .A2(n8999), .ZN(n9049) );
  NAND2_X1 U11440 ( .A1(n12826), .A2(n9013), .ZN(n9048) );
  NAND2_X1 U11441 ( .A1(n9049), .A2(n9048), .ZN(n9058) );
  AND2_X1 U11442 ( .A1(n9059), .A2(n9058), .ZN(n9050) );
  AND2_X1 U11443 ( .A1(n12827), .A2(n8999), .ZN(n9051) );
  AOI21_X1 U11444 ( .B1(n13002), .B2(n9013), .A(n9051), .ZN(n9057) );
  NAND2_X1 U11445 ( .A1(n13002), .A2(n6561), .ZN(n9053) );
  NAND2_X1 U11446 ( .A1(n12827), .A2(n9013), .ZN(n9052) );
  NAND2_X1 U11447 ( .A1(n9053), .A2(n9052), .ZN(n9056) );
  NAND2_X1 U11448 ( .A1(n9057), .A2(n9056), .ZN(n9054) );
  OR3_X1 U11449 ( .A1(n9060), .A2(n9059), .A3(n9058), .ZN(n9061) );
  INV_X1 U11450 ( .A(n9062), .ZN(n9065) );
  INV_X1 U11451 ( .A(n9063), .ZN(n9064) );
  NAND2_X1 U11452 ( .A1(n9065), .A2(n9064), .ZN(n9090) );
  NAND2_X1 U11453 ( .A1(n12960), .A2(n9013), .ZN(n9067) );
  OAI211_X1 U11454 ( .C1(n13134), .C2(n9013), .A(n9067), .B(n9096), .ZN(n9082)
         );
  NAND2_X1 U11455 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  INV_X1 U11456 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13256) );
  OR2_X1 U11457 ( .A1(n6567), .A2(n13256), .ZN(n9073) );
  OAI211_X1 U11458 ( .C1(n14749), .C2(n11288), .A(n9412), .B(n9130), .ZN(n9074) );
  INV_X1 U11459 ( .A(n9074), .ZN(n9075) );
  NAND2_X1 U11460 ( .A1(n12960), .A2(n8999), .ZN(n9095) );
  AOI21_X1 U11461 ( .B1(n9075), .B2(n9095), .A(n9077), .ZN(n9076) );
  AOI21_X1 U11462 ( .B1(n12956), .B2(n9013), .A(n9076), .ZN(n9094) );
  NAND2_X1 U11463 ( .A1(n12956), .A2(n6561), .ZN(n9079) );
  INV_X1 U11464 ( .A(n9077), .ZN(n12822) );
  NAND2_X1 U11465 ( .A1(n12822), .A2(n9013), .ZN(n9078) );
  NAND2_X1 U11466 ( .A1(n9079), .A2(n9078), .ZN(n9093) );
  INV_X1 U11467 ( .A(n9083), .ZN(n9087) );
  INV_X1 U11468 ( .A(n9084), .ZN(n9085) );
  NAND4_X1 U11469 ( .A1(n9099), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n9088)
         );
  OAI211_X1 U11470 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9088), .ZN(n9092)
         );
  NAND2_X1 U11471 ( .A1(n9093), .A2(n9094), .ZN(n9098) );
  OAI211_X1 U11472 ( .C1(n13134), .C2(n6561), .A(n9096), .B(n9095), .ZN(n9097)
         );
  INV_X1 U11473 ( .A(n9099), .ZN(n9123) );
  XNOR2_X1 U11474 ( .A(n12956), .B(n12822), .ZN(n9120) );
  NAND2_X1 U11475 ( .A1(n9101), .A2(n9100), .ZN(n12985) );
  NAND2_X1 U11476 ( .A1(n9103), .A2(n9102), .ZN(n13020) );
  XNOR2_X1 U11477 ( .A(n14410), .B(n14379), .ZN(n11216) );
  XNOR2_X1 U11478 ( .A(n10979), .B(n9104), .ZN(n10975) );
  OR2_X1 U11479 ( .A1(n8862), .A2(n9676), .ZN(n9105) );
  NAND2_X1 U11480 ( .A1(n10066), .A2(n9105), .ZN(n14756) );
  NAND2_X1 U11481 ( .A1(n14756), .A2(n14749), .ZN(n9106) );
  NOR2_X1 U11482 ( .A1(n9106), .A2(n9751), .ZN(n9108) );
  NOR2_X1 U11483 ( .A1(n10070), .A2(n8181), .ZN(n9107) );
  XNOR2_X1 U11484 ( .A(n10060), .B(n12847), .ZN(n10056) );
  NAND4_X1 U11485 ( .A1(n9108), .A2(n9107), .A3(n10056), .A4(n9943), .ZN(n9109) );
  NOR2_X1 U11486 ( .A1(n9109), .A2(n10026), .ZN(n9110) );
  NAND4_X1 U11487 ( .A1(n10813), .A2(n9110), .A3(n10675), .A4(n10546), .ZN(
        n9111) );
  OR4_X1 U11488 ( .A1(n11154), .A2(n11016), .A3(n10975), .A4(n9111), .ZN(n9112) );
  OR4_X1 U11489 ( .A1(n13102), .A2(n13119), .A3(n11216), .A4(n9112), .ZN(n9113) );
  XNOR2_X1 U11490 ( .A(n14396), .B(n11359), .ZN(n14395) );
  OR4_X1 U11491 ( .A1(n13083), .A2(n9113), .A3(n11364), .A4(n14395), .ZN(n9114) );
  NOR2_X1 U11492 ( .A1(n13071), .A2(n9114), .ZN(n9115) );
  NAND4_X1 U11493 ( .A1(n13020), .A2(n9115), .A3(n13043), .A4(n13060), .ZN(
        n9116) );
  NOR2_X1 U11494 ( .A1(n12985), .A2(n9117), .ZN(n9118) );
  NAND4_X1 U11495 ( .A1(n9120), .A2(n9119), .A3(n9118), .A4(n12976), .ZN(n9121) );
  OAI21_X1 U11496 ( .B1(n9125), .B2(n9124), .A(n11220), .ZN(n9129) );
  INV_X1 U11497 ( .A(n9125), .ZN(n9126) );
  NOR2_X1 U11498 ( .A1(n9126), .A2(n14748), .ZN(n9128) );
  MUX2_X1 U11499 ( .A(n11288), .B(n11220), .S(n14749), .Z(n9127) );
  OAI22_X1 U11500 ( .A1(n9129), .A2(n9128), .B1(n9127), .B2(n14748), .ZN(n9134) );
  NAND2_X1 U11501 ( .A1(n14748), .A2(n9130), .ZN(n9131) );
  OAI211_X1 U11502 ( .C1(n9409), .C2(n9136), .A(n9131), .B(n9412), .ZN(n9132)
         );
  AOI22_X1 U11503 ( .A1(n9135), .A2(n9134), .B1(n9133), .B2(n9132), .ZN(n9140)
         );
  OR2_X1 U11504 ( .A1(n9419), .A2(P2_U3088), .ZN(n11371) );
  NOR4_X1 U11505 ( .A1(n14764), .A2(n14378), .A3(n8140), .A4(n9412), .ZN(n9138) );
  OAI21_X1 U11506 ( .B1(n11371), .B2(n9136), .A(P2_B_REG_SCAN_IN), .ZN(n9137)
         );
  OR2_X1 U11507 ( .A1(n9138), .A2(n9137), .ZN(n9139) );
  OAI21_X1 U11508 ( .B1(n9140), .B2(n11371), .A(n9139), .ZN(P2_U3328) );
  AND2_X1 U11509 ( .A1(n9422), .A2(n9419), .ZN(n9175) );
  NAND2_X1 U11510 ( .A1(n9434), .A2(n9152), .ZN(n9220) );
  NAND2_X1 U11511 ( .A1(n9219), .A2(n15162), .ZN(n9167) );
  INV_X1 U11512 ( .A(n9167), .ZN(n9154) );
  INV_X1 U11513 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U11514 ( .A1(n9154), .A2(n9153), .ZN(n9162) );
  NOR2_X1 U11515 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n9159) );
  NOR2_X1 U11516 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9158) );
  NOR2_X1 U11517 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n9157) );
  NAND2_X1 U11518 ( .A1(n9223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9161) );
  OAI21_X2 U11519 ( .B1(n9162), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9164) );
  INV_X1 U11520 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9163) );
  INV_X1 U11521 ( .A(n9320), .ZN(n9165) );
  NAND2_X1 U11522 ( .A1(n9167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9168) );
  INV_X1 U11523 ( .A(n9325), .ZN(n9367) );
  OR2_X2 U11524 ( .A1(n10364), .A2(n9367), .ZN(n13695) );
  INV_X1 U11525 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n12858) );
  INV_X1 U11526 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9360) );
  AOI211_X1 U11527 ( .C1(n12857), .C2(n12858), .A(n12860), .B(n9360), .ZN(
        n9170) );
  INV_X1 U11528 ( .A(n12857), .ZN(n9182) );
  NAND2_X1 U11529 ( .A1(n9182), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11530 ( .A1(n9170), .A2(n9171), .ZN(n12862) );
  NAND2_X1 U11531 ( .A1(n12862), .A2(n9171), .ZN(n9299) );
  XNOR2_X1 U11532 ( .A(n9254), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9300) );
  INV_X1 U11533 ( .A(n9254), .ZN(n9307) );
  AOI22_X1 U11534 ( .A1(n9299), .A2(n9300), .B1(n9307), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n9178) );
  MUX2_X1 U11535 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9756), .S(n9333), .Z(n9177)
         );
  NOR2_X1 U11536 ( .A1(n9178), .A2(n9177), .ZN(n9344) );
  NAND2_X1 U11537 ( .A1(n9413), .A2(n9419), .ZN(n9172) );
  AND2_X1 U11538 ( .A1(n9173), .A2(n9172), .ZN(n9174) );
  OR2_X1 U11539 ( .A1(n9175), .A2(n9174), .ZN(n9188) );
  OR2_X1 U11540 ( .A1(n8131), .A2(P2_U3088), .ZN(n13262) );
  INV_X1 U11541 ( .A(n13262), .ZN(n9176) );
  NAND2_X1 U11542 ( .A1(n9188), .A2(n9176), .ZN(n9179) );
  AOI211_X1 U11544 ( .C1(n9178), .C2(n9177), .A(n9344), .B(n15310), .ZN(n9193)
         );
  INV_X1 U11545 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11546 ( .A1(n9180), .A2(n8140), .ZN(n11644) );
  MUX2_X1 U11547 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n7680), .S(n12857), .Z(
        n12854) );
  NOR3_X1 U11548 ( .A1(n12854), .A2(n12860), .A3(n9181), .ZN(n12853) );
  AOI21_X1 U11549 ( .B1(n9182), .B2(P2_REG1_REG_1__SCAN_IN), .A(n12853), .ZN(
        n9304) );
  MUX2_X1 U11550 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7699), .S(n9254), .Z(n9303)
         );
  OR2_X1 U11551 ( .A1(n9304), .A2(n9303), .ZN(n9301) );
  NAND2_X1 U11552 ( .A1(n9307), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9184) );
  MUX2_X1 U11553 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7716), .S(n9333), .Z(n9183)
         );
  AOI21_X1 U11554 ( .B1(n9301), .B2(n9184), .A(n9183), .ZN(n9334) );
  AND3_X1 U11555 ( .A1(n9301), .A2(n9184), .A3(n9183), .ZN(n9185) );
  NOR3_X1 U11556 ( .A1(n11644), .A2(n9334), .A3(n9185), .ZN(n9192) );
  NOR2_X2 U11557 ( .A1(n9188), .A2(P2_U3088), .ZN(n14718) );
  INV_X1 U11558 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9186) );
  NOR2_X1 U11559 ( .A1(n14706), .A2(n9186), .ZN(n9191) );
  AND2_X1 U11560 ( .A1(n8131), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11561 ( .A1(n9188), .A2(n9187), .ZN(n12925) );
  INV_X1 U11562 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9189) );
  OAI22_X1 U11563 ( .A1(n12925), .A2(n9333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9189), .ZN(n9190) );
  OR4_X1 U11564 ( .A1(n9193), .A2(n9192), .A3(n9191), .A4(n9190), .ZN(P2_U3217) );
  NOR2_X1 U11565 ( .A1(n9194), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9197) );
  NOR2_X1 U11566 ( .A1(n9197), .A2(n9479), .ZN(n9195) );
  MUX2_X1 U11567 ( .A(n9479), .B(n9195), .S(P1_IR_REG_5__SCAN_IN), .Z(n9198)
         );
  AND2_X1 U11568 ( .A1(n9197), .A2(n9196), .ZN(n9215) );
  OR2_X1 U11569 ( .A1(n9198), .A2(n9215), .ZN(n13756) );
  INV_X1 U11570 ( .A(n13756), .ZN(n13750) );
  NAND2_X1 U11571 ( .A1(n9194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9199) );
  XNOR2_X1 U11572 ( .A(n9199), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13732) );
  INV_X1 U11573 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9205) );
  NOR2_X1 U11574 ( .A1(n9200), .A2(n9479), .ZN(n9201) );
  MUX2_X1 U11575 ( .A(n9479), .B(n9201), .S(P1_IR_REG_2__SCAN_IN), .Z(n9204)
         );
  INV_X1 U11576 ( .A(n9202), .ZN(n9203) );
  MUX2_X1 U11577 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9205), .S(n13712), .Z(n9210) );
  NAND2_X1 U11578 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9206) );
  XNOR2_X1 U11579 ( .A(n9206), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9544) );
  INV_X1 U11580 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9207) );
  XNOR2_X1 U11581 ( .A(n9544), .B(n9207), .ZN(n9533) );
  AND2_X1 U11582 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9532) );
  NAND2_X1 U11583 ( .A1(n9533), .A2(n9532), .ZN(n9209) );
  NAND2_X1 U11584 ( .A1(n9544), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11585 ( .A1(n9209), .A2(n9208), .ZN(n13705) );
  NAND2_X1 U11586 ( .A1(n9210), .A2(n13705), .ZN(n13723) );
  NAND2_X1 U11587 ( .A1(n13712), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U11588 ( .A1(n13723), .A2(n13722), .ZN(n9214) );
  INV_X1 U11589 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11590 ( .A1(n9202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9211) );
  XNOR2_X1 U11591 ( .A(n9211), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13720) );
  MUX2_X1 U11592 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9212), .S(n13720), .Z(n9213) );
  NAND2_X1 U11593 ( .A1(n9214), .A2(n9213), .ZN(n13736) );
  NAND2_X1 U11594 ( .A1(n13720), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13735) );
  INV_X1 U11595 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15086) );
  MUX2_X1 U11596 ( .A(n15086), .B(P1_REG1_REG_4__SCAN_IN), .S(n13732), .Z(
        n13734) );
  AOI21_X1 U11597 ( .B1(n13732), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13733), .ZN(
        n13752) );
  INV_X1 U11598 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14667) );
  MUX2_X1 U11599 ( .A(n14667), .B(P1_REG1_REG_5__SCAN_IN), .S(n13756), .Z(
        n13753) );
  NAND2_X1 U11600 ( .A1(n13752), .A2(n13753), .ZN(n13751) );
  OAI21_X1 U11601 ( .B1(n13750), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13751), .ZN(
        n9229) );
  INV_X1 U11602 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14669) );
  NOR2_X1 U11603 ( .A1(n9215), .A2(n9479), .ZN(n9216) );
  MUX2_X1 U11604 ( .A(n9479), .B(n9216), .S(P1_IR_REG_6__SCAN_IN), .Z(n9218)
         );
  INV_X1 U11605 ( .A(n9217), .ZN(n10092) );
  MUX2_X1 U11606 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14669), .S(n10504), .Z(
        n9228) );
  OR2_X1 U11607 ( .A1(n10361), .A2(P1_U3086), .ZN(n13666) );
  INV_X1 U11608 ( .A(n13666), .ZN(n11368) );
  OR2_X1 U11609 ( .A1(n10231), .A2(n11368), .ZN(n9232) );
  NAND2_X1 U11610 ( .A1(n9220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9222) );
  INV_X1 U11611 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11612 ( .A1(n6847), .A2(n9461), .ZN(n13638) );
  INV_X1 U11613 ( .A(n13638), .ZN(n9227) );
  MUX2_X1 U11614 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9225), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9226) );
  AOI21_X1 U11615 ( .B1(n9227), .B2(n10361), .A(n6562), .ZN(n9230) );
  NAND2_X1 U11616 ( .A1(n9232), .A2(n9230), .ZN(n14528) );
  INV_X1 U11617 ( .A(n14142), .ZN(n14517) );
  NOR2_X2 U11618 ( .A1(n14528), .A2(n14517), .ZN(n13819) );
  AOI211_X1 U11619 ( .C1(n9229), .C2(n9228), .A(n13773), .B(n14536), .ZN(n9250) );
  INV_X1 U11620 ( .A(n9230), .ZN(n9231) );
  INV_X1 U11621 ( .A(n14525), .ZN(n14541) );
  OAI22_X1 U11622 ( .A1(n14541), .A2(n14164), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10367), .ZN(n9249) );
  INV_X1 U11623 ( .A(n14528), .ZN(n9235) );
  NOR2_X1 U11624 ( .A1(n9233), .A2(n14142), .ZN(n9234) );
  NAND2_X1 U11625 ( .A1(n9235), .A2(n9234), .ZN(n14534) );
  INV_X1 U11626 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9236) );
  MUX2_X1 U11627 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9236), .S(n13712), .Z(
        n13704) );
  INV_X1 U11628 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9237) );
  MUX2_X1 U11629 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9237), .S(n9544), .Z(n9537)
         );
  AND2_X1 U11630 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9238) );
  NAND2_X1 U11631 ( .A1(n9537), .A2(n9238), .ZN(n9536) );
  NAND2_X1 U11632 ( .A1(n9544), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11633 ( .A1(n9536), .A2(n9239), .ZN(n13703) );
  NAND2_X1 U11634 ( .A1(n13704), .A2(n13703), .ZN(n13718) );
  NAND2_X1 U11635 ( .A1(n13712), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13717) );
  NAND2_X1 U11636 ( .A1(n13718), .A2(n13717), .ZN(n9241) );
  INV_X1 U11637 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n15054) );
  MUX2_X1 U11638 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n15054), .S(n13720), .Z(
        n9240) );
  NAND2_X1 U11639 ( .A1(n9241), .A2(n9240), .ZN(n13742) );
  NAND2_X1 U11640 ( .A1(n13720), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13741) );
  INV_X1 U11641 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9242) );
  MUX2_X1 U11642 ( .A(n9242), .B(P1_REG2_REG_4__SCAN_IN), .S(n13732), .Z(
        n13740) );
  AOI21_X1 U11643 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13739) );
  INV_X1 U11644 ( .A(n13732), .ZN(n9262) );
  NOR2_X1 U11645 ( .A1(n9262), .A2(n9242), .ZN(n13755) );
  INV_X1 U11646 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10387) );
  MUX2_X1 U11647 ( .A(n10387), .B(P1_REG2_REG_5__SCAN_IN), .S(n13756), .Z(
        n9243) );
  OAI21_X1 U11648 ( .B1(n13739), .B2(n13755), .A(n9243), .ZN(n13761) );
  NAND2_X1 U11649 ( .A1(n13750), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9245) );
  INV_X1 U11650 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n15113) );
  MUX2_X1 U11651 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n15113), .S(n10504), .Z(
        n9244) );
  AOI21_X1 U11652 ( .B1(n13761), .B2(n9245), .A(n9244), .ZN(n13780) );
  AND3_X1 U11653 ( .A1(n13761), .A2(n9245), .A3(n9244), .ZN(n9246) );
  NOR3_X1 U11654 ( .A1(n14534), .A2(n13780), .A3(n9246), .ZN(n9248) );
  INV_X1 U11655 ( .A(n9233), .ZN(n13701) );
  NOR2_X1 U11656 ( .A1(n6779), .A2(n10504), .ZN(n9247) );
  OR4_X1 U11657 ( .A1(n9250), .A2(n9249), .A3(n9248), .A4(n9247), .ZN(P1_U3249) );
  INV_X1 U11658 ( .A(n9544), .ZN(n9252) );
  AND2_X1 U11659 ( .A1(n9020), .A2(P1_U3086), .ZN(n14136) );
  INV_X2 U11660 ( .A(n14136), .ZN(n14145) );
  OAI222_X1 U11661 ( .A1(P1_U3086), .A2(n9252), .B1(n14148), .B2(n9547), .C1(
        n7263), .C2(n14145), .ZN(P1_U3354) );
  AND2_X1 U11662 ( .A1(n7631), .A2(P2_U3088), .ZN(n13260) );
  INV_X2 U11663 ( .A(n13260), .ZN(n13272) );
  OAI222_X1 U11664 ( .A1(n13272), .A2(n9733), .B1(n9254), .B2(P2_U3088), .C1(
        n9253), .C2(n13269), .ZN(P2_U3325) );
  OAI222_X1 U11665 ( .A1(n13272), .A2(n9547), .B1(n12857), .B2(P2_U3088), .C1(
        n9255), .C2(n13269), .ZN(P2_U3326) );
  OAI222_X1 U11666 ( .A1(n13272), .A2(n10239), .B1(n9333), .B2(P2_U3088), .C1(
        n9256), .C2(n13269), .ZN(P2_U3324) );
  INV_X1 U11667 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9258) );
  INV_X1 U11668 ( .A(n13712), .ZN(n9257) );
  OAI222_X1 U11669 ( .A1(n14145), .A2(n9258), .B1(n14148), .B2(n9733), .C1(
        n9257), .C2(P1_U3086), .ZN(P1_U3353) );
  INV_X1 U11670 ( .A(n13720), .ZN(n9259) );
  OAI222_X1 U11671 ( .A1(n14145), .A2(n6842), .B1(n14148), .B2(n10239), .C1(
        n9259), .C2(P1_U3086), .ZN(P1_U3352) );
  NOR2_X1 U11672 ( .A1(n9020), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12602) );
  OAI222_X1 U11673 ( .A1(n12609), .A2(n9260), .B1(n12606), .B2(n7265), .C1(
        P3_U3151), .C2(n9601), .ZN(P3_U3294) );
  INV_X1 U11674 ( .A(n10241), .ZN(n9263) );
  INV_X1 U11675 ( .A(n9379), .ZN(n9346) );
  OAI222_X1 U11676 ( .A1(n13272), .A2(n9263), .B1(n9346), .B2(P2_U3088), .C1(
        n9261), .C2(n13269), .ZN(P2_U3323) );
  OAI222_X1 U11677 ( .A1(n14145), .A2(n6965), .B1(n14148), .B2(n9263), .C1(
        n9262), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U11678 ( .A(n9805), .ZN(n9810) );
  INV_X1 U11679 ( .A(n9264), .ZN(n9265) );
  INV_X1 U11680 ( .A(SI_3_), .ZN(n15242) );
  OAI222_X1 U11681 ( .A1(n9810), .A2(P3_U3151), .B1(n12609), .B2(n9265), .C1(
        n15242), .C2(n12606), .ZN(P3_U3292) );
  INV_X1 U11682 ( .A(n9836), .ZN(n9268) );
  INV_X1 U11683 ( .A(n9266), .ZN(n9267) );
  OAI222_X1 U11684 ( .A1(n9268), .A2(P3_U3151), .B1(n12609), .B2(n9267), .C1(
        n6729), .C2(n12606), .ZN(P3_U3291) );
  INV_X1 U11685 ( .A(n9269), .ZN(n9271) );
  INV_X1 U11686 ( .A(SI_5_), .ZN(n9270) );
  OAI222_X1 U11687 ( .A1(n9837), .A2(P3_U3151), .B1(n12609), .B2(n9271), .C1(
        n9270), .C2(n12606), .ZN(P3_U3290) );
  INV_X1 U11688 ( .A(n9782), .ZN(n9788) );
  INV_X1 U11689 ( .A(n9272), .ZN(n9274) );
  INV_X1 U11690 ( .A(SI_2_), .ZN(n9273) );
  OAI222_X1 U11691 ( .A1(n9788), .A2(P3_U3151), .B1(n12609), .B2(n9274), .C1(
        n9273), .C2(n12606), .ZN(P3_U3293) );
  OAI222_X1 U11692 ( .A1(P3_U3151), .A2(n9934), .B1(n12609), .B2(n9276), .C1(
        n9275), .C2(n12606), .ZN(P3_U3289) );
  INV_X1 U11693 ( .A(n12870), .ZN(n12867) );
  OAI222_X1 U11694 ( .A1(n13272), .A2(n10356), .B1(n12867), .B2(P2_U3088), 
        .C1(n9277), .C2(n13269), .ZN(P2_U3322) );
  INV_X1 U11695 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9278) );
  OAI222_X1 U11696 ( .A1(n14145), .A2(n9278), .B1(n14148), .B2(n10356), .C1(
        n13756), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U11697 ( .A1(n12606), .A2(n9280), .B1(n12609), .B2(n9279), .C1(
        n14856), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U11698 ( .A(n9347), .ZN(n12888) );
  OAI222_X1 U11699 ( .A1(n13272), .A2(n10503), .B1(n12888), .B2(P2_U3088), 
        .C1(n9281), .C2(n13269), .ZN(P2_U3321) );
  OAI222_X1 U11700 ( .A1(n14145), .A2(n9282), .B1(n14148), .B2(n10503), .C1(
        n10504), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U11701 ( .A(n9283), .ZN(n9284) );
  OAI222_X1 U11702 ( .A1(P3_U3151), .A2(n12194), .B1(n12606), .B2(n9285), .C1(
        n12609), .C2(n9284), .ZN(P3_U3285) );
  INV_X1 U11703 ( .A(n10110), .ZN(n10118) );
  INV_X1 U11704 ( .A(SI_7_), .ZN(n15224) );
  INV_X1 U11705 ( .A(n9286), .ZN(n9287) );
  OAI222_X1 U11706 ( .A1(P3_U3151), .A2(n10118), .B1(n12606), .B2(n15224), 
        .C1(n12609), .C2(n9287), .ZN(P3_U3288) );
  INV_X1 U11707 ( .A(n9288), .ZN(n9289) );
  OAI222_X1 U11708 ( .A1(P3_U3151), .A2(n12197), .B1(n12606), .B2(n9290), .C1(
        n12609), .C2(n9289), .ZN(P3_U3284) );
  INV_X1 U11709 ( .A(SI_9_), .ZN(n9293) );
  INV_X1 U11710 ( .A(n9291), .ZN(n9292) );
  OAI222_X1 U11711 ( .A1(P3_U3151), .A2(n10487), .B1(n12606), .B2(n9293), .C1(
        n12609), .C2(n9292), .ZN(P3_U3286) );
  OAI222_X1 U11712 ( .A1(n12609), .A2(n9295), .B1(n12606), .B2(n9294), .C1(
        P3_U3151), .C2(n10315), .ZN(P3_U3287) );
  INV_X1 U11713 ( .A(n12898), .ZN(n12906) );
  INV_X1 U11714 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9296) );
  OAI222_X1 U11715 ( .A1(n13272), .A2(n10511), .B1(n12906), .B2(P2_U3088), 
        .C1(n9296), .C2(n13269), .ZN(P2_U3320) );
  NAND2_X1 U11716 ( .A1(n10092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9297) );
  XNOR2_X1 U11717 ( .A(n9297), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13775) );
  INV_X1 U11718 ( .A(n13775), .ZN(n9487) );
  OAI222_X1 U11719 ( .A1(n14145), .A2(n9298), .B1(n14148), .B2(n10511), .C1(
        n9487), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U11720 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9310) );
  XOR2_X1 U11721 ( .A(n9300), .B(n9299), .Z(n9306) );
  INV_X1 U11722 ( .A(n9301), .ZN(n9302) );
  AOI211_X1 U11723 ( .C1(n9304), .C2(n9303), .A(n9302), .B(n11644), .ZN(n9305)
         );
  AOI21_X1 U11724 ( .B1(n6547), .B2(n9306), .A(n9305), .ZN(n9309) );
  INV_X1 U11725 ( .A(n12925), .ZN(n14720) );
  AOI22_X1 U11726 ( .A1(n14720), .A2(n9307), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3088), .ZN(n9308) );
  OAI211_X1 U11727 ( .C1(n14706), .C2(n9310), .A(n9309), .B(n9308), .ZN(
        P2_U3216) );
  INV_X1 U11728 ( .A(n9570), .ZN(n9343) );
  INV_X1 U11729 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9311) );
  OAI222_X1 U11730 ( .A1(n13272), .A2(n10622), .B1(n9343), .B2(P2_U3088), .C1(
        n9311), .C2(n13269), .ZN(P2_U3319) );
  INV_X1 U11731 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9314) );
  INV_X1 U11732 ( .A(n10283), .ZN(n9312) );
  NAND2_X1 U11733 ( .A1(n9312), .A2(n9319), .ZN(n9313) );
  OAI21_X1 U11734 ( .B1(n9319), .B2(n9314), .A(n9313), .ZN(P3_U3377) );
  NAND2_X1 U11735 ( .A1(n9478), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9357) );
  XNOR2_X1 U11736 ( .A(n9357), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10623) );
  INV_X1 U11737 ( .A(n10623), .ZN(n9492) );
  OAI222_X1 U11738 ( .A1(n14145), .A2(n9315), .B1(n14148), .B2(n10622), .C1(
        n9492), .C2(P1_U3086), .ZN(P1_U3347) );
  AND2_X1 U11739 ( .A1(n9329), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11740 ( .A1(n9329), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11741 ( .A1(n9329), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11742 ( .A1(n9329), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11743 ( .A1(n9329), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11744 ( .A1(n9329), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11745 ( .A1(n9329), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11746 ( .A1(n9329), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11747 ( .A1(n9329), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11748 ( .A1(n9329), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11749 ( .A1(n9329), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11750 ( .A1(n9329), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11751 ( .A1(n9329), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11752 ( .A1(n9329), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11753 ( .A1(n9329), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11754 ( .A1(n9329), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11755 ( .A1(n9329), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11756 ( .A1(n9329), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11757 ( .A1(n9329), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11758 ( .A1(n9329), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11759 ( .A1(n9329), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11760 ( .A1(n9329), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11761 ( .A1(n9329), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11762 ( .A1(n9329), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11763 ( .A1(n9329), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11764 ( .A1(n9329), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  INV_X1 U11765 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9318) );
  INV_X1 U11766 ( .A(n10040), .ZN(n9316) );
  NAND2_X1 U11767 ( .A1(n9316), .A2(n9319), .ZN(n9317) );
  OAI21_X1 U11768 ( .B1(n9319), .B2(n9318), .A(n9317), .ZN(P3_U3376) );
  NAND3_X1 U11769 ( .A1(n9320), .A2(P1_B_REG_SCAN_IN), .A3(n11952), .ZN(n9324)
         );
  INV_X1 U11770 ( .A(P1_B_REG_SCAN_IN), .ZN(n9321) );
  AOI21_X1 U11771 ( .B1(n9322), .B2(n9321), .A(n14149), .ZN(n9323) );
  NAND2_X1 U11772 ( .A1(n9324), .A2(n9323), .ZN(n9648) );
  NAND2_X1 U11773 ( .A1(n10231), .A2(n9648), .ZN(n14586) );
  INV_X1 U11774 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U11775 ( .A1(n9320), .A2(n14149), .ZN(n9649) );
  INV_X1 U11776 ( .A(n9649), .ZN(n9326) );
  AOI22_X1 U11777 ( .A1(n14586), .A2(n9645), .B1(n9326), .B2(n9325), .ZN(
        P1_U3446) );
  OAI222_X1 U11778 ( .A1(P3_U3151), .A2(n12201), .B1(n12606), .B2(n9328), .C1(
        n12609), .C2(n9327), .ZN(P3_U3282) );
  INV_X1 U11779 ( .A(n9329), .ZN(n9330) );
  INV_X1 U11780 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15009) );
  NOR2_X1 U11781 ( .A1(n9330), .A2(n15009), .ZN(P3_U3255) );
  INV_X1 U11782 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n15135) );
  NOR2_X1 U11783 ( .A1(n9330), .A2(n15135), .ZN(P3_U3248) );
  INV_X1 U11784 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n15251) );
  NOR2_X1 U11785 ( .A1(n9330), .A2(n15251), .ZN(P3_U3240) );
  INV_X1 U11786 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15153) );
  NOR2_X1 U11787 ( .A1(n9330), .A2(n15153), .ZN(P3_U3250) );
  INV_X1 U11788 ( .A(n14702), .ZN(n9332) );
  OAI222_X1 U11789 ( .A1(n13272), .A2(n10690), .B1(n9332), .B2(P2_U3088), .C1(
        n9331), .C2(n13269), .ZN(P2_U3318) );
  INV_X1 U11790 ( .A(n9333), .ZN(n9345) );
  AOI21_X1 U11791 ( .B1(n9345), .B2(P2_REG1_REG_3__SCAN_IN), .A(n9334), .ZN(
        n9374) );
  MUX2_X1 U11792 ( .A(n9335), .B(P2_REG1_REG_4__SCAN_IN), .S(n9379), .Z(n9373)
         );
  NOR2_X1 U11793 ( .A1(n9374), .A2(n9373), .ZN(n12874) );
  NOR2_X1 U11794 ( .A1(n9346), .A2(n9335), .ZN(n12869) );
  MUX2_X1 U11795 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9336), .S(n12870), .Z(n9337) );
  OAI21_X1 U11796 ( .B1(n12874), .B2(n12869), .A(n9337), .ZN(n12884) );
  NAND2_X1 U11797 ( .A1(n12870), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n12883) );
  INV_X1 U11798 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U11799 ( .A(n10226), .B(P2_REG1_REG_6__SCAN_IN), .S(n9347), .Z(
        n12882) );
  AOI21_X1 U11800 ( .B1(n12884), .B2(n12883), .A(n12882), .ZN(n12904) );
  NOR2_X1 U11801 ( .A1(n12888), .A2(n10226), .ZN(n12899) );
  INV_X1 U11802 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9338) );
  MUX2_X1 U11803 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9338), .S(n12898), .Z(n9339) );
  OAI21_X1 U11804 ( .B1(n12904), .B2(n12899), .A(n9339), .ZN(n12902) );
  NAND2_X1 U11805 ( .A1(n12898), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11806 ( .A(n7815), .B(P2_REG1_REG_8__SCAN_IN), .S(n9570), .Z(n9340)
         );
  AOI21_X1 U11807 ( .B1(n12902), .B2(n9341), .A(n9340), .ZN(n9566) );
  NAND3_X1 U11808 ( .A1(n12902), .A2(n9341), .A3(n9340), .ZN(n9342) );
  NAND2_X1 U11809 ( .A1(n9342), .A2(n14725), .ZN(n9355) );
  NAND2_X1 U11810 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10451) );
  OAI21_X1 U11811 ( .B1(n12925), .B2(n9343), .A(n10451), .ZN(n9353) );
  AOI21_X1 U11812 ( .B1(n9345), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9344), .ZN(
        n9371) );
  MUX2_X1 U11813 ( .A(n9951), .B(P2_REG2_REG_4__SCAN_IN), .S(n9379), .Z(n9370)
         );
  NOR2_X1 U11814 ( .A1(n9371), .A2(n9370), .ZN(n12877) );
  NOR2_X1 U11815 ( .A1(n9346), .A2(n9951), .ZN(n12876) );
  MUX2_X1 U11816 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10061), .S(n12870), .Z(
        n12875) );
  OAI21_X1 U11817 ( .B1(n12877), .B2(n12876), .A(n12875), .ZN(n12892) );
  NAND2_X1 U11818 ( .A1(n12870), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n12891) );
  MUX2_X1 U11819 ( .A(n7777), .B(P2_REG2_REG_6__SCAN_IN), .S(n9347), .Z(n12890) );
  AOI21_X1 U11820 ( .B1(n12892), .B2(n12891), .A(n12890), .ZN(n12910) );
  NOR2_X1 U11821 ( .A1(n12888), .A2(n7777), .ZN(n12909) );
  MUX2_X1 U11822 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9348), .S(n12898), .Z(
        n12908) );
  OAI21_X1 U11823 ( .B1(n12910), .B2(n12909), .A(n12908), .ZN(n12912) );
  NAND2_X1 U11824 ( .A1(n12898), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9350) );
  MUX2_X1 U11825 ( .A(n10678), .B(P2_REG2_REG_8__SCAN_IN), .S(n9570), .Z(n9349) );
  AOI21_X1 U11826 ( .B1(n12912), .B2(n9350), .A(n9349), .ZN(n9569) );
  AND3_X1 U11827 ( .A1(n12912), .A2(n9350), .A3(n9349), .ZN(n9351) );
  NOR3_X1 U11828 ( .A1(n9569), .A2(n9351), .A3(n15310), .ZN(n9352) );
  AOI211_X1 U11829 ( .C1(n14718), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9353), .B(
        n9352), .ZN(n9354) );
  OAI21_X1 U11830 ( .B1(n9566), .B2(n9355), .A(n9354), .ZN(P2_U3222) );
  INV_X1 U11831 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11832 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  NAND2_X1 U11833 ( .A1(n9358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9385) );
  XNOR2_X1 U11834 ( .A(n9385), .B(P1_IR_REG_9__SCAN_IN), .ZN(n13792) );
  INV_X1 U11835 ( .A(n13792), .ZN(n9359) );
  OAI222_X1 U11836 ( .A1(n14145), .A2(n15110), .B1(n14148), .B2(n10690), .C1(
        n9359), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U11837 ( .A1(n6547), .A2(n9360), .ZN(n9361) );
  OAI211_X1 U11838 ( .C1(n11644), .C2(P2_REG1_REG_0__SCAN_IN), .A(n9361), .B(
        n12925), .ZN(n9363) );
  OAI22_X1 U11839 ( .A1(n15310), .A2(n9360), .B1(n9181), .B2(n11644), .ZN(
        n9362) );
  MUX2_X1 U11840 ( .A(n9363), .B(n9362), .S(n12860), .Z(n9366) );
  INV_X1 U11841 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9364) );
  INV_X1 U11842 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14752) );
  OAI22_X1 U11843 ( .A1(n14706), .A2(n9364), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14752), .ZN(n9365) );
  OR2_X1 U11844 ( .A1(n9366), .A2(n9365), .ZN(P2_U3214) );
  INV_X1 U11845 ( .A(n14586), .ZN(n14585) );
  NAND2_X1 U11846 ( .A1(n11952), .A2(n14149), .ZN(n9454) );
  OAI22_X1 U11847 ( .A1(n14585), .A2(P1_D_REG_0__SCAN_IN), .B1(n9367), .B2(
        n9454), .ZN(n9368) );
  INV_X1 U11848 ( .A(n9368), .ZN(P1_U3445) );
  INV_X1 U11849 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U11850 ( .A1(n10720), .A2(P3_U3897), .ZN(n9369) );
  OAI21_X1 U11851 ( .B1(P3_U3897), .B2(n15174), .A(n9369), .ZN(P3_U3496) );
  INV_X1 U11852 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9381) );
  AOI211_X1 U11853 ( .C1(n9371), .C2(n9370), .A(n12877), .B(n15310), .ZN(n9372) );
  INV_X1 U11854 ( .A(n9372), .ZN(n9377) );
  AOI211_X1 U11855 ( .C1(n9374), .C2(n9373), .A(n12874), .B(n11644), .ZN(n9375) );
  INV_X1 U11856 ( .A(n9375), .ZN(n9376) );
  NAND2_X1 U11857 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  AND2_X1 U11858 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9695) );
  AOI211_X1 U11859 ( .C1(n14720), .C2(n9379), .A(n9378), .B(n9695), .ZN(n9380)
         );
  OAI21_X1 U11860 ( .B1(n14706), .B2(n9381), .A(n9380), .ZN(P2_U3218) );
  INV_X1 U11861 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n15249) );
  NAND2_X1 U11862 ( .A1(n12037), .A2(P3_U3897), .ZN(n9382) );
  OAI21_X1 U11863 ( .B1(P3_U3897), .B2(n15249), .A(n9382), .ZN(P3_U3498) );
  INV_X1 U11864 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U11865 ( .A1(n12437), .A2(P3_U3897), .ZN(n9383) );
  OAI21_X1 U11866 ( .B1(P3_U3897), .B2(n15019), .A(n9383), .ZN(P3_U3503) );
  NOR2_X1 U11867 ( .A1(n14525), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11868 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n15208) );
  INV_X1 U11869 ( .A(n10907), .ZN(n9388) );
  OAI222_X1 U11870 ( .A1(n13269), .A2(n15208), .B1(n13272), .B2(n9388), .C1(
        P2_U3088), .C2(n9888), .ZN(P2_U3317) );
  INV_X1 U11871 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11872 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U11873 ( .A1(n9386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U11874 ( .A(n9387), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10908) );
  INV_X1 U11875 ( .A(n10908), .ZN(n9496) );
  OAI222_X1 U11876 ( .A1(n14145), .A2(n9389), .B1(n14148), .B2(n9388), .C1(
        P1_U3086), .C2(n9496), .ZN(P1_U3345) );
  INV_X1 U11877 ( .A(n14905), .ZN(n9393) );
  INV_X1 U11878 ( .A(n9390), .ZN(n9391) );
  OAI222_X1 U11879 ( .A1(P3_U3151), .A2(n9393), .B1(n12606), .B2(n9392), .C1(
        n12609), .C2(n9391), .ZN(P3_U3281) );
  INV_X1 U11880 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15209) );
  NAND2_X1 U11881 ( .A1(n12423), .A2(P3_U3897), .ZN(n9394) );
  OAI21_X1 U11882 ( .B1(P3_U3897), .B2(n15209), .A(n9394), .ZN(P3_U3506) );
  INV_X1 U11883 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9396) );
  INV_X1 U11884 ( .A(n11808), .ZN(n9400) );
  AND2_X2 U11885 ( .A1(n9400), .A2(n9399), .ZN(n11731) );
  NAND2_X1 U11886 ( .A1(n11731), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9402) );
  NAND2_X2 U11887 ( .A1(n11808), .A2(n14139), .ZN(n11750) );
  NAND2_X1 U11888 ( .A1(n10244), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11889 ( .A1(P1_U4016), .A2(n6824), .ZN(n9403) );
  OAI21_X1 U11890 ( .B1(P1_U4016), .B2(n8252), .A(n9403), .ZN(P1_U3560) );
  NAND2_X1 U11891 ( .A1(n8862), .A2(n12800), .ZN(n9405) );
  NAND2_X1 U11892 ( .A1(n8876), .A2(n12801), .ZN(n9404) );
  AND2_X1 U11893 ( .A1(n9405), .A2(n9404), .ZN(n10072) );
  INV_X1 U11894 ( .A(n10134), .ZN(n10143) );
  NAND2_X1 U11895 ( .A1(n9406), .A2(n10143), .ZN(n9417) );
  NOR2_X1 U11896 ( .A1(n9417), .A2(n14764), .ZN(n9407) );
  NAND2_X1 U11897 ( .A1(n9408), .A2(n9407), .ZN(n9428) );
  NAND2_X1 U11898 ( .A1(n8178), .A2(n12664), .ZN(n9520) );
  XNOR2_X1 U11899 ( .A(n9520), .B(n9518), .ZN(n9517) );
  NAND2_X1 U11900 ( .A1(n8862), .A2(n12664), .ZN(n9410) );
  NAND2_X1 U11901 ( .A1(n9410), .A2(n9676), .ZN(n9682) );
  NAND2_X1 U11902 ( .A1(n14747), .A2(n12663), .ZN(n9411) );
  NAND2_X1 U11903 ( .A1(n9682), .A2(n9411), .ZN(n9516) );
  XNOR2_X1 U11904 ( .A(n9517), .B(n9516), .ZN(n9415) );
  OR2_X1 U11905 ( .A1(n14795), .A2(n9413), .ZN(n9414) );
  NAND2_X1 U11906 ( .A1(n9415), .A2(n14688), .ZN(n9431) );
  OR2_X1 U11907 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U11908 ( .A1(n9418), .A2(n10131), .ZN(n9425) );
  INV_X1 U11909 ( .A(n9419), .ZN(n9420) );
  OR2_X1 U11910 ( .A1(n9421), .A2(n9420), .ZN(n9423) );
  NOR2_X1 U11911 ( .A1(n9423), .A2(n9422), .ZN(n9424) );
  NAND2_X1 U11912 ( .A1(n9425), .A2(n9424), .ZN(n9698) );
  NOR2_X1 U11913 ( .A1(n9698), .A2(P2_U3088), .ZN(n9526) );
  INV_X1 U11914 ( .A(n9526), .ZN(n9679) );
  INV_X1 U11915 ( .A(n9426), .ZN(n9427) );
  OR2_X1 U11916 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  AOI22_X1 U11917 ( .A1(n9679), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8869), .B2(
        n14690), .ZN(n9430) );
  OAI211_X1 U11918 ( .C1(n10072), .C2(n12806), .A(n9431), .B(n9430), .ZN(
        P2_U3194) );
  INV_X1 U11919 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n15118) );
  NAND2_X1 U11920 ( .A1(n12385), .A2(P3_U3897), .ZN(n9432) );
  OAI21_X1 U11921 ( .B1(P3_U3897), .B2(n15118), .A(n9432), .ZN(P3_U3509) );
  OAI21_X1 U11922 ( .B1(n9648), .B2(P1_D_REG_1__SCAN_IN), .A(n9649), .ZN(n9453) );
  AND2_X1 U11923 ( .A1(n9433), .A2(n13464), .ZN(n9557) );
  NAND2_X1 U11924 ( .A1(n9439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U11925 ( .A1(n9437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U11926 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9438), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9440) );
  NAND2_X1 U11927 ( .A1(n14577), .A2(n13952), .ZN(n10229) );
  NOR4_X1 U11928 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9444) );
  NOR4_X1 U11929 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9443) );
  NOR4_X1 U11930 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9442) );
  NOR4_X1 U11931 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9441) );
  AND4_X1 U11932 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), .ZN(n9450)
         );
  NOR2_X1 U11933 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .ZN(
        n9448) );
  NOR4_X1 U11934 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9447) );
  NOR4_X1 U11935 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9446) );
  NOR4_X1 U11936 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9445) );
  AND4_X1 U11937 ( .A1(n9448), .A2(n9447), .A3(n9446), .A4(n9445), .ZN(n9449)
         );
  NAND2_X1 U11938 ( .A1(n9450), .A2(n9449), .ZN(n9646) );
  INV_X1 U11939 ( .A(n9646), .ZN(n9451) );
  OR2_X1 U11940 ( .A1(n9648), .A2(n9451), .ZN(n9452) );
  AND3_X1 U11941 ( .A1(n9453), .A2(n10229), .A3(n9452), .ZN(n9563) );
  INV_X1 U11942 ( .A(n10390), .ZN(n11783) );
  AND2_X1 U11943 ( .A1(n13636), .A2(n13965), .ZN(n9555) );
  OR2_X1 U11944 ( .A1(n13638), .A2(n9555), .ZN(n10362) );
  INV_X1 U11945 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9471) );
  INV_X1 U11946 ( .A(n9557), .ZN(n9469) );
  NOR2_X1 U11947 ( .A1(n8276), .A2(n9456), .ZN(n9458) );
  XNOR2_X1 U11948 ( .A(n9458), .B(n9457), .ZN(n14152) );
  INV_X1 U11949 ( .A(n9658), .ZN(n10442) );
  NAND2_X1 U11950 ( .A1(n9461), .A2(n13636), .ZN(n9652) );
  AND2_X2 U11951 ( .A1(n13463), .A2(n9652), .ZN(n11910) );
  NOR2_X1 U11952 ( .A1(n13463), .A2(n9652), .ZN(n9459) );
  INV_X1 U11953 ( .A(n10273), .ZN(n9460) );
  NAND2_X1 U11954 ( .A1(n9460), .A2(n13965), .ZN(n14628) );
  NAND2_X1 U11955 ( .A1(n9433), .A2(n13952), .ZN(n13462) );
  INV_X1 U11956 ( .A(n13636), .ZN(n10274) );
  OR2_X1 U11957 ( .A1(n9433), .A2(n13965), .ZN(n9462) );
  NAND2_X1 U11958 ( .A1(n9461), .A2(n10274), .ZN(n13615) );
  NAND2_X1 U11959 ( .A1(n10236), .A2(n9658), .ZN(n10265) );
  OR2_X1 U11960 ( .A1(n10236), .A2(n9658), .ZN(n9463) );
  INV_X1 U11961 ( .A(n13468), .ZN(n13416) );
  OAI21_X1 U11962 ( .B1(n14660), .B2(n14571), .A(n13416), .ZN(n9468) );
  NAND2_X1 U11963 ( .A1(n11731), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9467) );
  NAND2_X1 U11964 ( .A1(n10244), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U11965 ( .A1(n10245), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9464) );
  NAND4_X4 U11966 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n13696) );
  NAND2_X1 U11967 ( .A1(n13696), .A2(n13398), .ZN(n10441) );
  OAI211_X1 U11968 ( .C1(n9469), .C2(n10442), .A(n9468), .B(n10441), .ZN(
        n14116) );
  NAND2_X1 U11969 ( .A1(n14116), .A2(n14663), .ZN(n9470) );
  OAI21_X1 U11970 ( .B1(n14663), .B2(n9471), .A(n9470), .ZN(P1_U3459) );
  INV_X1 U11971 ( .A(n14323), .ZN(n12206) );
  INV_X1 U11972 ( .A(n9472), .ZN(n9473) );
  OAI222_X1 U11973 ( .A1(P3_U3151), .A2(n12206), .B1(n12606), .B2(n9474), .C1(
        n12609), .C2(n9473), .ZN(P3_U3280) );
  INV_X1 U11974 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9485) );
  INV_X1 U11975 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U11976 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  NOR2_X1 U11977 ( .A1(n9482), .A2(n9479), .ZN(n9480) );
  MUX2_X1 U11978 ( .A(n9479), .B(n9480), .S(P1_IR_REG_11__SCAN_IN), .Z(n9484)
         );
  INV_X1 U11979 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U11980 ( .A1(n9482), .A2(n9481), .ZN(n9629) );
  INV_X1 U11981 ( .A(n9629), .ZN(n9483) );
  MUX2_X1 U11982 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9485), .S(n9636), .Z(n9490) );
  INV_X1 U11983 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14677) );
  INV_X1 U11984 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14671) );
  NOR2_X1 U11985 ( .A1(n10504), .A2(n14669), .ZN(n13768) );
  MUX2_X1 U11986 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14671), .S(n13775), .Z(
        n9486) );
  OAI21_X1 U11987 ( .B1(n13773), .B2(n13768), .A(n9486), .ZN(n13771) );
  OAI21_X1 U11988 ( .B1(n14671), .B2(n9487), .A(n13771), .ZN(n9506) );
  INV_X1 U11989 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U11990 ( .A(n9488), .B(P1_REG1_REG_8__SCAN_IN), .S(n10623), .Z(n9507) );
  NOR2_X1 U11991 ( .A1(n9506), .A2(n9507), .ZN(n13787) );
  NOR2_X1 U11992 ( .A1(n10623), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13785) );
  INV_X1 U11993 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14674) );
  MUX2_X1 U11994 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14674), .S(n13792), .Z(
        n13786) );
  OAI21_X1 U11995 ( .B1(n13792), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13784), .ZN(
        n9615) );
  MUX2_X1 U11996 ( .A(n14677), .B(P1_REG1_REG_10__SCAN_IN), .S(n10908), .Z(
        n9614) );
  OAI21_X1 U11997 ( .B1(n14677), .B2(n9496), .A(n9616), .ZN(n9489) );
  NOR2_X1 U11998 ( .A1(n9489), .A2(n9490), .ZN(n9627) );
  AOI21_X1 U11999 ( .B1(n9490), .B2(n9489), .A(n9627), .ZN(n9505) );
  NOR2_X1 U12000 ( .A1(n10504), .A2(n15113), .ZN(n13774) );
  INV_X1 U12001 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10537) );
  MUX2_X1 U12002 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10537), .S(n13775), .Z(
        n9491) );
  OAI21_X1 U12003 ( .B1(n13780), .B2(n13774), .A(n9491), .ZN(n13778) );
  NAND2_X1 U12004 ( .A1(n13775), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9510) );
  INV_X1 U12005 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n15076) );
  MUX2_X1 U12006 ( .A(n15076), .B(P1_REG2_REG_8__SCAN_IN), .S(n10623), .Z(
        n9509) );
  AOI21_X1 U12007 ( .B1(n13778), .B2(n9510), .A(n9509), .ZN(n13798) );
  NOR2_X1 U12008 ( .A1(n9492), .A2(n15076), .ZN(n13793) );
  INV_X1 U12009 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U12010 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9493), .S(n13792), .Z(n9494) );
  OAI21_X1 U12011 ( .B1(n13798), .B2(n13793), .A(n9494), .ZN(n13796) );
  NAND2_X1 U12012 ( .A1(n13792), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9612) );
  INV_X1 U12013 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U12014 ( .A(n9495), .B(P1_REG2_REG_10__SCAN_IN), .S(n10908), .Z(
        n9611) );
  AOI21_X1 U12015 ( .B1(n13796), .B2(n9612), .A(n9611), .ZN(n9622) );
  NOR2_X1 U12016 ( .A1(n9496), .A2(n9495), .ZN(n9499) );
  INV_X1 U12017 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10932) );
  MUX2_X1 U12018 ( .A(n10932), .B(P1_REG2_REG_11__SCAN_IN), .S(n9636), .Z(
        n9498) );
  NOR3_X1 U12019 ( .A1(n9622), .A2(n9499), .A3(n9498), .ZN(n9497) );
  NOR2_X1 U12020 ( .A1(n9497), .A2(n14534), .ZN(n9503) );
  OAI21_X1 U12021 ( .B1(n9622), .B2(n9499), .A(n9498), .ZN(n9635) );
  INV_X1 U12022 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14177) );
  INV_X1 U12023 ( .A(n9636), .ZN(n10914) );
  NAND2_X1 U12024 ( .A1(n13817), .A2(n10914), .ZN(n9501) );
  NAND2_X1 U12025 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9500) );
  OAI211_X1 U12026 ( .C1(n14177), .C2(n14541), .A(n9501), .B(n9500), .ZN(n9502) );
  AOI21_X1 U12027 ( .B1(n9503), .B2(n9635), .A(n9502), .ZN(n9504) );
  OAI21_X1 U12028 ( .B1(n9505), .B2(n14536), .A(n9504), .ZN(P1_U3254) );
  AOI21_X1 U12029 ( .B1(n9507), .B2(n9506), .A(n13787), .ZN(n9515) );
  INV_X1 U12030 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14170) );
  NAND2_X1 U12031 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10805) );
  OAI21_X1 U12032 ( .B1(n14541), .B2(n14170), .A(n10805), .ZN(n9508) );
  AOI21_X1 U12033 ( .B1(n10623), .B2(n13817), .A(n9508), .ZN(n9514) );
  INV_X1 U12034 ( .A(n13798), .ZN(n9512) );
  NAND3_X1 U12035 ( .A1(n13778), .A2(n9510), .A3(n9509), .ZN(n9511) );
  NAND3_X1 U12036 ( .A1(n13813), .A2(n9512), .A3(n9511), .ZN(n9513) );
  OAI211_X1 U12037 ( .C1(n9515), .C2(n14536), .A(n9514), .B(n9513), .ZN(
        P1_U3251) );
  INV_X1 U12038 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U12039 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  NAND2_X1 U12040 ( .A1(n8876), .A2(n13104), .ZN(n9687) );
  XNOR2_X1 U12041 ( .A(n9765), .B(n12663), .ZN(n9685) );
  XNOR2_X1 U12042 ( .A(n9687), .B(n9685), .ZN(n9683) );
  XOR2_X1 U12043 ( .A(n9683), .B(n9684), .Z(n9529) );
  INV_X1 U12044 ( .A(n12806), .ZN(n14685) );
  NAND2_X1 U12045 ( .A1(n8178), .A2(n12800), .ZN(n9524) );
  NAND2_X1 U12046 ( .A1(n12849), .A2(n12801), .ZN(n9523) );
  NAND2_X1 U12047 ( .A1(n9524), .A2(n9523), .ZN(n9773) );
  OAI22_X1 U12048 ( .A1(n12821), .A2(n14780), .B1(n9526), .B2(n9525), .ZN(
        n9527) );
  AOI21_X1 U12049 ( .B1(n14685), .B2(n9773), .A(n9527), .ZN(n9528) );
  OAI21_X1 U12050 ( .B1(n9529), .B2(n12792), .A(n9528), .ZN(P2_U3209) );
  INV_X1 U12051 ( .A(n14326), .ZN(n12165) );
  OAI222_X1 U12052 ( .A1(n12606), .A2(n9531), .B1(n12609), .B2(n9530), .C1(
        n12165), .C2(P3_U3151), .ZN(P3_U3279) );
  XNOR2_X1 U12053 ( .A(n9533), .B(n9532), .ZN(n9540) );
  INV_X1 U12054 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9534) );
  OAI22_X1 U12055 ( .A1(n14541), .A2(n6736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9534), .ZN(n9535) );
  AOI21_X1 U12056 ( .B1(n9544), .B2(n13817), .A(n9535), .ZN(n9539) );
  NAND2_X1 U12057 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13698) );
  OAI211_X1 U12058 ( .C1(n9238), .C2(n9537), .A(n13813), .B(n9536), .ZN(n9538)
         );
  OAI211_X1 U12059 ( .C1(n14536), .C2(n9540), .A(n9539), .B(n9538), .ZN(
        P1_U3244) );
  INV_X1 U12060 ( .A(n10913), .ZN(n9542) );
  INV_X1 U12061 ( .A(n12917), .ZN(n12924) );
  OAI222_X1 U12062 ( .A1(n13272), .A2(n9542), .B1(n12924), .B2(P2_U3088), .C1(
        n9541), .C2(n13269), .ZN(P2_U3316) );
  OAI222_X1 U12063 ( .A1(n14145), .A2(n9543), .B1(n14148), .B2(n9542), .C1(
        n9636), .C2(P1_U3086), .ZN(P1_U3344) );
  NAND2_X1 U12064 ( .A1(n11702), .A2(n9544), .ZN(n9545) );
  AOI21_X1 U12065 ( .B1(n13417), .B2(n6824), .A(n14550), .ZN(n9548) );
  OR2_X1 U12066 ( .A1(n13638), .A2(n9233), .ZN(n13387) );
  NOR2_X1 U12067 ( .A1(n9548), .A2(n13662), .ZN(n10461) );
  NOR2_X1 U12068 ( .A1(n13473), .A2(n9658), .ZN(n14579) );
  INV_X1 U12069 ( .A(n14579), .ZN(n9550) );
  NAND2_X1 U12070 ( .A1(n13473), .A2(n9658), .ZN(n9549) );
  NAND2_X1 U12071 ( .A1(n9550), .A2(n9549), .ZN(n9558) );
  XNOR2_X1 U12072 ( .A(n9558), .B(n7412), .ZN(n10460) );
  NOR3_X1 U12073 ( .A1(n10461), .A2(n14550), .A3(n10460), .ZN(n9562) );
  NAND2_X1 U12074 ( .A1(n10245), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U12075 ( .A1(n11731), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9553) );
  INV_X2 U12076 ( .A(n11750), .ZN(n11778) );
  NAND2_X1 U12077 ( .A1(n11778), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U12078 ( .A1(n10244), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U12079 ( .A1(n13694), .A2(n13398), .ZN(n9670) );
  OAI21_X1 U12080 ( .B1(n10461), .B2(n9671), .A(n9670), .ZN(n10464) );
  INV_X1 U12081 ( .A(n9555), .ZN(n9556) );
  NOR2_X1 U12082 ( .A1(n9558), .A2(n6570), .ZN(n10458) );
  INV_X1 U12083 ( .A(n10458), .ZN(n9559) );
  OAI21_X1 U12084 ( .B1(n10237), .B2(n14655), .A(n9559), .ZN(n9561) );
  XNOR2_X1 U12085 ( .A(n10265), .B(n13417), .ZN(n10467) );
  AOI21_X1 U12086 ( .B1(n14628), .B2(n14642), .A(n10467), .ZN(n9560) );
  NOR4_X1 U12087 ( .A1(n9562), .A2(n10464), .A3(n9561), .A4(n9560), .ZN(n14588) );
  NAND2_X1 U12088 ( .A1(n14676), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9565) );
  OAI21_X1 U12089 ( .B1(n14588), .B2(n14676), .A(n9565), .ZN(P1_U3529) );
  AOI21_X1 U12090 ( .B1(n9570), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9566), .ZN(
        n14697) );
  MUX2_X1 U12091 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7832), .S(n14702), .Z(
        n14696) );
  NAND2_X1 U12092 ( .A1(n14697), .A2(n14696), .ZN(n14695) );
  OAI21_X1 U12093 ( .B1(n14702), .B2(P2_REG1_REG_9__SCAN_IN), .A(n14695), .ZN(
        n9568) );
  INV_X1 U12094 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14831) );
  MUX2_X1 U12095 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14831), .S(n9888), .Z(
        n9567) );
  NOR2_X1 U12096 ( .A1(n9568), .A2(n9567), .ZN(n12922) );
  AOI211_X1 U12097 ( .C1(n9568), .C2(n9567), .A(n11644), .B(n12922), .ZN(n9576) );
  AOI21_X1 U12098 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9570), .A(n9569), .ZN(
        n14700) );
  MUX2_X1 U12099 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10821), .S(n14702), .Z(
        n14699) );
  NAND2_X1 U12100 ( .A1(n14700), .A2(n14699), .ZN(n14698) );
  OAI21_X1 U12101 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n14702), .A(n14698), .ZN(
        n9572) );
  MUX2_X1 U12102 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10981), .S(n9888), .Z(
        n9571) );
  NOR2_X1 U12103 ( .A1(n9572), .A2(n9571), .ZN(n9895) );
  AOI211_X1 U12104 ( .C1(n9572), .C2(n9571), .A(n15310), .B(n9895), .ZN(n9575)
         );
  NAND2_X1 U12105 ( .A1(n14718), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U12106 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10765)
         );
  OAI211_X1 U12107 ( .C1(n12925), .C2(n9888), .A(n9573), .B(n10765), .ZN(n9574) );
  OR3_X1 U12108 ( .A1(n9576), .A2(n9575), .A3(n9574), .ZN(P2_U3224) );
  INV_X1 U12109 ( .A(n9982), .ZN(n9577) );
  OR2_X1 U12110 ( .A1(n9962), .A2(P3_U3151), .ZN(n11622) );
  NAND2_X1 U12111 ( .A1(n9577), .A2(n11622), .ZN(n9589) );
  NAND2_X1 U12112 ( .A1(n11569), .A2(n9962), .ZN(n9578) );
  AND2_X1 U12113 ( .A1(n9579), .A2(n9578), .ZN(n9587) );
  INV_X1 U12114 ( .A(n9593), .ZN(n9580) );
  MUX2_X1 U12115 ( .A(n12140), .B(n9580), .S(n6831), .Z(n14357) );
  INV_X4 U12116 ( .A(n12223), .ZN(n12164) );
  NAND2_X1 U12117 ( .A1(n9593), .A2(n12164), .ZN(n14313) );
  INV_X1 U12118 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9581) );
  MUX2_X1 U12119 ( .A(n9581), .B(P3_REG1_REG_2__SCAN_IN), .S(n9782), .Z(n9586)
         );
  INV_X1 U12120 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U12121 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9582), .ZN(n9583) );
  INV_X1 U12122 ( .A(n9583), .ZN(n9995) );
  OR2_X1 U12123 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9583), .ZN(n9584) );
  OAI21_X1 U12124 ( .B1(n9601), .B2(n9995), .A(n9584), .ZN(n9851) );
  OR2_X1 U12125 ( .A1(n9851), .A2(n8259), .ZN(n9849) );
  NAND2_X1 U12126 ( .A1(n9849), .A2(n9584), .ZN(n9585) );
  OAI21_X1 U12127 ( .B1(n9586), .B2(n9585), .A(n9787), .ZN(n9600) );
  INV_X1 U12128 ( .A(n9587), .ZN(n9588) );
  AND2_X1 U12129 ( .A1(n9589), .A2(n9588), .ZN(n14899) );
  INV_X1 U12130 ( .A(n14899), .ZN(n14878) );
  INV_X1 U12131 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9590) );
  INV_X1 U12132 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n14917) );
  OAI22_X1 U12133 ( .A1(n14878), .A2(n9590), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14917), .ZN(n9599) );
  INV_X1 U12134 ( .A(n9591), .ZN(n9592) );
  INV_X1 U12135 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15262) );
  INV_X1 U12136 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9603) );
  NOR2_X1 U12137 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n9603), .ZN(n9994) );
  NAND2_X1 U12138 ( .A1(n8245), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9594) );
  OAI21_X1 U12139 ( .B1(n9601), .B2(n9994), .A(n9594), .ZN(n9854) );
  INV_X1 U12140 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n14948) );
  OR2_X1 U12141 ( .A1(n9854), .A2(n14948), .ZN(n9856) );
  OAI21_X1 U12142 ( .B1(n9596), .B2(n9595), .A(n9790), .ZN(n9597) );
  AND2_X1 U12143 ( .A1(n14843), .A2(n9597), .ZN(n9598) );
  AOI211_X1 U12144 ( .C1(n14895), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9610)
         );
  MUX2_X1 U12145 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12164), .Z(n9604) );
  INV_X1 U12146 ( .A(n9601), .ZN(n9859) );
  XNOR2_X1 U12147 ( .A(n9604), .B(n9859), .ZN(n9848) );
  INV_X1 U12148 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9602) );
  MUX2_X1 U12149 ( .A(n9603), .B(n9602), .S(n12164), .Z(n9999) );
  AND2_X1 U12150 ( .A1(n9999), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U12151 ( .A1(n9848), .A2(n10004), .ZN(n9607) );
  INV_X1 U12152 ( .A(n9604), .ZN(n9605) );
  NAND2_X1 U12153 ( .A1(n9605), .A2(n9859), .ZN(n9606) );
  NAND2_X1 U12154 ( .A1(n9607), .A2(n9606), .ZN(n9780) );
  MUX2_X1 U12155 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12164), .Z(n9781) );
  XNOR2_X1 U12156 ( .A(n9781), .B(n9782), .ZN(n9779) );
  XNOR2_X1 U12157 ( .A(n9780), .B(n9779), .ZN(n9608) );
  AND2_X1 U12158 ( .A1(P3_U3897), .A2(n6831), .ZN(n14903) );
  NAND2_X1 U12159 ( .A1(n9608), .A2(n14903), .ZN(n9609) );
  OAI211_X1 U12160 ( .C1(n14357), .C2(n9788), .A(n9610), .B(n9609), .ZN(
        P3_U3184) );
  NAND3_X1 U12161 ( .A1(n13796), .A2(n9612), .A3(n9611), .ZN(n9613) );
  NAND2_X1 U12162 ( .A1(n9613), .A2(n13813), .ZN(n9621) );
  AOI21_X1 U12163 ( .B1(n9615), .B2(n9614), .A(n14536), .ZN(n9617) );
  NAND2_X1 U12164 ( .A1(n9617), .A2(n9616), .ZN(n9620) );
  INV_X1 U12165 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U12166 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14438)
         );
  OAI21_X1 U12167 ( .B1(n14541), .B2(n15010), .A(n14438), .ZN(n9618) );
  AOI21_X1 U12168 ( .B1(n10908), .B2(n13817), .A(n9618), .ZN(n9619) );
  OAI211_X1 U12169 ( .C1(n9622), .C2(n9621), .A(n9620), .B(n9619), .ZN(
        P1_U3253) );
  INV_X1 U12170 ( .A(n11055), .ZN(n9643) );
  INV_X1 U12171 ( .A(n9897), .ZN(n10997) );
  OAI222_X1 U12172 ( .A1(n13272), .A2(n9643), .B1(n10997), .B2(P2_U3088), .C1(
        n9623), .C2(n13269), .ZN(P2_U3315) );
  INV_X1 U12173 ( .A(n12210), .ZN(n14356) );
  INV_X1 U12174 ( .A(n9624), .ZN(n9626) );
  INV_X1 U12175 ( .A(SI_17_), .ZN(n9625) );
  OAI222_X1 U12176 ( .A1(n14356), .A2(P3_U3151), .B1(n12609), .B2(n9626), .C1(
        n9625), .C2(n12606), .ZN(P3_U3278) );
  NAND2_X1 U12177 ( .A1(n9629), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9628) );
  MUX2_X1 U12178 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9628), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n9630) );
  INV_X1 U12179 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14290) );
  INV_X1 U12180 ( .A(n11056), .ZN(n10152) );
  AOI22_X1 U12181 ( .A1(n11056), .A2(n14290), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n10152), .ZN(n9631) );
  NOR2_X1 U12182 ( .A1(n9632), .A2(n9631), .ZN(n10151) );
  AOI21_X1 U12183 ( .B1(n9632), .B2(n9631), .A(n10151), .ZN(n9642) );
  INV_X1 U12184 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n15137) );
  NOR2_X1 U12185 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15137), .ZN(n9634) );
  NOR2_X1 U12186 ( .A1(n6779), .A2(n10152), .ZN(n9633) );
  AOI211_X1 U12187 ( .C1(n14525), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9634), .B(
        n9633), .ZN(n9641) );
  OAI21_X1 U12188 ( .B1(n10932), .B2(n9636), .A(n9635), .ZN(n9638) );
  INV_X1 U12189 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U12190 ( .A1(n11056), .A2(n15154), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10152), .ZN(n9637) );
  NOR2_X1 U12191 ( .A1(n9637), .A2(n9638), .ZN(n10148) );
  AOI21_X1 U12192 ( .B1(n9638), .B2(n9637), .A(n10148), .ZN(n9639) );
  OR2_X1 U12193 ( .A1(n9639), .A2(n14534), .ZN(n9640) );
  OAI211_X1 U12194 ( .C1(n9642), .C2(n14536), .A(n9641), .B(n9640), .ZN(
        P1_U3255) );
  OAI222_X1 U12195 ( .A1(n14145), .A2(n9644), .B1(n14148), .B2(n9643), .C1(
        n10152), .C2(P1_U3086), .ZN(P1_U3343) );
  NOR2_X1 U12196 ( .A1(n9646), .A2(n9645), .ZN(n9647) );
  OR2_X1 U12197 ( .A1(n9648), .A2(n9647), .ZN(n9650) );
  AND2_X1 U12198 ( .A1(n9650), .A2(n9649), .ZN(n9669) );
  NAND2_X1 U12199 ( .A1(n10390), .A2(n9669), .ZN(n9651) );
  NAND2_X1 U12200 ( .A1(n9651), .A2(n10229), .ZN(n10365) );
  INV_X1 U12201 ( .A(n9652), .ZN(n13639) );
  AND2_X2 U12202 ( .A1(n9653), .A2(n13639), .ZN(n9654) );
  INV_X4 U12203 ( .A(n11910), .ZN(n11941) );
  XNOR2_X1 U12204 ( .A(n9655), .B(n11941), .ZN(n9734) );
  XNOR2_X1 U12205 ( .A(n9734), .B(n9737), .ZN(n9664) );
  INV_X1 U12206 ( .A(n10364), .ZN(n9657) );
  INV_X1 U12207 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12208 ( .A1(n9707), .A2(n9662), .ZN(n9663) );
  NAND2_X1 U12209 ( .A1(n9664), .A2(n9663), .ZN(n9735) );
  OAI21_X1 U12210 ( .B1(n9664), .B2(n9663), .A(n9735), .ZN(n9668) );
  INV_X1 U12211 ( .A(n10231), .ZN(n9666) );
  NAND2_X1 U12212 ( .A1(n14655), .A2(n13638), .ZN(n9665) );
  NOR2_X1 U12213 ( .A1(n9666), .A2(n9665), .ZN(n9667) );
  NAND3_X1 U12214 ( .A1(n10390), .A2(n9669), .A3(n9667), .ZN(n14458) );
  NAND2_X1 U12215 ( .A1(n9668), .A2(n14440), .ZN(n9675) );
  OAI21_X1 U12216 ( .B1(n9671), .B2(n13387), .A(n9670), .ZN(n9673) );
  NAND2_X1 U12217 ( .A1(n10365), .A2(n9672), .ZN(n9745) );
  AOI22_X1 U12218 ( .A1(n14433), .A2(n9673), .B1(n9745), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9674) );
  OAI211_X1 U12219 ( .C1(n10237), .C2(n13414), .A(n9675), .B(n9674), .ZN(
        P1_U3222) );
  NAND2_X1 U12220 ( .A1(n14688), .A2(n12619), .ZN(n12794) );
  INV_X1 U12221 ( .A(n12794), .ZN(n12813) );
  NAND2_X1 U12222 ( .A1(n12813), .A2(n8862), .ZN(n9677) );
  MUX2_X1 U12223 ( .A(n9677), .B(n12821), .S(n9676), .Z(n9681) );
  NOR2_X1 U12224 ( .A1(n12806), .A2(n14754), .ZN(n9678) );
  AOI22_X1 U12225 ( .A1(n9679), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n9678), .B2(
        n8178), .ZN(n9680) );
  OAI211_X1 U12226 ( .C1(n12792), .C2(n9682), .A(n9681), .B(n9680), .ZN(
        P2_U3204) );
  NAND2_X1 U12227 ( .A1(n12848), .A2(n12664), .ZN(n9906) );
  XNOR2_X1 U12228 ( .A(n9913), .B(n9906), .ZN(n9702) );
  INV_X1 U12229 ( .A(n9685), .ZN(n9686) );
  NAND2_X1 U12230 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  XNOR2_X1 U12231 ( .A(n9757), .B(n12673), .ZN(n9693) );
  NAND2_X1 U12232 ( .A1(n9689), .A2(n9693), .ZN(n9690) );
  NAND2_X1 U12233 ( .A1(n9691), .A2(n9690), .ZN(n9723) );
  AND2_X1 U12234 ( .A1(n9702), .A2(n9691), .ZN(n9692) );
  OAI21_X1 U12235 ( .B1(n9702), .B2(n9721), .A(n9912), .ZN(n9705) );
  INV_X1 U12236 ( .A(n9693), .ZN(n9694) );
  NAND3_X1 U12237 ( .A1(n12813), .A2(n12849), .A3(n9694), .ZN(n9703) );
  AOI21_X1 U12238 ( .B1(n14690), .B2(n14794), .A(n9695), .ZN(n9701) );
  NAND2_X1 U12239 ( .A1(n12849), .A2(n12800), .ZN(n9697) );
  NAND2_X1 U12240 ( .A1(n12847), .A2(n12801), .ZN(n9696) );
  NAND2_X1 U12241 ( .A1(n9697), .A2(n9696), .ZN(n9949) );
  INV_X1 U12242 ( .A(n14694), .ZN(n12803) );
  INV_X1 U12243 ( .A(n9955), .ZN(n9699) );
  AOI22_X1 U12244 ( .A1(n14685), .A2(n9949), .B1(n12803), .B2(n9699), .ZN(
        n9700) );
  OAI211_X1 U12245 ( .C1(n9703), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9704)
         );
  AOI21_X1 U12246 ( .B1(n9705), .B2(n14688), .A(n9704), .ZN(n9706) );
  INV_X1 U12247 ( .A(n9706), .ZN(P2_U3202) );
  OAI21_X1 U12248 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(n13697) );
  NAND2_X1 U12249 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9745), .ZN(n9710) );
  OAI21_X1 U12250 ( .B1(n14456), .B2(n10441), .A(n9710), .ZN(n9711) );
  AOI21_X1 U12251 ( .B1(n13697), .B2(n14440), .A(n9711), .ZN(n9712) );
  OAI21_X1 U12252 ( .B1(n10442), .B2(n13414), .A(n9712), .ZN(P1_U3232) );
  INV_X1 U12253 ( .A(n12226), .ZN(n12231) );
  INV_X1 U12254 ( .A(n9713), .ZN(n9715) );
  INV_X1 U12255 ( .A(SI_18_), .ZN(n9714) );
  OAI222_X1 U12256 ( .A1(n12231), .A2(P3_U3151), .B1(n12609), .B2(n9715), .C1(
        n9714), .C2(n12606), .ZN(P3_U3277) );
  INV_X1 U12257 ( .A(n11061), .ZN(n9719) );
  NAND2_X1 U12258 ( .A1(n10103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9716) );
  INV_X1 U12259 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n15078) );
  XNOR2_X1 U12260 ( .A(n9716), .B(n15078), .ZN(n11064) );
  OAI222_X1 U12261 ( .A1(n14145), .A2(n11062), .B1(n14148), .B2(n9719), .C1(
        n11064), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U12262 ( .A1(n12609), .A2(n9718), .B1(n12606), .B2(n9717), .C1(
        P3_U3151), .C2(n12237), .ZN(P3_U3276) );
  OAI222_X1 U12263 ( .A1(n13269), .A2(n9720), .B1(n10999), .B2(P2_U3088), .C1(
        n13272), .C2(n9719), .ZN(P2_U3314) );
  INV_X1 U12264 ( .A(n9721), .ZN(n9722) );
  AOI211_X1 U12265 ( .C1(n9724), .C2(n9723), .A(n12792), .B(n9722), .ZN(n9730)
         );
  AOI22_X1 U12266 ( .A1(n14694), .A2(n9189), .B1(P2_STATE_REG_SCAN_IN), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n9729) );
  INV_X1 U12267 ( .A(n12848), .ZN(n9725) );
  OAI22_X1 U12268 ( .A1(n9726), .A2(n14378), .B1(n9725), .B2(n14754), .ZN(
        n9754) );
  INV_X1 U12269 ( .A(n9754), .ZN(n9727) );
  OAI22_X1 U12270 ( .A1(n9727), .A2(n12806), .B1(n14789), .B2(n12821), .ZN(
        n9728) );
  OR3_X1 U12271 ( .A1(n9730), .A2(n9729), .A3(n9728), .ZN(P2_U3190) );
  NAND2_X1 U12272 ( .A1(n6551), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12273 ( .A1(n6562), .A2(n13712), .ZN(n9731) );
  INV_X1 U12274 ( .A(n9734), .ZN(n9736) );
  OAI21_X1 U12275 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n10344) );
  AOI22_X1 U12276 ( .A1(n6559), .A2(n13694), .B1(n11821), .B2(n14573), .ZN(
        n9738) );
  XNOR2_X1 U12277 ( .A(n9738), .B(n11941), .ZN(n10342) );
  INV_X1 U12278 ( .A(n6565), .ZN(n9739) );
  INV_X1 U12279 ( .A(n13694), .ZN(n10436) );
  OAI22_X1 U12280 ( .A1(n9656), .A2(n10436), .B1(n14590), .B2(n11884), .ZN(
        n10340) );
  XNOR2_X1 U12281 ( .A(n10342), .B(n10340), .ZN(n10343) );
  XNOR2_X1 U12282 ( .A(n10344), .B(n10343), .ZN(n9740) );
  NAND2_X1 U12283 ( .A1(n9740), .A2(n14440), .ZN(n9747) );
  NAND2_X1 U12284 ( .A1(n10245), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9744) );
  INV_X4 U12285 ( .A(n11731), .ZN(n11769) );
  NAND2_X1 U12286 ( .A1(n11778), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U12287 ( .A1(n10244), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9741) );
  OAI22_X1 U12288 ( .A1(n7412), .A2(n13387), .B1(n10271), .B2(n13388), .ZN(
        n14569) );
  AOI22_X1 U12289 ( .A1(n14433), .A2(n14569), .B1(n9745), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9746) );
  OAI211_X1 U12290 ( .C1(n14590), .C2(n13414), .A(n9747), .B(n9746), .ZN(
        P1_U3237) );
  XNOR2_X1 U12291 ( .A(n9749), .B(n9748), .ZN(n14785) );
  NAND3_X1 U12292 ( .A1(n9772), .A2(n9752), .A3(n9751), .ZN(n9753) );
  AOI21_X1 U12293 ( .B1(n9750), .B2(n9753), .A(n13189), .ZN(n9755) );
  NOR2_X1 U12294 ( .A1(n9755), .A2(n9754), .ZN(n14788) );
  MUX2_X1 U12295 ( .A(n9756), .B(n14788), .S(n6558), .Z(n9762) );
  NAND2_X1 U12296 ( .A1(n9766), .A2(n9757), .ZN(n9758) );
  NAND2_X1 U12297 ( .A1(n9758), .A2(n10011), .ZN(n9759) );
  NOR2_X1 U12298 ( .A1(n9952), .A2(n9759), .ZN(n14786) );
  OAI22_X1 U12299 ( .A1(n14739), .A2(n14789), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14751), .ZN(n9760) );
  AOI21_X1 U12300 ( .B1(n14786), .B2(n14731), .A(n9760), .ZN(n9761) );
  OAI211_X1 U12301 ( .C1(n14785), .C2(n13114), .A(n9762), .B(n9761), .ZN(
        P2_U3262) );
  XNOR2_X1 U12302 ( .A(n9764), .B(n9763), .ZN(n14777) );
  AOI21_X1 U12303 ( .B1(n10074), .B2(n9765), .A(n13104), .ZN(n9767) );
  NAND2_X1 U12304 ( .A1(n9767), .A2(n9766), .ZN(n14778) );
  INV_X1 U12305 ( .A(n14778), .ZN(n9777) );
  NAND2_X1 U12306 ( .A1(n14736), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9769) );
  NAND2_X1 U12307 ( .A1(n14734), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9768) );
  OAI211_X1 U12308 ( .C1(n14739), .C2(n14780), .A(n9769), .B(n9768), .ZN(n9776) );
  NAND3_X1 U12309 ( .A1(n10067), .A2(n9770), .A3(n8181), .ZN(n9771) );
  AOI21_X1 U12310 ( .B1(n9772), .B2(n9771), .A(n13189), .ZN(n9774) );
  NOR2_X1 U12311 ( .A1(n9774), .A2(n9773), .ZN(n14779) );
  NOR2_X1 U12312 ( .A1(n14779), .A2(n14736), .ZN(n9775) );
  AOI211_X1 U12313 ( .C1(n9777), .C2(n14731), .A(n9776), .B(n9775), .ZN(n9778)
         );
  OAI21_X1 U12314 ( .B1(n13114), .B2(n14777), .A(n9778), .ZN(P2_U3263) );
  MUX2_X1 U12315 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12164), .Z(n9804) );
  XNOR2_X1 U12316 ( .A(n9804), .B(n9805), .ZN(n9802) );
  NAND2_X1 U12317 ( .A1(n9780), .A2(n9779), .ZN(n9785) );
  INV_X1 U12318 ( .A(n9781), .ZN(n9783) );
  NAND2_X1 U12319 ( .A1(n9783), .A2(n9782), .ZN(n9784) );
  NAND2_X1 U12320 ( .A1(n9785), .A2(n9784), .ZN(n9803) );
  XOR2_X1 U12321 ( .A(n9802), .B(n9803), .Z(n9801) );
  NAND2_X1 U12322 ( .A1(n9788), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U12323 ( .A1(n9787), .A2(n9786), .ZN(n9811) );
  XNOR2_X1 U12324 ( .A(n9811), .B(n9805), .ZN(n9809) );
  XOR2_X1 U12325 ( .A(n9809), .B(P3_REG1_REG_3__SCAN_IN), .Z(n9798) );
  NAND2_X1 U12326 ( .A1(n9788), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U12327 ( .A1(n9792), .A2(n9810), .ZN(n9817) );
  INV_X1 U12328 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15066) );
  OAI21_X1 U12329 ( .B1(n9794), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9818), .ZN(
        n9795) );
  NAND2_X1 U12330 ( .A1(n14843), .A2(n9795), .ZN(n9797) );
  NOR2_X1 U12331 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8295), .ZN(n10166) );
  AOI21_X1 U12332 ( .B1(n14899), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10166), .ZN(
        n9796) );
  OAI211_X1 U12333 ( .C1(n9798), .C2(n14313), .A(n9797), .B(n9796), .ZN(n9799)
         );
  AOI21_X1 U12334 ( .B1(n14906), .B2(n9805), .A(n9799), .ZN(n9800) );
  OAI21_X1 U12335 ( .B1(n9801), .B2(n14882), .A(n9800), .ZN(P3_U3185) );
  MUX2_X1 U12336 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12164), .Z(n9830) );
  XNOR2_X1 U12337 ( .A(n9830), .B(n9836), .ZN(n9828) );
  NAND2_X1 U12338 ( .A1(n9803), .A2(n9802), .ZN(n9808) );
  INV_X1 U12339 ( .A(n9804), .ZN(n9806) );
  NAND2_X1 U12340 ( .A1(n9806), .A2(n9805), .ZN(n9807) );
  NAND2_X1 U12341 ( .A1(n9808), .A2(n9807), .ZN(n9829) );
  XOR2_X1 U12342 ( .A(n9828), .B(n9829), .Z(n9827) );
  MUX2_X1 U12343 ( .A(n10329), .B(P3_REG1_REG_4__SCAN_IN), .S(n9836), .Z(n9815) );
  NAND2_X1 U12344 ( .A1(n9809), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U12345 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  NAND2_X1 U12346 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U12347 ( .A1(n9814), .A2(n9815), .ZN(n9834) );
  OAI21_X1 U12348 ( .B1(n9815), .B2(n9814), .A(n9834), .ZN(n9816) );
  INV_X1 U12349 ( .A(n9816), .ZN(n9824) );
  INV_X1 U12350 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15258) );
  MUX2_X1 U12351 ( .A(n15258), .B(P3_REG2_REG_4__SCAN_IN), .S(n9836), .Z(n9820) );
  OAI21_X1 U12352 ( .B1(n9820), .B2(n9819), .A(n9835), .ZN(n9821) );
  NAND2_X1 U12353 ( .A1(n14843), .A2(n9821), .ZN(n9823) );
  AND2_X1 U12354 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10409) );
  AOI21_X1 U12355 ( .B1(n14899), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10409), .ZN(
        n9822) );
  OAI211_X1 U12356 ( .C1(n9824), .C2(n14313), .A(n9823), .B(n9822), .ZN(n9825)
         );
  AOI21_X1 U12357 ( .B1(n14906), .B2(n9836), .A(n9825), .ZN(n9826) );
  OAI21_X1 U12358 ( .B1(n9827), .B2(n14882), .A(n9826), .ZN(P3_U3186) );
  MUX2_X1 U12359 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12164), .Z(n9864) );
  XNOR2_X1 U12360 ( .A(n9864), .B(n9874), .ZN(n9862) );
  NAND2_X1 U12361 ( .A1(n9829), .A2(n9828), .ZN(n9833) );
  INV_X1 U12362 ( .A(n9830), .ZN(n9831) );
  NAND2_X1 U12363 ( .A1(n9831), .A2(n9836), .ZN(n9832) );
  NAND2_X1 U12364 ( .A1(n9833), .A2(n9832), .ZN(n9863) );
  XOR2_X1 U12365 ( .A(n9862), .B(n9863), .Z(n9847) );
  INV_X1 U12366 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10329) );
  XNOR2_X1 U12367 ( .A(n9876), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n9844) );
  AND2_X1 U12368 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10605) );
  INV_X1 U12369 ( .A(n14843), .ZN(n14912) );
  INV_X1 U12370 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9840) );
  AOI21_X1 U12371 ( .B1(n9840), .B2(n9839), .A(n9871), .ZN(n9841) );
  NOR2_X1 U12372 ( .A1(n14912), .A2(n9841), .ZN(n9842) );
  AOI211_X1 U12373 ( .C1(n14899), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10605), .B(
        n9842), .ZN(n9843) );
  OAI21_X1 U12374 ( .B1(n9844), .B2(n14313), .A(n9843), .ZN(n9845) );
  AOI21_X1 U12375 ( .B1(n9874), .B2(n14906), .A(n9845), .ZN(n9846) );
  OAI21_X1 U12376 ( .B1(n9847), .B2(n14882), .A(n9846), .ZN(P3_U3187) );
  XOR2_X1 U12377 ( .A(n10004), .B(n9848), .Z(n9861) );
  INV_X1 U12378 ( .A(n9849), .ZN(n9850) );
  AOI21_X1 U12379 ( .B1(n8259), .B2(n9851), .A(n9850), .ZN(n9853) );
  AOI22_X1 U12380 ( .A1(n14899), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9852) );
  OAI21_X1 U12381 ( .B1(n9853), .B2(n14313), .A(n9852), .ZN(n9858) );
  NAND2_X1 U12382 ( .A1(n9854), .A2(n14948), .ZN(n9855) );
  AOI21_X1 U12383 ( .B1(n9856), .B2(n9855), .A(n14912), .ZN(n9857) );
  AOI211_X1 U12384 ( .C1(n14906), .C2(n9859), .A(n9858), .B(n9857), .ZN(n9860)
         );
  OAI21_X1 U12385 ( .B1(n14882), .B2(n9861), .A(n9860), .ZN(P3_U3183) );
  MUX2_X1 U12386 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12164), .Z(n9922) );
  XNOR2_X1 U12387 ( .A(n9922), .B(n6555), .ZN(n9920) );
  NAND2_X1 U12388 ( .A1(n9863), .A2(n9862), .ZN(n9867) );
  INV_X1 U12389 ( .A(n9864), .ZN(n9865) );
  NAND2_X1 U12390 ( .A1(n9865), .A2(n9874), .ZN(n9866) );
  NAND2_X1 U12391 ( .A1(n9867), .A2(n9866), .ZN(n9921) );
  XOR2_X1 U12392 ( .A(n9920), .B(n9921), .Z(n9886) );
  INV_X1 U12393 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U12394 ( .A1(n6555), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n9868), .B2(
        n9934), .ZN(n9933) );
  INV_X1 U12395 ( .A(n9869), .ZN(n9870) );
  XOR2_X1 U12396 ( .A(n9933), .B(n6722), .Z(n9883) );
  INV_X1 U12397 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U12398 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9872), .ZN(n10662) );
  AOI21_X1 U12399 ( .B1(n14899), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10662), .ZN(
        n9882) );
  INV_X1 U12400 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9877) );
  INV_X1 U12401 ( .A(n9873), .ZN(n9875) );
  OAI22_X1 U12402 ( .A1(n9877), .A2(n9876), .B1(n9875), .B2(n9874), .ZN(n9879)
         );
  INV_X1 U12403 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U12404 ( .A1(n6555), .A2(n10726), .B1(P3_REG1_REG_6__SCAN_IN), .B2(
        n9934), .ZN(n9878) );
  OAI21_X1 U12405 ( .B1(n9879), .B2(n9878), .A(n9927), .ZN(n9880) );
  NAND2_X1 U12406 ( .A1(n14895), .A2(n9880), .ZN(n9881) );
  OAI211_X1 U12407 ( .C1(n14912), .C2(n9883), .A(n9882), .B(n9881), .ZN(n9884)
         );
  AOI21_X1 U12408 ( .B1(n6555), .B2(n14906), .A(n9884), .ZN(n9885) );
  OAI21_X1 U12409 ( .B1(n9886), .B2(n14882), .A(n9885), .ZN(P3_U3188) );
  NOR2_X1 U12410 ( .A1(n9897), .A2(n9891), .ZN(n9887) );
  AOI21_X1 U12411 ( .B1(n9891), .B2(n9897), .A(n9887), .ZN(n9893) );
  INV_X1 U12412 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15047) );
  NOR2_X1 U12413 ( .A1(n9888), .A2(n14831), .ZN(n12916) );
  MUX2_X1 U12414 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15047), .S(n12917), .Z(
        n9889) );
  OAI21_X1 U12415 ( .B1(n12922), .B2(n12916), .A(n9889), .ZN(n12920) );
  OAI21_X1 U12416 ( .B1(n15047), .B2(n12924), .A(n12920), .ZN(n9892) );
  NOR2_X1 U12417 ( .A1(n10997), .A2(n9891), .ZN(n9890) );
  AOI211_X1 U12418 ( .C1(n10997), .C2(n9891), .A(n9890), .B(n9892), .ZN(n10986) );
  AOI21_X1 U12419 ( .B1(n9893), .B2(n9892), .A(n10986), .ZN(n9905) );
  NAND2_X1 U12420 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14691)
         );
  OAI21_X1 U12421 ( .B1(n12925), .B2(n10997), .A(n14691), .ZN(n9894) );
  AOI21_X1 U12422 ( .B1(n14718), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n9894), .ZN(
        n9904) );
  AOI21_X1 U12423 ( .B1(n9896), .B2(P2_REG2_REG_10__SCAN_IN), .A(n9895), .ZN(
        n12929) );
  MUX2_X1 U12424 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11024), .S(n12917), .Z(
        n12928) );
  NAND2_X1 U12425 ( .A1(n12929), .A2(n12928), .ZN(n12927) );
  NAND2_X1 U12426 ( .A1(n12924), .A2(n11024), .ZN(n9900) );
  OR2_X1 U12427 ( .A1(n9897), .A2(n15207), .ZN(n9899) );
  INV_X1 U12428 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n15207) );
  NAND2_X1 U12429 ( .A1(n9897), .A2(n15207), .ZN(n9898) );
  AND2_X1 U12430 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  AOI21_X1 U12431 ( .B1(n12927), .B2(n9900), .A(n9901), .ZN(n10996) );
  AND3_X1 U12432 ( .A1(n12927), .A2(n9901), .A3(n9900), .ZN(n9902) );
  OAI21_X1 U12433 ( .B1(n10996), .B2(n9902), .A(n6547), .ZN(n9903) );
  OAI211_X1 U12434 ( .C1(n9905), .C2(n11644), .A(n9904), .B(n9903), .ZN(
        P2_U3226) );
  INV_X1 U12435 ( .A(n9913), .ZN(n9907) );
  NAND2_X1 U12436 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  NAND2_X1 U12437 ( .A1(n9912), .A2(n9908), .ZN(n9909) );
  NAND2_X1 U12438 ( .A1(n12847), .A2(n12664), .ZN(n10007) );
  XNOR2_X1 U12439 ( .A(n10006), .B(n10007), .ZN(n9914) );
  AOI22_X1 U12440 ( .A1(n12800), .A2(n12848), .B1(n12846), .B2(n12801), .ZN(
        n10135) );
  NAND2_X1 U12441 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n12866) );
  INV_X1 U12442 ( .A(n9910), .ZN(n10059) );
  NAND2_X1 U12443 ( .A1(n12803), .A2(n10059), .ZN(n9911) );
  OAI211_X1 U12444 ( .C1(n10135), .C2(n12806), .A(n12866), .B(n9911), .ZN(
        n9918) );
  INV_X1 U12445 ( .A(n9912), .ZN(n9916) );
  AOI22_X1 U12446 ( .A1(n12813), .A2(n12848), .B1(n14688), .B2(n9913), .ZN(
        n9915) );
  NOR3_X1 U12447 ( .A1(n9916), .A2(n9915), .A3(n9914), .ZN(n9917) );
  AOI211_X1 U12448 ( .C1(n10060), .C2(n14690), .A(n9918), .B(n9917), .ZN(n9919) );
  OAI21_X1 U12449 ( .B1(n10010), .B2(n12792), .A(n9919), .ZN(P2_U3199) );
  MUX2_X1 U12450 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12164), .Z(n10109) );
  XNOR2_X1 U12451 ( .A(n10109), .B(n10110), .ZN(n10107) );
  NAND2_X1 U12452 ( .A1(n9921), .A2(n9920), .ZN(n9925) );
  INV_X1 U12453 ( .A(n9922), .ZN(n9923) );
  NAND2_X1 U12454 ( .A1(n9923), .A2(n6555), .ZN(n9924) );
  NAND2_X1 U12455 ( .A1(n9925), .A2(n9924), .ZN(n10108) );
  XOR2_X1 U12456 ( .A(n10107), .B(n10108), .Z(n9942) );
  OR2_X1 U12457 ( .A1(n6555), .A2(n10726), .ZN(n9928) );
  XNOR2_X1 U12458 ( .A(n10117), .B(n10110), .ZN(n9929) );
  NAND2_X1 U12459 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n9929), .ZN(n10119) );
  OAI21_X1 U12460 ( .B1(n9929), .B2(P3_REG1_REG_7__SCAN_IN), .A(n10119), .ZN(
        n9930) );
  INV_X1 U12461 ( .A(n9930), .ZN(n9932) );
  AND2_X1 U12462 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n10734) );
  AOI21_X1 U12463 ( .B1(n14899), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10734), .ZN(
        n9931) );
  OAI21_X1 U12464 ( .B1(n14313), .B2(n9932), .A(n9931), .ZN(n9940) );
  INV_X1 U12465 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9936) );
  AOI21_X1 U12466 ( .B1(n9937), .B2(n9936), .A(n10114), .ZN(n9938) );
  NOR2_X1 U12467 ( .A1(n14912), .A2(n9938), .ZN(n9939) );
  AOI211_X1 U12468 ( .C1(n14906), .C2(n10110), .A(n9940), .B(n9939), .ZN(n9941) );
  OAI21_X1 U12469 ( .B1(n9942), .B2(n14882), .A(n9941), .ZN(P3_U3189) );
  XNOR2_X1 U12470 ( .A(n9944), .B(n9943), .ZN(n14798) );
  NAND3_X1 U12471 ( .A1(n9750), .A2(n9946), .A3(n9945), .ZN(n9947) );
  AOI21_X1 U12472 ( .B1(n9948), .B2(n9947), .A(n13189), .ZN(n9950) );
  NOR2_X1 U12473 ( .A1(n9950), .A2(n9949), .ZN(n14796) );
  MUX2_X1 U12474 ( .A(n9951), .B(n14796), .S(n6558), .Z(n9959) );
  INV_X1 U12475 ( .A(n9952), .ZN(n9954) );
  INV_X1 U12476 ( .A(n9953), .ZN(n10058) );
  AOI211_X1 U12477 ( .C1(n14794), .C2(n9954), .A(n13104), .B(n10058), .ZN(
        n14793) );
  OAI22_X1 U12478 ( .A1(n14739), .A2(n9956), .B1(n14751), .B2(n9955), .ZN(
        n9957) );
  AOI21_X1 U12479 ( .B1(n14793), .B2(n14731), .A(n9957), .ZN(n9958) );
  OAI211_X1 U12480 ( .C1(n13114), .C2(n14798), .A(n9959), .B(n9958), .ZN(
        P2_U3261) );
  INV_X1 U12481 ( .A(n9974), .ZN(n9960) );
  NAND2_X1 U12482 ( .A1(n9979), .A2(n9960), .ZN(n9966) );
  NAND3_X1 U12483 ( .A1(n9963), .A2(n9962), .A3(n9961), .ZN(n9964) );
  AOI21_X1 U12484 ( .B1(n9984), .B2(n9972), .A(n9964), .ZN(n9965) );
  NAND2_X1 U12485 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  NAND2_X1 U12486 ( .A1(n9967), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9971) );
  INV_X1 U12487 ( .A(n9988), .ZN(n9968) );
  NAND2_X1 U12488 ( .A1(n9982), .A2(n9968), .ZN(n11618) );
  INV_X1 U12489 ( .A(n11618), .ZN(n9969) );
  NAND2_X1 U12490 ( .A1(n9979), .A2(n9969), .ZN(n9970) );
  NOR2_X1 U12491 ( .A1(n12124), .A2(P3_U3151), .ZN(n10090) );
  INV_X1 U12492 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15223) );
  NAND2_X1 U12493 ( .A1(n9972), .A2(n14971), .ZN(n9973) );
  OAI22_X1 U12494 ( .A1(n9979), .A2(n9974), .B1(n9984), .B2(n9973), .ZN(n9975)
         );
  NAND2_X1 U12495 ( .A1(n8751), .A2(n10100), .ZN(n11429) );
  INV_X1 U12496 ( .A(n11429), .ZN(n9976) );
  NOR2_X1 U12497 ( .A1(n14930), .A2(n9976), .ZN(n11587) );
  INV_X1 U12498 ( .A(n11587), .ZN(n9986) );
  INV_X1 U12499 ( .A(n11580), .ZN(n9977) );
  NAND2_X1 U12500 ( .A1(n9982), .A2(n9977), .ZN(n9978) );
  OR2_X1 U12501 ( .A1(n9979), .A2(n9978), .ZN(n10049) );
  INV_X1 U12502 ( .A(n10049), .ZN(n9980) );
  NAND2_X1 U12503 ( .A1(n9982), .A2(n14966), .ZN(n9983) );
  NOR2_X1 U12504 ( .A1(n11613), .A2(n14971), .ZN(n9981) );
  OAI22_X1 U12505 ( .A1(n12120), .A2(n14922), .B1(n12121), .B2(n10100), .ZN(
        n9985) );
  AOI21_X1 U12506 ( .B1(n12058), .B2(n9986), .A(n9985), .ZN(n9987) );
  OAI21_X1 U12507 ( .B1(n10090), .B2(n15223), .A(n9987), .ZN(P3_U3172) );
  INV_X1 U12508 ( .A(n12544), .ZN(n12525) );
  NAND2_X1 U12509 ( .A1(n9988), .A2(n14971), .ZN(n9989) );
  OR2_X1 U12510 ( .A1(n11587), .A2(n9989), .ZN(n9991) );
  NAND2_X1 U12511 ( .A1(n12139), .A2(n12453), .ZN(n9990) );
  NAND2_X1 U12512 ( .A1(n9991), .A2(n9990), .ZN(n10471) );
  MUX2_X1 U12513 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n10471), .S(n14989), .Z(
        n9992) );
  AOI21_X1 U12514 ( .B1(n12525), .B2(n10474), .A(n9992), .ZN(n9993) );
  INV_X1 U12515 ( .A(n9993), .ZN(P3_U3459) );
  NAND3_X1 U12516 ( .A1(n14912), .A2(n14882), .A3(n14313), .ZN(n10003) );
  INV_X1 U12517 ( .A(n9994), .ZN(n9998) );
  AOI22_X1 U12518 ( .A1(n14899), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9997) );
  NAND2_X1 U12519 ( .A1(n14895), .A2(n9995), .ZN(n9996) );
  OAI211_X1 U12520 ( .C1(n14912), .C2(n9998), .A(n9997), .B(n9996), .ZN(n10002) );
  NOR2_X1 U12521 ( .A1(n14882), .A2(n9999), .ZN(n10000) );
  MUX2_X1 U12522 ( .A(n10000), .B(n14906), .S(P3_IR_REG_0__SCAN_IN), .Z(n10001) );
  AOI211_X1 U12523 ( .C1(n10004), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10005) );
  INV_X1 U12524 ( .A(n10005), .ZN(P3_U3182) );
  INV_X1 U12525 ( .A(n10219), .ZN(n10035) );
  INV_X1 U12526 ( .A(n10006), .ZN(n10008) );
  NAND2_X1 U12527 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  XNOR2_X1 U12528 ( .A(n10219), .B(n12663), .ZN(n10012) );
  AND2_X1 U12529 ( .A1(n12846), .A2(n12664), .ZN(n10013) );
  NAND2_X1 U12530 ( .A1(n10012), .A2(n10013), .ZN(n10187) );
  INV_X1 U12531 ( .A(n10012), .ZN(n10186) );
  INV_X1 U12532 ( .A(n10013), .ZN(n10014) );
  NAND2_X1 U12533 ( .A1(n10186), .A2(n10014), .ZN(n10015) );
  NAND2_X1 U12534 ( .A1(n10187), .A2(n10015), .ZN(n10016) );
  AOI21_X1 U12535 ( .B1(n10017), .B2(n10016), .A(n12792), .ZN(n10018) );
  NAND2_X1 U12536 ( .A1(n10018), .A2(n10188), .ZN(n10023) );
  NAND2_X1 U12537 ( .A1(n12847), .A2(n12800), .ZN(n10020) );
  NAND2_X1 U12538 ( .A1(n12845), .A2(n12801), .ZN(n10019) );
  NAND2_X1 U12539 ( .A1(n10020), .A2(n10019), .ZN(n10218) );
  NAND2_X1 U12540 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n12887) );
  OAI21_X1 U12541 ( .B1(n14694), .B2(n10030), .A(n12887), .ZN(n10021) );
  AOI21_X1 U12542 ( .B1(n14685), .B2(n10218), .A(n10021), .ZN(n10022) );
  OAI211_X1 U12543 ( .C1(n10035), .C2(n12821), .A(n10023), .B(n10022), .ZN(
        P2_U3211) );
  XNOR2_X1 U12544 ( .A(n10024), .B(n10026), .ZN(n10222) );
  INV_X1 U12545 ( .A(n13131), .ZN(n13058) );
  OAI21_X1 U12546 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(n10216) );
  INV_X1 U12547 ( .A(n13114), .ZN(n10037) );
  NAND2_X1 U12548 ( .A1(n10057), .A2(n10219), .ZN(n10028) );
  NAND2_X1 U12549 ( .A1(n10028), .A2(n10011), .ZN(n10029) );
  NOR2_X1 U12550 ( .A1(n10550), .A2(n10029), .ZN(n10217) );
  NAND2_X1 U12551 ( .A1(n10217), .A2(n14731), .ZN(n10034) );
  INV_X1 U12552 ( .A(n10030), .ZN(n10032) );
  MUX2_X1 U12553 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10218), .S(n6558), .Z(
        n10031) );
  AOI21_X1 U12554 ( .B1(n14734), .B2(n10032), .A(n10031), .ZN(n10033) );
  OAI211_X1 U12555 ( .C1(n10035), .C2(n14739), .A(n10034), .B(n10033), .ZN(
        n10036) );
  AOI21_X1 U12556 ( .B1(n10216), .B2(n10037), .A(n10036), .ZN(n10038) );
  OAI21_X1 U12557 ( .B1(n10222), .B2(n13058), .A(n10038), .ZN(P2_U3259) );
  INV_X1 U12558 ( .A(n10039), .ZN(n11616) );
  XNOR2_X1 U12559 ( .A(n10160), .B(n6553), .ZN(n10047) );
  XNOR2_X1 U12560 ( .A(n12139), .B(n6756), .ZN(n10041) );
  INV_X1 U12561 ( .A(n10086), .ZN(n14936) );
  AOI21_X1 U12562 ( .B1(n10042), .B2(n11968), .A(n14936), .ZN(n10043) );
  XNOR2_X1 U12563 ( .A(n11032), .B(n6756), .ZN(n10044) );
  NAND2_X1 U12564 ( .A1(n10044), .A2(n14922), .ZN(n10045) );
  NAND2_X1 U12565 ( .A1(n10084), .A2(n10045), .ZN(n10046) );
  OAI21_X1 U12566 ( .B1(n10047), .B2(n10046), .A(n10162), .ZN(n10048) );
  NAND2_X1 U12567 ( .A1(n10048), .A2(n12058), .ZN(n10053) );
  INV_X1 U12568 ( .A(n12120), .ZN(n12109) );
  OAI22_X1 U12569 ( .A1(n12112), .A2(n14922), .B1(n12121), .B2(n10050), .ZN(
        n10051) );
  AOI21_X1 U12570 ( .B1(n12109), .B2(n12138), .A(n10051), .ZN(n10052) );
  OAI211_X1 U12571 ( .C1(n10090), .C2(n14917), .A(n10053), .B(n10052), .ZN(
        P3_U3177) );
  XOR2_X1 U12572 ( .A(n10056), .B(n10054), .Z(n10141) );
  XOR2_X1 U12573 ( .A(n10056), .B(n10055), .Z(n10139) );
  OAI211_X1 U12574 ( .C1(n10058), .C2(n10137), .A(n10011), .B(n10057), .ZN(
        n10136) );
  AOI22_X1 U12575 ( .A1(n14393), .A2(n10060), .B1(n10059), .B2(n14734), .ZN(
        n10063) );
  MUX2_X1 U12576 ( .A(n10061), .B(n10135), .S(n6558), .Z(n10062) );
  OAI211_X1 U12577 ( .C1(n10136), .C2(n13129), .A(n10063), .B(n10062), .ZN(
        n10064) );
  AOI21_X1 U12578 ( .B1(n10139), .B2(n10037), .A(n10064), .ZN(n10065) );
  OAI21_X1 U12579 ( .B1(n10141), .B2(n13058), .A(n10065), .ZN(P2_U3260) );
  XNOR2_X1 U12580 ( .A(n10070), .B(n10066), .ZN(n14775) );
  INV_X1 U12581 ( .A(n14775), .ZN(n10079) );
  NAND2_X1 U12582 ( .A1(n6558), .A2(n6720), .ZN(n10826) );
  INV_X1 U12583 ( .A(n10067), .ZN(n10068) );
  AOI21_X1 U12584 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10073) );
  NAND2_X1 U12585 ( .A1(n14775), .A2(n14816), .ZN(n10071) );
  OAI211_X1 U12586 ( .C1(n10073), .C2(n13189), .A(n10072), .B(n10071), .ZN(
        n14773) );
  NAND2_X1 U12587 ( .A1(n14773), .A2(n6558), .ZN(n10078) );
  OAI22_X1 U12588 ( .A1(n6558), .A2(n12858), .B1(n12851), .B2(n14751), .ZN(
        n10076) );
  OAI211_X1 U12589 ( .C1(n14772), .C2(n14747), .A(n10011), .B(n10074), .ZN(
        n14771) );
  NOR2_X1 U12590 ( .A1(n13129), .A2(n14771), .ZN(n10075) );
  AOI211_X1 U12591 ( .C1(n14393), .C2(n8869), .A(n10076), .B(n10075), .ZN(
        n10077) );
  OAI211_X1 U12592 ( .C1(n10079), .C2(n10826), .A(n10078), .B(n10077), .ZN(
        P2_U3264) );
  INV_X1 U12593 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n14933) );
  INV_X1 U12594 ( .A(n8751), .ZN(n14940) );
  OAI22_X1 U12595 ( .A1(n12112), .A2(n14940), .B1(n6756), .B2(n12121), .ZN(
        n10080) );
  AOI21_X1 U12596 ( .B1(n12109), .B2(n6553), .A(n10080), .ZN(n10089) );
  INV_X1 U12597 ( .A(n14930), .ZN(n10082) );
  NAND3_X1 U12598 ( .A1(n10082), .A2(n11968), .A3(n14937), .ZN(n10083) );
  OAI211_X1 U12599 ( .C1(n10086), .C2(n10085), .A(n10084), .B(n10083), .ZN(
        n10087) );
  NAND2_X1 U12600 ( .A1(n10087), .A2(n12058), .ZN(n10088) );
  OAI211_X1 U12601 ( .C1(n10090), .C2(n14933), .A(n10089), .B(n10088), .ZN(
        P3_U3162) );
  INV_X1 U12602 ( .A(n11290), .ZN(n10102) );
  OR2_X1 U12603 ( .A1(n10092), .A2(n10091), .ZN(n10333) );
  NOR2_X1 U12604 ( .A1(n10333), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n10335) );
  OR2_X1 U12605 ( .A1(n10335), .A2(n9479), .ZN(n10093) );
  MUX2_X1 U12606 ( .A(n10093), .B(P1_IR_REG_31__SCAN_IN), .S(n10094), .Z(
        n10095) );
  NAND2_X1 U12607 ( .A1(n10335), .A2(n10094), .ZN(n10649) );
  AND2_X1 U12608 ( .A1(n10095), .A2(n10649), .ZN(n11291) );
  INV_X1 U12609 ( .A(n11291), .ZN(n11269) );
  OAI222_X1 U12610 ( .A1(n14145), .A2(n10096), .B1(n14148), .B2(n10102), .C1(
        n11269), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12611 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10097) );
  NOR2_X1 U12612 ( .A1(n14979), .A2(n10097), .ZN(n10098) );
  AOI21_X1 U12613 ( .B1(n14979), .B2(n10471), .A(n10098), .ZN(n10099) );
  OAI21_X1 U12614 ( .B1(n10100), .B2(n12597), .A(n10099), .ZN(P3_U3390) );
  INV_X1 U12615 ( .A(n11171), .ZN(n10105) );
  INV_X1 U12616 ( .A(n12938), .ZN(n11002) );
  OAI222_X1 U12617 ( .A1(n13272), .A2(n10105), .B1(n11002), .B2(P2_U3088), 
        .C1(n10101), .C2(n13269), .ZN(P2_U3313) );
  INV_X1 U12618 ( .A(n11133), .ZN(n11007) );
  OAI222_X1 U12619 ( .A1(n13269), .A2(n15273), .B1(n11007), .B2(P2_U3088), 
        .C1(n13272), .C2(n10102), .ZN(P2_U3311) );
  OAI21_X1 U12620 ( .B1(n10103), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10104) );
  XNOR2_X1 U12621 ( .A(n10104), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11172) );
  INV_X1 U12622 ( .A(n11172), .ZN(n10877) );
  OAI222_X1 U12623 ( .A1(n14145), .A2(n10106), .B1(n14148), .B2(n10105), .C1(
        n10877), .C2(P1_U3086), .ZN(P1_U3341) );
  MUX2_X1 U12624 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12164), .Z(n10304) );
  XNOR2_X1 U12625 ( .A(n10304), .B(n10309), .ZN(n10302) );
  NAND2_X1 U12626 ( .A1(n10108), .A2(n10107), .ZN(n10113) );
  INV_X1 U12627 ( .A(n10109), .ZN(n10111) );
  NAND2_X1 U12628 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  NAND2_X1 U12629 ( .A1(n10113), .A2(n10112), .ZN(n10303) );
  XOR2_X1 U12630 ( .A(n10302), .B(n10303), .Z(n10130) );
  INV_X1 U12631 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U12632 ( .A1(n10309), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n10116), 
        .B2(n10315), .ZN(n10312) );
  XNOR2_X1 U12633 ( .A(n10313), .B(n10312), .ZN(n10128) );
  INV_X1 U12634 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U12635 ( .A1(n10309), .A2(n14982), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n10315), .ZN(n10122) );
  NAND2_X1 U12636 ( .A1(n10118), .A2(n10117), .ZN(n10120) );
  NAND2_X1 U12637 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  NAND2_X1 U12638 ( .A1(n10122), .A2(n10121), .ZN(n10308) );
  OAI21_X1 U12639 ( .B1(n10122), .B2(n10121), .A(n10308), .ZN(n10123) );
  NAND2_X1 U12640 ( .A1(n10123), .A2(n14895), .ZN(n10126) );
  INV_X1 U12641 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U12642 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10124), .ZN(n12035) );
  AOI21_X1 U12643 ( .B1(n14899), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12035), .ZN(
        n10125) );
  OAI211_X1 U12644 ( .C1(n14357), .C2(n10315), .A(n10126), .B(n10125), .ZN(
        n10127) );
  AOI21_X1 U12645 ( .B1(n14843), .B2(n10128), .A(n10127), .ZN(n10129) );
  OAI21_X1 U12646 ( .B1(n10130), .B2(n14882), .A(n10129), .ZN(P3_U3190) );
  NAND2_X1 U12647 ( .A1(n10131), .A2(n14766), .ZN(n10132) );
  INV_X1 U12648 ( .A(n8861), .ZN(n14809) );
  OAI211_X1 U12649 ( .C1(n10137), .C2(n14819), .A(n10136), .B(n10135), .ZN(
        n10138) );
  AOI21_X1 U12650 ( .B1(n10139), .B2(n7116), .A(n10138), .ZN(n10140) );
  OAI21_X1 U12651 ( .B1(n10141), .B2(n13189), .A(n10140), .ZN(n10145) );
  NAND2_X1 U12652 ( .A1(n10145), .A2(n14833), .ZN(n10142) );
  OAI21_X1 U12653 ( .B1(n14833), .B2(n9336), .A(n10142), .ZN(P2_U3504) );
  INV_X1 U12654 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10147) );
  NAND2_X1 U12655 ( .A1(n10145), .A2(n14814), .ZN(n10146) );
  OAI21_X1 U12656 ( .B1(n14814), .B2(n10147), .A(n10146), .ZN(P2_U3445) );
  AOI21_X1 U12657 ( .B1(n10152), .B2(n15154), .A(n10148), .ZN(n10150) );
  MUX2_X1 U12658 ( .A(n11083), .B(P1_REG2_REG_13__SCAN_IN), .S(n11064), .Z(
        n10149) );
  NAND2_X1 U12659 ( .A1(n10149), .A2(n10150), .ZN(n10208) );
  OAI211_X1 U12660 ( .C1(n10150), .C2(n10149), .A(n13813), .B(n10208), .ZN(
        n10159) );
  NAND2_X1 U12661 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13370)
         );
  INV_X1 U12662 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U12663 ( .A(n10153), .B(P1_REG1_REG_13__SCAN_IN), .S(n11064), .Z(
        n10154) );
  NAND2_X1 U12664 ( .A1(n10155), .A2(n10154), .ZN(n10203) );
  OAI211_X1 U12665 ( .C1(n10155), .C2(n10154), .A(n10203), .B(n13819), .ZN(
        n10156) );
  NAND2_X1 U12666 ( .A1(n13370), .A2(n10156), .ZN(n10157) );
  AOI21_X1 U12667 ( .B1(n14525), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10157), 
        .ZN(n10158) );
  OAI211_X1 U12668 ( .C1(n6779), .C2(n11064), .A(n10159), .B(n10158), .ZN(
        P1_U3256) );
  INV_X1 U12669 ( .A(n6553), .ZN(n14942) );
  NAND2_X1 U12670 ( .A1(n10160), .A2(n14942), .ZN(n10161) );
  XNOR2_X1 U12671 ( .A(n11032), .B(n10298), .ZN(n10397) );
  XNOR2_X1 U12672 ( .A(n10397), .B(n12138), .ZN(n10163) );
  OAI211_X1 U12673 ( .C1(n10164), .C2(n10163), .A(n10400), .B(n12058), .ZN(
        n10168) );
  INV_X1 U12674 ( .A(n12137), .ZN(n10745) );
  OAI22_X1 U12675 ( .A1(n12112), .A2(n14942), .B1(n10745), .B2(n12120), .ZN(
        n10165) );
  AOI211_X1 U12676 ( .C1(n12469), .C2(n6545), .A(n10166), .B(n10165), .ZN(
        n10167) );
  OAI211_X1 U12677 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11042), .A(n10168), .B(
        n10167), .ZN(P3_U3158) );
  OR2_X1 U12678 ( .A1(n10169), .A2(n11595), .ZN(n10170) );
  NAND2_X1 U12679 ( .A1(n10171), .A2(n10170), .ZN(n12472) );
  INV_X1 U12680 ( .A(n12472), .ZN(n10177) );
  OAI211_X1 U12681 ( .C1(n10174), .C2(n10173), .A(n10172), .B(n12450), .ZN(
        n10176) );
  AOI22_X1 U12682 ( .A1(n12456), .A2(n6553), .B1(n12137), .B2(n12453), .ZN(
        n10175) );
  AND2_X1 U12683 ( .A1(n10176), .A2(n10175), .ZN(n12467) );
  OAI21_X1 U12684 ( .B1(n10177), .B2(n14973), .A(n12467), .ZN(n10300) );
  INV_X1 U12685 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10178) );
  OAI22_X1 U12686 ( .A1(n12544), .A2(n10298), .B1(n14989), .B2(n10178), .ZN(
        n10179) );
  AOI21_X1 U12687 ( .B1(n10300), .B2(n14989), .A(n10179), .ZN(n10180) );
  INV_X1 U12688 ( .A(n10180), .ZN(P3_U3462) );
  XNOR2_X1 U12689 ( .A(n10552), .B(n12663), .ZN(n10447) );
  AND2_X1 U12690 ( .A1(n12845), .A2(n12664), .ZN(n10181) );
  NAND2_X1 U12691 ( .A1(n10447), .A2(n10181), .ZN(n10416) );
  INV_X1 U12692 ( .A(n10447), .ZN(n10183) );
  INV_X1 U12693 ( .A(n10181), .ZN(n10182) );
  NAND2_X1 U12694 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  AND2_X1 U12695 ( .A1(n10416), .A2(n10184), .ZN(n10189) );
  INV_X1 U12696 ( .A(n10189), .ZN(n10185) );
  AOI21_X1 U12697 ( .B1(n10188), .B2(n10185), .A(n12792), .ZN(n10192) );
  NOR3_X1 U12698 ( .A1(n10186), .A2(n10193), .A3(n12794), .ZN(n10191) );
  OAI21_X1 U12699 ( .B1(n10192), .B2(n10191), .A(n10449), .ZN(n10196) );
  OAI22_X1 U12700 ( .A1(n10193), .A2(n14378), .B1(n10424), .B2(n14754), .ZN(
        n10548) );
  NAND2_X1 U12701 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n12905) );
  OAI21_X1 U12702 ( .B1(n14694), .B2(n14733), .A(n12905), .ZN(n10194) );
  AOI21_X1 U12703 ( .B1(n10548), .B2(n14685), .A(n10194), .ZN(n10195) );
  OAI211_X1 U12704 ( .C1(n14740), .C2(n12821), .A(n10196), .B(n10195), .ZN(
        P2_U3185) );
  INV_X1 U12705 ( .A(n11689), .ZN(n10227) );
  NAND2_X1 U12706 ( .A1(n10649), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10197) );
  XNOR2_X1 U12707 ( .A(n10197), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11690) );
  INV_X1 U12708 ( .A(n11690), .ZN(n11377) );
  OAI222_X1 U12709 ( .A1(n14145), .A2(n10198), .B1(n14148), .B2(n10227), .C1(
        n11377), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12710 ( .A(n10199), .ZN(n10200) );
  OAI222_X1 U12711 ( .A1(P3_U3151), .A2(n10202), .B1(n12606), .B2(n10201), 
        .C1(n12609), .C2(n10200), .ZN(P3_U3275) );
  INV_X1 U12712 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U12713 ( .A1(n11172), .A2(n14472), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10877), .ZN(n10205) );
  OAI21_X1 U12714 ( .B1(n11064), .B2(n10153), .A(n10203), .ZN(n10204) );
  NOR2_X1 U12715 ( .A1(n10205), .A2(n10204), .ZN(n10876) );
  AOI21_X1 U12716 ( .B1(n10205), .B2(n10204), .A(n10876), .ZN(n10215) );
  NAND2_X1 U12717 ( .A1(n14525), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U12718 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14435)
         );
  NAND2_X1 U12719 ( .A1(n10206), .A2(n14435), .ZN(n10207) );
  AOI21_X1 U12720 ( .B1(n11172), .B2(n13817), .A(n10207), .ZN(n10214) );
  INV_X1 U12721 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11083) );
  OAI21_X1 U12722 ( .B1(n11064), .B2(n11083), .A(n10208), .ZN(n10212) );
  INV_X1 U12723 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10209) );
  MUX2_X1 U12724 ( .A(n10209), .B(P1_REG2_REG_14__SCAN_IN), .S(n11172), .Z(
        n10210) );
  INV_X1 U12725 ( .A(n10210), .ZN(n10211) );
  NAND2_X1 U12726 ( .A1(n10211), .A2(n10212), .ZN(n10882) );
  OAI211_X1 U12727 ( .C1(n10212), .C2(n10211), .A(n13813), .B(n10882), .ZN(
        n10213) );
  OAI211_X1 U12728 ( .C1(n10215), .C2(n14536), .A(n10214), .B(n10213), .ZN(
        P1_U3257) );
  NAND2_X1 U12729 ( .A1(n10216), .A2(n7116), .ZN(n10221) );
  AOI211_X1 U12730 ( .C1(n14795), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        n10220) );
  OAI211_X1 U12731 ( .C1(n10222), .C2(n13189), .A(n10221), .B(n10220), .ZN(
        n10224) );
  NAND2_X1 U12732 ( .A1(n10224), .A2(n14814), .ZN(n10223) );
  OAI21_X1 U12733 ( .B1(n14814), .B2(n7774), .A(n10223), .ZN(P2_U3448) );
  NAND2_X1 U12734 ( .A1(n10224), .A2(n14833), .ZN(n10225) );
  OAI21_X1 U12735 ( .B1(n14833), .B2(n10226), .A(n10225), .ZN(P2_U3505) );
  INV_X1 U12736 ( .A(n11636), .ZN(n11011) );
  OAI222_X1 U12737 ( .A1(n13269), .A2(n10228), .B1(n11011), .B2(P2_U3088), 
        .C1(n13272), .C2(n10227), .ZN(P2_U3310) );
  INV_X1 U12738 ( .A(n10229), .ZN(n10230) );
  INV_X1 U12739 ( .A(n10251), .ZN(n10235) );
  INV_X1 U12740 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10233) );
  INV_X1 U12741 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U12742 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12743 ( .A1(n10235), .A2(n10234), .ZN(n10611) );
  NAND2_X1 U12744 ( .A1(n13694), .A2(n14590), .ZN(n13478) );
  NAND2_X1 U12745 ( .A1(n14564), .A2(n13479), .ZN(n10435) );
  AOI22_X1 U12746 ( .A1(n6551), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6562), .B2(
        n13720), .ZN(n10238) );
  NAND2_X1 U12747 ( .A1(n10348), .A2(n13693), .ZN(n13486) );
  NAND2_X1 U12748 ( .A1(n10435), .A2(n13486), .ZN(n10240) );
  NAND2_X1 U12749 ( .A1(n10271), .A2(n14596), .ZN(n13487) );
  NAND2_X1 U12750 ( .A1(n10240), .A2(n13487), .ZN(n10382) );
  NAND2_X1 U12751 ( .A1(n10241), .A2(n13444), .ZN(n10243) );
  AOI22_X1 U12752 ( .A1(n13455), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6562), 
        .B2(n13732), .ZN(n10242) );
  NAND2_X1 U12753 ( .A1(n13448), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10250) );
  INV_X1 U12754 ( .A(n10245), .ZN(n11738) );
  OR2_X1 U12755 ( .A1(n11738), .A2(n15086), .ZN(n10249) );
  OR2_X1 U12756 ( .A1(n11769), .A2(n10611), .ZN(n10248) );
  INV_X1 U12757 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10246) );
  OR2_X1 U12758 ( .A1(n11750), .A2(n10246), .ZN(n10247) );
  XNOR2_X1 U12759 ( .A(n10382), .B(n13419), .ZN(n10259) );
  NAND2_X1 U12760 ( .A1(n13693), .A2(n13662), .ZN(n10258) );
  NAND2_X1 U12761 ( .A1(n10245), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U12762 ( .A1(n10251), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10516) );
  OAI21_X1 U12763 ( .B1(n10251), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10516), .ZN(
        n10392) );
  OR2_X1 U12764 ( .A1(n11769), .A2(n10392), .ZN(n10255) );
  NAND2_X1 U12765 ( .A1(n13448), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U12766 ( .A1(n11778), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U12767 ( .A1(n13691), .A2(n13398), .ZN(n10257) );
  NAND2_X1 U12768 ( .A1(n10258), .A2(n10257), .ZN(n10609) );
  AOI21_X1 U12769 ( .B1(n10259), .B2(n14571), .A(n10609), .ZN(n14609) );
  NAND2_X1 U12770 ( .A1(n14579), .A2(n14590), .ZN(n14578) );
  NAND2_X1 U12771 ( .A1(n10431), .A2(n13491), .ZN(n10260) );
  NAND2_X1 U12772 ( .A1(n10260), .A2(n14577), .ZN(n10261) );
  NOR2_X1 U12773 ( .A1(n10388), .A2(n10261), .ZN(n14605) );
  NAND2_X1 U12774 ( .A1(n14605), .A2(n13965), .ZN(n10262) );
  OAI211_X1 U12775 ( .C1(n14010), .C2(n10611), .A(n14609), .B(n10262), .ZN(
        n10264) );
  NAND2_X1 U12776 ( .A1(n11784), .A2(n11783), .ZN(n10263) );
  MUX2_X1 U12777 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10264), .S(n14002), .Z(
        n10277) );
  INV_X1 U12778 ( .A(n10265), .ZN(n10266) );
  NOR2_X1 U12779 ( .A1(n13696), .A2(n13473), .ZN(n13472) );
  INV_X1 U12780 ( .A(n13472), .ZN(n10267) );
  INV_X1 U12781 ( .A(n14566), .ZN(n13415) );
  NAND2_X1 U12782 ( .A1(n14567), .A2(n13415), .ZN(n10270) );
  OR2_X1 U12783 ( .A1(n13694), .A2(n14573), .ZN(n10269) );
  NAND2_X1 U12784 ( .A1(n13487), .A2(n13486), .ZN(n13482) );
  NAND2_X1 U12785 ( .A1(n10271), .A2(n10348), .ZN(n10272) );
  XNOR2_X1 U12786 ( .A(n10379), .B(n13419), .ZN(n14606) );
  NAND2_X1 U12787 ( .A1(n13464), .A2(n10274), .ZN(n13644) );
  INV_X1 U12788 ( .A(n13644), .ZN(n13660) );
  NAND2_X1 U12789 ( .A1(n13660), .A2(n9433), .ZN(n10275) );
  OAI22_X1 U12790 ( .A1(n14606), .A2(n14020), .B1(n14603), .B2(n14012), .ZN(
        n10276) );
  OR2_X1 U12791 ( .A1(n10277), .A2(n10276), .ZN(P1_U3289) );
  OAI21_X1 U12792 ( .B1(n10279), .B2(n11447), .A(n10278), .ZN(n10280) );
  INV_X1 U12793 ( .A(n10280), .ZN(n10325) );
  INV_X1 U12794 ( .A(n10281), .ZN(n10284) );
  OAI22_X1 U12795 ( .A1(n10284), .A2(n10283), .B1(n10040), .B2(n10282), .ZN(
        n10286) );
  OR2_X1 U12796 ( .A1(n11613), .A2(n11433), .ZN(n12265) );
  NAND2_X1 U12797 ( .A1(n14920), .A2(n12265), .ZN(n14945) );
  OAI211_X1 U12798 ( .C1(n10288), .C2(n11590), .A(n10287), .B(n12450), .ZN(
        n10290) );
  AOI22_X1 U12799 ( .A1(n12453), .A2(n10720), .B1(n12138), .B2(n12456), .ZN(
        n10289) );
  AND2_X1 U12800 ( .A1(n10290), .A2(n10289), .ZN(n10324) );
  MUX2_X1 U12801 ( .A(n15258), .B(n10324), .S(n14946), .Z(n10293) );
  INV_X1 U12802 ( .A(n11613), .ZN(n14935) );
  NOR2_X1 U12803 ( .A1(n10291), .A2(n14935), .ZN(n12461) );
  AOI22_X1 U12804 ( .A1(n12470), .A2(n10410), .B1(n12468), .B2(n10396), .ZN(
        n10292) );
  OAI211_X1 U12805 ( .C1(n10325), .C2(n12431), .A(n10293), .B(n10292), .ZN(
        P3_U3229) );
  INV_X1 U12806 ( .A(n10294), .ZN(n10296) );
  OAI222_X1 U12807 ( .A1(n12609), .A2(n10296), .B1(n12606), .B2(n10295), .C1(
        P3_U3151), .C2(n11433), .ZN(P3_U3274) );
  INV_X1 U12808 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10297) );
  OAI22_X1 U12809 ( .A1(n12597), .A2(n10298), .B1(n14979), .B2(n10297), .ZN(
        n10299) );
  AOI21_X1 U12810 ( .B1(n10300), .B2(n14979), .A(n10299), .ZN(n10301) );
  INV_X1 U12811 ( .A(n10301), .ZN(P3_U3399) );
  MUX2_X1 U12812 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12164), .Z(n10478) );
  XNOR2_X1 U12813 ( .A(n10478), .B(n10483), .ZN(n10476) );
  NAND2_X1 U12814 ( .A1(n10303), .A2(n10302), .ZN(n10307) );
  INV_X1 U12815 ( .A(n10304), .ZN(n10305) );
  NAND2_X1 U12816 ( .A1(n10305), .A2(n10309), .ZN(n10306) );
  NAND2_X1 U12817 ( .A1(n10307), .A2(n10306), .ZN(n10477) );
  XOR2_X1 U12818 ( .A(n10476), .B(n10477), .Z(n10323) );
  OAI21_X1 U12819 ( .B1(n10309), .B2(n14982), .A(n10308), .ZN(n10486) );
  OAI21_X1 U12820 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n10310), .A(n10488), .ZN(
        n10321) );
  AND2_X1 U12821 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n10791) );
  AOI21_X1 U12822 ( .B1(n14899), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10791), .ZN(
        n10311) );
  OAI21_X1 U12823 ( .B1(n14357), .B2(n10487), .A(n10311), .ZN(n10320) );
  NOR2_X1 U12824 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  XNOR2_X1 U12825 ( .A(n10483), .B(n10482), .ZN(n10317) );
  INV_X1 U12826 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10316) );
  AOI21_X1 U12827 ( .B1(n10317), .B2(n10316), .A(n10484), .ZN(n10318) );
  NOR2_X1 U12828 ( .A1(n10318), .A2(n14912), .ZN(n10319) );
  AOI211_X1 U12829 ( .C1(n14895), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10322) );
  OAI21_X1 U12830 ( .B1(n10323), .B2(n14882), .A(n10322), .ZN(P3_U3191) );
  OAI21_X1 U12831 ( .B1(n10325), .B2(n14973), .A(n10324), .ZN(n10331) );
  INV_X1 U12832 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10326) );
  OAI22_X1 U12833 ( .A1(n12597), .A2(n10401), .B1(n14979), .B2(n10326), .ZN(
        n10327) );
  AOI21_X1 U12834 ( .B1(n10331), .B2(n14979), .A(n10327), .ZN(n10328) );
  INV_X1 U12835 ( .A(n10328), .ZN(P3_U3402) );
  OAI22_X1 U12836 ( .A1(n12544), .A2(n10401), .B1(n14989), .B2(n10329), .ZN(
        n10330) );
  AOI21_X1 U12837 ( .B1(n10331), .B2(n14989), .A(n10330), .ZN(n10332) );
  INV_X1 U12838 ( .A(n10332), .ZN(P3_U3463) );
  INV_X1 U12839 ( .A(n11243), .ZN(n10414) );
  NAND2_X1 U12840 ( .A1(n10333), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10334) );
  MUX2_X1 U12841 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10334), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n10337) );
  INV_X1 U12842 ( .A(n10335), .ZN(n10336) );
  AND2_X1 U12843 ( .A1(n10337), .A2(n10336), .ZN(n11244) );
  INV_X1 U12844 ( .A(n11244), .ZN(n14537) );
  OAI222_X1 U12845 ( .A1(n14145), .A2(n10338), .B1(n14148), .B2(n10414), .C1(
        n14537), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U12846 ( .A(n13490), .ZN(n13692) );
  AOI22_X1 U12847 ( .A1(n11821), .A2(n13491), .B1(n11931), .B2(n13692), .ZN(
        n10339) );
  XNOR2_X1 U12848 ( .A(n10339), .B(n11941), .ZN(n10613) );
  INV_X1 U12849 ( .A(n10340), .ZN(n10341) );
  NAND2_X1 U12850 ( .A1(n11821), .A2(n14596), .ZN(n10346) );
  NAND2_X1 U12851 ( .A1(n6559), .A2(n13693), .ZN(n10345) );
  NAND2_X1 U12852 ( .A1(n10346), .A2(n10345), .ZN(n10347) );
  XNOR2_X1 U12853 ( .A(n10347), .B(n11910), .ZN(n10351) );
  NOR2_X1 U12854 ( .A1(n11884), .A2(n10348), .ZN(n10349) );
  AOI21_X1 U12855 ( .B1(n6565), .B2(n13693), .A(n10349), .ZN(n10350) );
  NOR2_X1 U12856 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  AOI21_X1 U12857 ( .B1(n10351), .B2(n10350), .A(n10352), .ZN(n13293) );
  INV_X1 U12858 ( .A(n10352), .ZN(n10353) );
  OAI22_X1 U12859 ( .A1(n13490), .A2(n9739), .B1(n14603), .B2(n11884), .ZN(
        n10354) );
  OR2_X1 U12860 ( .A1(n10356), .A2(n13453), .ZN(n10358) );
  AOI22_X1 U12861 ( .A1(n13455), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6562), 
        .B2(n13750), .ZN(n10357) );
  NAND2_X1 U12862 ( .A1(n10358), .A2(n10357), .ZN(n13497) );
  AOI22_X1 U12863 ( .A1(n13497), .A2(n11930), .B1(n11931), .B2(n13691), .ZN(
        n10359) );
  XOR2_X1 U12864 ( .A(n11941), .B(n10359), .Z(n10560) );
  AOI22_X1 U12865 ( .A1(n11931), .A2(n13497), .B1(n6565), .B2(n13691), .ZN(
        n10558) );
  INV_X1 U12866 ( .A(n10558), .ZN(n10559) );
  XNOR2_X1 U12867 ( .A(n10560), .B(n10559), .ZN(n10360) );
  XNOR2_X1 U12868 ( .A(n10562), .B(n10360), .ZN(n10376) );
  AND2_X1 U12869 ( .A1(n10362), .A2(n10361), .ZN(n10363) );
  AND2_X1 U12870 ( .A1(n10364), .A2(n10363), .ZN(n13663) );
  NAND2_X1 U12871 ( .A1(n10365), .A2(n13663), .ZN(n10366) );
  NAND2_X1 U12872 ( .A1(n13448), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10371) );
  INV_X1 U12873 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10367) );
  XNOR2_X1 U12874 ( .A(n10516), .B(n10367), .ZN(n14552) );
  OR2_X1 U12875 ( .A1(n11769), .A2(n14552), .ZN(n10370) );
  NAND2_X1 U12876 ( .A1(n10245), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U12877 ( .A1(n11778), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U12878 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n13690) );
  NAND2_X1 U12879 ( .A1(n13690), .A2(n13398), .ZN(n10372) );
  OAI21_X1 U12880 ( .B1(n13490), .B2(n13387), .A(n10372), .ZN(n14611) );
  AOI22_X1 U12881 ( .A1(n14433), .A2(n14611), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10374) );
  AND2_X1 U12882 ( .A1(n13497), .A2(n14636), .ZN(n14613) );
  NAND2_X1 U12883 ( .A1(n14451), .A2(n14613), .ZN(n10373) );
  OAI211_X1 U12884 ( .C1(n14463), .C2(n10392), .A(n10374), .B(n10373), .ZN(
        n10375) );
  AOI21_X1 U12885 ( .B1(n10376), .B2(n14440), .A(n10375), .ZN(n10377) );
  INV_X1 U12886 ( .A(n10377), .ZN(P1_U3227) );
  INV_X1 U12887 ( .A(n13419), .ZN(n10378) );
  NAND2_X1 U12888 ( .A1(n14603), .A2(n13490), .ZN(n10380) );
  NAND2_X1 U12889 ( .A1(n10381), .A2(n10380), .ZN(n10500) );
  INV_X1 U12890 ( .A(n13691), .ZN(n10523) );
  XNOR2_X1 U12891 ( .A(n13497), .B(n10523), .ZN(n13422) );
  XOR2_X1 U12892 ( .A(n10500), .B(n13422), .Z(n14610) );
  NAND2_X1 U12893 ( .A1(n10382), .A2(n13419), .ZN(n10384) );
  NAND2_X1 U12894 ( .A1(n13491), .A2(n13490), .ZN(n10383) );
  XNOR2_X1 U12895 ( .A(n10522), .B(n13422), .ZN(n10385) );
  NOR2_X1 U12896 ( .A1(n10385), .A2(n14550), .ZN(n14614) );
  NOR2_X1 U12897 ( .A1(n14614), .A2(n14611), .ZN(n10386) );
  MUX2_X1 U12898 ( .A(n10387), .B(n10386), .S(n14002), .Z(n10395) );
  INV_X1 U12899 ( .A(n10388), .ZN(n10389) );
  INV_X1 U12900 ( .A(n13497), .ZN(n10524) );
  AOI211_X1 U12901 ( .C1(n13497), .C2(n10389), .A(n6570), .B(n14554), .ZN(
        n14612) );
  NOR2_X1 U12902 ( .A1(n10390), .A2(n13952), .ZN(n10391) );
  OAI22_X1 U12903 ( .A1(n14012), .A2(n10524), .B1(n14010), .B2(n10392), .ZN(
        n10393) );
  AOI21_X1 U12904 ( .B1(n14612), .B2(n14581), .A(n10393), .ZN(n10394) );
  OAI211_X1 U12905 ( .C1(n14020), .C2(n14610), .A(n10395), .B(n10394), .ZN(
        P1_U3288) );
  INV_X1 U12906 ( .A(n10396), .ZN(n10413) );
  INV_X1 U12907 ( .A(n10397), .ZN(n10398) );
  NAND2_X1 U12908 ( .A1(n10398), .A2(n12138), .ZN(n10399) );
  XNOR2_X1 U12909 ( .A(n11032), .B(n10401), .ZN(n10402) );
  NAND2_X1 U12910 ( .A1(n10402), .A2(n10745), .ZN(n10598) );
  INV_X1 U12911 ( .A(n10402), .ZN(n10403) );
  NAND2_X1 U12912 ( .A1(n10403), .A2(n12137), .ZN(n10404) );
  AND2_X1 U12913 ( .A1(n10598), .A2(n10404), .ZN(n10405) );
  OAI21_X1 U12914 ( .B1(n10406), .B2(n10405), .A(n10599), .ZN(n10407) );
  NAND2_X1 U12915 ( .A1(n10407), .A2(n12058), .ZN(n10412) );
  INV_X1 U12916 ( .A(n12138), .ZN(n14921) );
  OAI22_X1 U12917 ( .A1(n12112), .A2(n14921), .B1(n10660), .B2(n12120), .ZN(
        n10408) );
  AOI211_X1 U12918 ( .C1(n10410), .C2(n6545), .A(n10409), .B(n10408), .ZN(
        n10411) );
  OAI211_X1 U12919 ( .C1(n10413), .C2(n11042), .A(n10412), .B(n10411), .ZN(
        P3_U3170) );
  INV_X1 U12920 ( .A(n14719), .ZN(n11006) );
  OAI222_X1 U12921 ( .A1(n13269), .A2(n10415), .B1(n11006), .B2(P2_U3088), 
        .C1(n13272), .C2(n10414), .ZN(P2_U3312) );
  XNOR2_X1 U12922 ( .A(n10680), .B(n6554), .ZN(n10418) );
  NAND2_X1 U12923 ( .A1(n12844), .A2(n12664), .ZN(n10419) );
  XNOR2_X1 U12924 ( .A(n10418), .B(n10419), .ZN(n10457) );
  INV_X1 U12925 ( .A(n10418), .ZN(n10425) );
  NAND2_X1 U12926 ( .A1(n10425), .A2(n10419), .ZN(n10420) );
  XNOR2_X1 U12927 ( .A(n6569), .B(n6554), .ZN(n10752) );
  NAND2_X1 U12928 ( .A1(n12843), .A2(n12619), .ZN(n10753) );
  XNOR2_X1 U12929 ( .A(n10752), .B(n10753), .ZN(n10423) );
  AOI22_X1 U12930 ( .A1(n12800), .A2(n12844), .B1(n12842), .B2(n12801), .ZN(
        n10816) );
  NOR2_X1 U12931 ( .A1(n10816), .A2(n12806), .ZN(n10422) );
  NAND2_X1 U12932 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14704) );
  OAI21_X1 U12933 ( .B1(n14694), .B2(n10820), .A(n14704), .ZN(n10421) );
  AOI211_X1 U12934 ( .C1(n6569), .C2(n14690), .A(n10422), .B(n10421), .ZN(
        n10429) );
  INV_X1 U12935 ( .A(n10423), .ZN(n10427) );
  OAI22_X1 U12936 ( .A1(n10425), .A2(n12792), .B1(n10424), .B2(n12794), .ZN(
        n10426) );
  NAND3_X1 U12937 ( .A1(n10448), .A2(n10427), .A3(n10426), .ZN(n10428) );
  OAI211_X1 U12938 ( .C1(n10755), .C2(n12792), .A(n10429), .B(n10428), .ZN(
        P2_U3203) );
  INV_X1 U12939 ( .A(n13482), .ZN(n13418) );
  XNOR2_X1 U12940 ( .A(n10430), .B(n13418), .ZN(n14599) );
  INV_X1 U12941 ( .A(n10431), .ZN(n10432) );
  AOI211_X1 U12942 ( .C1(n14596), .C2(n14578), .A(n6570), .B(n10432), .ZN(
        n14595) );
  INV_X1 U12943 ( .A(n14595), .ZN(n10433) );
  OAI22_X1 U12944 ( .A1(n10433), .A2(n14016), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14010), .ZN(n10434) );
  AOI21_X1 U12945 ( .B1(n14572), .B2(n14596), .A(n10434), .ZN(n10439) );
  XNOR2_X1 U12946 ( .A(n10435), .B(n13418), .ZN(n10437) );
  OAI22_X1 U12947 ( .A1(n10436), .A2(n13387), .B1(n13490), .B2(n13388), .ZN(
        n13295) );
  AOI21_X1 U12948 ( .B1(n10437), .B2(n14571), .A(n13295), .ZN(n14597) );
  MUX2_X1 U12949 ( .A(n14597), .B(n15054), .S(n14276), .Z(n10438) );
  OAI211_X1 U12950 ( .C1(n14020), .C2(n14599), .A(n10439), .B(n10438), .ZN(
        P1_U3290) );
  INV_X1 U12951 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10440) );
  OAI22_X1 U12952 ( .A1(n14575), .A2(n10441), .B1(n10440), .B2(n14010), .ZN(
        n10444) );
  NOR2_X1 U12953 ( .A1(n14016), .A2(n6570), .ZN(n13825) );
  INV_X1 U12954 ( .A(n13825), .ZN(n11096) );
  AOI21_X1 U12955 ( .B1(n11096), .B2(n14012), .A(n10442), .ZN(n10443) );
  AOI211_X1 U12956 ( .C1(n14276), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10444), .B(
        n10443), .ZN(n10446) );
  NAND2_X1 U12957 ( .A1(n14002), .A2(n14571), .ZN(n13924) );
  INV_X1 U12958 ( .A(n13924), .ZN(n14018) );
  INV_X1 U12959 ( .A(n14020), .ZN(n13922) );
  OAI21_X1 U12960 ( .B1(n14018), .B2(n13922), .A(n13416), .ZN(n10445) );
  NAND2_X1 U12961 ( .A1(n10446), .A2(n10445), .ZN(P1_U3293) );
  NAND3_X1 U12962 ( .A1(n10447), .A2(n12813), .A3(n12845), .ZN(n10456) );
  OAI21_X1 U12963 ( .B1(n10457), .B2(n10449), .A(n10448), .ZN(n10450) );
  NAND2_X1 U12964 ( .A1(n10450), .A2(n14688), .ZN(n10455) );
  OAI21_X1 U12965 ( .B1(n14694), .B2(n10677), .A(n10451), .ZN(n10453) );
  AOI22_X1 U12966 ( .A1(n12800), .A2(n12845), .B1(n12843), .B2(n12801), .ZN(
        n10670) );
  NOR2_X1 U12967 ( .A1(n10670), .A2(n12806), .ZN(n10452) );
  AOI211_X1 U12968 ( .C1(n10680), .C2(n14690), .A(n10453), .B(n10452), .ZN(
        n10454) );
  OAI211_X1 U12969 ( .C1(n10457), .C2(n10456), .A(n10455), .B(n10454), .ZN(
        P2_U3193) );
  INV_X1 U12970 ( .A(n14010), .ZN(n14574) );
  AOI22_X1 U12971 ( .A1(n14581), .A2(n10458), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14574), .ZN(n10459) );
  OAI21_X1 U12972 ( .B1(n14002), .B2(n9237), .A(n10459), .ZN(n10463) );
  NOR3_X1 U12973 ( .A1(n13924), .A2(n10461), .A3(n10460), .ZN(n10462) );
  AOI211_X1 U12974 ( .C1(n14572), .C2(n13473), .A(n10463), .B(n10462), .ZN(
        n10466) );
  NAND2_X1 U12975 ( .A1(n10464), .A2(n14002), .ZN(n10465) );
  OAI211_X1 U12976 ( .C1(n14020), .C2(n10467), .A(n10466), .B(n10465), .ZN(
        P1_U3292) );
  INV_X1 U12977 ( .A(n10468), .ZN(n10470) );
  OAI22_X1 U12978 ( .A1(n11619), .A2(P3_U3151), .B1(SI_22_), .B2(n12606), .ZN(
        n10469) );
  AOI21_X1 U12979 ( .B1(n10470), .B2(n12602), .A(n10469), .ZN(P3_U3273) );
  NOR2_X1 U12980 ( .A1(n14934), .A2(n15223), .ZN(n10473) );
  INV_X2 U12981 ( .A(n14946), .ZN(n14949) );
  MUX2_X1 U12982 ( .A(n10471), .B(P3_REG2_REG_0__SCAN_IN), .S(n14949), .Z(
        n10472) );
  AOI211_X1 U12983 ( .C1(n12470), .C2(n10474), .A(n10473), .B(n10472), .ZN(
        n10475) );
  INV_X1 U12984 ( .A(n10475), .ZN(P3_U3233) );
  MUX2_X1 U12985 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12164), .Z(n12143) );
  XNOR2_X1 U12986 ( .A(n12143), .B(n12144), .ZN(n12141) );
  NAND2_X1 U12987 ( .A1(n10477), .A2(n10476), .ZN(n10481) );
  INV_X1 U12988 ( .A(n10478), .ZN(n10479) );
  NAND2_X1 U12989 ( .A1(n10479), .A2(n10483), .ZN(n10480) );
  NAND2_X1 U12990 ( .A1(n10481), .A2(n10480), .ZN(n12142) );
  XOR2_X1 U12991 ( .A(n12141), .B(n12142), .Z(n10499) );
  NAND2_X1 U12992 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n12194), .ZN(n10485) );
  OAI21_X1 U12993 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12194), .A(n10485), 
        .ZN(n12174) );
  XNOR2_X1 U12994 ( .A(n12175), .B(n12174), .ZN(n10497) );
  INV_X1 U12995 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U12996 ( .A1(n12144), .A2(n14987), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n12194), .ZN(n10491) );
  NAND2_X1 U12997 ( .A1(n10487), .A2(n10486), .ZN(n10489) );
  NAND2_X1 U12998 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  OAI21_X1 U12999 ( .B1(n10491), .B2(n10490), .A(n12195), .ZN(n10492) );
  NAND2_X1 U13000 ( .A1(n10492), .A2(n14895), .ZN(n10495) );
  INV_X1 U13001 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n10493) );
  NOR2_X1 U13002 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10493), .ZN(n11039) );
  AOI21_X1 U13003 ( .B1(n14899), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11039), 
        .ZN(n10494) );
  OAI211_X1 U13004 ( .C1(n14357), .C2(n12194), .A(n10495), .B(n10494), .ZN(
        n10496) );
  AOI21_X1 U13005 ( .B1(n14843), .B2(n10497), .A(n10496), .ZN(n10498) );
  OAI21_X1 U13006 ( .B1(n10499), .B2(n14882), .A(n10498), .ZN(P3_U3192) );
  NAND2_X1 U13007 ( .A1(n10500), .A2(n13422), .ZN(n10502) );
  NAND2_X1 U13008 ( .A1(n10524), .A2(n10523), .ZN(n10501) );
  NAND2_X1 U13009 ( .A1(n10502), .A2(n10501), .ZN(n14543) );
  OR2_X1 U13010 ( .A1(n10503), .A2(n13453), .ZN(n10507) );
  INV_X1 U13011 ( .A(n10504), .ZN(n10505) );
  AOI22_X1 U13012 ( .A1(n13455), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6562), 
        .B2(n10505), .ZN(n10506) );
  NAND2_X1 U13013 ( .A1(n10507), .A2(n10506), .ZN(n14559) );
  INV_X1 U13014 ( .A(n13690), .ZN(n10566) );
  NAND2_X1 U13015 ( .A1(n14559), .A2(n10566), .ZN(n10526) );
  OR2_X1 U13016 ( .A1(n14559), .A2(n10566), .ZN(n10508) );
  NAND2_X1 U13017 ( .A1(n10526), .A2(n10508), .ZN(n14547) );
  NAND2_X1 U13018 ( .A1(n14543), .A2(n14547), .ZN(n10510) );
  OR2_X1 U13019 ( .A1(n14559), .A2(n13690), .ZN(n10509) );
  OR2_X1 U13020 ( .A1(n10511), .A2(n13453), .ZN(n10513) );
  AOI22_X1 U13021 ( .A1(n13455), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6562), 
        .B2(n13775), .ZN(n10512) );
  NAND2_X1 U13022 ( .A1(n10513), .A2(n10512), .ZN(n13506) );
  NAND2_X1 U13023 ( .A1(n13448), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10521) );
  INV_X1 U13024 ( .A(n10516), .ZN(n10514) );
  AOI21_X1 U13025 ( .B1(n10514), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U13026 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n10515) );
  OR2_X1 U13027 ( .A1(n10517), .A2(n10528), .ZN(n10591) );
  OR2_X1 U13028 ( .A1(n11769), .A2(n10591), .ZN(n10520) );
  NAND2_X1 U13029 ( .A1(n10245), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10519) );
  NAND2_X1 U13030 ( .A1(n11778), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13031 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n13689) );
  XNOR2_X1 U13032 ( .A(n13506), .B(n13689), .ZN(n13423) );
  XNOR2_X1 U13033 ( .A(n10620), .B(n13423), .ZN(n14627) );
  NAND2_X1 U13034 ( .A1(n10524), .A2(n13691), .ZN(n10525) );
  NAND2_X1 U13035 ( .A1(n14544), .A2(n10526), .ZN(n10527) );
  OAI21_X1 U13036 ( .B1(n10527), .B2(n13423), .A(n10632), .ZN(n10536) );
  NAND2_X1 U13037 ( .A1(n13690), .A2(n13662), .ZN(n10535) );
  NAND2_X1 U13038 ( .A1(n10245), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13039 ( .A1(n10528), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10634) );
  OR2_X1 U13040 ( .A1(n10528), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U13041 ( .A1(n10634), .A2(n10529), .ZN(n10806) );
  OR2_X1 U13042 ( .A1(n11769), .A2(n10806), .ZN(n10532) );
  NAND2_X1 U13043 ( .A1(n11778), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10531) );
  NAND2_X1 U13044 ( .A1(n13448), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13045 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n13688) );
  NAND2_X1 U13046 ( .A1(n13688), .A2(n13398), .ZN(n10534) );
  NAND2_X1 U13047 ( .A1(n10535), .A2(n10534), .ZN(n10589) );
  AOI21_X1 U13048 ( .B1(n10536), .B2(n14571), .A(n10589), .ZN(n14626) );
  MUX2_X1 U13049 ( .A(n14626), .B(n10537), .S(n14276), .Z(n10542) );
  INV_X1 U13050 ( .A(n14559), .ZN(n10538) );
  INV_X1 U13051 ( .A(n10645), .ZN(n10539) );
  AOI211_X1 U13052 ( .C1(n13506), .C2(n14555), .A(n6570), .B(n10539), .ZN(
        n14624) );
  INV_X1 U13053 ( .A(n13506), .ZN(n10588) );
  OAI22_X1 U13054 ( .A1(n14012), .A2(n10588), .B1(n14010), .B2(n10591), .ZN(
        n10540) );
  AOI21_X1 U13055 ( .B1(n14624), .B2(n14581), .A(n10540), .ZN(n10541) );
  OAI211_X1 U13056 ( .C1(n14020), .C2(n14627), .A(n10542), .B(n10541), .ZN(
        P1_U3286) );
  OAI21_X1 U13057 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(n14742) );
  INV_X1 U13058 ( .A(n14742), .ZN(n10554) );
  XNOR2_X1 U13059 ( .A(n10547), .B(n10546), .ZN(n10549) );
  AOI21_X1 U13060 ( .B1(n10549), .B2(n14753), .A(n10548), .ZN(n14744) );
  INV_X1 U13061 ( .A(n10550), .ZN(n10551) );
  AOI211_X1 U13062 ( .C1(n10552), .C2(n10551), .A(n13104), .B(n10676), .ZN(
        n14732) );
  AOI21_X1 U13063 ( .B1(n14795), .B2(n10552), .A(n14732), .ZN(n10553) );
  OAI211_X1 U13064 ( .C1(n10554), .C2(n14799), .A(n14744), .B(n10553), .ZN(
        n10556) );
  NAND2_X1 U13065 ( .A1(n10556), .A2(n14833), .ZN(n10555) );
  OAI21_X1 U13066 ( .B1(n14833), .B2(n9338), .A(n10555), .ZN(P2_U3506) );
  NAND2_X1 U13067 ( .A1(n10556), .A2(n14814), .ZN(n10557) );
  OAI21_X1 U13068 ( .B1(n14814), .B2(n7793), .A(n10557), .ZN(P2_U3451) );
  NAND2_X1 U13069 ( .A1(n6752), .A2(n10558), .ZN(n10561) );
  NAND2_X1 U13070 ( .A1(n14559), .A2(n11930), .ZN(n10564) );
  NAND2_X1 U13071 ( .A1(n11931), .A2(n13690), .ZN(n10563) );
  NAND2_X1 U13072 ( .A1(n10564), .A2(n10563), .ZN(n10565) );
  XNOR2_X1 U13073 ( .A(n10565), .B(n11910), .ZN(n10571) );
  INV_X1 U13074 ( .A(n10571), .ZN(n10569) );
  NOR2_X1 U13075 ( .A1(n9739), .A2(n10566), .ZN(n10567) );
  AOI21_X1 U13076 ( .B1(n14559), .B2(n11931), .A(n10567), .ZN(n10570) );
  INV_X1 U13077 ( .A(n10570), .ZN(n10568) );
  NAND2_X1 U13078 ( .A1(n10569), .A2(n10568), .ZN(n10582) );
  INV_X1 U13079 ( .A(n10582), .ZN(n10572) );
  AND2_X1 U13080 ( .A1(n10571), .A2(n10570), .ZN(n10581) );
  NOR2_X1 U13081 ( .A1(n10572), .A2(n10581), .ZN(n10573) );
  XNOR2_X1 U13082 ( .A(n10583), .B(n10573), .ZN(n10579) );
  NAND2_X1 U13083 ( .A1(n13691), .A2(n13662), .ZN(n10575) );
  NAND2_X1 U13084 ( .A1(n13689), .A2(n13398), .ZN(n10574) );
  NAND2_X1 U13085 ( .A1(n10575), .A2(n10574), .ZN(n14548) );
  AOI22_X1 U13086 ( .A1(n14433), .A2(n14548), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10577) );
  AND2_X1 U13087 ( .A1(n14559), .A2(n14636), .ZN(n14620) );
  NAND2_X1 U13088 ( .A1(n14620), .A2(n14451), .ZN(n10576) );
  OAI211_X1 U13089 ( .C1(n14463), .C2(n14552), .A(n10577), .B(n10576), .ZN(
        n10578) );
  AOI21_X1 U13090 ( .B1(n10579), .B2(n14440), .A(n10578), .ZN(n10580) );
  INV_X1 U13091 ( .A(n10580), .ZN(P1_U3239) );
  INV_X1 U13092 ( .A(n13689), .ZN(n10628) );
  NOR2_X1 U13093 ( .A1(n9739), .A2(n10628), .ZN(n10584) );
  AOI21_X1 U13094 ( .B1(n13506), .B2(n11931), .A(n10584), .ZN(n10800) );
  AOI22_X1 U13095 ( .A1(n13506), .A2(n11930), .B1(n11931), .B2(n13689), .ZN(
        n10585) );
  XNOR2_X1 U13096 ( .A(n10585), .B(n11941), .ZN(n10799) );
  XOR2_X1 U13097 ( .A(n10800), .B(n10799), .Z(n10586) );
  OAI211_X1 U13098 ( .C1(n10587), .C2(n10586), .A(n10798), .B(n14440), .ZN(
        n10594) );
  NOR2_X1 U13099 ( .A1(n10588), .A2(n14655), .ZN(n14623) );
  NAND2_X1 U13100 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U13101 ( .A1(n14433), .A2(n10589), .ZN(n10590) );
  OAI211_X1 U13102 ( .C1(n14463), .C2(n10591), .A(n13765), .B(n10590), .ZN(
        n10592) );
  AOI21_X1 U13103 ( .B1(n14623), .B2(n14451), .A(n10592), .ZN(n10593) );
  NAND2_X1 U13104 ( .A1(n10594), .A2(n10593), .ZN(P1_U3213) );
  INV_X1 U13105 ( .A(n10595), .ZN(n10861) );
  INV_X1 U13106 ( .A(n10599), .ZN(n10597) );
  INV_X1 U13107 ( .A(n10598), .ZN(n10596) );
  XNOR2_X1 U13108 ( .A(n11032), .B(n10862), .ZN(n10655) );
  XNOR2_X1 U13109 ( .A(n10655), .B(n10720), .ZN(n10600) );
  NOR3_X1 U13110 ( .A1(n10597), .A2(n10596), .A3(n10600), .ZN(n10603) );
  INV_X1 U13111 ( .A(n10785), .ZN(n10602) );
  OAI21_X1 U13112 ( .B1(n10603), .B2(n10602), .A(n12058), .ZN(n10608) );
  INV_X1 U13113 ( .A(n10862), .ZN(n10606) );
  INV_X1 U13114 ( .A(n12136), .ZN(n10775) );
  OAI22_X1 U13115 ( .A1(n12112), .A2(n10745), .B1(n10775), .B2(n12120), .ZN(
        n10604) );
  AOI211_X1 U13116 ( .C1(n10606), .C2(n6545), .A(n10605), .B(n10604), .ZN(
        n10607) );
  OAI211_X1 U13117 ( .C1(n10861), .C2(n11042), .A(n10608), .B(n10607), .ZN(
        P3_U3167) );
  NAND2_X1 U13118 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U13119 ( .A1(n14433), .A2(n10609), .ZN(n10610) );
  OAI211_X1 U13120 ( .C1(n14463), .C2(n10611), .A(n13729), .B(n10610), .ZN(
        n10617) );
  NAND2_X1 U13121 ( .A1(n6598), .A2(n10612), .ZN(n10614) );
  XNOR2_X1 U13122 ( .A(n10614), .B(n10613), .ZN(n10615) );
  NOR2_X1 U13123 ( .A1(n10615), .A2(n14458), .ZN(n10616) );
  AOI211_X1 U13124 ( .C1(n14447), .C2(n13491), .A(n10617), .B(n10616), .ZN(
        n10618) );
  INV_X1 U13125 ( .A(n10618), .ZN(P1_U3230) );
  INV_X1 U13126 ( .A(n13423), .ZN(n10619) );
  OR2_X1 U13127 ( .A1(n13506), .A2(n13689), .ZN(n10621) );
  OR2_X1 U13128 ( .A1(n10622), .A2(n13453), .ZN(n10625) );
  AOI22_X1 U13129 ( .A1(n13455), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6562), 
        .B2(n10623), .ZN(n10624) );
  INV_X1 U13130 ( .A(n13688), .ZN(n10626) );
  OR2_X1 U13131 ( .A1(n14635), .A2(n10626), .ZN(n10693) );
  NAND2_X1 U13132 ( .A1(n14635), .A2(n10626), .ZN(n10627) );
  XNOR2_X1 U13133 ( .A(n10687), .B(n13425), .ZN(n14638) );
  NAND2_X1 U13134 ( .A1(n13506), .A2(n10628), .ZN(n10630) );
  NAND2_X1 U13135 ( .A1(n10632), .A2(n10630), .ZN(n10629) );
  INV_X1 U13136 ( .A(n13425), .ZN(n10686) );
  NAND2_X1 U13137 ( .A1(n10629), .A2(n10686), .ZN(n10633) );
  AND2_X1 U13138 ( .A1(n13425), .A2(n10630), .ZN(n10631) );
  NAND3_X1 U13139 ( .A1(n10633), .A2(n14571), .A3(n10694), .ZN(n10643) );
  NAND2_X1 U13140 ( .A1(n13689), .A2(n13662), .ZN(n10641) );
  NAND2_X1 U13141 ( .A1(n10245), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10639) );
  NAND2_X1 U13142 ( .A1(n10634), .A2(n10950), .ZN(n10635) );
  NAND2_X1 U13143 ( .A1(n10697), .A2(n10635), .ZN(n10949) );
  OR2_X1 U13144 ( .A1(n11769), .A2(n10949), .ZN(n10638) );
  NAND2_X1 U13145 ( .A1(n11778), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U13146 ( .A1(n13448), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13147 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n13687) );
  NAND2_X1 U13148 ( .A1(n13687), .A2(n13398), .ZN(n10640) );
  NAND2_X1 U13149 ( .A1(n10641), .A2(n10640), .ZN(n10803) );
  INV_X1 U13150 ( .A(n10803), .ZN(n10642) );
  NAND2_X1 U13151 ( .A1(n10643), .A2(n10642), .ZN(n14633) );
  MUX2_X1 U13152 ( .A(n14633), .B(P1_REG2_REG_8__SCAN_IN), .S(n14276), .Z(
        n10644) );
  INV_X1 U13153 ( .A(n10644), .ZN(n10648) );
  AOI211_X1 U13154 ( .C1(n14635), .C2(n10645), .A(n6570), .B(n7543), .ZN(
        n14634) );
  OAI22_X1 U13155 ( .A1(n7080), .A2(n14012), .B1(n10806), .B2(n14010), .ZN(
        n10646) );
  AOI21_X1 U13156 ( .B1(n14634), .B2(n14581), .A(n10646), .ZN(n10647) );
  OAI211_X1 U13157 ( .C1(n14638), .C2(n14020), .A(n10648), .B(n10647), .ZN(
        P1_U3285) );
  INV_X1 U13158 ( .A(n11693), .ZN(n10652) );
  OAI21_X1 U13159 ( .B1(n10649), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10650) );
  XNOR2_X1 U13160 ( .A(n10650), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13808) );
  INV_X1 U13161 ( .A(n13808), .ZN(n11386) );
  OAI222_X1 U13162 ( .A1(n14145), .A2(n10651), .B1(n14148), .B2(n10652), .C1(
        P1_U3086), .C2(n11386), .ZN(P1_U3337) );
  INV_X1 U13163 ( .A(n12949), .ZN(n11639) );
  OAI222_X1 U13164 ( .A1(n13269), .A2(n10653), .B1(n13272), .B2(n10652), .C1(
        P2_U3088), .C2(n11639), .ZN(P2_U3309) );
  INV_X1 U13165 ( .A(n10654), .ZN(n10854) );
  NAND2_X1 U13166 ( .A1(n10655), .A2(n10660), .ZN(n10773) );
  AND2_X1 U13167 ( .A1(n10785), .A2(n10773), .ZN(n10658) );
  XNOR2_X1 U13168 ( .A(n11032), .B(n10855), .ZN(n10776) );
  XNOR2_X1 U13169 ( .A(n10776), .B(n12136), .ZN(n10657) );
  AND2_X1 U13170 ( .A1(n10657), .A2(n10773), .ZN(n10656) );
  NAND2_X1 U13171 ( .A1(n10785), .A2(n10656), .ZN(n10732) );
  OAI211_X1 U13172 ( .C1(n10658), .C2(n10657), .A(n12058), .B(n10732), .ZN(
        n10665) );
  INV_X1 U13173 ( .A(n12037), .ZN(n10659) );
  OAI22_X1 U13174 ( .A1(n12112), .A2(n10660), .B1(n10659), .B2(n12120), .ZN(
        n10661) );
  AOI211_X1 U13175 ( .C1(n10663), .C2(n6545), .A(n10662), .B(n10661), .ZN(
        n10664) );
  OAI211_X1 U13176 ( .C1(n10854), .C2(n11042), .A(n10665), .B(n10664), .ZN(
        P3_U3179) );
  INV_X1 U13177 ( .A(n10666), .ZN(n10667) );
  AOI21_X1 U13178 ( .B1(n10669), .B2(n10668), .A(n10667), .ZN(n10671) );
  OAI21_X1 U13179 ( .B1(n10671), .B2(n13189), .A(n10670), .ZN(n14804) );
  INV_X1 U13180 ( .A(n14804), .ZN(n10684) );
  INV_X1 U13181 ( .A(n10672), .ZN(n10673) );
  AOI21_X1 U13182 ( .B1(n10675), .B2(n10674), .A(n10673), .ZN(n14806) );
  OAI211_X1 U13183 ( .C1(n10676), .C2(n14803), .A(n10011), .B(n10818), .ZN(
        n14802) );
  OAI22_X1 U13184 ( .A1(n6558), .A2(n10678), .B1(n10677), .B2(n14751), .ZN(
        n10679) );
  AOI21_X1 U13185 ( .B1(n10680), .B2(n14393), .A(n10679), .ZN(n10681) );
  OAI21_X1 U13186 ( .B1(n14802), .B2(n13129), .A(n10681), .ZN(n10682) );
  AOI21_X1 U13187 ( .B1(n14806), .B2(n10037), .A(n10682), .ZN(n10683) );
  OAI21_X1 U13188 ( .B1(n10684), .B2(n14736), .A(n10683), .ZN(P2_U3257) );
  NAND2_X1 U13189 ( .A1(n12140), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10685) );
  OAI21_X1 U13190 ( .B1(n12261), .B2(n12140), .A(n10685), .ZN(P3_U3519) );
  OR2_X1 U13191 ( .A1(n14635), .A2(n13688), .ZN(n10688) );
  NAND2_X1 U13192 ( .A1(n10689), .A2(n10688), .ZN(n10904) );
  OR2_X1 U13193 ( .A1(n10690), .A2(n13453), .ZN(n10692) );
  AOI22_X1 U13194 ( .A1(n13455), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6562), 
        .B2(n13792), .ZN(n10691) );
  XNOR2_X1 U13195 ( .A(n10904), .B(n13426), .ZN(n14643) );
  OAI21_X1 U13196 ( .B1(n10695), .B2(n13426), .A(n10923), .ZN(n10704) );
  NAND2_X1 U13197 ( .A1(n13448), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10702) );
  INV_X1 U13198 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10696) );
  AND2_X1 U13199 ( .A1(n10697), .A2(n10696), .ZN(n10698) );
  OR2_X1 U13200 ( .A1(n10698), .A2(n10917), .ZN(n14449) );
  OR2_X1 U13201 ( .A1(n11769), .A2(n14449), .ZN(n10701) );
  NAND2_X1 U13202 ( .A1(n10245), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10700) );
  NAND2_X1 U13203 ( .A1(n11778), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10699) );
  NAND4_X1 U13204 ( .A1(n10702), .A2(n10701), .A3(n10700), .A4(n10699), .ZN(
        n13686) );
  AOI22_X1 U13205 ( .A1(n13662), .A2(n13688), .B1(n13686), .B2(n13398), .ZN(
        n10951) );
  INV_X1 U13206 ( .A(n10951), .ZN(n10703) );
  AOI21_X1 U13207 ( .B1(n10704), .B2(n14571), .A(n10703), .ZN(n14645) );
  INV_X1 U13208 ( .A(n14645), .ZN(n10710) );
  XNOR2_X1 U13209 ( .A(n7543), .B(n13514), .ZN(n10705) );
  NAND2_X1 U13210 ( .A1(n10705), .A2(n14577), .ZN(n14644) );
  NAND2_X1 U13211 ( .A1(n14575), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10706) );
  OAI21_X1 U13212 ( .B1(n14010), .B2(n10949), .A(n10706), .ZN(n10707) );
  AOI21_X1 U13213 ( .B1(n13514), .B2(n14572), .A(n10707), .ZN(n10708) );
  OAI21_X1 U13214 ( .B1(n14644), .B2(n14016), .A(n10708), .ZN(n10709) );
  AOI21_X1 U13215 ( .B1(n10710), .B2(n14002), .A(n10709), .ZN(n10711) );
  OAI21_X1 U13216 ( .B1(n14020), .B2(n14643), .A(n10711), .ZN(P1_U3284) );
  NAND2_X1 U13217 ( .A1(n10712), .A2(n12602), .ZN(n10713) );
  OAI211_X1 U13218 ( .C1(n10714), .C2(n12606), .A(n10713), .B(n11622), .ZN(
        P3_U3272) );
  OAI21_X1 U13219 ( .B1(n10716), .B2(n11594), .A(n10715), .ZN(n10859) );
  NAND2_X1 U13220 ( .A1(n10717), .A2(n11594), .ZN(n10718) );
  NAND3_X1 U13221 ( .A1(n10719), .A2(n12450), .A3(n10718), .ZN(n10722) );
  AOI22_X1 U13222 ( .A1(n12453), .A2(n12037), .B1(n10720), .B2(n12456), .ZN(
        n10721) );
  NAND2_X1 U13223 ( .A1(n10722), .A2(n10721), .ZN(n10856) );
  AOI21_X1 U13224 ( .B1(n14963), .B2(n10859), .A(n10856), .ZN(n10729) );
  INV_X1 U13225 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n10723) );
  OAI22_X1 U13226 ( .A1(n12597), .A2(n10855), .B1(n14979), .B2(n10723), .ZN(
        n10724) );
  INV_X1 U13227 ( .A(n10724), .ZN(n10725) );
  OAI21_X1 U13228 ( .B1(n10729), .B2(n14977), .A(n10725), .ZN(P3_U3408) );
  OAI22_X1 U13229 ( .A1(n12544), .A2(n10855), .B1(n14989), .B2(n10726), .ZN(
        n10727) );
  INV_X1 U13230 ( .A(n10727), .ZN(n10728) );
  OAI21_X1 U13231 ( .B1(n10729), .B2(n14986), .A(n10728), .ZN(P3_U3465) );
  INV_X1 U13232 ( .A(n10776), .ZN(n10730) );
  AND2_X1 U13233 ( .A1(n10730), .A2(n12136), .ZN(n10778) );
  INV_X1 U13234 ( .A(n10778), .ZN(n10731) );
  NAND2_X1 U13235 ( .A1(n10732), .A2(n10731), .ZN(n12031) );
  XNOR2_X1 U13236 ( .A(n12031), .B(n12030), .ZN(n10737) );
  OAI22_X1 U13237 ( .A1(n12112), .A2(n10775), .B1(n10789), .B2(n12120), .ZN(
        n10733) );
  AOI211_X1 U13238 ( .C1(n10872), .C2(n6545), .A(n10734), .B(n10733), .ZN(
        n10736) );
  NAND2_X1 U13239 ( .A1(n12124), .A2(n10871), .ZN(n10735) );
  OAI211_X1 U13240 ( .C1(n10737), .C2(n12126), .A(n10736), .B(n10735), .ZN(
        P3_U3153) );
  NAND2_X1 U13241 ( .A1(n12140), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10738) );
  OAI21_X1 U13242 ( .B1(n12026), .B2(n12140), .A(n10738), .ZN(P3_U3520) );
  OAI21_X1 U13243 ( .B1(n10740), .B2(n11588), .A(n10739), .ZN(n10866) );
  INV_X1 U13244 ( .A(n10741), .ZN(n10742) );
  AOI21_X1 U13245 ( .B1(n11588), .B2(n10743), .A(n10742), .ZN(n10744) );
  OAI222_X1 U13246 ( .A1(n14941), .A2(n10745), .B1(n14943), .B2(n10775), .C1(
        n14939), .C2(n10744), .ZN(n10863) );
  AOI21_X1 U13247 ( .B1(n14963), .B2(n10866), .A(n10863), .ZN(n10751) );
  OAI22_X1 U13248 ( .A1(n12544), .A2(n10862), .B1(n14989), .B2(n9877), .ZN(
        n10746) );
  INV_X1 U13249 ( .A(n10746), .ZN(n10747) );
  OAI21_X1 U13250 ( .B1(n10751), .B2(n14986), .A(n10747), .ZN(P3_U3464) );
  INV_X1 U13251 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10748) );
  OAI22_X1 U13252 ( .A1(n12597), .A2(n10862), .B1(n14979), .B2(n10748), .ZN(
        n10749) );
  INV_X1 U13253 ( .A(n10749), .ZN(n10750) );
  OAI21_X1 U13254 ( .B1(n10751), .B2(n14977), .A(n10750), .ZN(P3_U3405) );
  INV_X1 U13255 ( .A(n10752), .ZN(n10754) );
  XNOR2_X1 U13256 ( .A(n10979), .B(n12663), .ZN(n10842) );
  AND2_X1 U13257 ( .A1(n12842), .A2(n12664), .ZN(n10756) );
  NAND2_X1 U13258 ( .A1(n10842), .A2(n10756), .ZN(n10843) );
  INV_X1 U13259 ( .A(n10842), .ZN(n10758) );
  INV_X1 U13260 ( .A(n10756), .ZN(n10757) );
  NAND2_X1 U13261 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  NAND2_X1 U13262 ( .A1(n10843), .A2(n10759), .ZN(n10761) );
  AOI21_X1 U13263 ( .B1(n10760), .B2(n10761), .A(n12792), .ZN(n10764) );
  INV_X1 U13264 ( .A(n10760), .ZN(n10763) );
  INV_X1 U13265 ( .A(n10761), .ZN(n10762) );
  NAND2_X1 U13266 ( .A1(n10764), .A2(n10844), .ZN(n10769) );
  AOI22_X1 U13267 ( .A1(n12800), .A2(n12843), .B1(n12841), .B2(n12801), .ZN(
        n10976) );
  INV_X1 U13268 ( .A(n10976), .ZN(n10767) );
  OAI21_X1 U13269 ( .B1(n14694), .B2(n10980), .A(n10765), .ZN(n10766) );
  AOI21_X1 U13270 ( .B1(n10767), .B2(n14685), .A(n10766), .ZN(n10768) );
  OAI211_X1 U13271 ( .C1(n7148), .C2(n12821), .A(n10769), .B(n10768), .ZN(
        P2_U3189) );
  INV_X1 U13272 ( .A(n11701), .ZN(n10771) );
  OAI222_X1 U13273 ( .A1(n13269), .A2(n10770), .B1(n13272), .B2(n10771), .C1(
        P2_U3088), .C2(n14748), .ZN(P2_U3308) );
  OAI222_X1 U13274 ( .A1(n14145), .A2(n10772), .B1(n14148), .B2(n10771), .C1(
        P1_U3086), .C2(n13965), .ZN(P1_U3336) );
  INV_X1 U13275 ( .A(n11050), .ZN(n10794) );
  XNOR2_X1 U13276 ( .A(n11032), .B(n14959), .ZN(n10780) );
  XNOR2_X1 U13277 ( .A(n10780), .B(n10789), .ZN(n12032) );
  NAND2_X1 U13278 ( .A1(n12030), .A2(n10773), .ZN(n10774) );
  AOI211_X1 U13279 ( .C1(n10776), .C2(n10775), .A(n12032), .B(n10774), .ZN(
        n10784) );
  INV_X1 U13280 ( .A(n12032), .ZN(n10779) );
  AOI21_X1 U13281 ( .B1(n10779), .B2(n12037), .A(n12030), .ZN(n10782) );
  INV_X1 U13282 ( .A(n12030), .ZN(n10777) );
  AOI21_X1 U13283 ( .B1(n10779), .B2(n10778), .A(n10777), .ZN(n10781) );
  OAI22_X1 U13284 ( .A1(n10782), .A2(n10781), .B1(n10789), .B2(n10780), .ZN(
        n10783) );
  XNOR2_X1 U13285 ( .A(n11032), .B(n14967), .ZN(n11034) );
  XNOR2_X1 U13286 ( .A(n11034), .B(n11473), .ZN(n10786) );
  OAI21_X1 U13287 ( .B1(n10787), .B2(n10786), .A(n11033), .ZN(n10788) );
  NAND2_X1 U13288 ( .A1(n10788), .A2(n12058), .ZN(n10793) );
  INV_X1 U13289 ( .A(n12133), .ZN(n11317) );
  OAI22_X1 U13290 ( .A1(n12112), .A2(n10789), .B1(n11317), .B2(n12120), .ZN(
        n10790) );
  AOI211_X1 U13291 ( .C1(n14967), .C2(n6545), .A(n10791), .B(n10790), .ZN(
        n10792) );
  OAI211_X1 U13292 ( .C1(n10794), .C2(n11042), .A(n10793), .B(n10792), .ZN(
        P3_U3171) );
  AOI22_X1 U13293 ( .A1(n14635), .A2(n11931), .B1(n6565), .B2(n13688), .ZN(
        n10941) );
  NAND2_X1 U13294 ( .A1(n14635), .A2(n11930), .ZN(n10796) );
  NAND2_X1 U13295 ( .A1(n11931), .A2(n13688), .ZN(n10795) );
  NAND2_X1 U13296 ( .A1(n10796), .A2(n10795), .ZN(n10797) );
  XNOR2_X1 U13297 ( .A(n10797), .B(n11941), .ZN(n10938) );
  XOR2_X1 U13298 ( .A(n10941), .B(n10938), .Z(n10802) );
  AOI21_X1 U13299 ( .B1(n10802), .B2(n10801), .A(n10939), .ZN(n10809) );
  NAND2_X1 U13300 ( .A1(n14433), .A2(n10803), .ZN(n10804) );
  OAI211_X1 U13301 ( .C1(n14463), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n10807) );
  AOI21_X1 U13302 ( .B1(n14635), .B2(n14447), .A(n10807), .ZN(n10808) );
  OAI21_X1 U13303 ( .B1(n10809), .B2(n14458), .A(n10808), .ZN(P1_U3221) );
  XNOR2_X1 U13304 ( .A(n10811), .B(n10810), .ZN(n10898) );
  OAI211_X1 U13305 ( .C1(n10814), .C2(n10813), .A(n10812), .B(n14753), .ZN(
        n10815) );
  OAI211_X1 U13306 ( .C1(n10898), .C2(n6774), .A(n10816), .B(n10815), .ZN(
        n10893) );
  NAND2_X1 U13307 ( .A1(n10893), .A2(n6558), .ZN(n10825) );
  INV_X1 U13308 ( .A(n10978), .ZN(n10817) );
  AOI211_X1 U13309 ( .C1(n6569), .C2(n10818), .A(n12664), .B(n10817), .ZN(
        n10894) );
  INV_X1 U13310 ( .A(n6569), .ZN(n10819) );
  NOR2_X1 U13311 ( .A1(n10819), .A2(n14739), .ZN(n10823) );
  OAI22_X1 U13312 ( .A1(n6558), .A2(n10821), .B1(n10820), .B2(n14751), .ZN(
        n10822) );
  AOI211_X1 U13313 ( .C1(n10894), .C2(n14731), .A(n10823), .B(n10822), .ZN(
        n10824) );
  OAI211_X1 U13314 ( .C1(n10898), .C2(n10826), .A(n10825), .B(n10824), .ZN(
        P2_U3256) );
  OAI21_X1 U13315 ( .B1(n10828), .B2(n11589), .A(n10827), .ZN(n10868) );
  OAI211_X1 U13316 ( .C1(n10831), .C2(n10830), .A(n10829), .B(n12450), .ZN(
        n10833) );
  AOI22_X1 U13317 ( .A1(n12456), .A2(n12136), .B1(n12135), .B2(n12453), .ZN(
        n10832) );
  NAND2_X1 U13318 ( .A1(n10833), .A2(n10832), .ZN(n10869) );
  AOI21_X1 U13319 ( .B1(n14963), .B2(n10868), .A(n10869), .ZN(n10841) );
  INV_X1 U13320 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n10834) );
  OAI22_X1 U13321 ( .A1(n12597), .A2(n10838), .B1(n14979), .B2(n10834), .ZN(
        n10835) );
  INV_X1 U13322 ( .A(n10835), .ZN(n10836) );
  OAI21_X1 U13323 ( .B1(n10841), .B2(n14977), .A(n10836), .ZN(P3_U3411) );
  INV_X1 U13324 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10837) );
  OAI22_X1 U13325 ( .A1(n12544), .A2(n10838), .B1(n14989), .B2(n10837), .ZN(
        n10839) );
  INV_X1 U13326 ( .A(n10839), .ZN(n10840) );
  OAI21_X1 U13327 ( .B1(n10841), .B2(n14986), .A(n10840), .ZN(P3_U3466) );
  XNOR2_X1 U13328 ( .A(n11027), .B(n6554), .ZN(n11111) );
  NAND2_X1 U13329 ( .A1(n12841), .A2(n12619), .ZN(n11112) );
  XNOR2_X1 U13330 ( .A(n11111), .B(n11112), .ZN(n10853) );
  NAND3_X1 U13331 ( .A1(n10842), .A2(n12813), .A3(n12842), .ZN(n10852) );
  OAI21_X1 U13332 ( .B1(n10844), .B2(n10853), .A(n11115), .ZN(n10845) );
  NAND2_X1 U13333 ( .A1(n10845), .A2(n14688), .ZN(n10851) );
  NAND2_X1 U13334 ( .A1(n12842), .A2(n12800), .ZN(n10847) );
  NAND2_X1 U13335 ( .A1(n12840), .A2(n12801), .ZN(n10846) );
  AND2_X1 U13336 ( .A1(n10847), .A2(n10846), .ZN(n11021) );
  NOR2_X1 U13337 ( .A1(n11021), .A2(n12806), .ZN(n10849) );
  NAND2_X1 U13338 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12923)
         );
  OAI21_X1 U13339 ( .B1(n14694), .B2(n11023), .A(n12923), .ZN(n10848) );
  AOI211_X1 U13340 ( .C1(n11027), .C2(n14690), .A(n10849), .B(n10848), .ZN(
        n10850) );
  OAI211_X1 U13341 ( .C1(n10853), .C2(n10852), .A(n10851), .B(n10850), .ZN(
        P2_U3208) );
  OAI22_X1 U13342 ( .A1(n12428), .A2(n10855), .B1(n10854), .B2(n14934), .ZN(
        n10858) );
  MUX2_X1 U13343 ( .A(n10856), .B(P3_REG2_REG_6__SCAN_IN), .S(n14949), .Z(
        n10857) );
  AOI211_X1 U13344 ( .C1(n12471), .C2(n10859), .A(n10858), .B(n10857), .ZN(
        n10860) );
  INV_X1 U13345 ( .A(n10860), .ZN(P3_U3227) );
  OAI22_X1 U13346 ( .A1(n12428), .A2(n10862), .B1(n10861), .B2(n14934), .ZN(
        n10865) );
  MUX2_X1 U13347 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n10863), .S(n14946), .Z(
        n10864) );
  AOI211_X1 U13348 ( .C1(n12471), .C2(n10866), .A(n10865), .B(n10864), .ZN(
        n10867) );
  INV_X1 U13349 ( .A(n10867), .ZN(P3_U3228) );
  INV_X1 U13350 ( .A(n10868), .ZN(n10875) );
  MUX2_X1 U13351 ( .A(n10869), .B(P3_REG2_REG_7__SCAN_IN), .S(n14949), .Z(
        n10870) );
  INV_X1 U13352 ( .A(n10870), .ZN(n10874) );
  AOI22_X1 U13353 ( .A1(n12470), .A2(n10872), .B1(n12468), .B2(n10871), .ZN(
        n10873) );
  OAI211_X1 U13354 ( .C1(n12431), .C2(n10875), .A(n10874), .B(n10873), .ZN(
        P3_U3226) );
  INV_X1 U13355 ( .A(n10878), .ZN(n10879) );
  XNOR2_X1 U13356 ( .A(n10878), .B(n11244), .ZN(n14530) );
  NOR2_X1 U13357 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14530), .ZN(n14529) );
  XOR2_X1 U13358 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11291), .Z(n10880) );
  NAND2_X1 U13359 ( .A1(n10880), .A2(n10881), .ZN(n11270) );
  OAI211_X1 U13360 ( .C1(n10881), .C2(n10880), .A(n13819), .B(n11270), .ZN(
        n10892) );
  NAND2_X1 U13361 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13332)
         );
  NAND2_X1 U13362 ( .A1(n11172), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13363 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  INV_X1 U13364 ( .A(n10884), .ZN(n10885) );
  XNOR2_X1 U13365 ( .A(n10884), .B(n11244), .ZN(n14532) );
  NOR2_X1 U13366 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14532), .ZN(n14531) );
  AOI21_X1 U13367 ( .B1(n14537), .B2(n10885), .A(n14531), .ZN(n10888) );
  INV_X1 U13368 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11268) );
  NOR2_X1 U13369 ( .A1(n11268), .A2(n11269), .ZN(n10886) );
  AOI21_X1 U13370 ( .B1(n11268), .B2(n11269), .A(n10886), .ZN(n10887) );
  NAND2_X1 U13371 ( .A1(n10887), .A2(n10888), .ZN(n11267) );
  OAI211_X1 U13372 ( .C1(n10888), .C2(n10887), .A(n13813), .B(n11267), .ZN(
        n10889) );
  NAND2_X1 U13373 ( .A1(n13332), .A2(n10889), .ZN(n10890) );
  AOI21_X1 U13374 ( .B1(n14525), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10890), 
        .ZN(n10891) );
  OAI211_X1 U13375 ( .C1(n6779), .C2(n11269), .A(n10892), .B(n10891), .ZN(
        P1_U3259) );
  INV_X1 U13376 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10900) );
  INV_X1 U13377 ( .A(n10893), .ZN(n10897) );
  AOI21_X1 U13378 ( .B1(n14795), .B2(n6569), .A(n10894), .ZN(n10896) );
  OAI211_X1 U13379 ( .C1(n10898), .C2(n14809), .A(n10897), .B(n10896), .ZN(
        n10901) );
  NAND2_X1 U13380 ( .A1(n10901), .A2(n14814), .ZN(n10899) );
  OAI21_X1 U13381 ( .B1(n14814), .B2(n10900), .A(n10899), .ZN(P2_U3457) );
  NAND2_X1 U13382 ( .A1(n10901), .A2(n14833), .ZN(n10902) );
  OAI21_X1 U13383 ( .B1(n14833), .B2(n7832), .A(n10902), .ZN(P2_U3508) );
  INV_X1 U13384 ( .A(n13426), .ZN(n10903) );
  NAND2_X1 U13385 ( .A1(n10904), .A2(n10903), .ZN(n10906) );
  OR2_X1 U13386 ( .A1(n13514), .A2(n13687), .ZN(n10905) );
  NAND2_X1 U13387 ( .A1(n10907), .A2(n13444), .ZN(n10910) );
  AOI22_X1 U13388 ( .A1(n10908), .A2(n6562), .B1(n13455), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10909) );
  INV_X1 U13389 ( .A(n13686), .ZN(n11334) );
  OR2_X1 U13390 ( .A1(n14653), .A2(n11334), .ZN(n10924) );
  NAND2_X1 U13391 ( .A1(n14653), .A2(n11334), .ZN(n10911) );
  NAND2_X1 U13392 ( .A1(n10924), .A2(n10911), .ZN(n13428) );
  OR2_X1 U13393 ( .A1(n14653), .A2(n13686), .ZN(n10912) );
  NAND2_X1 U13394 ( .A1(n10913), .A2(n13444), .ZN(n10916) );
  AOI22_X1 U13395 ( .A1(n10914), .A2(n6562), .B1(n13455), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U13396 ( .A1(n10245), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10922) );
  NOR2_X1 U13397 ( .A1(n10917), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10918) );
  OR2_X1 U13398 ( .A1(n10925), .A2(n10918), .ZN(n14464) );
  OR2_X1 U13399 ( .A1(n11769), .A2(n14464), .ZN(n10921) );
  NAND2_X1 U13400 ( .A1(n11778), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13401 ( .A1(n13448), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10919) );
  NAND4_X1 U13402 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n13685) );
  INV_X1 U13403 ( .A(n13685), .ZN(n11077) );
  XNOR2_X1 U13404 ( .A(n14450), .B(n11077), .ZN(n13429) );
  INV_X1 U13405 ( .A(n13429), .ZN(n11075) );
  XNOR2_X1 U13406 ( .A(n11054), .B(n11075), .ZN(n14484) );
  INV_X1 U13407 ( .A(n13687), .ZN(n10945) );
  NAND2_X1 U13408 ( .A1(n10960), .A2(n10924), .ZN(n11076) );
  XNOR2_X1 U13409 ( .A(n11076), .B(n11075), .ZN(n10931) );
  NAND2_X1 U13410 ( .A1(n13448), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10930) );
  OR2_X1 U13411 ( .A1(n10925), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13412 ( .A1(n11069), .A2(n10926), .ZN(n11351) );
  OR2_X1 U13413 ( .A1(n11769), .A2(n11351), .ZN(n10929) );
  NAND2_X1 U13414 ( .A1(n10245), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U13415 ( .A1(n11778), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U13416 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n13684) );
  AOI22_X1 U13417 ( .A1(n13662), .A2(n13686), .B1(n13684), .B2(n13398), .ZN(
        n14457) );
  OAI21_X1 U13418 ( .B1(n10931), .B2(n14550), .A(n14457), .ZN(n14486) );
  NAND2_X1 U13419 ( .A1(n14486), .A2(n14002), .ZN(n10937) );
  OAI22_X1 U13420 ( .A1(n14002), .A2(n10932), .B1(n14464), .B2(n14010), .ZN(
        n10935) );
  INV_X1 U13421 ( .A(n14450), .ZN(n10933) );
  INV_X1 U13422 ( .A(n13514), .ZN(n14646) );
  NAND2_X1 U13423 ( .A1(n10933), .A2(n10963), .ZN(n14277) );
  OAI211_X1 U13424 ( .C1(n10933), .C2(n10963), .A(n14577), .B(n14277), .ZN(
        n14482) );
  NOR2_X1 U13425 ( .A1(n14482), .A2(n14016), .ZN(n10934) );
  AOI211_X1 U13426 ( .C1(n14572), .C2(n14450), .A(n10935), .B(n10934), .ZN(
        n10936) );
  OAI211_X1 U13427 ( .C1(n14484), .C2(n14020), .A(n10937), .B(n10936), .ZN(
        P1_U3282) );
  INV_X1 U13428 ( .A(n10938), .ZN(n10940) );
  NAND2_X1 U13429 ( .A1(n13514), .A2(n11930), .ZN(n10943) );
  NAND2_X1 U13430 ( .A1(n11931), .A2(n13687), .ZN(n10942) );
  NAND2_X1 U13431 ( .A1(n10943), .A2(n10942), .ZN(n10944) );
  XNOR2_X1 U13432 ( .A(n10944), .B(n11941), .ZN(n11329) );
  NOR2_X1 U13433 ( .A1(n9739), .A2(n10945), .ZN(n10946) );
  AOI21_X1 U13434 ( .B1(n13514), .B2(n11931), .A(n10946), .ZN(n11330) );
  XNOR2_X1 U13435 ( .A(n11329), .B(n11330), .ZN(n10947) );
  OAI211_X1 U13436 ( .C1(n10948), .C2(n10947), .A(n11333), .B(n14440), .ZN(
        n10955) );
  INV_X1 U13437 ( .A(n10949), .ZN(n10953) );
  INV_X1 U13438 ( .A(n14463), .ZN(n13410) );
  OAI22_X1 U13439 ( .A1(n14456), .A2(n10951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10950), .ZN(n10952) );
  AOI21_X1 U13440 ( .B1(n10953), .B2(n13410), .A(n10952), .ZN(n10954) );
  OAI211_X1 U13441 ( .C1(n14646), .C2(n13414), .A(n10955), .B(n10954), .ZN(
        P1_U3231) );
  INV_X1 U13442 ( .A(n10956), .ZN(n10958) );
  OAI222_X1 U13443 ( .A1(P3_U3151), .A2(n8777), .B1(n12609), .B2(n10958), .C1(
        n10957), .C2(n12606), .ZN(P3_U3271) );
  XOR2_X1 U13444 ( .A(n13428), .B(n10959), .Z(n14652) );
  INV_X1 U13445 ( .A(n10960), .ZN(n10961) );
  AOI211_X1 U13446 ( .C1(n13428), .C2(n10962), .A(n14550), .B(n10961), .ZN(
        n14657) );
  AOI211_X1 U13447 ( .C1(n14653), .C2(n10964), .A(n6570), .B(n10963), .ZN(
        n10968) );
  NAND2_X1 U13448 ( .A1(n13687), .A2(n13662), .ZN(n10966) );
  NAND2_X1 U13449 ( .A1(n13685), .A2(n13398), .ZN(n10965) );
  AND2_X1 U13450 ( .A1(n10966), .A2(n10965), .ZN(n14439) );
  INV_X1 U13451 ( .A(n14439), .ZN(n10967) );
  NOR2_X1 U13452 ( .A1(n10968), .A2(n10967), .ZN(n14654) );
  NOR2_X1 U13453 ( .A1(n14654), .A2(n13952), .ZN(n10969) );
  OAI21_X1 U13454 ( .B1(n14657), .B2(n10969), .A(n14002), .ZN(n10972) );
  OAI22_X1 U13455 ( .A1(n14002), .A2(n9495), .B1(n14449), .B2(n14010), .ZN(
        n10970) );
  AOI21_X1 U13456 ( .B1(n14653), .B2(n14572), .A(n10970), .ZN(n10971) );
  OAI211_X1 U13457 ( .C1(n14652), .C2(n14020), .A(n10972), .B(n10971), .ZN(
        P1_U3283) );
  XNOR2_X1 U13458 ( .A(n10973), .B(n10975), .ZN(n14807) );
  XOR2_X1 U13459 ( .A(n10975), .B(n10974), .Z(n10977) );
  OAI21_X1 U13460 ( .B1(n10977), .B2(n13189), .A(n10976), .ZN(n14813) );
  NAND2_X1 U13461 ( .A1(n14813), .A2(n6558), .ZN(n10985) );
  AOI211_X1 U13462 ( .C1(n10979), .C2(n10978), .A(n12664), .B(n6712), .ZN(
        n14811) );
  NOR2_X1 U13463 ( .A1(n7148), .A2(n14739), .ZN(n10983) );
  OAI22_X1 U13464 ( .A1(n6558), .A2(n10981), .B1(n10980), .B2(n14751), .ZN(
        n10982) );
  AOI211_X1 U13465 ( .C1(n14811), .C2(n14731), .A(n10983), .B(n10982), .ZN(
        n10984) );
  OAI211_X1 U13466 ( .C1(n13114), .C2(n14807), .A(n10985), .B(n10984), .ZN(
        P2_U3255) );
  NAND2_X1 U13467 ( .A1(n11133), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10993) );
  XNOR2_X1 U13468 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11007), .ZN(n11130) );
  AOI21_X1 U13469 ( .B1(n9891), .B2(n10997), .A(n10986), .ZN(n14713) );
  MUX2_X1 U13470 ( .A(n10987), .B(P2_REG1_REG_13__SCAN_IN), .S(n10999), .Z(
        n14712) );
  NAND2_X1 U13471 ( .A1(n14713), .A2(n14712), .ZN(n14711) );
  OAI21_X1 U13472 ( .B1(n10987), .B2(n10999), .A(n14711), .ZN(n12936) );
  NAND2_X1 U13473 ( .A1(n12938), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10988) );
  OAI21_X1 U13474 ( .B1(n12938), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10988), 
        .ZN(n10989) );
  INV_X1 U13475 ( .A(n10989), .ZN(n12935) );
  NAND2_X1 U13476 ( .A1(n12936), .A2(n12935), .ZN(n12934) );
  OAI21_X1 U13477 ( .B1(n7910), .B2(n11002), .A(n12934), .ZN(n10990) );
  INV_X1 U13478 ( .A(n10990), .ZN(n10992) );
  XNOR2_X1 U13479 ( .A(n10990), .B(n14719), .ZN(n14724) );
  INV_X1 U13480 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10991) );
  OAI22_X1 U13481 ( .A1(n10992), .A2(n11006), .B1(n14724), .B2(n10991), .ZN(
        n11129) );
  NAND2_X1 U13482 ( .A1(n11130), .A2(n11129), .ZN(n11128) );
  NAND2_X1 U13483 ( .A1(n10993), .A2(n11128), .ZN(n11635) );
  INV_X1 U13484 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10994) );
  XNOR2_X1 U13485 ( .A(n11636), .B(n10994), .ZN(n11634) );
  XNOR2_X1 U13486 ( .A(n11635), .B(n11634), .ZN(n11015) );
  NAND2_X1 U13487 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12751)
         );
  NAND2_X1 U13488 ( .A1(n11636), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11630) );
  INV_X1 U13489 ( .A(n11630), .ZN(n10995) );
  AOI21_X1 U13490 ( .B1(n13107), .B2(n11011), .A(n10995), .ZN(n11009) );
  MUX2_X1 U13491 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13125), .S(n11133), .Z(
        n11126) );
  NAND2_X1 U13492 ( .A1(n14710), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11000) );
  AOI21_X1 U13493 ( .B1(n10997), .B2(n15207), .A(n10996), .ZN(n14709) );
  INV_X1 U13494 ( .A(n11000), .ZN(n10998) );
  AOI21_X1 U13495 ( .B1(n7896), .B2(n10999), .A(n10998), .ZN(n14708) );
  NAND2_X1 U13496 ( .A1(n14709), .A2(n14708), .ZN(n14707) );
  NAND2_X1 U13497 ( .A1(n11000), .A2(n14707), .ZN(n11001) );
  NAND2_X1 U13498 ( .A1(n12938), .A2(n11001), .ZN(n11003) );
  XNOR2_X1 U13499 ( .A(n11002), .B(n11001), .ZN(n12940) );
  NAND2_X1 U13500 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n12940), .ZN(n12939) );
  NAND2_X1 U13501 ( .A1(n11003), .A2(n12939), .ZN(n11004) );
  XNOR2_X1 U13502 ( .A(n11004), .B(n14719), .ZN(n14721) );
  INV_X1 U13503 ( .A(n11004), .ZN(n11005) );
  OAI22_X1 U13504 ( .A1(n14721), .A2(n11360), .B1(n11006), .B2(n11005), .ZN(
        n11127) );
  NAND2_X1 U13505 ( .A1(n11126), .A2(n11127), .ZN(n11125) );
  OAI21_X1 U13506 ( .B1(n11007), .B2(n13125), .A(n11125), .ZN(n11008) );
  NAND2_X1 U13507 ( .A1(n11008), .A2(n11009), .ZN(n11629) );
  OAI211_X1 U13508 ( .C1(n11009), .C2(n11008), .A(n6547), .B(n11629), .ZN(
        n11010) );
  NAND2_X1 U13509 ( .A1(n12751), .A2(n11010), .ZN(n11013) );
  NOR2_X1 U13510 ( .A1(n12925), .A2(n11011), .ZN(n11012) );
  AOI211_X1 U13511 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n14718), .A(n11013), 
        .B(n11012), .ZN(n11014) );
  OAI21_X1 U13512 ( .B1(n11015), .B2(n11644), .A(n11014), .ZN(P2_U3231) );
  XNOR2_X1 U13513 ( .A(n11017), .B(n11016), .ZN(n14815) );
  INV_X1 U13514 ( .A(n14815), .ZN(n11030) );
  XNOR2_X1 U13515 ( .A(n11019), .B(n11018), .ZN(n11020) );
  NAND2_X1 U13516 ( .A1(n11020), .A2(n14753), .ZN(n11022) );
  NAND2_X1 U13517 ( .A1(n11022), .A2(n11021), .ZN(n14823) );
  NAND2_X1 U13518 ( .A1(n14823), .A2(n6558), .ZN(n11029) );
  OAI22_X1 U13519 ( .A1(n6558), .A2(n11024), .B1(n11023), .B2(n14751), .ZN(
        n11026) );
  OAI211_X1 U13520 ( .C1(n14820), .C2(n6712), .A(n10011), .B(n11160), .ZN(
        n14818) );
  NOR2_X1 U13521 ( .A1(n14818), .A2(n13129), .ZN(n11025) );
  AOI211_X1 U13522 ( .C1(n14393), .C2(n11027), .A(n11026), .B(n11025), .ZN(
        n11028) );
  OAI211_X1 U13523 ( .C1(n13114), .C2(n11030), .A(n11029), .B(n11028), .ZN(
        P2_U3254) );
  INV_X1 U13524 ( .A(n11031), .ZN(n11148) );
  XNOR2_X1 U13525 ( .A(n11032), .B(n11150), .ZN(n11101) );
  XNOR2_X1 U13526 ( .A(n11101), .B(n12133), .ZN(n11036) );
  AOI211_X1 U13527 ( .C1(n11036), .C2(n11035), .A(n12126), .B(n11100), .ZN(
        n11037) );
  INV_X1 U13528 ( .A(n11037), .ZN(n11041) );
  OAI22_X1 U13529 ( .A1(n12112), .A2(n11473), .B1(n11231), .B2(n12120), .ZN(
        n11038) );
  AOI211_X1 U13530 ( .C1(n11150), .C2(n6545), .A(n11039), .B(n11038), .ZN(
        n11040) );
  OAI211_X1 U13531 ( .C1(n11148), .C2(n11042), .A(n11041), .B(n11040), .ZN(
        P3_U3157) );
  INV_X1 U13532 ( .A(n11712), .ZN(n11109) );
  OAI222_X1 U13533 ( .A1(n13272), .A2(n11109), .B1(n11044), .B2(P2_U3088), 
        .C1(n11043), .C2(n13269), .ZN(P2_U3307) );
  XNOR2_X1 U13534 ( .A(n11045), .B(n11468), .ZN(n14969) );
  OAI211_X1 U13535 ( .C1(n11047), .C2(n11468), .A(n11046), .B(n12450), .ZN(
        n11049) );
  AOI22_X1 U13536 ( .A1(n12456), .A2(n12135), .B1(n12133), .B2(n12453), .ZN(
        n11048) );
  NAND2_X1 U13537 ( .A1(n11049), .A2(n11048), .ZN(n14965) );
  AOI22_X1 U13538 ( .A1(n14949), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n12468), 
        .B2(n11050), .ZN(n11051) );
  OAI21_X1 U13539 ( .B1(n12428), .B2(n11474), .A(n11051), .ZN(n11052) );
  AOI21_X1 U13540 ( .B1(n14965), .B2(n14946), .A(n11052), .ZN(n11053) );
  OAI21_X1 U13541 ( .B1(n12431), .B2(n14969), .A(n11053), .ZN(P3_U3224) );
  NAND2_X1 U13542 ( .A1(n11055), .A2(n13444), .ZN(n11058) );
  AOI22_X1 U13543 ( .A1(n11056), .A2(n6562), .B1(n13455), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11057) );
  INV_X1 U13544 ( .A(n13684), .ZN(n11348) );
  XNOR2_X1 U13545 ( .A(n14274), .B(n11348), .ZN(n14266) );
  NAND2_X1 U13546 ( .A1(n14267), .A2(n14266), .ZN(n11060) );
  OR2_X1 U13547 ( .A1(n14274), .A2(n13684), .ZN(n11059) );
  NAND2_X1 U13548 ( .A1(n11060), .A2(n11059), .ZN(n11187) );
  NAND2_X1 U13549 ( .A1(n11061), .A2(n13444), .ZN(n11067) );
  OAI22_X1 U13550 ( .A1(n11064), .A2(n11671), .B1(n11063), .B2(n11062), .ZN(
        n11065) );
  INV_X1 U13551 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13552 ( .A1(n13448), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11074) );
  INV_X1 U13553 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U13554 ( .A1(n11069), .A2(n11068), .ZN(n11070) );
  NAND2_X1 U13555 ( .A1(n11085), .A2(n11070), .ZN(n13369) );
  OR2_X1 U13556 ( .A1(n11769), .A2(n13369), .ZN(n11073) );
  NAND2_X1 U13557 ( .A1(n10245), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U13558 ( .A1(n13449), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U13559 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n13683) );
  INV_X1 U13560 ( .A(n13683), .ZN(n13534) );
  XNOR2_X1 U13561 ( .A(n14476), .B(n13534), .ZN(n13431) );
  XNOR2_X1 U13562 ( .A(n11187), .B(n13431), .ZN(n14481) );
  INV_X1 U13563 ( .A(n14481), .ZN(n11099) );
  NAND2_X1 U13564 ( .A1(n11076), .A2(n11075), .ZN(n11079) );
  OR2_X1 U13565 ( .A1(n14450), .A2(n11077), .ZN(n11078) );
  NAND2_X1 U13566 ( .A1(n11079), .A2(n11078), .ZN(n14269) );
  INV_X1 U13567 ( .A(n14266), .ZN(n14268) );
  NAND2_X1 U13568 ( .A1(n14269), .A2(n14268), .ZN(n11081) );
  OR2_X1 U13569 ( .A1(n14274), .A2(n11348), .ZN(n11080) );
  NAND2_X1 U13570 ( .A1(n11081), .A2(n11080), .ZN(n11168) );
  XNOR2_X1 U13571 ( .A(n11168), .B(n13431), .ZN(n14473) );
  NAND2_X1 U13572 ( .A1(n14476), .A2(n14278), .ZN(n11082) );
  NAND2_X1 U13573 ( .A1(n11175), .A2(n11082), .ZN(n14479) );
  NOR2_X1 U13574 ( .A1(n14002), .A2(n11083), .ZN(n11094) );
  INV_X1 U13575 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U13576 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  NAND2_X1 U13577 ( .A1(n11178), .A2(n11086), .ZN(n14437) );
  OR2_X1 U13578 ( .A1(n11769), .A2(n14437), .ZN(n11090) );
  NAND2_X1 U13579 ( .A1(n10245), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11089) );
  NAND2_X1 U13580 ( .A1(n13449), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U13581 ( .A1(n13448), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11087) );
  NAND4_X1 U13582 ( .A1(n11090), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n13682) );
  NAND2_X1 U13583 ( .A1(n13682), .A2(n13398), .ZN(n11092) );
  NAND2_X1 U13584 ( .A1(n13684), .A2(n13662), .ZN(n11091) );
  AND2_X1 U13585 ( .A1(n11092), .A2(n11091), .ZN(n14474) );
  OAI22_X1 U13586 ( .A1(n14575), .A2(n14474), .B1(n13369), .B2(n14010), .ZN(
        n11093) );
  AOI211_X1 U13587 ( .C1(n14476), .C2(n14572), .A(n11094), .B(n11093), .ZN(
        n11095) );
  OAI21_X1 U13588 ( .B1(n14479), .B2(n11096), .A(n11095), .ZN(n11097) );
  AOI21_X1 U13589 ( .B1(n14473), .B2(n14018), .A(n11097), .ZN(n11098) );
  OAI21_X1 U13590 ( .B1(n14020), .B2(n11099), .A(n11098), .ZN(P1_U3280) );
  XNOR2_X1 U13591 ( .A(n11032), .B(n11105), .ZN(n11224) );
  XNOR2_X1 U13592 ( .A(n11224), .B(n12455), .ZN(n11102) );
  XNOR2_X1 U13593 ( .A(n11227), .B(n11102), .ZN(n11108) );
  NAND2_X1 U13594 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14847)
         );
  INV_X1 U13595 ( .A(n14847), .ZN(n11104) );
  INV_X1 U13596 ( .A(n12437), .ZN(n11318) );
  OAI22_X1 U13597 ( .A1(n12112), .A2(n11317), .B1(n11318), .B2(n12120), .ZN(
        n11103) );
  AOI211_X1 U13598 ( .C1(n11105), .C2(n6545), .A(n11104), .B(n11103), .ZN(
        n11107) );
  NAND2_X1 U13599 ( .A1(n12124), .A2(n11320), .ZN(n11106) );
  OAI211_X1 U13600 ( .C1(n11108), .C2(n12126), .A(n11107), .B(n11106), .ZN(
        P3_U3176) );
  OAI222_X1 U13601 ( .A1(n14145), .A2(n11110), .B1(n14148), .B2(n11109), .C1(
        n13636), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13602 ( .A(n11111), .ZN(n11113) );
  NAND2_X1 U13603 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  XNOR2_X1 U13604 ( .A(n14689), .B(n12673), .ZN(n11116) );
  NAND2_X1 U13605 ( .A1(n12840), .A2(n12619), .ZN(n11117) );
  AND2_X1 U13606 ( .A1(n11116), .A2(n11117), .ZN(n14681) );
  INV_X1 U13607 ( .A(n11116), .ZN(n11119) );
  INV_X1 U13608 ( .A(n11117), .ZN(n11118) );
  NAND2_X1 U13609 ( .A1(n11119), .A2(n11118), .ZN(n14680) );
  XNOR2_X1 U13610 ( .A(n14410), .B(n6554), .ZN(n12616) );
  NAND2_X1 U13611 ( .A1(n12839), .A2(n12619), .ZN(n12614) );
  XNOR2_X1 U13612 ( .A(n12616), .B(n12614), .ZN(n12612) );
  XNOR2_X1 U13613 ( .A(n12613), .B(n12612), .ZN(n11124) );
  OAI22_X1 U13614 ( .A1(n11359), .A2(n14754), .B1(n11120), .B2(n14378), .ZN(
        n14409) );
  INV_X1 U13615 ( .A(n14409), .ZN(n11211) );
  NOR2_X1 U13616 ( .A1(n11211), .A2(n12806), .ZN(n11122) );
  OAI22_X1 U13617 ( .A1(n14694), .A2(n11208), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7893), .ZN(n11121) );
  AOI211_X1 U13618 ( .C1(n14410), .C2(n14690), .A(n11122), .B(n11121), .ZN(
        n11123) );
  OAI21_X1 U13619 ( .B1(n11124), .B2(n12792), .A(n11123), .ZN(P2_U3206) );
  OAI211_X1 U13620 ( .C1(n11127), .C2(n11126), .A(n6547), .B(n11125), .ZN(
        n11135) );
  NAND2_X1 U13621 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12740)
         );
  OAI211_X1 U13622 ( .C1(n11130), .C2(n11129), .A(n11128), .B(n14725), .ZN(
        n11131) );
  NAND2_X1 U13623 ( .A1(n12740), .A2(n11131), .ZN(n11132) );
  AOI21_X1 U13624 ( .B1(n14720), .B2(n11133), .A(n11132), .ZN(n11134) );
  OAI211_X1 U13625 ( .C1(n14706), .C2(n15017), .A(n11135), .B(n11134), .ZN(
        P2_U3230) );
  INV_X1 U13626 ( .A(n11136), .ZN(n11139) );
  INV_X1 U13627 ( .A(SI_25_), .ZN(n11138) );
  OAI222_X1 U13628 ( .A1(n12609), .A2(n11139), .B1(n12606), .B2(n11138), .C1(
        n11137), .C2(P3_U3151), .ZN(P3_U3270) );
  INV_X1 U13629 ( .A(n11140), .ZN(n11142) );
  OAI21_X1 U13630 ( .B1(n11142), .B2(n6754), .A(n11141), .ZN(n14974) );
  OAI211_X1 U13631 ( .C1(n11145), .C2(n11144), .A(n11143), .B(n12450), .ZN(
        n11147) );
  AOI22_X1 U13632 ( .A1(n12453), .A2(n12455), .B1(n12134), .B2(n12456), .ZN(
        n11146) );
  NAND2_X1 U13633 ( .A1(n11147), .A2(n11146), .ZN(n14975) );
  NAND2_X1 U13634 ( .A1(n14975), .A2(n14946), .ZN(n11152) );
  OAI22_X1 U13635 ( .A1(n14946), .A2(n7022), .B1(n11148), .B2(n14934), .ZN(
        n11149) );
  AOI21_X1 U13636 ( .B1(n12470), .B2(n11150), .A(n11149), .ZN(n11151) );
  OAI211_X1 U13637 ( .C1(n14974), .C2(n12431), .A(n11152), .B(n11151), .ZN(
        P3_U3223) );
  XOR2_X1 U13638 ( .A(n11153), .B(n11154), .Z(n14422) );
  INV_X1 U13639 ( .A(n14422), .ZN(n14416) );
  AOI21_X1 U13640 ( .B1(n11155), .B2(n11154), .A(n13189), .ZN(n11159) );
  NAND2_X1 U13641 ( .A1(n12841), .A2(n12800), .ZN(n11157) );
  NAND2_X1 U13642 ( .A1(n12839), .A2(n12801), .ZN(n11156) );
  NAND2_X1 U13643 ( .A1(n11157), .A2(n11156), .ZN(n14686) );
  AOI21_X1 U13644 ( .B1(n11159), .B2(n11158), .A(n14686), .ZN(n14418) );
  INV_X1 U13645 ( .A(n14418), .ZN(n11165) );
  AOI21_X1 U13646 ( .B1(n11160), .B2(n14689), .A(n13104), .ZN(n11161) );
  NAND2_X1 U13647 ( .A1(n11161), .A2(n11212), .ZN(n14417) );
  OAI22_X1 U13648 ( .A1(n6558), .A2(n15207), .B1(n14693), .B2(n14751), .ZN(
        n11162) );
  AOI21_X1 U13649 ( .B1(n14689), .B2(n14393), .A(n11162), .ZN(n11163) );
  OAI21_X1 U13650 ( .B1(n14417), .B2(n13129), .A(n11163), .ZN(n11164) );
  AOI21_X1 U13651 ( .B1(n11165), .B2(n6558), .A(n11164), .ZN(n11166) );
  OAI21_X1 U13652 ( .B1(n13114), .B2(n14416), .A(n11166), .ZN(P2_U3253) );
  INV_X1 U13653 ( .A(n13431), .ZN(n11167) );
  NAND2_X1 U13654 ( .A1(n11168), .A2(n11167), .ZN(n11170) );
  OR2_X1 U13655 ( .A1(n14476), .A2(n13534), .ZN(n11169) );
  NAND2_X1 U13656 ( .A1(n11171), .A2(n13444), .ZN(n11174) );
  AOI22_X1 U13657 ( .A1(n11172), .A2(n6562), .B1(n13455), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11173) );
  NAND2_X2 U13658 ( .A1(n11174), .A2(n11173), .ZN(n14431) );
  INV_X1 U13659 ( .A(n13545), .ZN(n13436) );
  XNOR2_X1 U13660 ( .A(n11242), .B(n13436), .ZN(n14471) );
  AOI21_X1 U13661 ( .B1(n14431), .B2(n11175), .A(n6570), .ZN(n11176) );
  NAND2_X1 U13662 ( .A1(n11176), .A2(n11260), .ZN(n14466) );
  INV_X1 U13663 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11177) );
  NOR2_X1 U13664 ( .A1(n11248), .A2(n7537), .ZN(n13411) );
  NAND2_X1 U13665 ( .A1(n13411), .A2(n11731), .ZN(n11182) );
  NAND2_X1 U13666 ( .A1(n13448), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U13667 ( .A1(n10245), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U13668 ( .A1(n13449), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11179) );
  NAND4_X1 U13669 ( .A1(n11182), .A2(n11181), .A3(n11180), .A4(n11179), .ZN(
        n13681) );
  NAND2_X1 U13670 ( .A1(n13681), .A2(n13398), .ZN(n11184) );
  NAND2_X1 U13671 ( .A1(n13683), .A2(n13662), .ZN(n11183) );
  NAND2_X1 U13672 ( .A1(n11184), .A2(n11183), .ZN(n14434) );
  INV_X1 U13673 ( .A(n14434), .ZN(n14465) );
  OAI22_X1 U13674 ( .A1(n14575), .A2(n14465), .B1(n14437), .B2(n14010), .ZN(
        n11186) );
  INV_X1 U13675 ( .A(n14431), .ZN(n14467) );
  NOR2_X1 U13676 ( .A1(n14467), .A2(n14012), .ZN(n11185) );
  AOI211_X1 U13677 ( .C1(n14276), .C2(P1_REG2_REG_14__SCAN_IN), .A(n11186), 
        .B(n11185), .ZN(n11192) );
  NAND2_X1 U13678 ( .A1(n11187), .A2(n13431), .ZN(n11189) );
  OR2_X1 U13679 ( .A1(n14476), .A2(n13683), .ZN(n11188) );
  NAND2_X1 U13680 ( .A1(n11189), .A2(n11188), .ZN(n11190) );
  NAND2_X1 U13681 ( .A1(n13545), .A2(n11190), .ZN(n14468) );
  NAND3_X1 U13682 ( .A1(n11256), .A2(n14468), .A3(n13922), .ZN(n11191) );
  OAI211_X1 U13683 ( .C1(n14466), .C2(n14016), .A(n11192), .B(n11191), .ZN(
        n11193) );
  AOI21_X1 U13684 ( .B1(n14018), .B2(n14471), .A(n11193), .ZN(n11194) );
  INV_X1 U13685 ( .A(n11194), .ZN(P1_U3279) );
  OAI21_X1 U13686 ( .B1(n11196), .B2(n11586), .A(n11195), .ZN(n14962) );
  INV_X1 U13687 ( .A(n12038), .ZN(n11197) );
  OAI22_X1 U13688 ( .A1(n12428), .A2(n14959), .B1(n11197), .B2(n14934), .ZN(
        n11205) );
  NAND2_X1 U13689 ( .A1(n11199), .A2(n11586), .ZN(n11200) );
  NAND2_X1 U13690 ( .A1(n11198), .A2(n11200), .ZN(n11201) );
  NAND2_X1 U13691 ( .A1(n11201), .A2(n12450), .ZN(n11203) );
  AOI22_X1 U13692 ( .A1(n12456), .A2(n12037), .B1(n12134), .B2(n12453), .ZN(
        n11202) );
  NAND2_X1 U13693 ( .A1(n11203), .A2(n11202), .ZN(n14960) );
  MUX2_X1 U13694 ( .A(n14960), .B(P3_REG2_REG_8__SCAN_IN), .S(n14949), .Z(
        n11204) );
  AOI211_X1 U13695 ( .C1(n12471), .C2(n14962), .A(n11205), .B(n11204), .ZN(
        n11206) );
  INV_X1 U13696 ( .A(n11206), .ZN(P3_U3225) );
  XOR2_X1 U13697 ( .A(n11207), .B(n11216), .Z(n14413) );
  INV_X1 U13698 ( .A(n11208), .ZN(n11209) );
  AOI22_X1 U13699 ( .A1(n14736), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11209), 
        .B2(n14734), .ZN(n11210) );
  OAI21_X1 U13700 ( .B1(n11211), .B2(n14736), .A(n11210), .ZN(n11215) );
  NAND2_X1 U13701 ( .A1(n14410), .A2(n11212), .ZN(n11213) );
  NAND3_X1 U13702 ( .A1(n14397), .A2(n10011), .A3(n11213), .ZN(n14411) );
  NOR2_X1 U13703 ( .A1(n14411), .A2(n13129), .ZN(n11214) );
  AOI211_X1 U13704 ( .C1(n14393), .C2(n14410), .A(n11215), .B(n11214), .ZN(
        n11219) );
  XNOR2_X1 U13705 ( .A(n11217), .B(n11216), .ZN(n14415) );
  NAND2_X1 U13706 ( .A1(n14415), .A2(n13131), .ZN(n11218) );
  OAI211_X1 U13707 ( .C1(n14413), .C2(n13114), .A(n11219), .B(n11218), .ZN(
        P2_U3252) );
  INV_X1 U13708 ( .A(n11685), .ZN(n11222) );
  OAI222_X1 U13709 ( .A1(n13269), .A2(n11221), .B1(n13272), .B2(n11222), .C1(
        P2_U3088), .C2(n11220), .ZN(P2_U3306) );
  OAI222_X1 U13710 ( .A1(n14145), .A2(n11223), .B1(n14148), .B2(n11222), .C1(
        P1_U3086), .C2(n13464), .ZN(P1_U3334) );
  XNOR2_X1 U13711 ( .A(n11032), .B(n11233), .ZN(n11278) );
  XNOR2_X1 U13712 ( .A(n11278), .B(n12437), .ZN(n11229) );
  NOR2_X1 U13713 ( .A1(n11224), .A2(n12455), .ZN(n11226) );
  INV_X1 U13714 ( .A(n11224), .ZN(n11225) );
  AOI21_X1 U13715 ( .B1(n11229), .B2(n11228), .A(n6717), .ZN(n11236) );
  NOR2_X1 U13716 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11230), .ZN(n14858) );
  OAI22_X1 U13717 ( .A1(n12112), .A2(n11231), .B1(n11964), .B2(n12120), .ZN(
        n11232) );
  AOI211_X1 U13718 ( .C1(n11233), .C2(n6545), .A(n14858), .B(n11232), .ZN(
        n11235) );
  NAND2_X1 U13719 ( .A1(n12124), .A2(n12460), .ZN(n11234) );
  OAI211_X1 U13720 ( .C1(n11236), .C2(n12126), .A(n11235), .B(n11234), .ZN(
        P3_U3164) );
  INV_X1 U13721 ( .A(n11237), .ZN(n11239) );
  OAI222_X1 U13722 ( .A1(P3_U3151), .A2(n11240), .B1(n12609), .B2(n11239), 
        .C1(n11238), .C2(n12606), .ZN(P3_U3269) );
  INV_X1 U13723 ( .A(n13682), .ZN(n13538) );
  OR2_X1 U13724 ( .A1(n14431), .A2(n13538), .ZN(n13537) );
  INV_X1 U13725 ( .A(n13537), .ZN(n11241) );
  AOI21_X2 U13726 ( .B1(n11242), .B2(n13545), .A(n11241), .ZN(n11294) );
  NAND2_X1 U13727 ( .A1(n11243), .A2(n13444), .ZN(n11246) );
  AOI22_X1 U13728 ( .A1(n13455), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6562), 
        .B2(n11244), .ZN(n11245) );
  INV_X1 U13729 ( .A(n13681), .ZN(n11838) );
  NAND2_X1 U13730 ( .A1(n11837), .A2(n11838), .ZN(n13550) );
  NAND2_X1 U13731 ( .A1(n13549), .A2(n13550), .ZN(n13433) );
  XNOR2_X1 U13732 ( .A(n11294), .B(n11258), .ZN(n11247) );
  NAND2_X1 U13733 ( .A1(n11247), .A2(n14571), .ZN(n11254) );
  NAND2_X1 U13734 ( .A1(n11248), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11300) );
  OR2_X1 U13735 ( .A1(n11248), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U13736 ( .A1(n11300), .A2(n11249), .ZN(n13333) );
  NAND2_X1 U13737 ( .A1(n13448), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11251) );
  NAND2_X1 U13738 ( .A1(n10245), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11250) );
  AND2_X1 U13739 ( .A1(n11251), .A2(n11250), .ZN(n11253) );
  NAND2_X1 U13740 ( .A1(n13449), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11252) );
  OAI211_X1 U13741 ( .C1(n11769), .C2(n13333), .A(n11253), .B(n11252), .ZN(
        n13680) );
  AOI22_X1 U13742 ( .A1(n13680), .A2(n13398), .B1(n13682), .B2(n13662), .ZN(
        n13408) );
  NAND2_X1 U13743 ( .A1(n11254), .A2(n13408), .ZN(n14115) );
  INV_X1 U13744 ( .A(n14115), .ZN(n11266) );
  NAND2_X1 U13745 ( .A1(n14431), .A2(n13682), .ZN(n11255) );
  NAND2_X1 U13746 ( .A1(n11258), .A2(n11257), .ZN(n11259) );
  NAND2_X1 U13747 ( .A1(n11310), .A2(n11259), .ZN(n14111) );
  AOI21_X1 U13748 ( .B1(n11837), .B2(n11260), .A(n6570), .ZN(n11261) );
  NAND2_X1 U13749 ( .A1(n11261), .A2(n11296), .ZN(n14112) );
  AOI22_X1 U13750 ( .A1(n14276), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13411), 
        .B2(n14574), .ZN(n11263) );
  NAND2_X1 U13751 ( .A1(n11837), .A2(n14572), .ZN(n11262) );
  OAI211_X1 U13752 ( .C1(n14112), .C2(n14016), .A(n11263), .B(n11262), .ZN(
        n11264) );
  AOI21_X1 U13753 ( .B1(n14111), .B2(n13922), .A(n11264), .ZN(n11265) );
  OAI21_X1 U13754 ( .B1(n11266), .B2(n14575), .A(n11265), .ZN(P1_U3278) );
  XNOR2_X1 U13755 ( .A(n11377), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n11375) );
  OAI21_X1 U13756 ( .B1(n11269), .B2(n11268), .A(n11267), .ZN(n11374) );
  XNOR2_X1 U13757 ( .A(n11375), .B(n11374), .ZN(n11277) );
  NAND2_X1 U13758 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13343)
         );
  INV_X1 U13759 ( .A(n11270), .ZN(n11271) );
  AOI21_X1 U13760 ( .B1(n11291), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11271), 
        .ZN(n11379) );
  XNOR2_X1 U13761 ( .A(n11690), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11380) );
  XOR2_X1 U13762 ( .A(n11379), .B(n11380), .Z(n11272) );
  NAND2_X1 U13763 ( .A1(n13819), .A2(n11272), .ZN(n11273) );
  NAND2_X1 U13764 ( .A1(n13343), .A2(n11273), .ZN(n11275) );
  NOR2_X1 U13765 ( .A1(n6779), .A2(n11377), .ZN(n11274) );
  AOI211_X1 U13766 ( .C1(n14525), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n11275), 
        .B(n11274), .ZN(n11276) );
  OAI21_X1 U13767 ( .B1(n11277), .B2(n14534), .A(n11276), .ZN(P1_U3260) );
  INV_X1 U13768 ( .A(n11278), .ZN(n11279) );
  XNOR2_X1 U13769 ( .A(n12596), .B(n11032), .ZN(n11963) );
  XNOR2_X1 U13770 ( .A(n11963), .B(n12454), .ZN(n11280) );
  OAI211_X1 U13771 ( .C1(n11281), .C2(n11280), .A(n11962), .B(n12058), .ZN(
        n11286) );
  NOR2_X1 U13772 ( .A1(n12121), .A2(n12596), .ZN(n11284) );
  NAND2_X1 U13773 ( .A1(n12118), .A2(n12437), .ZN(n11282) );
  NAND2_X1 U13774 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n14876)
         );
  OAI211_X1 U13775 ( .C1(n12120), .C2(n12409), .A(n11282), .B(n14876), .ZN(
        n11283) );
  AOI211_X1 U13776 ( .C1(n12440), .C2(n12124), .A(n11284), .B(n11283), .ZN(
        n11285) );
  NAND2_X1 U13777 ( .A1(n11286), .A2(n11285), .ZN(P3_U3174) );
  INV_X1 U13778 ( .A(n11287), .ZN(n11289) );
  OAI222_X1 U13779 ( .A1(n13269), .A2(n15202), .B1(n13272), .B2(n11289), .C1(
        P2_U3088), .C2(n11288), .ZN(P2_U3305) );
  NAND2_X1 U13780 ( .A1(n11290), .A2(n13444), .ZN(n11293) );
  AOI22_X1 U13781 ( .A1(n13455), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11291), 
        .B2(n6562), .ZN(n11292) );
  INV_X1 U13782 ( .A(n13680), .ZN(n13341) );
  XNOR2_X1 U13783 ( .A(n14106), .B(n13341), .ZN(n13432) );
  AOI21_X1 U13784 ( .B1(n13432), .B2(n11295), .A(n6705), .ZN(n14110) );
  NAND2_X1 U13785 ( .A1(n11296), .A2(n14106), .ZN(n11297) );
  NAND2_X1 U13786 ( .A1(n11297), .A2(n14577), .ZN(n11298) );
  NOR2_X1 U13787 ( .A1(n14008), .A2(n11298), .ZN(n14104) );
  INV_X1 U13788 ( .A(n14106), .ZN(n11688) );
  INV_X1 U13789 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U13790 ( .A1(n11300), .A2(n11299), .ZN(n11301) );
  NAND2_X1 U13791 ( .A1(n11697), .A2(n11301), .ZN(n14011) );
  AOI22_X1 U13792 ( .A1(n13448), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10245), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U13793 ( .A1(n13449), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11302) );
  OAI211_X1 U13794 ( .C1(n14011), .C2(n11769), .A(n11303), .B(n11302), .ZN(
        n13679) );
  NAND2_X1 U13795 ( .A1(n13679), .A2(n13398), .ZN(n11305) );
  NAND2_X1 U13796 ( .A1(n13681), .A2(n13662), .ZN(n11304) );
  NAND2_X1 U13797 ( .A1(n11305), .A2(n11304), .ZN(n14105) );
  INV_X1 U13798 ( .A(n14105), .ZN(n11306) );
  OAI22_X1 U13799 ( .A1(n14575), .A2(n11306), .B1(n13333), .B2(n14010), .ZN(
        n11307) );
  AOI21_X1 U13800 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14276), .A(n11307), 
        .ZN(n11308) );
  OAI21_X1 U13801 ( .B1(n11688), .B2(n14012), .A(n11308), .ZN(n11309) );
  AOI21_X1 U13802 ( .B1(n14104), .B2(n14581), .A(n11309), .ZN(n11312) );
  XNOR2_X1 U13803 ( .A(n11790), .B(n13432), .ZN(n14107) );
  NAND2_X1 U13804 ( .A1(n14107), .A2(n13922), .ZN(n11311) );
  OAI211_X1 U13805 ( .C1(n14110), .C2(n13924), .A(n11312), .B(n11311), .ZN(
        P1_U3277) );
  INV_X1 U13806 ( .A(n11313), .ZN(n11314) );
  AOI21_X1 U13807 ( .B1(n11481), .B2(n11315), .A(n11314), .ZN(n11316) );
  OAI222_X1 U13808 ( .A1(n14943), .A2(n11318), .B1(n14941), .B2(n11317), .C1(
        n14939), .C2(n11316), .ZN(n14369) );
  INV_X1 U13809 ( .A(n14369), .ZN(n11325) );
  OAI21_X1 U13810 ( .B1(n6716), .B2(n11481), .A(n11319), .ZN(n14371) );
  INV_X1 U13811 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11322) );
  NOR2_X1 U13812 ( .A1(n11486), .A2(n14971), .ZN(n14370) );
  AOI22_X1 U13813 ( .A1(n12461), .A2(n14370), .B1(n12468), .B2(n11320), .ZN(
        n11321) );
  OAI21_X1 U13814 ( .B1(n11322), .B2(n14946), .A(n11321), .ZN(n11323) );
  AOI21_X1 U13815 ( .B1(n14371), .B2(n12471), .A(n11323), .ZN(n11324) );
  OAI21_X1 U13816 ( .B1(n11325), .B2(n14949), .A(n11324), .ZN(P3_U3222) );
  INV_X1 U13817 ( .A(n14274), .ZN(n14284) );
  AOI22_X1 U13818 ( .A1(n14450), .A2(n11931), .B1(n6565), .B2(n13685), .ZN(
        n11344) );
  NAND2_X1 U13819 ( .A1(n14450), .A2(n11930), .ZN(n11327) );
  NAND2_X1 U13820 ( .A1(n11931), .A2(n13685), .ZN(n11326) );
  NAND2_X1 U13821 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  XNOR2_X1 U13822 ( .A(n11328), .B(n11941), .ZN(n11342) );
  INV_X1 U13823 ( .A(n11342), .ZN(n11343) );
  NOR2_X1 U13824 ( .A1(n9739), .A2(n11334), .ZN(n11335) );
  AOI21_X1 U13825 ( .B1(n14653), .B2(n11931), .A(n11335), .ZN(n11338) );
  AOI22_X1 U13826 ( .A1(n14653), .A2(n11930), .B1(n11931), .B2(n13686), .ZN(
        n11336) );
  XNOR2_X1 U13827 ( .A(n11336), .B(n11941), .ZN(n11337) );
  XOR2_X1 U13828 ( .A(n11338), .B(n11337), .Z(n14442) );
  INV_X1 U13829 ( .A(n11337), .ZN(n11340) );
  INV_X1 U13830 ( .A(n11338), .ZN(n11339) );
  NAND2_X1 U13831 ( .A1(n11340), .A2(n11339), .ZN(n11341) );
  XOR2_X1 U13832 ( .A(n11344), .B(n11342), .Z(n14455) );
  NAND2_X1 U13833 ( .A1(n14274), .A2(n11930), .ZN(n11346) );
  NAND2_X1 U13834 ( .A1(n11931), .A2(n13684), .ZN(n11345) );
  NAND2_X1 U13835 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  XNOR2_X1 U13836 ( .A(n11347), .B(n11941), .ZN(n11815) );
  NOR2_X1 U13837 ( .A1(n9739), .A2(n11348), .ZN(n11349) );
  AOI21_X1 U13838 ( .B1(n14274), .B2(n11931), .A(n11349), .ZN(n11816) );
  XNOR2_X1 U13839 ( .A(n11815), .B(n11816), .ZN(n11350) );
  OAI211_X1 U13840 ( .C1(n6708), .C2(n11350), .A(n11819), .B(n14440), .ZN(
        n11356) );
  INV_X1 U13841 ( .A(n11351), .ZN(n14273) );
  NAND2_X1 U13842 ( .A1(n13685), .A2(n13662), .ZN(n11353) );
  NAND2_X1 U13843 ( .A1(n13683), .A2(n13398), .ZN(n11352) );
  AND2_X1 U13844 ( .A1(n11353), .A2(n11352), .ZN(n14270) );
  OAI22_X1 U13845 ( .A1(n14456), .A2(n14270), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15137), .ZN(n11354) );
  AOI21_X1 U13846 ( .B1(n14273), .B2(n13410), .A(n11354), .ZN(n11355) );
  OAI211_X1 U13847 ( .C1(n14284), .C2(n13414), .A(n11356), .B(n11355), .ZN(
        P1_U3224) );
  XOR2_X1 U13848 ( .A(n11357), .B(n11364), .Z(n13232) );
  AOI21_X1 U13849 ( .B1(n13228), .B2(n14398), .A(n12664), .ZN(n11358) );
  AND2_X1 U13850 ( .A1(n11358), .A2(n6700), .ZN(n13226) );
  OAI22_X1 U13851 ( .A1(n12749), .A2(n14754), .B1(n11359), .B2(n14378), .ZN(
        n13227) );
  OAI22_X1 U13852 ( .A1(n6558), .A2(n11360), .B1(n12817), .B2(n14751), .ZN(
        n11361) );
  AOI21_X1 U13853 ( .B1(n13227), .B2(n6558), .A(n11361), .ZN(n11362) );
  OAI21_X1 U13854 ( .B1(n7146), .B2(n14739), .A(n11362), .ZN(n11363) );
  AOI21_X1 U13855 ( .B1(n14731), .B2(n13226), .A(n11363), .ZN(n11367) );
  NAND2_X1 U13856 ( .A1(n11365), .A2(n11364), .ZN(n13229) );
  NAND3_X1 U13857 ( .A1(n6699), .A2(n13131), .A3(n13229), .ZN(n11366) );
  OAI211_X1 U13858 ( .C1(n13232), .C2(n13114), .A(n11367), .B(n11366), .ZN(
        P2_U3250) );
  INV_X1 U13859 ( .A(n11726), .ZN(n11370) );
  AOI21_X1 U13860 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n14136), .A(n11368), 
        .ZN(n11369) );
  OAI21_X1 U13861 ( .B1(n11370), .B2(n14148), .A(n11369), .ZN(P1_U3332) );
  NAND2_X1 U13862 ( .A1(n11726), .A2(n13260), .ZN(n11372) );
  OAI211_X1 U13863 ( .C1(n11373), .C2(n13269), .A(n11372), .B(n11371), .ZN(
        P2_U3304) );
  AOI22_X1 U13864 ( .A1(n11375), .A2(n11374), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n11690), .ZN(n13802) );
  XNOR2_X1 U13865 ( .A(n13802), .B(n13808), .ZN(n11376) );
  NAND2_X1 U13866 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11376), .ZN(n13805) );
  OAI211_X1 U13867 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11376), .A(n13813), 
        .B(n13805), .ZN(n11385) );
  NAND2_X1 U13868 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13389)
         );
  INV_X1 U13869 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11378) );
  XNOR2_X1 U13870 ( .A(n11386), .B(n13807), .ZN(n11381) );
  NAND2_X1 U13871 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11381), .ZN(n13810) );
  OAI211_X1 U13872 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11381), .A(n13819), 
        .B(n13810), .ZN(n11382) );
  NAND2_X1 U13873 ( .A1(n13389), .A2(n11382), .ZN(n11383) );
  AOI21_X1 U13874 ( .B1(n14525), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11383), 
        .ZN(n11384) );
  OAI211_X1 U13875 ( .C1(n6779), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        P1_U3261) );
  INV_X1 U13876 ( .A(n11661), .ZN(n11953) );
  OAI222_X1 U13877 ( .A1(n13269), .A2(n11388), .B1(n13272), .B2(n11953), .C1(
        P2_U3088), .C2(n11387), .ZN(P2_U3303) );
  INV_X1 U13878 ( .A(n13261), .ZN(n11389) );
  OAI222_X1 U13879 ( .A1(n14145), .A2(n11390), .B1(n14148), .B2(n11389), .C1(
        P1_U3086), .C2(n9233), .ZN(P1_U3327) );
  INV_X1 U13880 ( .A(n11392), .ZN(n11393) );
  NAND2_X1 U13881 ( .A1(n11394), .A2(n11393), .ZN(n11396) );
  NAND2_X1 U13882 ( .A1(n14141), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11395) );
  XNOR2_X1 U13883 ( .A(n13256), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11407) );
  INV_X1 U13884 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11807) );
  XNOR2_X1 U13885 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11397) );
  XNOR2_X1 U13886 ( .A(n11398), .B(n11397), .ZN(n12603) );
  NAND2_X1 U13887 ( .A1(n12603), .A2(n11409), .ZN(n11400) );
  INV_X1 U13888 ( .A(SI_31_), .ZN(n12599) );
  OR2_X1 U13889 ( .A1(n11411), .A2(n12599), .ZN(n11399) );
  NAND2_X1 U13890 ( .A1(n8711), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11404) );
  NAND2_X1 U13891 ( .A1(n8819), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11403) );
  NAND2_X1 U13892 ( .A1(n11401), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11402) );
  AND3_X1 U13893 ( .A1(n11404), .A2(n11403), .A3(n11402), .ZN(n11405) );
  XNOR2_X1 U13894 ( .A(n11408), .B(n11407), .ZN(n11811) );
  NAND2_X1 U13895 ( .A1(n11811), .A2(n11409), .ZN(n11413) );
  INV_X1 U13896 ( .A(SI_30_), .ZN(n11410) );
  OR2_X1 U13897 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  NAND2_X1 U13898 ( .A1(n11415), .A2(n11417), .ZN(n11414) );
  INV_X1 U13899 ( .A(n12243), .ZN(n12128) );
  OAI21_X1 U13900 ( .B1(n14364), .B2(n12128), .A(n11572), .ZN(n11416) );
  NOR2_X1 U13901 ( .A1(n11608), .A2(n11416), .ZN(n11420) );
  INV_X1 U13902 ( .A(n11417), .ZN(n12129) );
  XNOR2_X1 U13903 ( .A(n11422), .B(n12237), .ZN(n11617) );
  INV_X1 U13904 ( .A(n11423), .ZN(n11556) );
  INV_X1 U13905 ( .A(n11424), .ZN(n11425) );
  MUX2_X1 U13906 ( .A(n11426), .B(n11425), .S(n11569), .Z(n11427) );
  NOR2_X1 U13907 ( .A1(n12275), .A2(n11427), .ZN(n11560) );
  NAND2_X1 U13908 ( .A1(n11429), .A2(n11619), .ZN(n11432) );
  NAND2_X1 U13909 ( .A1(n11429), .A2(n11428), .ZN(n11430) );
  NAND3_X1 U13910 ( .A1(n11437), .A2(n11430), .A3(n11577), .ZN(n11431) );
  OAI21_X1 U13911 ( .B1(n14937), .B2(n11432), .A(n11431), .ZN(n11435) );
  NAND2_X1 U13912 ( .A1(n14930), .A2(n11433), .ZN(n11434) );
  AOI21_X1 U13913 ( .B1(n11435), .B2(n11434), .A(n11591), .ZN(n11444) );
  MUX2_X1 U13914 ( .A(n11437), .B(n11436), .S(n11577), .Z(n11443) );
  NAND2_X1 U13915 ( .A1(n11446), .A2(n11438), .ZN(n11441) );
  NAND2_X1 U13916 ( .A1(n11445), .A2(n11439), .ZN(n11440) );
  MUX2_X1 U13917 ( .A(n11441), .B(n11440), .S(n11569), .Z(n11442) );
  AOI21_X1 U13918 ( .B1(n11444), .B2(n11443), .A(n11442), .ZN(n11453) );
  MUX2_X1 U13919 ( .A(n11446), .B(n11445), .S(n11577), .Z(n11448) );
  NAND2_X1 U13920 ( .A1(n11448), .A2(n11447), .ZN(n11452) );
  MUX2_X1 U13921 ( .A(n11450), .B(n11449), .S(n11569), .Z(n11451) );
  OAI211_X1 U13922 ( .C1(n11453), .C2(n11452), .A(n11588), .B(n11451), .ZN(
        n11457) );
  NAND2_X1 U13923 ( .A1(n11462), .A2(n11454), .ZN(n11455) );
  NAND2_X1 U13924 ( .A1(n11455), .A2(n11569), .ZN(n11456) );
  NAND2_X1 U13925 ( .A1(n11457), .A2(n11456), .ZN(n11461) );
  AOI21_X1 U13926 ( .B1(n11460), .B2(n11458), .A(n11569), .ZN(n11459) );
  AOI21_X1 U13927 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n11467) );
  OAI21_X1 U13928 ( .B1(n11569), .B2(n11462), .A(n11589), .ZN(n11466) );
  MUX2_X1 U13929 ( .A(n11464), .B(n11463), .S(n11577), .Z(n11465) );
  OAI211_X1 U13930 ( .C1(n11467), .C2(n11466), .A(n11586), .B(n11465), .ZN(
        n11472) );
  INV_X1 U13931 ( .A(n11468), .ZN(n11596) );
  MUX2_X1 U13932 ( .A(n11470), .B(n11469), .S(n11569), .Z(n11471) );
  NAND3_X1 U13933 ( .A1(n11472), .A2(n11596), .A3(n11471), .ZN(n11478) );
  NAND2_X1 U13934 ( .A1(n11473), .A2(n11569), .ZN(n11476) );
  NAND2_X1 U13935 ( .A1(n12134), .A2(n11577), .ZN(n11475) );
  MUX2_X1 U13936 ( .A(n11476), .B(n11475), .S(n11474), .Z(n11477) );
  NAND2_X1 U13937 ( .A1(n11478), .A2(n11477), .ZN(n11484) );
  MUX2_X1 U13938 ( .A(n11480), .B(n11479), .S(n11569), .Z(n11482) );
  NAND2_X1 U13939 ( .A1(n11482), .A2(n11481), .ZN(n11483) );
  AOI21_X1 U13940 ( .B1(n11484), .B2(n6754), .A(n11483), .ZN(n11494) );
  NAND2_X1 U13941 ( .A1(n11491), .A2(n11485), .ZN(n11489) );
  NAND2_X1 U13942 ( .A1(n12455), .A2(n11486), .ZN(n11487) );
  NAND2_X1 U13943 ( .A1(n11490), .A2(n11487), .ZN(n11488) );
  MUX2_X1 U13944 ( .A(n11489), .B(n11488), .S(n11569), .Z(n11493) );
  INV_X1 U13945 ( .A(n12434), .ZN(n12444) );
  MUX2_X1 U13946 ( .A(n11491), .B(n11490), .S(n11577), .Z(n11492) );
  OAI211_X1 U13947 ( .C1(n11494), .C2(n11493), .A(n12444), .B(n11492), .ZN(
        n11499) );
  INV_X1 U13948 ( .A(n12421), .ZN(n11495) );
  AND2_X1 U13949 ( .A1(n12412), .A2(n11495), .ZN(n11600) );
  MUX2_X1 U13950 ( .A(n11497), .B(n11496), .S(n11569), .Z(n11498) );
  NAND3_X1 U13951 ( .A1(n11499), .A2(n11600), .A3(n11498), .ZN(n11506) );
  INV_X1 U13952 ( .A(n11500), .ZN(n11501) );
  NAND2_X1 U13953 ( .A1(n12412), .A2(n11501), .ZN(n11503) );
  NAND3_X1 U13954 ( .A1(n11503), .A2(n11502), .A3(n11513), .ZN(n11504) );
  NAND2_X1 U13955 ( .A1(n11504), .A2(n11577), .ZN(n11505) );
  AOI21_X1 U13956 ( .B1(n11506), .B2(n11505), .A(n7032), .ZN(n11515) );
  INV_X1 U13957 ( .A(n11507), .ZN(n11510) );
  INV_X1 U13958 ( .A(n11508), .ZN(n11509) );
  AOI21_X1 U13959 ( .B1(n12412), .B2(n11510), .A(n11509), .ZN(n11512) );
  AOI21_X1 U13960 ( .B1(n11512), .B2(n11511), .A(n11577), .ZN(n11514) );
  OAI22_X1 U13961 ( .A1(n11515), .A2(n11514), .B1(n11577), .B2(n11513), .ZN(
        n11529) );
  NOR2_X1 U13962 ( .A1(n12373), .A2(n7034), .ZN(n11528) );
  INV_X1 U13963 ( .A(n11516), .ZN(n11520) );
  INV_X1 U13964 ( .A(n11517), .ZN(n11518) );
  AND2_X1 U13965 ( .A1(n11523), .A2(n11518), .ZN(n11519) );
  OR3_X1 U13966 ( .A1(n11521), .A2(n11520), .A3(n11519), .ZN(n11526) );
  OAI211_X1 U13967 ( .C1(n12373), .C2(n11524), .A(n11523), .B(n11522), .ZN(
        n11525) );
  MUX2_X1 U13968 ( .A(n11526), .B(n11525), .S(n11577), .Z(n11527) );
  AOI21_X1 U13969 ( .B1(n11529), .B2(n11528), .A(n11527), .ZN(n11533) );
  INV_X1 U13970 ( .A(n11584), .ZN(n11531) );
  MUX2_X1 U13971 ( .A(n12370), .B(n12572), .S(n11569), .Z(n11530) );
  NOR2_X1 U13972 ( .A1(n11531), .A2(n11530), .ZN(n11532) );
  OR3_X1 U13973 ( .A1(n11533), .A2(n12351), .A3(n11532), .ZN(n11537) );
  XNOR2_X1 U13974 ( .A(n12338), .B(n12345), .ZN(n12337) );
  NAND2_X1 U13975 ( .A1(n12509), .A2(n12360), .ZN(n11535) );
  MUX2_X1 U13976 ( .A(n11535), .B(n11534), .S(n11569), .Z(n11536) );
  NAND3_X1 U13977 ( .A1(n11537), .A2(n12337), .A3(n11536), .ZN(n11541) );
  MUX2_X1 U13978 ( .A(n11539), .B(n11538), .S(n11577), .Z(n11540) );
  NAND3_X1 U13979 ( .A1(n11541), .A2(n12326), .A3(n11540), .ZN(n11545) );
  MUX2_X1 U13980 ( .A(n11543), .B(n11542), .S(n11569), .Z(n11544) );
  NAND3_X1 U13981 ( .A1(n11545), .A2(n12316), .A3(n11544), .ZN(n11547) );
  NAND3_X1 U13982 ( .A1(n12496), .A2(n12324), .A3(n11569), .ZN(n11546) );
  AND2_X1 U13983 ( .A1(n11547), .A2(n11546), .ZN(n11555) );
  INV_X1 U13984 ( .A(n11548), .ZN(n11549) );
  NAND2_X1 U13985 ( .A1(n11553), .A2(n11549), .ZN(n11551) );
  AND2_X1 U13986 ( .A1(n11551), .A2(n11550), .ZN(n11552) );
  MUX2_X1 U13987 ( .A(n11553), .B(n11552), .S(n11577), .Z(n11554) );
  OAI211_X1 U13988 ( .C1(n11555), .C2(n12303), .A(n11554), .B(n12291), .ZN(
        n11559) );
  MUX2_X1 U13989 ( .A(n11557), .B(n11556), .S(n11569), .Z(n11558) );
  AOI21_X1 U13990 ( .B1(n11560), .B2(n11559), .A(n11558), .ZN(n11562) );
  NAND2_X1 U13991 ( .A1(n12130), .A2(n11577), .ZN(n11561) );
  OAI22_X1 U13992 ( .A1(n11562), .A2(n8717), .B1(n12477), .B2(n11561), .ZN(
        n11564) );
  INV_X1 U13993 ( .A(n11563), .ZN(n12021) );
  NAND2_X1 U13994 ( .A1(n11564), .A2(n12021), .ZN(n11571) );
  NAND2_X1 U13995 ( .A1(n11566), .A2(n11565), .ZN(n11568) );
  INV_X1 U13996 ( .A(n11576), .ZN(n11573) );
  NAND2_X1 U13997 ( .A1(n11573), .A2(n11572), .ZN(n11579) );
  INV_X1 U13998 ( .A(n11574), .ZN(n11575) );
  NOR2_X1 U13999 ( .A1(n11576), .A2(n11575), .ZN(n11578) );
  INV_X1 U14000 ( .A(n11614), .ZN(n11581) );
  INV_X1 U14001 ( .A(n12291), .ZN(n11604) );
  INV_X1 U14002 ( .A(n11583), .ZN(n11585) );
  NAND4_X1 U14003 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11592) );
  NOR4_X1 U14004 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n14937), .ZN(
        n11593) );
  NAND2_X1 U14005 ( .A1(n11593), .A2(n12449), .ZN(n11598) );
  NAND4_X1 U14006 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n6754), .ZN(
        n11597) );
  NOR4_X1 U14007 ( .A1(n11598), .A2(n8444), .A3(n12434), .A4(n11597), .ZN(
        n11599) );
  NAND4_X1 U14008 ( .A1(n12400), .A2(n12391), .A3(n11600), .A4(n11599), .ZN(
        n11601) );
  NOR4_X1 U14009 ( .A1(n12351), .A2(n12361), .A3(n12373), .A4(n11601), .ZN(
        n11602) );
  NAND4_X1 U14010 ( .A1(n12316), .A2(n12326), .A3(n11602), .A4(n12337), .ZN(
        n11603) );
  NOR4_X1 U14011 ( .A1(n12275), .A2(n11604), .A3(n12303), .A4(n11603), .ZN(
        n11606) );
  XNOR2_X1 U14012 ( .A(n11610), .B(n12222), .ZN(n11612) );
  OAI22_X1 U14013 ( .A1(n11614), .A2(n11613), .B1(n11612), .B2(n11611), .ZN(
        n11615) );
  NOR3_X1 U14014 ( .A1(n11618), .A2(n12223), .A3(n6831), .ZN(n11621) );
  OAI21_X1 U14015 ( .B1(n11622), .B2(n11619), .A(P3_B_REG_SCAN_IN), .ZN(n11620) );
  INV_X1 U14016 ( .A(n11653), .ZN(n13271) );
  OAI222_X1 U14017 ( .A1(n14145), .A2(n11624), .B1(n14148), .B2(n13271), .C1(
        P1_U3086), .C2(n9320), .ZN(P1_U3330) );
  INV_X1 U14018 ( .A(n11625), .ZN(n11628) );
  OAI222_X1 U14019 ( .A1(n12609), .A2(n11628), .B1(P3_U3151), .B2(n11627), 
        .C1(n11626), .C2(n12606), .ZN(P3_U3266) );
  NAND2_X1 U14020 ( .A1(n11630), .A2(n11629), .ZN(n11631) );
  XOR2_X1 U14021 ( .A(n11639), .B(n11631), .Z(n12945) );
  NOR2_X1 U14022 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12945), .ZN(n12944) );
  NOR2_X1 U14023 ( .A1(n12949), .A2(n11631), .ZN(n11632) );
  NOR2_X1 U14024 ( .A1(n12944), .A2(n11632), .ZN(n11633) );
  XOR2_X1 U14025 ( .A(n11633), .B(P2_REG2_REG_19__SCAN_IN), .Z(n11648) );
  INV_X1 U14026 ( .A(n11648), .ZN(n11646) );
  NAND2_X1 U14027 ( .A1(n11635), .A2(n11634), .ZN(n11638) );
  NAND2_X1 U14028 ( .A1(n11636), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n11637) );
  NAND2_X1 U14029 ( .A1(n11638), .A2(n11637), .ZN(n11640) );
  XNOR2_X1 U14030 ( .A(n11640), .B(n11639), .ZN(n12951) );
  NAND2_X1 U14031 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n12951), .ZN(n12950) );
  NAND2_X1 U14032 ( .A1(n12949), .A2(n11640), .ZN(n11641) );
  NAND2_X1 U14033 ( .A1(n12950), .A2(n11641), .ZN(n11643) );
  XNOR2_X1 U14034 ( .A(n11643), .B(n11642), .ZN(n11647) );
  OAI21_X1 U14035 ( .B1(n11647), .B2(n11644), .A(n12925), .ZN(n11645) );
  AOI21_X1 U14036 ( .B1(n11646), .B2(n6547), .A(n11645), .ZN(n11650) );
  AOI22_X1 U14037 ( .A1(n11648), .A2(n6547), .B1(n14725), .B2(n11647), .ZN(
        n11649) );
  MUX2_X1 U14038 ( .A(n11650), .B(n11649), .S(n14748), .Z(n11651) );
  NAND2_X1 U14039 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12696)
         );
  OAI211_X1 U14040 ( .C1(n11652), .C2(n14706), .A(n11651), .B(n12696), .ZN(
        P2_U3233) );
  NAND2_X1 U14041 ( .A1(n11653), .A2(n13444), .ZN(n11655) );
  NAND2_X1 U14042 ( .A1(n13455), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11654) );
  INV_X1 U14043 ( .A(n14051), .ZN(n13886) );
  NAND2_X1 U14044 ( .A1(n13448), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11660) );
  INV_X1 U14045 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11696) );
  INV_X1 U14046 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U14047 ( .A1(n11729), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11664) );
  INV_X1 U14048 ( .A(n11664), .ZN(n11656) );
  NAND2_X1 U14049 ( .A1(n11656), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11739) );
  OAI21_X1 U14050 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11656), .A(n11739), 
        .ZN(n13882) );
  OR2_X1 U14051 ( .A1(n11769), .A2(n13882), .ZN(n11659) );
  NAND2_X1 U14052 ( .A1(n10245), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U14053 ( .A1(n13449), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14054 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n13672) );
  NAND2_X1 U14055 ( .A1(n11661), .A2(n13444), .ZN(n11663) );
  NAND2_X1 U14056 ( .A1(n13455), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14057 ( .A1(n13448), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11668) );
  OAI21_X1 U14058 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11729), .A(n11664), 
        .ZN(n13903) );
  OR2_X1 U14059 ( .A1(n11769), .A2(n13903), .ZN(n11667) );
  NAND2_X1 U14060 ( .A1(n10245), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14061 ( .A1(n13449), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11665) );
  NAND4_X1 U14062 ( .A1(n11668), .A2(n11667), .A3(n11666), .A4(n11665), .ZN(
        n13673) );
  NAND2_X2 U14063 ( .A1(n14150), .A2(n11671), .ZN(n13937) );
  INV_X1 U14064 ( .A(n13937), .ZN(n14072) );
  OR2_X1 U14065 ( .A1(n11680), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11672) );
  AND2_X1 U14066 ( .A1(n11672), .A2(n11730), .ZN(n13935) );
  NAND2_X1 U14067 ( .A1(n13935), .A2(n11731), .ZN(n11678) );
  INV_X1 U14068 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14069 ( .A1(n13449), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11674) );
  NAND2_X1 U14070 ( .A1(n10245), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n11673) );
  OAI211_X1 U14071 ( .C1(n10252), .C2(n11675), .A(n11674), .B(n11673), .ZN(
        n11676) );
  INV_X1 U14072 ( .A(n11676), .ZN(n11677) );
  NOR2_X1 U14073 ( .A1(n11717), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11679) );
  OR2_X1 U14074 ( .A1(n11680), .A2(n11679), .ZN(n13948) );
  INV_X1 U14075 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U14076 ( .A1(n13448), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14077 ( .A1(n13449), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11681) );
  OAI211_X1 U14078 ( .C1(n11738), .C2(n15259), .A(n11682), .B(n11681), .ZN(
        n11683) );
  INV_X1 U14079 ( .A(n11683), .ZN(n11684) );
  OAI21_X1 U14080 ( .B1(n13948), .B2(n11769), .A(n11684), .ZN(n13675) );
  INV_X1 U14081 ( .A(n13675), .ZN(n11725) );
  NAND2_X1 U14082 ( .A1(n11685), .A2(n13444), .ZN(n11687) );
  NAND2_X1 U14083 ( .A1(n13455), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11686) );
  NAND2_X1 U14084 ( .A1(n11689), .A2(n13444), .ZN(n11692) );
  AOI22_X1 U14085 ( .A1(n6562), .A2(n11690), .B1(n13455), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n11691) );
  INV_X1 U14086 ( .A(n13679), .ZN(n13434) );
  OR2_X1 U14087 ( .A1(n13435), .A2(n13434), .ZN(n13560) );
  NAND2_X1 U14088 ( .A1(n13435), .A2(n13434), .ZN(n13561) );
  NAND2_X1 U14089 ( .A1(n11693), .A2(n13444), .ZN(n11695) );
  AOI22_X1 U14090 ( .A1(n13808), .A2(n6562), .B1(n13455), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n11694) );
  AND2_X1 U14091 ( .A1(n11697), .A2(n11696), .ZN(n11698) );
  OR2_X1 U14092 ( .A1(n11698), .A2(n11705), .ZN(n13997) );
  AOI22_X1 U14093 ( .A1(n13448), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10245), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14094 ( .A1(n13449), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11699) );
  OAI211_X1 U14095 ( .C1(n13997), .C2(n11769), .A(n11700), .B(n11699), .ZN(
        n13678) );
  INV_X1 U14096 ( .A(n13678), .ZN(n13342) );
  OR2_X1 U14097 ( .A1(n14094), .A2(n13342), .ZN(n13563) );
  NAND2_X1 U14098 ( .A1(n14094), .A2(n13342), .ZN(n13564) );
  NAND2_X1 U14099 ( .A1(n13991), .A2(n13990), .ZN(n13989) );
  NAND2_X1 U14100 ( .A1(n11701), .A2(n13444), .ZN(n11704) );
  AOI22_X1 U14101 ( .A1(n13455), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13952), 
        .B2(n6562), .ZN(n11703) );
  NOR2_X1 U14102 ( .A1(n11705), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11706) );
  OR2_X1 U14103 ( .A1(n11715), .A2(n11706), .ZN(n13982) );
  INV_X1 U14104 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13811) );
  NAND2_X1 U14105 ( .A1(n13448), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14106 ( .A1(n13449), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11707) );
  OAI211_X1 U14107 ( .C1(n11738), .C2(n13811), .A(n11708), .B(n11707), .ZN(
        n11709) );
  INV_X1 U14108 ( .A(n11709), .ZN(n11710) );
  OAI21_X1 U14109 ( .B1(n13982), .B2(n11769), .A(n11710), .ZN(n13677) );
  XNOR2_X1 U14110 ( .A(n14089), .B(n13677), .ZN(n13566) );
  INV_X1 U14111 ( .A(n13677), .ZN(n13568) );
  NAND2_X1 U14112 ( .A1(n14089), .A2(n13568), .ZN(n13569) );
  INV_X1 U14113 ( .A(n13569), .ZN(n11711) );
  NAND2_X1 U14114 ( .A1(n11712), .A2(n13444), .ZN(n11714) );
  NAND2_X1 U14115 ( .A1(n13455), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11713) );
  NOR2_X1 U14116 ( .A1(n11715), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11716) );
  OR2_X1 U14117 ( .A1(n11717), .A2(n11716), .ZN(n13967) );
  INV_X1 U14118 ( .A(n13967), .ZN(n11722) );
  INV_X1 U14119 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U14120 ( .A1(n13449), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14121 ( .A1(n10245), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11718) );
  OAI211_X1 U14122 ( .C1(n10252), .C2(n11720), .A(n11719), .B(n11718), .ZN(
        n11721) );
  AOI21_X1 U14123 ( .B1(n11722), .B2(n11731), .A(n11721), .ZN(n13573) );
  INV_X1 U14124 ( .A(n13573), .ZN(n13676) );
  NAND2_X1 U14125 ( .A1(n13962), .A2(n13676), .ZN(n11724) );
  OR2_X1 U14126 ( .A1(n13962), .A2(n13676), .ZN(n11723) );
  NAND2_X1 U14127 ( .A1(n11724), .A2(n11723), .ZN(n13958) );
  NAND2_X1 U14128 ( .A1(n13960), .A2(n11724), .ZN(n13947) );
  XNOR2_X1 U14129 ( .A(n13954), .B(n11725), .ZN(n13439) );
  NAND2_X1 U14130 ( .A1(n13947), .A2(n13946), .ZN(n13945) );
  INV_X1 U14131 ( .A(n15203), .ZN(n13582) );
  NAND2_X1 U14132 ( .A1(n11726), .A2(n13444), .ZN(n11728) );
  NAND2_X1 U14133 ( .A1(n13455), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11727) );
  NAND2_X2 U14134 ( .A1(n11728), .A2(n11727), .ZN(n13919) );
  NAND2_X1 U14135 ( .A1(n13448), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11735) );
  INV_X1 U14136 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15176) );
  OR2_X1 U14137 ( .A1(n11750), .A2(n15176), .ZN(n11734) );
  NAND2_X1 U14138 ( .A1(n10245), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11733) );
  AOI21_X1 U14139 ( .B1(n15150), .B2(n11730), .A(n11729), .ZN(n13916) );
  NAND2_X1 U14140 ( .A1(n11731), .A2(n13916), .ZN(n11732) );
  NAND4_X1 U14141 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n13674) );
  XNOR2_X1 U14142 ( .A(n13919), .B(n13674), .ZN(n13909) );
  INV_X1 U14143 ( .A(n13909), .ZN(n13911) );
  INV_X1 U14144 ( .A(n13919), .ZN(n14065) );
  XNOR2_X1 U14145 ( .A(n13900), .B(n13673), .ZN(n13895) );
  INV_X1 U14146 ( .A(n13895), .ZN(n13899) );
  NOR2_X1 U14147 ( .A1(n13898), .A2(n13899), .ZN(n13897) );
  XNOR2_X1 U14148 ( .A(n14051), .B(n13672), .ZN(n13890) );
  NAND2_X1 U14149 ( .A1(n13267), .A2(n13444), .ZN(n11737) );
  NAND2_X1 U14150 ( .A1(n13455), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11736) );
  INV_X1 U14151 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15260) );
  OR2_X1 U14152 ( .A1(n11738), .A2(n15260), .ZN(n11744) );
  INV_X1 U14153 ( .A(n11739), .ZN(n11740) );
  NAND2_X1 U14154 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n11740), .ZN(n11747) );
  OAI21_X1 U14155 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n11740), .A(n11747), 
        .ZN(n13868) );
  OR2_X1 U14156 ( .A1(n11769), .A2(n13868), .ZN(n11743) );
  NAND2_X1 U14157 ( .A1(n13448), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U14158 ( .A1(n13449), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11741) );
  NAND4_X1 U14159 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n13671) );
  INV_X1 U14160 ( .A(n13671), .ZN(n11745) );
  XNOR2_X1 U14161 ( .A(n14045), .B(n11745), .ZN(n13871) );
  INV_X1 U14162 ( .A(n11747), .ZN(n11746) );
  NAND2_X1 U14163 ( .A1(n11746), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11761) );
  INV_X1 U14164 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14165 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND2_X1 U14166 ( .A1(n11761), .A2(n11749), .ZN(n13852) );
  OR2_X1 U14167 ( .A1(n11769), .A2(n13852), .ZN(n11754) );
  INV_X1 U14168 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15129) );
  OR2_X1 U14169 ( .A1(n11750), .A2(n15129), .ZN(n11753) );
  NAND2_X1 U14170 ( .A1(n13448), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14171 ( .A1(n10245), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U14172 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n13670) );
  NAND2_X1 U14173 ( .A1(n13265), .A2(n13444), .ZN(n11756) );
  NAND2_X1 U14174 ( .A1(n13455), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11755) );
  INV_X1 U14175 ( .A(n14040), .ZN(n13855) );
  NAND2_X1 U14176 ( .A1(n13261), .A2(n13444), .ZN(n11758) );
  NAND2_X1 U14177 ( .A1(n13455), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14178 ( .A1(n13448), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11766) );
  INV_X1 U14179 ( .A(n11761), .ZN(n11759) );
  NAND2_X1 U14180 ( .A1(n11759), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11786) );
  INV_X1 U14181 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14182 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  NAND2_X1 U14183 ( .A1(n11786), .A2(n11762), .ZN(n13839) );
  NAND2_X1 U14184 ( .A1(n10245), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U14185 ( .A1(n13449), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U14186 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n13669) );
  INV_X1 U14187 ( .A(n13669), .ZN(n11803) );
  NAND2_X1 U14188 ( .A1(n13258), .A2(n13444), .ZN(n11768) );
  NAND2_X1 U14189 ( .A1(n13455), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U14190 ( .A1(n13448), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11773) );
  OR2_X1 U14191 ( .A1(n11769), .A2(n11786), .ZN(n11772) );
  NAND2_X1 U14192 ( .A1(n10245), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U14193 ( .A1(n11778), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11770) );
  NAND4_X1 U14194 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n13668) );
  XNOR2_X1 U14195 ( .A(n14029), .B(n13668), .ZN(n13459) );
  INV_X1 U14196 ( .A(n13459), .ZN(n11774) );
  XNOR2_X1 U14197 ( .A(n11775), .B(n11774), .ZN(n11777) );
  INV_X1 U14198 ( .A(n13435), .ZN(n14099) );
  NAND2_X1 U14199 ( .A1(n14008), .A2(n14099), .ZN(n14007) );
  NAND2_X1 U14200 ( .A1(n13937), .A2(n13944), .ZN(n13913) );
  NAND2_X1 U14201 ( .A1(n10245), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U14202 ( .A1(n13448), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U14203 ( .A1(n11778), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11779) );
  NAND3_X1 U14204 ( .A1(n11781), .A2(n11780), .A3(n11779), .ZN(n13667) );
  INV_X1 U14205 ( .A(n13667), .ZN(n13611) );
  NAND2_X1 U14206 ( .A1(n14517), .A2(P1_B_REG_SCAN_IN), .ZN(n11782) );
  NAND2_X1 U14207 ( .A1(n13398), .A2(n11782), .ZN(n13826) );
  NOR2_X1 U14208 ( .A1(n13611), .A2(n13826), .ZN(n14028) );
  NAND3_X1 U14209 ( .A1(n11784), .A2(n14028), .A3(n11783), .ZN(n11785) );
  OAI21_X1 U14210 ( .B1(n14010), .B2(n11786), .A(n11785), .ZN(n11787) );
  AOI21_X1 U14211 ( .B1(n14575), .B2(P1_REG2_REG_29__SCAN_IN), .A(n11787), 
        .ZN(n11788) );
  OAI21_X1 U14212 ( .B1(n13619), .B2(n14012), .A(n11788), .ZN(n11806) );
  NOR2_X1 U14213 ( .A1(n14106), .A2(n13680), .ZN(n11789) );
  NAND2_X1 U14214 ( .A1(n14106), .A2(n13680), .ZN(n11791) );
  AND2_X1 U14215 ( .A1(n13435), .A2(n13679), .ZN(n11793) );
  OR2_X1 U14216 ( .A1(n13435), .A2(n13679), .ZN(n11792) );
  NAND2_X1 U14217 ( .A1(n14094), .A2(n13678), .ZN(n11794) );
  OR2_X1 U14218 ( .A1(n13954), .A2(n13675), .ZN(n11796) );
  NAND2_X1 U14219 ( .A1(n13937), .A2(n15203), .ZN(n11797) );
  NAND2_X1 U14220 ( .A1(n13919), .A2(n13674), .ZN(n11798) );
  NAND2_X1 U14221 ( .A1(n13896), .A2(n13899), .ZN(n11800) );
  OR2_X1 U14222 ( .A1(n13900), .A2(n13673), .ZN(n11799) );
  NAND2_X1 U14223 ( .A1(n11800), .A2(n11799), .ZN(n13891) );
  NAND2_X1 U14224 ( .A1(n14051), .A2(n13672), .ZN(n11801) );
  NOR2_X1 U14225 ( .A1(n13841), .A2(n11803), .ZN(n11804) );
  AOI21_X1 U14226 ( .B1(n13841), .B2(n11803), .A(n11804), .ZN(n13443) );
  INV_X1 U14227 ( .A(n13443), .ZN(n13845) );
  OAI222_X1 U14228 ( .A1(n11808), .A2(P1_U3086), .B1(n14148), .B2(n13454), 
        .C1(n11807), .C2(n14145), .ZN(P1_U3325) );
  INV_X1 U14229 ( .A(n11809), .ZN(n11810) );
  OAI222_X1 U14230 ( .A1(n12609), .A2(n11810), .B1(n12606), .B2(n15059), .C1(
        P3_U3151), .C2(n12164), .ZN(P3_U3268) );
  INV_X1 U14231 ( .A(n11811), .ZN(n11813) );
  OAI222_X1 U14232 ( .A1(n12609), .A2(n11813), .B1(n12606), .B2(n11410), .C1(
        n11812), .C2(P3_U3151), .ZN(P3_U3265) );
  AOI22_X1 U14233 ( .A1(n14106), .A2(n11931), .B1(n6565), .B2(n13680), .ZN(
        n11842) );
  AOI22_X1 U14234 ( .A1(n14106), .A2(n11821), .B1(n11931), .B2(n13680), .ZN(
        n11814) );
  XNOR2_X1 U14235 ( .A(n11814), .B(n11941), .ZN(n11843) );
  INV_X1 U14236 ( .A(n11816), .ZN(n11817) );
  NAND2_X1 U14237 ( .A1(n11815), .A2(n11817), .ZN(n11818) );
  NOR2_X1 U14238 ( .A1(n9739), .A2(n13534), .ZN(n11820) );
  AOI21_X1 U14239 ( .B1(n14476), .B2(n11931), .A(n11820), .ZN(n11824) );
  AOI22_X1 U14240 ( .A1(n14476), .A2(n11930), .B1(n11931), .B2(n13683), .ZN(
        n11822) );
  XNOR2_X1 U14241 ( .A(n11822), .B(n11941), .ZN(n11823) );
  XOR2_X1 U14242 ( .A(n11824), .B(n11823), .Z(n13367) );
  INV_X1 U14243 ( .A(n11823), .ZN(n11826) );
  INV_X1 U14244 ( .A(n11824), .ZN(n11825) );
  AOI22_X1 U14245 ( .A1(n14431), .A2(n11931), .B1(n6565), .B2(n13682), .ZN(
        n11831) );
  NAND2_X1 U14246 ( .A1(n14431), .A2(n11930), .ZN(n11829) );
  NAND2_X1 U14247 ( .A1(n11931), .A2(n13682), .ZN(n11828) );
  NAND2_X1 U14248 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  XNOR2_X1 U14249 ( .A(n11830), .B(n11941), .ZN(n11833) );
  XOR2_X1 U14250 ( .A(n11831), .B(n11833), .Z(n14427) );
  INV_X1 U14251 ( .A(n11831), .ZN(n11832) );
  NAND2_X1 U14252 ( .A1(n11837), .A2(n11930), .ZN(n11835) );
  NAND2_X1 U14253 ( .A1(n11931), .A2(n13681), .ZN(n11834) );
  NAND2_X1 U14254 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  XNOR2_X1 U14255 ( .A(n11836), .B(n11941), .ZN(n11839) );
  XNOR2_X1 U14256 ( .A(n11841), .B(n11839), .ZN(n13407) );
  OAI22_X1 U14257 ( .A1(n7089), .A2(n11884), .B1(n11838), .B2(n9739), .ZN(
        n13406) );
  INV_X1 U14258 ( .A(n11839), .ZN(n11840) );
  NAND2_X1 U14259 ( .A1(n13405), .A2(n7536), .ZN(n13329) );
  INV_X1 U14260 ( .A(n13329), .ZN(n11845) );
  XNOR2_X1 U14261 ( .A(n11843), .B(n11842), .ZN(n13330) );
  NAND2_X1 U14262 ( .A1(n13435), .A2(n11930), .ZN(n11847) );
  NAND2_X1 U14263 ( .A1(n13679), .A2(n11931), .ZN(n11846) );
  NAND2_X1 U14264 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  XNOR2_X1 U14265 ( .A(n11848), .B(n11941), .ZN(n13338) );
  NAND2_X1 U14266 ( .A1(n13435), .A2(n11931), .ZN(n11850) );
  NAND2_X1 U14267 ( .A1(n6565), .A2(n13679), .ZN(n11849) );
  NAND2_X1 U14268 ( .A1(n11850), .A2(n11849), .ZN(n13337) );
  NOR2_X1 U14269 ( .A1(n13338), .A2(n13337), .ZN(n11853) );
  INV_X1 U14270 ( .A(n13338), .ZN(n11852) );
  INV_X1 U14271 ( .A(n13337), .ZN(n11851) );
  AOI22_X1 U14272 ( .A1(n14094), .A2(n11931), .B1(n6565), .B2(n13678), .ZN(
        n11861) );
  NAND2_X1 U14273 ( .A1(n14094), .A2(n11930), .ZN(n11855) );
  NAND2_X1 U14274 ( .A1(n13678), .A2(n11931), .ZN(n11854) );
  NAND2_X1 U14275 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  XNOR2_X1 U14276 ( .A(n11856), .B(n11941), .ZN(n11863) );
  XOR2_X1 U14277 ( .A(n11861), .B(n11863), .Z(n13386) );
  NAND2_X1 U14278 ( .A1(n14089), .A2(n11930), .ZN(n11858) );
  NAND2_X1 U14279 ( .A1(n13677), .A2(n11931), .ZN(n11857) );
  NAND2_X1 U14280 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  XNOR2_X1 U14281 ( .A(n11859), .B(n11910), .ZN(n11864) );
  AND2_X1 U14282 ( .A1(n13677), .A2(n6565), .ZN(n11860) );
  AOI21_X1 U14283 ( .B1(n14089), .B2(n11931), .A(n11860), .ZN(n11865) );
  XNOR2_X1 U14284 ( .A(n11864), .B(n11865), .ZN(n13299) );
  INV_X1 U14285 ( .A(n11861), .ZN(n11862) );
  NOR2_X1 U14286 ( .A1(n11863), .A2(n11862), .ZN(n13300) );
  INV_X1 U14287 ( .A(n11864), .ZN(n11867) );
  INV_X1 U14288 ( .A(n11865), .ZN(n11866) );
  NAND2_X1 U14289 ( .A1(n11867), .A2(n11866), .ZN(n11868) );
  OAI22_X1 U14290 ( .A1(n13962), .A2(n11882), .B1(n13573), .B2(n11884), .ZN(
        n11869) );
  XNOR2_X1 U14291 ( .A(n11869), .B(n11941), .ZN(n11873) );
  AND2_X1 U14292 ( .A1(n13676), .A2(n6565), .ZN(n11870) );
  AOI21_X1 U14293 ( .B1(n14083), .B2(n11931), .A(n11870), .ZN(n11871) );
  XNOR2_X1 U14294 ( .A(n11873), .B(n11871), .ZN(n13358) );
  INV_X1 U14295 ( .A(n11871), .ZN(n11872) );
  NAND2_X1 U14296 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  NAND2_X1 U14297 ( .A1(n13954), .A2(n11930), .ZN(n11876) );
  NAND2_X1 U14298 ( .A1(n13675), .A2(n11931), .ZN(n11875) );
  NAND2_X1 U14299 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  XNOR2_X1 U14300 ( .A(n11877), .B(n11910), .ZN(n11880) );
  AND2_X1 U14301 ( .A1(n13675), .A2(n6565), .ZN(n11878) );
  AOI21_X1 U14302 ( .B1(n13954), .B2(n11931), .A(n11878), .ZN(n11879) );
  NAND2_X1 U14303 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  OAI21_X1 U14304 ( .B1(n11880), .B2(n11879), .A(n11881), .ZN(n13308) );
  OAI22_X1 U14305 ( .A1(n13937), .A2(n11882), .B1(n15203), .B2(n11884), .ZN(
        n11883) );
  XNOR2_X1 U14306 ( .A(n11883), .B(n11941), .ZN(n11888) );
  OR2_X1 U14307 ( .A1(n13937), .A2(n11884), .ZN(n11886) );
  NAND2_X1 U14308 ( .A1(n13582), .A2(n6565), .ZN(n11885) );
  NAND2_X1 U14309 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  NOR2_X1 U14310 ( .A1(n11888), .A2(n11887), .ZN(n11889) );
  AOI21_X1 U14311 ( .B1(n11888), .B2(n11887), .A(n11889), .ZN(n13377) );
  INV_X1 U14312 ( .A(n11889), .ZN(n11890) );
  NAND2_X1 U14313 ( .A1(n13919), .A2(n11930), .ZN(n11892) );
  NAND2_X1 U14314 ( .A1(n11931), .A2(n13674), .ZN(n11891) );
  NAND2_X1 U14315 ( .A1(n11892), .A2(n11891), .ZN(n11893) );
  XNOR2_X1 U14316 ( .A(n11893), .B(n11941), .ZN(n11897) );
  NAND2_X1 U14317 ( .A1(n13919), .A2(n11931), .ZN(n11895) );
  NAND2_X1 U14318 ( .A1(n6565), .A2(n13674), .ZN(n11894) );
  NAND2_X1 U14319 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  NOR2_X1 U14320 ( .A1(n11897), .A2(n11896), .ZN(n13348) );
  AOI21_X1 U14321 ( .B1(n11897), .B2(n11896), .A(n13348), .ZN(n13286) );
  NAND2_X1 U14322 ( .A1(n13900), .A2(n11930), .ZN(n11899) );
  NAND2_X1 U14323 ( .A1(n11931), .A2(n13673), .ZN(n11898) );
  NAND2_X1 U14324 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  XNOR2_X1 U14325 ( .A(n11900), .B(n11910), .ZN(n11903) );
  INV_X1 U14326 ( .A(n13673), .ZN(n11901) );
  NOR2_X1 U14327 ( .A1(n9739), .A2(n11901), .ZN(n11902) );
  AOI21_X1 U14328 ( .B1(n13900), .B2(n11931), .A(n11902), .ZN(n11904) );
  NAND2_X1 U14329 ( .A1(n11903), .A2(n11904), .ZN(n13321) );
  INV_X1 U14330 ( .A(n11903), .ZN(n11906) );
  INV_X1 U14331 ( .A(n11904), .ZN(n11905) );
  NAND2_X1 U14332 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  NAND2_X1 U14333 ( .A1(n13318), .A2(n13321), .ZN(n11919) );
  NAND2_X1 U14334 ( .A1(n14051), .A2(n11930), .ZN(n11909) );
  NAND2_X1 U14335 ( .A1(n11931), .A2(n13672), .ZN(n11908) );
  NAND2_X1 U14336 ( .A1(n11909), .A2(n11908), .ZN(n11911) );
  XNOR2_X1 U14337 ( .A(n11911), .B(n11910), .ZN(n11914) );
  INV_X1 U14338 ( .A(n13672), .ZN(n11912) );
  NOR2_X1 U14339 ( .A1(n9739), .A2(n11912), .ZN(n11913) );
  AOI21_X1 U14340 ( .B1(n14051), .B2(n6559), .A(n11913), .ZN(n11915) );
  NAND2_X1 U14341 ( .A1(n11914), .A2(n11915), .ZN(n11920) );
  INV_X1 U14342 ( .A(n11914), .ZN(n11917) );
  INV_X1 U14343 ( .A(n11915), .ZN(n11916) );
  NAND2_X1 U14344 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  NAND2_X1 U14345 ( .A1(n14045), .A2(n11930), .ZN(n11922) );
  NAND2_X1 U14346 ( .A1(n11931), .A2(n13671), .ZN(n11921) );
  NAND2_X1 U14347 ( .A1(n11922), .A2(n11921), .ZN(n11923) );
  XNOR2_X1 U14348 ( .A(n11923), .B(n11941), .ZN(n11927) );
  NAND2_X1 U14349 ( .A1(n14045), .A2(n11931), .ZN(n11925) );
  NAND2_X1 U14350 ( .A1(n6565), .A2(n13671), .ZN(n11924) );
  NAND2_X1 U14351 ( .A1(n11925), .A2(n11924), .ZN(n11926) );
  NOR2_X1 U14352 ( .A1(n11927), .A2(n11926), .ZN(n11928) );
  AOI21_X1 U14353 ( .B1(n11927), .B2(n11926), .A(n11928), .ZN(n13396) );
  INV_X1 U14354 ( .A(n11928), .ZN(n11929) );
  NAND2_X1 U14355 ( .A1(n14040), .A2(n11930), .ZN(n11933) );
  NAND2_X1 U14356 ( .A1(n11931), .A2(n13670), .ZN(n11932) );
  NAND2_X1 U14357 ( .A1(n11933), .A2(n11932), .ZN(n11934) );
  XNOR2_X1 U14358 ( .A(n11934), .B(n11941), .ZN(n11938) );
  NAND2_X1 U14359 ( .A1(n14040), .A2(n11931), .ZN(n11936) );
  NAND2_X1 U14360 ( .A1(n6565), .A2(n13670), .ZN(n11935) );
  NAND2_X1 U14361 ( .A1(n11936), .A2(n11935), .ZN(n11937) );
  NOR2_X1 U14362 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  AOI21_X1 U14363 ( .B1(n11938), .B2(n11937), .A(n11939), .ZN(n13278) );
  AOI22_X1 U14364 ( .A1(n14033), .A2(n11931), .B1(n6565), .B2(n13669), .ZN(
        n11942) );
  XNOR2_X1 U14365 ( .A(n11942), .B(n11941), .ZN(n11944) );
  AOI22_X1 U14366 ( .A1(n14033), .A2(n11930), .B1(n6559), .B2(n13669), .ZN(
        n11943) );
  XNOR2_X1 U14367 ( .A(n11944), .B(n11943), .ZN(n11945) );
  NAND2_X1 U14368 ( .A1(n13668), .A2(n13398), .ZN(n11947) );
  NAND2_X1 U14369 ( .A1(n13670), .A2(n13662), .ZN(n11946) );
  NAND2_X1 U14370 ( .A1(n11947), .A2(n11946), .ZN(n13837) );
  AOI22_X1 U14371 ( .A1(n14433), .A2(n13837), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11948) );
  OAI21_X1 U14372 ( .B1(n13839), .B2(n14463), .A(n11948), .ZN(n11949) );
  AOI21_X1 U14373 ( .B1(n14033), .B2(n14447), .A(n11949), .ZN(n11950) );
  OAI21_X1 U14374 ( .B1(n11951), .B2(n14458), .A(n11950), .ZN(P1_U3220) );
  OAI222_X1 U14375 ( .A1(n14145), .A2(n11954), .B1(n14148), .B2(n11953), .C1(
        P1_U3086), .C2(n11952), .ZN(P1_U3331) );
  INV_X1 U14376 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n11956) );
  NAND2_X1 U14377 ( .A1(n11955), .A2(n12468), .ZN(n12244) );
  OAI21_X1 U14378 ( .B1(n14946), .B2(n11956), .A(n12244), .ZN(n11958) );
  XNOR2_X1 U14379 ( .A(n12477), .B(n11032), .ZN(n12019) );
  XNOR2_X1 U14380 ( .A(n12019), .B(n12130), .ZN(n12020) );
  XNOR2_X1 U14381 ( .A(n12509), .B(n11032), .ZN(n11975) );
  XNOR2_X1 U14382 ( .A(n11961), .B(n11032), .ZN(n11967) );
  XNOR2_X1 U14383 ( .A(n12592), .B(n11032), .ZN(n11998) );
  NOR2_X1 U14384 ( .A1(n11998), .A2(n12409), .ZN(n11965) );
  XNOR2_X1 U14385 ( .A(n11966), .B(n12423), .ZN(n12117) );
  XNOR2_X1 U14386 ( .A(n11967), .B(n12410), .ZN(n12060) );
  XNOR2_X1 U14387 ( .A(n12579), .B(n11968), .ZN(n12066) );
  NAND2_X1 U14388 ( .A1(n12066), .A2(n12397), .ZN(n11970) );
  INV_X1 U14389 ( .A(n12066), .ZN(n11969) );
  XNOR2_X1 U14390 ( .A(n12101), .B(n11032), .ZN(n12097) );
  NAND2_X1 U14391 ( .A1(n12097), .A2(n12385), .ZN(n11972) );
  INV_X1 U14392 ( .A(n12097), .ZN(n11971) );
  XNOR2_X1 U14393 ( .A(n12572), .B(n11032), .ZN(n11973) );
  XNOR2_X1 U14394 ( .A(n11973), .B(n12346), .ZN(n12013) );
  NAND2_X1 U14395 ( .A1(n12014), .A2(n12013), .ZN(n12012) );
  XNOR2_X1 U14396 ( .A(n11975), .B(n12131), .ZN(n12084) );
  XNOR2_X1 U14397 ( .A(n12338), .B(n11032), .ZN(n11976) );
  XNOR2_X1 U14398 ( .A(n11976), .B(n12323), .ZN(n12044) );
  XNOR2_X1 U14399 ( .A(n12327), .B(n11032), .ZN(n11979) );
  XNOR2_X2 U14400 ( .A(n11978), .B(n11979), .ZN(n12091) );
  NAND2_X1 U14401 ( .A1(n12091), .A2(n12335), .ZN(n11982) );
  XNOR2_X1 U14402 ( .A(n12496), .B(n11032), .ZN(n11985) );
  NAND2_X1 U14403 ( .A1(n12006), .A2(n12324), .ZN(n11984) );
  XNOR2_X1 U14404 ( .A(n12492), .B(n11032), .ZN(n11986) );
  XNOR2_X1 U14405 ( .A(n11986), .B(n12054), .ZN(n12075) );
  INV_X1 U14406 ( .A(n11986), .ZN(n11987) );
  NAND2_X1 U14407 ( .A1(n11987), .A2(n12054), .ZN(n11988) );
  XNOR2_X1 U14408 ( .A(n12486), .B(n11032), .ZN(n11990) );
  XNOR2_X1 U14409 ( .A(n11990), .B(n12274), .ZN(n12051) );
  INV_X1 U14410 ( .A(n11990), .ZN(n11991) );
  NAND2_X1 U14411 ( .A1(n11991), .A2(n12274), .ZN(n11992) );
  XNOR2_X1 U14412 ( .A(n12277), .B(n11032), .ZN(n11993) );
  XNOR2_X1 U14413 ( .A(n11993), .B(n12260), .ZN(n12107) );
  AOI22_X1 U14414 ( .A1(n12285), .A2(n12118), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11995) );
  NAND2_X1 U14415 ( .A1(n12266), .A2(n12124), .ZN(n11994) );
  OAI211_X1 U14416 ( .C1(n12261), .C2(n12120), .A(n11995), .B(n11994), .ZN(
        n11996) );
  AOI21_X1 U14417 ( .B1(n12477), .B2(n6545), .A(n11996), .ZN(n11997) );
  XNOR2_X1 U14418 ( .A(n11998), .B(n12436), .ZN(n11999) );
  XNOR2_X1 U14419 ( .A(n12000), .B(n11999), .ZN(n12005) );
  NOR2_X1 U14420 ( .A1(n12592), .A2(n12121), .ZN(n12003) );
  NAND2_X1 U14421 ( .A1(n12118), .A2(n12454), .ZN(n12001) );
  NAND2_X1 U14422 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n14897)
         );
  OAI211_X1 U14423 ( .C1(n12120), .C2(n12398), .A(n12001), .B(n14897), .ZN(
        n12002) );
  AOI211_X1 U14424 ( .C1(n12426), .C2(n12124), .A(n12003), .B(n12002), .ZN(
        n12004) );
  OAI21_X1 U14425 ( .B1(n12005), .B2(n12126), .A(n12004), .ZN(P3_U3155) );
  XNOR2_X1 U14426 ( .A(n12006), .B(n12297), .ZN(n12011) );
  AOI22_X1 U14427 ( .A1(n12118), .A2(n12310), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12008) );
  NAND2_X1 U14428 ( .A1(n12124), .A2(n12312), .ZN(n12007) );
  OAI211_X1 U14429 ( .C1(n12054), .C2(n12120), .A(n12008), .B(n12007), .ZN(
        n12009) );
  AOI21_X1 U14430 ( .B1(n12496), .B2(n6545), .A(n12009), .ZN(n12010) );
  OAI21_X1 U14431 ( .B1(n12011), .B2(n12126), .A(n12010), .ZN(P3_U3156) );
  OAI211_X1 U14432 ( .C1(n12014), .C2(n12013), .A(n12012), .B(n12058), .ZN(
        n12018) );
  NAND2_X1 U14433 ( .A1(n12118), .A2(n12385), .ZN(n12015) );
  NAND2_X1 U14434 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12236)
         );
  OAI211_X1 U14435 ( .C1(n12120), .C2(n12360), .A(n12015), .B(n12236), .ZN(
        n12016) );
  AOI21_X1 U14436 ( .B1(n12363), .B2(n12124), .A(n12016), .ZN(n12017) );
  OAI211_X1 U14437 ( .C1(n12121), .C2(n12572), .A(n12018), .B(n12017), .ZN(
        P3_U3159) );
  XNOR2_X1 U14438 ( .A(n12021), .B(n11032), .ZN(n12022) );
  XNOR2_X1 U14439 ( .A(n12023), .B(n12022), .ZN(n12029) );
  AOI22_X1 U14440 ( .A1(n12130), .A2(n12118), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12025) );
  NAND2_X1 U14441 ( .A1(n12249), .A2(n12124), .ZN(n12024) );
  OAI211_X1 U14442 ( .C1(n12026), .C2(n12120), .A(n12025), .B(n12024), .ZN(
        n12027) );
  AOI21_X1 U14443 ( .B1(n12253), .B2(n6545), .A(n12027), .ZN(n12028) );
  OAI21_X1 U14444 ( .B1(n12029), .B2(n12126), .A(n12028), .ZN(P3_U3160) );
  MUX2_X1 U14445 ( .A(n12037), .B(n12031), .S(n12030), .Z(n12033) );
  XNOR2_X1 U14446 ( .A(n12033), .B(n12032), .ZN(n12034) );
  NAND2_X1 U14447 ( .A1(n12034), .A2(n12058), .ZN(n12042) );
  INV_X1 U14448 ( .A(n14959), .ZN(n12036) );
  AOI21_X1 U14449 ( .B1(n6545), .B2(n12036), .A(n12035), .ZN(n12041) );
  AOI22_X1 U14450 ( .A1(n12109), .A2(n12134), .B1(n12118), .B2(n12037), .ZN(
        n12040) );
  NAND2_X1 U14451 ( .A1(n12124), .A2(n12038), .ZN(n12039) );
  NAND4_X1 U14452 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        P3_U3161) );
  XOR2_X1 U14453 ( .A(n12043), .B(n12044), .Z(n12049) );
  AOI22_X1 U14454 ( .A1(n12118), .A2(n12131), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12046) );
  NAND2_X1 U14455 ( .A1(n12124), .A2(n12339), .ZN(n12045) );
  OAI211_X1 U14456 ( .C1(n12335), .C2(n12120), .A(n12046), .B(n12045), .ZN(
        n12047) );
  AOI21_X1 U14457 ( .B1(n12338), .B2(n6545), .A(n12047), .ZN(n12048) );
  OAI21_X1 U14458 ( .B1(n12049), .B2(n12126), .A(n12048), .ZN(P3_U3163) );
  XOR2_X1 U14459 ( .A(n12051), .B(n12050), .Z(n12057) );
  AOI22_X1 U14460 ( .A1(n12285), .A2(n12109), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12053) );
  NAND2_X1 U14461 ( .A1(n12124), .A2(n12287), .ZN(n12052) );
  OAI211_X1 U14462 ( .C1(n12054), .C2(n12112), .A(n12053), .B(n12052), .ZN(
        n12055) );
  AOI21_X1 U14463 ( .B1(n12486), .B2(n6545), .A(n12055), .ZN(n12056) );
  OAI21_X1 U14464 ( .B1(n12057), .B2(n12126), .A(n12056), .ZN(P3_U3165) );
  OAI211_X1 U14465 ( .C1(n12061), .C2(n12060), .A(n12059), .B(n12058), .ZN(
        n12065) );
  AND2_X1 U14466 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14335) );
  AOI21_X1 U14467 ( .B1(n12109), .B2(n12132), .A(n14335), .ZN(n12062) );
  OAI21_X1 U14468 ( .B1(n12398), .B2(n12112), .A(n12062), .ZN(n12063) );
  AOI21_X1 U14469 ( .B1(n12402), .B2(n12124), .A(n12063), .ZN(n12064) );
  OAI211_X1 U14470 ( .C1(n12584), .C2(n12121), .A(n12065), .B(n12064), .ZN(
        P3_U3166) );
  XNOR2_X1 U14471 ( .A(n12066), .B(n12132), .ZN(n12067) );
  XNOR2_X1 U14472 ( .A(n12068), .B(n12067), .ZN(n12073) );
  AND2_X1 U14473 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14354) );
  AOI21_X1 U14474 ( .B1(n12109), .B2(n12385), .A(n14354), .ZN(n12070) );
  NAND2_X1 U14475 ( .A1(n12124), .A2(n12388), .ZN(n12069) );
  OAI211_X1 U14476 ( .C1(n12410), .C2(n12112), .A(n12070), .B(n12069), .ZN(
        n12071) );
  AOI21_X1 U14477 ( .B1(n12579), .B2(n6545), .A(n12071), .ZN(n12072) );
  OAI21_X1 U14478 ( .B1(n12073), .B2(n12126), .A(n12072), .ZN(P3_U3168) );
  XOR2_X1 U14479 ( .A(n12075), .B(n12074), .Z(n12080) );
  AOI22_X1 U14480 ( .A1(n12296), .A2(n12109), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12077) );
  NAND2_X1 U14481 ( .A1(n12124), .A2(n12298), .ZN(n12076) );
  OAI211_X1 U14482 ( .C1(n12324), .C2(n12112), .A(n12077), .B(n12076), .ZN(
        n12078) );
  AOI21_X1 U14483 ( .B1(n12492), .B2(n6545), .A(n12078), .ZN(n12079) );
  OAI21_X1 U14484 ( .B1(n12080), .B2(n12126), .A(n12079), .ZN(P3_U3169) );
  INV_X1 U14485 ( .A(n12081), .ZN(n12082) );
  AOI21_X1 U14486 ( .B1(n12084), .B2(n12083), .A(n12082), .ZN(n12090) );
  AOI22_X1 U14487 ( .A1(n12109), .A2(n12345), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12086) );
  NAND2_X1 U14488 ( .A1(n12124), .A2(n12352), .ZN(n12085) );
  OAI211_X1 U14489 ( .C1(n12370), .C2(n12112), .A(n12086), .B(n12085), .ZN(
        n12087) );
  AOI21_X1 U14490 ( .B1(n12509), .B2(n6545), .A(n12087), .ZN(n12089) );
  OAI21_X1 U14491 ( .B1(n12090), .B2(n12126), .A(n12089), .ZN(P3_U3173) );
  XNOR2_X1 U14492 ( .A(n12091), .B(n12310), .ZN(n12096) );
  AOI22_X1 U14493 ( .A1(n12118), .A2(n12345), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12093) );
  NAND2_X1 U14494 ( .A1(n12124), .A2(n12328), .ZN(n12092) );
  OAI211_X1 U14495 ( .C1(n12324), .C2(n12120), .A(n12093), .B(n12092), .ZN(
        n12094) );
  AOI21_X1 U14496 ( .B1(n12327), .B2(n6545), .A(n12094), .ZN(n12095) );
  OAI21_X1 U14497 ( .B1(n12096), .B2(n12126), .A(n12095), .ZN(P3_U3175) );
  XNOR2_X1 U14498 ( .A(n12097), .B(n12385), .ZN(n12098) );
  XNOR2_X1 U14499 ( .A(n12099), .B(n12098), .ZN(n12105) );
  NAND2_X1 U14500 ( .A1(n12118), .A2(n12132), .ZN(n12100) );
  NAND2_X1 U14501 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12190)
         );
  OAI211_X1 U14502 ( .C1(n12120), .C2(n12370), .A(n12100), .B(n12190), .ZN(
        n12103) );
  INV_X1 U14503 ( .A(n12101), .ZN(n12576) );
  NOR2_X1 U14504 ( .A1(n12576), .A2(n12121), .ZN(n12102) );
  AOI211_X1 U14505 ( .C1(n12376), .C2(n12124), .A(n12103), .B(n12102), .ZN(
        n12104) );
  OAI21_X1 U14506 ( .B1(n12105), .B2(n12126), .A(n12104), .ZN(P3_U3178) );
  XOR2_X1 U14507 ( .A(n12107), .B(n12106), .Z(n12115) );
  AOI22_X1 U14508 ( .A1(n12130), .A2(n12109), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12111) );
  NAND2_X1 U14509 ( .A1(n12278), .A2(n12124), .ZN(n12110) );
  OAI211_X1 U14510 ( .C1(n12274), .C2(n12112), .A(n12111), .B(n12110), .ZN(
        n12113) );
  AOI21_X1 U14511 ( .B1(n12277), .B2(n6545), .A(n12113), .ZN(n12114) );
  OAI21_X1 U14512 ( .B1(n12115), .B2(n12126), .A(n12114), .ZN(P3_U3180) );
  XOR2_X1 U14513 ( .A(n12117), .B(n12116), .Z(n12127) );
  NAND2_X1 U14514 ( .A1(n12118), .A2(n12436), .ZN(n12119) );
  NAND2_X1 U14515 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14314)
         );
  OAI211_X1 U14516 ( .C1(n12120), .C2(n12410), .A(n12119), .B(n14314), .ZN(
        n12123) );
  NOR2_X1 U14517 ( .A1(n12588), .A2(n12121), .ZN(n12122) );
  AOI211_X1 U14518 ( .C1(n12414), .C2(n12124), .A(n12123), .B(n12122), .ZN(
        n12125) );
  OAI21_X1 U14519 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(P3_U3181) );
  MUX2_X1 U14520 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12128), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14521 ( .A(n12129), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12140), .Z(
        P3_U3521) );
  MUX2_X1 U14522 ( .A(n12130), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12140), .Z(
        P3_U3518) );
  MUX2_X1 U14523 ( .A(n12285), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12140), .Z(
        P3_U3517) );
  MUX2_X1 U14524 ( .A(n12296), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12140), .Z(
        P3_U3516) );
  MUX2_X1 U14525 ( .A(n12309), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12140), .Z(
        P3_U3515) );
  MUX2_X1 U14526 ( .A(n12297), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12140), .Z(
        P3_U3514) );
  MUX2_X1 U14527 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12310), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14528 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12345), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14529 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12131), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14530 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12346), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14531 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12132), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14532 ( .A(n12384), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12140), .Z(
        P3_U3507) );
  MUX2_X1 U14533 ( .A(n12436), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12140), .Z(
        P3_U3505) );
  MUX2_X1 U14534 ( .A(n12454), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12140), .Z(
        P3_U3504) );
  MUX2_X1 U14535 ( .A(n12455), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12140), .Z(
        P3_U3502) );
  MUX2_X1 U14536 ( .A(n12133), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12140), .Z(
        P3_U3501) );
  MUX2_X1 U14537 ( .A(n12134), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12140), .Z(
        P3_U3500) );
  MUX2_X1 U14538 ( .A(n12135), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12140), .Z(
        P3_U3499) );
  MUX2_X1 U14539 ( .A(n12136), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12140), .Z(
        P3_U3497) );
  MUX2_X1 U14540 ( .A(n12137), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12140), .Z(
        P3_U3495) );
  MUX2_X1 U14541 ( .A(n12138), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12140), .Z(
        P3_U3494) );
  MUX2_X1 U14542 ( .A(n6553), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12140), .Z(
        P3_U3493) );
  MUX2_X1 U14543 ( .A(n12139), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12140), .Z(
        P3_U3492) );
  MUX2_X1 U14544 ( .A(n8751), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12140), .Z(
        P3_U3491) );
  MUX2_X1 U14545 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12164), .Z(n12171) );
  MUX2_X1 U14546 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12164), .Z(n12169) );
  NAND2_X1 U14547 ( .A1(n12142), .A2(n12141), .ZN(n12147) );
  INV_X1 U14548 ( .A(n12143), .ZN(n12145) );
  NAND2_X1 U14549 ( .A1(n12145), .A2(n12144), .ZN(n12146) );
  NAND2_X1 U14550 ( .A1(n12147), .A2(n12146), .ZN(n14838) );
  MUX2_X1 U14551 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12164), .Z(n12148) );
  XNOR2_X1 U14552 ( .A(n12148), .B(n14836), .ZN(n14837) );
  NAND2_X1 U14553 ( .A1(n14838), .A2(n14837), .ZN(n12151) );
  INV_X1 U14554 ( .A(n12148), .ZN(n12149) );
  NAND2_X1 U14555 ( .A1(n12149), .A2(n14836), .ZN(n12150) );
  NAND2_X1 U14556 ( .A1(n12151), .A2(n12150), .ZN(n14863) );
  MUX2_X1 U14557 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12164), .Z(n12152) );
  XNOR2_X1 U14558 ( .A(n12152), .B(n14856), .ZN(n14862) );
  NAND2_X1 U14559 ( .A1(n12152), .A2(n14856), .ZN(n12153) );
  NAND2_X1 U14560 ( .A1(n12154), .A2(n12153), .ZN(n14881) );
  MUX2_X1 U14561 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12164), .Z(n12155) );
  XNOR2_X1 U14562 ( .A(n12155), .B(n12201), .ZN(n14880) );
  INV_X1 U14563 ( .A(n12155), .ZN(n12156) );
  INV_X1 U14564 ( .A(n12201), .ZN(n14875) );
  NAND2_X1 U14565 ( .A1(n12156), .A2(n14875), .ZN(n12157) );
  NAND2_X1 U14566 ( .A1(n14884), .A2(n12157), .ZN(n14901) );
  INV_X1 U14567 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12158) );
  OR2_X1 U14568 ( .A1(n14905), .A2(n12158), .ZN(n12173) );
  NAND2_X1 U14569 ( .A1(n14905), .A2(n12158), .ZN(n12159) );
  NAND2_X1 U14570 ( .A1(n12173), .A2(n12159), .ZN(n14891) );
  INV_X1 U14571 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12537) );
  OR2_X1 U14572 ( .A1(n14905), .A2(n12537), .ZN(n12205) );
  NAND2_X1 U14573 ( .A1(n14905), .A2(n12537), .ZN(n12160) );
  NAND2_X1 U14574 ( .A1(n12205), .A2(n12160), .ZN(n12192) );
  MUX2_X1 U14575 ( .A(n14891), .B(n12192), .S(n12164), .Z(n14900) );
  MUX2_X1 U14576 ( .A(n12173), .B(n12205), .S(n12164), .Z(n12161) );
  NAND2_X1 U14577 ( .A1(n14904), .A2(n12161), .ZN(n12162) );
  XNOR2_X1 U14578 ( .A(n12162), .B(n14323), .ZN(n14319) );
  MUX2_X1 U14579 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12164), .Z(n14318) );
  NAND2_X1 U14580 ( .A1(n14319), .A2(n14318), .ZN(n14317) );
  NAND2_X1 U14581 ( .A1(n12162), .A2(n12206), .ZN(n12163) );
  NAND2_X1 U14582 ( .A1(n14317), .A2(n12163), .ZN(n14330) );
  MUX2_X1 U14583 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12164), .Z(n12166) );
  XNOR2_X1 U14584 ( .A(n12166), .B(n12165), .ZN(n14329) );
  INV_X1 U14585 ( .A(n12166), .ZN(n12167) );
  NAND2_X1 U14586 ( .A1(n12167), .A2(n14326), .ZN(n12168) );
  NAND2_X1 U14587 ( .A1(n14332), .A2(n12168), .ZN(n14350) );
  XNOR2_X1 U14588 ( .A(n12169), .B(n14356), .ZN(n14349) );
  NOR2_X1 U14589 ( .A1(n14350), .A2(n14349), .ZN(n14353) );
  AOI21_X1 U14590 ( .B1(n12169), .B2(n14356), .A(n14353), .ZN(n12227) );
  XNOR2_X1 U14591 ( .A(n12227), .B(n12226), .ZN(n12170) );
  NOR2_X1 U14592 ( .A1(n12170), .A2(n12171), .ZN(n12225) );
  AOI21_X1 U14593 ( .B1(n12171), .B2(n12170), .A(n12225), .ZN(n12219) );
  INV_X1 U14594 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12172) );
  NOR2_X1 U14595 ( .A1(n12226), .A2(n12172), .ZN(n12220) );
  AOI21_X1 U14596 ( .B1(n12226), .B2(n12172), .A(n12220), .ZN(n12188) );
  INV_X1 U14597 ( .A(n12173), .ZN(n12181) );
  NOR2_X1 U14598 ( .A1(n14836), .A2(n12176), .ZN(n12177) );
  XOR2_X1 U14599 ( .A(n12176), .B(n12197), .Z(n14844) );
  NAND2_X1 U14600 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n14856), .ZN(n12178) );
  OAI21_X1 U14601 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n14856), .A(n12178), 
        .ZN(n14851) );
  NOR2_X1 U14602 ( .A1(n14875), .A2(n12179), .ZN(n12180) );
  INV_X1 U14603 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14872) );
  NOR2_X1 U14604 ( .A1(n12181), .A2(n14890), .ZN(n12182) );
  NOR2_X1 U14605 ( .A1(n14323), .A2(n12182), .ZN(n12183) );
  INV_X1 U14606 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14308) );
  INV_X1 U14607 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12184) );
  MUX2_X1 U14608 ( .A(P3_REG2_REG_16__SCAN_IN), .B(n12184), .S(n14326), .Z(
        n14337) );
  OR2_X1 U14609 ( .A1(n14326), .A2(n12184), .ZN(n12185) );
  INV_X1 U14610 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14346) );
  OAI21_X1 U14611 ( .B1(n12188), .B2(n12187), .A(n12221), .ZN(n12189) );
  INV_X1 U14612 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12191) );
  OAI21_X1 U14613 ( .B1(n14878), .B2(n12191), .A(n12190), .ZN(n12217) );
  INV_X1 U14614 ( .A(n12192), .ZN(n14893) );
  NAND2_X1 U14615 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14856), .ZN(n12200) );
  INV_X1 U14616 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12193) );
  MUX2_X1 U14617 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12193), .S(n14856), .Z(
        n14854) );
  NAND2_X1 U14618 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12194), .ZN(n12196) );
  NAND2_X1 U14619 ( .A1(n12197), .A2(n12198), .ZN(n12199) );
  XNOR2_X1 U14620 ( .A(n12198), .B(n14836), .ZN(n14840) );
  NAND2_X1 U14621 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14840), .ZN(n14839) );
  NAND2_X1 U14622 ( .A1(n12199), .A2(n14839), .ZN(n14855) );
  NAND2_X1 U14623 ( .A1(n14854), .A2(n14855), .ZN(n14853) );
  NAND2_X1 U14624 ( .A1(n12200), .A2(n14853), .ZN(n12202) );
  NAND2_X1 U14625 ( .A1(n12201), .A2(n12202), .ZN(n12203) );
  XNOR2_X1 U14626 ( .A(n12202), .B(n14875), .ZN(n14874) );
  NAND2_X1 U14627 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n14874), .ZN(n14873) );
  NAND2_X1 U14628 ( .A1(n12203), .A2(n14873), .ZN(n14894) );
  NAND2_X1 U14629 ( .A1(n14893), .A2(n14894), .ZN(n12204) );
  NAND2_X1 U14630 ( .A1(n12205), .A2(n12204), .ZN(n12207) );
  NAND2_X1 U14631 ( .A1(n12206), .A2(n12207), .ZN(n12208) );
  XNOR2_X1 U14632 ( .A(n14323), .B(n12207), .ZN(n14310) );
  NAND2_X1 U14633 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14310), .ZN(n14309) );
  NAND2_X1 U14634 ( .A1(n12208), .A2(n14309), .ZN(n14328) );
  XNOR2_X1 U14635 ( .A(n14326), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14327) );
  INV_X1 U14636 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12529) );
  NOR2_X1 U14637 ( .A1(n14326), .A2(n12529), .ZN(n12209) );
  AOI21_X1 U14638 ( .B1(n14328), .B2(n14327), .A(n12209), .ZN(n12211) );
  OR2_X1 U14639 ( .A1(n12211), .A2(n12210), .ZN(n12213) );
  XNOR2_X1 U14640 ( .A(n12211), .B(n14356), .ZN(n14348) );
  NAND2_X1 U14641 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14348), .ZN(n14347) );
  INV_X1 U14642 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12519) );
  XNOR2_X1 U14643 ( .A(n12226), .B(n12519), .ZN(n12212) );
  INV_X1 U14644 ( .A(n12230), .ZN(n12215) );
  NAND3_X1 U14645 ( .A1(n12213), .A2(n14347), .A3(n12212), .ZN(n12214) );
  AOI21_X1 U14646 ( .B1(n12215), .B2(n12214), .A(n14313), .ZN(n12216) );
  AOI211_X1 U14647 ( .C1(n14906), .C2(n12226), .A(n12217), .B(n12216), .ZN(
        n12218) );
  XNOR2_X1 U14648 ( .A(n12222), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12224) );
  XNOR2_X1 U14649 ( .A(n12222), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12232) );
  MUX2_X1 U14650 ( .A(n12232), .B(n12224), .S(n12223), .Z(n12229) );
  AOI21_X1 U14651 ( .B1(n12227), .B2(n12226), .A(n12225), .ZN(n12228) );
  XOR2_X1 U14652 ( .A(n12229), .B(n12228), .Z(n12240) );
  XNOR2_X1 U14653 ( .A(n12233), .B(n12232), .ZN(n12234) );
  NOR2_X1 U14654 ( .A1(n12234), .A2(n14313), .ZN(n12239) );
  NAND2_X1 U14655 ( .A1(n14899), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12235) );
  OAI211_X1 U14656 ( .C1(n14357), .C2(n12237), .A(n12236), .B(n12235), .ZN(
        n12238) );
  AOI21_X1 U14657 ( .B1(n12244), .B2(n14363), .A(n14949), .ZN(n12246) );
  AOI21_X1 U14658 ( .B1(n14949), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12246), 
        .ZN(n12245) );
  OAI21_X1 U14659 ( .B1(n12547), .B2(n12428), .A(n12245), .ZN(P3_U3202) );
  AOI21_X1 U14660 ( .B1(n14949), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12246), 
        .ZN(n12247) );
  OAI21_X1 U14661 ( .B1(n14364), .B2(n12428), .A(n12247), .ZN(P3_U3203) );
  INV_X1 U14662 ( .A(n12249), .ZN(n12251) );
  INV_X1 U14663 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12250) );
  OAI22_X1 U14664 ( .A1(n12251), .A2(n14934), .B1(n14946), .B2(n12250), .ZN(
        n12252) );
  AOI21_X1 U14665 ( .B1(n12253), .B2(n12470), .A(n12252), .ZN(n12256) );
  NAND2_X1 U14666 ( .A1(n12254), .A2(n12471), .ZN(n12255) );
  OAI211_X1 U14667 ( .C1(n12248), .C2(n14949), .A(n12256), .B(n12255), .ZN(
        P3_U3205) );
  OAI22_X1 U14668 ( .A1(n12261), .A2(n14943), .B1(n12260), .B2(n14941), .ZN(
        n12262) );
  INV_X1 U14669 ( .A(n12265), .ZN(n14928) );
  NAND2_X1 U14670 ( .A1(n14946), .A2(n14928), .ZN(n12269) );
  AOI22_X1 U14671 ( .A1(n12266), .A2(n12468), .B1(n14949), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12268) );
  NAND2_X1 U14672 ( .A1(n12477), .A2(n12470), .ZN(n12267) );
  OAI211_X1 U14673 ( .C1(n12479), .C2(n12269), .A(n12268), .B(n12267), .ZN(
        n12270) );
  AOI21_X1 U14674 ( .B1(n12480), .B2(n14946), .A(n12270), .ZN(n12271) );
  INV_X1 U14675 ( .A(n12271), .ZN(P3_U3206) );
  INV_X1 U14676 ( .A(n12482), .ZN(n12282) );
  XNOR2_X1 U14677 ( .A(n12276), .B(n12275), .ZN(n12483) );
  INV_X1 U14678 ( .A(n12277), .ZN(n12554) );
  AOI22_X1 U14679 ( .A1(n12278), .A2(n12468), .B1(n14949), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12279) );
  OAI21_X1 U14680 ( .B1(n12554), .B2(n12428), .A(n12279), .ZN(n12280) );
  AOI21_X1 U14681 ( .B1(n12483), .B2(n12471), .A(n12280), .ZN(n12281) );
  OAI21_X1 U14682 ( .B1(n12282), .B2(n14949), .A(n12281), .ZN(P3_U3207) );
  NAND2_X1 U14683 ( .A1(n12283), .A2(n12291), .ZN(n12284) );
  AOI22_X1 U14684 ( .A1(n12285), .A2(n12453), .B1(n12456), .B2(n12309), .ZN(
        n12286) );
  INV_X1 U14685 ( .A(n12287), .ZN(n12289) );
  INV_X1 U14686 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12288) );
  OAI22_X1 U14687 ( .A1(n12289), .A2(n14934), .B1(n14946), .B2(n12288), .ZN(
        n12290) );
  AOI21_X1 U14688 ( .B1(n12486), .B2(n12470), .A(n12290), .ZN(n12294) );
  XNOR2_X1 U14689 ( .A(n12292), .B(n12291), .ZN(n12487) );
  NAND2_X1 U14690 ( .A1(n12487), .A2(n12471), .ZN(n12293) );
  OAI211_X1 U14691 ( .C1(n12489), .C2(n14949), .A(n12294), .B(n12293), .ZN(
        P3_U3208) );
  INV_X1 U14692 ( .A(n12298), .ZN(n12300) );
  OAI22_X1 U14693 ( .A1(n12300), .A2(n14934), .B1(n14946), .B2(n12299), .ZN(
        n12306) );
  INV_X1 U14694 ( .A(n12301), .ZN(n12302) );
  AOI21_X1 U14695 ( .B1(n12304), .B2(n12303), .A(n12302), .ZN(n12495) );
  NOR2_X1 U14696 ( .A1(n12495), .A2(n12431), .ZN(n12305) );
  AOI211_X1 U14697 ( .C1(n12470), .C2(n12492), .A(n12306), .B(n12305), .ZN(
        n12307) );
  OAI21_X1 U14698 ( .B1(n12494), .B2(n14949), .A(n12307), .ZN(P3_U3209) );
  XNOR2_X1 U14699 ( .A(n12308), .B(n12316), .ZN(n12311) );
  AOI222_X1 U14700 ( .A1(n12450), .A2(n12311), .B1(n12310), .B2(n12456), .C1(
        n12309), .C2(n12453), .ZN(n12499) );
  INV_X1 U14701 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12314) );
  INV_X1 U14702 ( .A(n12312), .ZN(n12313) );
  OAI22_X1 U14703 ( .A1(n14946), .A2(n12314), .B1(n12313), .B2(n14934), .ZN(
        n12315) );
  AOI21_X1 U14704 ( .B1(n12496), .B2(n12470), .A(n12315), .ZN(n12320) );
  OR2_X1 U14705 ( .A1(n12317), .A2(n12316), .ZN(n12497) );
  NAND3_X1 U14706 ( .A1(n12497), .A2(n12318), .A3(n12471), .ZN(n12319) );
  OAI211_X1 U14707 ( .C1(n12499), .C2(n14949), .A(n12320), .B(n12319), .ZN(
        P3_U3210) );
  XNOR2_X1 U14708 ( .A(n12321), .B(n12326), .ZN(n12322) );
  OAI222_X1 U14709 ( .A1(n14943), .A2(n12324), .B1(n14941), .B2(n12323), .C1(
        n14939), .C2(n12322), .ZN(n12501) );
  INV_X1 U14710 ( .A(n12501), .ZN(n12332) );
  XOR2_X1 U14711 ( .A(n12325), .B(n12326), .Z(n12502) );
  INV_X1 U14712 ( .A(n12327), .ZN(n12564) );
  AOI22_X1 U14713 ( .A1(n14949), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n12468), 
        .B2(n12328), .ZN(n12329) );
  OAI21_X1 U14714 ( .B1(n12564), .B2(n12428), .A(n12329), .ZN(n12330) );
  AOI21_X1 U14715 ( .B1(n12502), .B2(n12471), .A(n12330), .ZN(n12331) );
  OAI21_X1 U14716 ( .B1(n12332), .B2(n14949), .A(n12331), .ZN(P3_U3211) );
  XOR2_X1 U14717 ( .A(n12333), .B(n12337), .Z(n12334) );
  OAI222_X1 U14718 ( .A1(n14943), .A2(n12335), .B1(n14941), .B2(n12360), .C1(
        n14939), .C2(n12334), .ZN(n12505) );
  INV_X1 U14719 ( .A(n12505), .ZN(n12343) );
  XOR2_X1 U14720 ( .A(n12337), .B(n12336), .Z(n12506) );
  INV_X1 U14721 ( .A(n12338), .ZN(n12567) );
  AOI22_X1 U14722 ( .A1(n14949), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12468), 
        .B2(n12339), .ZN(n12340) );
  OAI21_X1 U14723 ( .B1(n12567), .B2(n12428), .A(n12340), .ZN(n12341) );
  AOI21_X1 U14724 ( .B1(n12506), .B2(n12471), .A(n12341), .ZN(n12342) );
  OAI21_X1 U14725 ( .B1(n12343), .B2(n14949), .A(n12342), .ZN(P3_U3212) );
  XOR2_X1 U14726 ( .A(n12344), .B(n12351), .Z(n12347) );
  AOI222_X1 U14727 ( .A1(n12450), .A2(n12347), .B1(n12346), .B2(n12456), .C1(
        n12345), .C2(n12453), .ZN(n12512) );
  INV_X1 U14728 ( .A(n12348), .ZN(n12349) );
  AOI21_X1 U14729 ( .B1(n12351), .B2(n12350), .A(n12349), .ZN(n12510) );
  INV_X1 U14730 ( .A(n12509), .ZN(n12354) );
  AOI22_X1 U14731 ( .A1(n14949), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n12468), 
        .B2(n12352), .ZN(n12353) );
  OAI21_X1 U14732 ( .B1(n12354), .B2(n12428), .A(n12353), .ZN(n12355) );
  AOI21_X1 U14733 ( .B1(n12510), .B2(n12471), .A(n12355), .ZN(n12356) );
  OAI21_X1 U14734 ( .B1(n12512), .B2(n14949), .A(n12356), .ZN(P3_U3213) );
  XOR2_X1 U14735 ( .A(n12357), .B(n12361), .Z(n12358) );
  OAI222_X1 U14736 ( .A1(n14943), .A2(n12360), .B1(n14941), .B2(n12359), .C1(
        n12358), .C2(n14939), .ZN(n12513) );
  INV_X1 U14737 ( .A(n12513), .ZN(n12367) );
  XNOR2_X1 U14738 ( .A(n12362), .B(n12361), .ZN(n12514) );
  AOI22_X1 U14739 ( .A1(n14949), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n12468), 
        .B2(n12363), .ZN(n12364) );
  OAI21_X1 U14740 ( .B1(n12572), .B2(n12428), .A(n12364), .ZN(n12365) );
  AOI21_X1 U14741 ( .B1(n12514), .B2(n12471), .A(n12365), .ZN(n12366) );
  OAI21_X1 U14742 ( .B1(n12367), .B2(n14949), .A(n12366), .ZN(P3_U3214) );
  OAI21_X1 U14743 ( .B1(n12369), .B2(n12373), .A(n12368), .ZN(n12372) );
  OAI22_X1 U14744 ( .A1(n12397), .A2(n14941), .B1(n12370), .B2(n14943), .ZN(
        n12371) );
  AOI21_X1 U14745 ( .B1(n12372), .B2(n12450), .A(n12371), .ZN(n12518) );
  INV_X1 U14746 ( .A(n12373), .ZN(n12374) );
  XNOR2_X1 U14747 ( .A(n12375), .B(n12374), .ZN(n12516) );
  AOI22_X1 U14748 ( .A1(n14949), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n12468), 
        .B2(n12376), .ZN(n12377) );
  OAI21_X1 U14749 ( .B1(n12576), .B2(n12428), .A(n12377), .ZN(n12378) );
  AOI21_X1 U14750 ( .B1(n12516), .B2(n12471), .A(n12378), .ZN(n12379) );
  OAI21_X1 U14751 ( .B1(n12518), .B2(n14949), .A(n12379), .ZN(P3_U3215) );
  NAND2_X1 U14752 ( .A1(n12381), .A2(n12391), .ZN(n12382) );
  NAND3_X1 U14753 ( .A1(n12383), .A2(n12450), .A3(n12382), .ZN(n12387) );
  AOI22_X1 U14754 ( .A1(n12385), .A2(n12453), .B1(n12456), .B2(n12384), .ZN(
        n12386) );
  INV_X1 U14755 ( .A(n12388), .ZN(n12389) );
  OAI22_X1 U14756 ( .A1(n14946), .A2(n14346), .B1(n12389), .B2(n14934), .ZN(
        n12390) );
  AOI21_X1 U14757 ( .B1(n12579), .B2(n12470), .A(n12390), .ZN(n12394) );
  XNOR2_X1 U14758 ( .A(n12392), .B(n12391), .ZN(n12521) );
  NAND2_X1 U14759 ( .A1(n12521), .A2(n12471), .ZN(n12393) );
  OAI211_X1 U14760 ( .C1(n12523), .C2(n14949), .A(n12394), .B(n12393), .ZN(
        P3_U3216) );
  XOR2_X1 U14761 ( .A(n12395), .B(n12400), .Z(n12396) );
  OAI222_X1 U14762 ( .A1(n14941), .A2(n12398), .B1(n14943), .B2(n12397), .C1(
        n12396), .C2(n14939), .ZN(n12527) );
  INV_X1 U14763 ( .A(n12527), .ZN(n12406) );
  OAI21_X1 U14764 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12528) );
  AOI22_X1 U14765 ( .A1(n14949), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12468), 
        .B2(n12402), .ZN(n12403) );
  OAI21_X1 U14766 ( .B1(n12584), .B2(n12428), .A(n12403), .ZN(n12404) );
  AOI21_X1 U14767 ( .B1(n12528), .B2(n12471), .A(n12404), .ZN(n12405) );
  OAI21_X1 U14768 ( .B1(n12406), .B2(n14949), .A(n12405), .ZN(P3_U3217) );
  XOR2_X1 U14769 ( .A(n12407), .B(n12412), .Z(n12408) );
  OAI222_X1 U14770 ( .A1(n14943), .A2(n12410), .B1(n14941), .B2(n12409), .C1(
        n12408), .C2(n14939), .ZN(n12531) );
  INV_X1 U14771 ( .A(n12531), .ZN(n12418) );
  OAI21_X1 U14772 ( .B1(n12413), .B2(n12412), .A(n12411), .ZN(n12532) );
  AOI22_X1 U14773 ( .A1(n14949), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12468), 
        .B2(n12414), .ZN(n12415) );
  OAI21_X1 U14774 ( .B1(n12428), .B2(n12588), .A(n12415), .ZN(n12416) );
  AOI21_X1 U14775 ( .B1(n12532), .B2(n12471), .A(n12416), .ZN(n12417) );
  OAI21_X1 U14776 ( .B1(n12418), .B2(n14949), .A(n12417), .ZN(P3_U3218) );
  XNOR2_X1 U14777 ( .A(n12419), .B(n12421), .ZN(n12536) );
  INV_X1 U14778 ( .A(n12536), .ZN(n12432) );
  OAI211_X1 U14779 ( .C1(n12422), .C2(n12421), .A(n12420), .B(n12450), .ZN(
        n12425) );
  AOI22_X1 U14780 ( .A1(n12423), .A2(n12453), .B1(n12456), .B2(n12454), .ZN(
        n12424) );
  NAND2_X1 U14781 ( .A1(n12425), .A2(n12424), .ZN(n12535) );
  AOI22_X1 U14782 ( .A1(n14949), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n12468), 
        .B2(n12426), .ZN(n12427) );
  OAI21_X1 U14783 ( .B1(n12428), .B2(n12592), .A(n12427), .ZN(n12429) );
  AOI21_X1 U14784 ( .B1(n12535), .B2(n14946), .A(n12429), .ZN(n12430) );
  OAI21_X1 U14785 ( .B1(n12432), .B2(n12431), .A(n12430), .ZN(P3_U3219) );
  OAI211_X1 U14786 ( .C1(n12435), .C2(n12434), .A(n12433), .B(n12450), .ZN(
        n12439) );
  AOI22_X1 U14787 ( .A1(n12456), .A2(n12437), .B1(n12436), .B2(n12453), .ZN(
        n12438) );
  AND2_X1 U14788 ( .A1(n12439), .A2(n12438), .ZN(n12541) );
  INV_X1 U14789 ( .A(n12596), .ZN(n12443) );
  INV_X1 U14790 ( .A(n12440), .ZN(n12441) );
  OAI22_X1 U14791 ( .A1(n14946), .A2(n14872), .B1(n12441), .B2(n14934), .ZN(
        n12442) );
  AOI21_X1 U14792 ( .B1(n12470), .B2(n12443), .A(n12442), .ZN(n12447) );
  XNOR2_X1 U14793 ( .A(n12445), .B(n12444), .ZN(n12539) );
  NAND2_X1 U14794 ( .A1(n12539), .A2(n12471), .ZN(n12446) );
  OAI211_X1 U14795 ( .C1(n12541), .C2(n14949), .A(n12447), .B(n12446), .ZN(
        P3_U3220) );
  XNOR2_X1 U14796 ( .A(n12448), .B(n12449), .ZN(n14368) );
  INV_X1 U14797 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12464) );
  OAI211_X1 U14798 ( .C1(n6709), .C2(n12452), .A(n12451), .B(n12450), .ZN(
        n12458) );
  AOI22_X1 U14799 ( .A1(n12456), .A2(n12455), .B1(n12454), .B2(n12453), .ZN(
        n12457) );
  NAND2_X1 U14800 ( .A1(n12458), .A2(n12457), .ZN(n14366) );
  NAND2_X1 U14801 ( .A1(n14366), .A2(n14946), .ZN(n12463) );
  NOR2_X1 U14802 ( .A1(n12459), .A2(n14971), .ZN(n14367) );
  AOI22_X1 U14803 ( .A1(n12461), .A2(n14367), .B1(n12468), .B2(n12460), .ZN(
        n12462) );
  OAI211_X1 U14804 ( .C1(n14946), .C2(n12464), .A(n12463), .B(n12462), .ZN(
        n12465) );
  AOI21_X1 U14805 ( .B1(n12471), .B2(n14368), .A(n12465), .ZN(n12466) );
  INV_X1 U14806 ( .A(n12466), .ZN(P3_U3221) );
  MUX2_X1 U14807 ( .A(n15066), .B(n12467), .S(n14946), .Z(n12475) );
  AOI22_X1 U14808 ( .A1(n12470), .A2(n12469), .B1(n12468), .B2(n8295), .ZN(
        n12474) );
  NAND2_X1 U14809 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  NAND3_X1 U14810 ( .A1(n12475), .A2(n12474), .A3(n12473), .ZN(P3_U3230) );
  INV_X1 U14811 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n15183) );
  MUX2_X1 U14812 ( .A(n14363), .B(n15183), .S(n14986), .Z(n12476) );
  OAI21_X1 U14813 ( .B1(n12547), .B2(n12544), .A(n12476), .ZN(P3_U3490) );
  INV_X1 U14814 ( .A(n12477), .ZN(n12550) );
  INV_X1 U14815 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12481) );
  INV_X1 U14816 ( .A(n12478), .ZN(n14958) );
  INV_X1 U14817 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12484) );
  AOI21_X1 U14818 ( .B1(n14963), .B2(n12483), .A(n12482), .ZN(n12551) );
  MUX2_X1 U14819 ( .A(n12484), .B(n12551), .S(n14989), .Z(n12485) );
  OAI21_X1 U14820 ( .B1(n12554), .B2(n12544), .A(n12485), .ZN(P3_U3485) );
  INV_X1 U14821 ( .A(n12486), .ZN(n12558) );
  INV_X1 U14822 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U14823 ( .A1(n12487), .A2(n14963), .ZN(n12488) );
  MUX2_X1 U14824 ( .A(n12490), .B(n12555), .S(n14989), .Z(n12491) );
  NAND2_X1 U14825 ( .A1(n12492), .A2(n14966), .ZN(n12493) );
  OAI211_X1 U14826 ( .C1(n14973), .C2(n12495), .A(n12494), .B(n12493), .ZN(
        n12559) );
  MUX2_X1 U14827 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12559), .S(n14989), .Z(
        P3_U3483) );
  INV_X1 U14828 ( .A(n12496), .ZN(n12500) );
  NAND3_X1 U14829 ( .A1(n12497), .A2(n12318), .A3(n14963), .ZN(n12498) );
  OAI211_X1 U14830 ( .C1(n12500), .C2(n14971), .A(n12499), .B(n12498), .ZN(
        n12560) );
  MUX2_X1 U14831 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12560), .S(n14989), .Z(
        P3_U3482) );
  AOI21_X1 U14832 ( .B1(n14963), .B2(n12502), .A(n12501), .ZN(n12561) );
  MUX2_X1 U14833 ( .A(n12503), .B(n12561), .S(n14989), .Z(n12504) );
  OAI21_X1 U14834 ( .B1(n12564), .B2(n12544), .A(n12504), .ZN(P3_U3481) );
  INV_X1 U14835 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12507) );
  AOI21_X1 U14836 ( .B1(n12506), .B2(n14963), .A(n12505), .ZN(n12565) );
  MUX2_X1 U14837 ( .A(n12507), .B(n12565), .S(n14989), .Z(n12508) );
  OAI21_X1 U14838 ( .B1(n12567), .B2(n12544), .A(n12508), .ZN(P3_U3480) );
  AOI22_X1 U14839 ( .A1(n12510), .A2(n14963), .B1(n14966), .B2(n12509), .ZN(
        n12511) );
  NAND2_X1 U14840 ( .A1(n12512), .A2(n12511), .ZN(n12568) );
  MUX2_X1 U14841 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12568), .S(n14989), .Z(
        P3_U3479) );
  INV_X1 U14842 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n15015) );
  AOI21_X1 U14843 ( .B1(n12514), .B2(n14963), .A(n12513), .ZN(n12569) );
  MUX2_X1 U14844 ( .A(n15015), .B(n12569), .S(n14989), .Z(n12515) );
  OAI21_X1 U14845 ( .B1(n12544), .B2(n12572), .A(n12515), .ZN(P3_U3478) );
  NAND2_X1 U14846 ( .A1(n12516), .A2(n14963), .ZN(n12517) );
  AND2_X1 U14847 ( .A1(n12518), .A2(n12517), .ZN(n12573) );
  MUX2_X1 U14848 ( .A(n12519), .B(n12573), .S(n14989), .Z(n12520) );
  OAI21_X1 U14849 ( .B1(n12576), .B2(n12544), .A(n12520), .ZN(P3_U3477) );
  NAND2_X1 U14850 ( .A1(n12521), .A2(n14963), .ZN(n12522) );
  NAND2_X1 U14851 ( .A1(n12523), .A2(n12522), .ZN(n12577) );
  MUX2_X1 U14852 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12577), .S(n14989), .Z(
        n12524) );
  AOI21_X1 U14853 ( .B1(n12525), .B2(n12579), .A(n12524), .ZN(n12526) );
  INV_X1 U14854 ( .A(n12526), .ZN(P3_U3476) );
  AOI21_X1 U14855 ( .B1(n14963), .B2(n12528), .A(n12527), .ZN(n12581) );
  MUX2_X1 U14856 ( .A(n12529), .B(n12581), .S(n14989), .Z(n12530) );
  OAI21_X1 U14857 ( .B1(n12584), .B2(n12544), .A(n12530), .ZN(P3_U3475) );
  INV_X1 U14858 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12533) );
  AOI21_X1 U14859 ( .B1(n14963), .B2(n12532), .A(n12531), .ZN(n12585) );
  MUX2_X1 U14860 ( .A(n12533), .B(n12585), .S(n14989), .Z(n12534) );
  OAI21_X1 U14861 ( .B1(n12588), .B2(n12544), .A(n12534), .ZN(P3_U3474) );
  AOI21_X1 U14862 ( .B1(n14963), .B2(n12536), .A(n12535), .ZN(n12589) );
  MUX2_X1 U14863 ( .A(n12537), .B(n12589), .S(n14989), .Z(n12538) );
  OAI21_X1 U14864 ( .B1(n12592), .B2(n12544), .A(n12538), .ZN(P3_U3473) );
  INV_X1 U14865 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U14866 ( .A1(n12539), .A2(n14963), .ZN(n12540) );
  MUX2_X1 U14867 ( .A(n12542), .B(n12593), .S(n14989), .Z(n12543) );
  OAI21_X1 U14868 ( .B1(n12544), .B2(n12596), .A(n12543), .ZN(P3_U3472) );
  INV_X1 U14869 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12545) );
  MUX2_X1 U14870 ( .A(n14363), .B(n12545), .S(n14977), .Z(n12546) );
  OAI21_X1 U14871 ( .B1(n12547), .B2(n12597), .A(n12546), .ZN(P3_U3458) );
  MUX2_X1 U14872 ( .A(n12552), .B(n12551), .S(n14979), .Z(n12553) );
  OAI21_X1 U14873 ( .B1(n12554), .B2(n12597), .A(n12553), .ZN(P3_U3453) );
  MUX2_X1 U14874 ( .A(n12556), .B(n12555), .S(n14979), .Z(n12557) );
  OAI21_X1 U14875 ( .B1(n12558), .B2(n12597), .A(n12557), .ZN(P3_U3452) );
  MUX2_X1 U14876 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12559), .S(n14979), .Z(
        P3_U3451) );
  MUX2_X1 U14877 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12560), .S(n14979), .Z(
        P3_U3450) );
  INV_X1 U14878 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12562) );
  MUX2_X1 U14879 ( .A(n12562), .B(n12561), .S(n14979), .Z(n12563) );
  OAI21_X1 U14880 ( .B1(n12564), .B2(n12597), .A(n12563), .ZN(P3_U3449) );
  INV_X1 U14881 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n15244) );
  MUX2_X1 U14882 ( .A(n15244), .B(n12565), .S(n14979), .Z(n12566) );
  OAI21_X1 U14883 ( .B1(n12567), .B2(n12597), .A(n12566), .ZN(P3_U3448) );
  MUX2_X1 U14884 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12568), .S(n14979), .Z(
        P3_U3447) );
  INV_X1 U14885 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12570) );
  MUX2_X1 U14886 ( .A(n12570), .B(n12569), .S(n14979), .Z(n12571) );
  OAI21_X1 U14887 ( .B1(n12597), .B2(n12572), .A(n12571), .ZN(P3_U3446) );
  INV_X1 U14888 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12574) );
  MUX2_X1 U14889 ( .A(n12574), .B(n12573), .S(n14979), .Z(n12575) );
  OAI21_X1 U14890 ( .B1(n12576), .B2(n12597), .A(n12575), .ZN(P3_U3444) );
  MUX2_X1 U14891 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12577), .S(n14979), .Z(
        n12578) );
  AOI21_X1 U14892 ( .B1(n8834), .B2(n12579), .A(n12578), .ZN(n12580) );
  INV_X1 U14893 ( .A(n12580), .ZN(P3_U3441) );
  INV_X1 U14894 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12582) );
  MUX2_X1 U14895 ( .A(n12582), .B(n12581), .S(n14979), .Z(n12583) );
  OAI21_X1 U14896 ( .B1(n12584), .B2(n12597), .A(n12583), .ZN(P3_U3438) );
  INV_X1 U14897 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12586) );
  MUX2_X1 U14898 ( .A(n12586), .B(n12585), .S(n14979), .Z(n12587) );
  OAI21_X1 U14899 ( .B1(n12588), .B2(n12597), .A(n12587), .ZN(P3_U3435) );
  INV_X1 U14900 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12590) );
  MUX2_X1 U14901 ( .A(n12590), .B(n12589), .S(n14979), .Z(n12591) );
  OAI21_X1 U14902 ( .B1(n12592), .B2(n12597), .A(n12591), .ZN(P3_U3432) );
  INV_X1 U14903 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12594) );
  MUX2_X1 U14904 ( .A(n12594), .B(n12593), .S(n14979), .Z(n12595) );
  OAI21_X1 U14905 ( .B1(n12597), .B2(n12596), .A(n12595), .ZN(P3_U3429) );
  NAND4_X1 U14906 ( .A1(n7434), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .A4(n15270), .ZN(n12600) );
  OAI22_X1 U14907 ( .A1(n12598), .A2(n12600), .B1(n12599), .B2(n12606), .ZN(
        n12601) );
  AOI21_X1 U14908 ( .B1(n12603), .B2(n12602), .A(n12601), .ZN(n12604) );
  INV_X1 U14909 ( .A(n12604), .ZN(P3_U3264) );
  INV_X1 U14910 ( .A(n12605), .ZN(n12608) );
  OAI222_X1 U14911 ( .A1(P3_U3151), .A2(n6831), .B1(n12609), .B2(n12608), .C1(
        n12607), .C2(n12606), .ZN(P3_U3267) );
  MUX2_X1 U14912 ( .A(n12611), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U14913 ( .A(n12991), .B(n12673), .ZN(n12672) );
  NAND2_X1 U14914 ( .A1(n12826), .A2(n12619), .ZN(n12671) );
  XNOR2_X1 U14915 ( .A(n13053), .B(n12663), .ZN(n12651) );
  NAND2_X1 U14916 ( .A1(n12831), .A2(n12619), .ZN(n12652) );
  XNOR2_X1 U14917 ( .A(n13194), .B(n12663), .ZN(n12647) );
  INV_X1 U14918 ( .A(n12647), .ZN(n12650) );
  NAND2_X1 U14919 ( .A1(n12832), .A2(n12619), .ZN(n12649) );
  XNOR2_X1 U14920 ( .A(n13078), .B(n6554), .ZN(n12764) );
  NAND2_X1 U14921 ( .A1(n12613), .A2(n12612), .ZN(n12618) );
  INV_X1 U14922 ( .A(n12614), .ZN(n12615) );
  NAND2_X1 U14923 ( .A1(n12616), .A2(n12615), .ZN(n12617) );
  NAND2_X1 U14924 ( .A1(n12618), .A2(n12617), .ZN(n14382) );
  XNOR2_X1 U14925 ( .A(n14396), .B(n12673), .ZN(n12620) );
  NAND2_X1 U14926 ( .A1(n12838), .A2(n12619), .ZN(n12621) );
  NAND2_X1 U14927 ( .A1(n12620), .A2(n12621), .ZN(n12625) );
  INV_X1 U14928 ( .A(n12620), .ZN(n12623) );
  INV_X1 U14929 ( .A(n12621), .ZN(n12622) );
  NAND2_X1 U14930 ( .A1(n12623), .A2(n12622), .ZN(n12624) );
  NAND2_X1 U14931 ( .A1(n12625), .A2(n12624), .ZN(n14381) );
  XNOR2_X1 U14932 ( .A(n13228), .B(n12663), .ZN(n12627) );
  AND2_X1 U14933 ( .A1(n12837), .A2(n12664), .ZN(n12628) );
  XNOR2_X1 U14934 ( .A(n13219), .B(n12663), .ZN(n12630) );
  AND2_X1 U14935 ( .A1(n12836), .A2(n12664), .ZN(n12631) );
  AND2_X1 U14936 ( .A1(n12630), .A2(n12631), .ZN(n12735) );
  AOI21_X1 U14937 ( .B1(n12627), .B2(n12628), .A(n12735), .ZN(n12626) );
  INV_X1 U14938 ( .A(n12627), .ZN(n12733) );
  INV_X1 U14939 ( .A(n12735), .ZN(n12629) );
  INV_X1 U14940 ( .A(n12628), .ZN(n12812) );
  AND2_X1 U14941 ( .A1(n12629), .A2(n12812), .ZN(n12634) );
  INV_X1 U14942 ( .A(n12630), .ZN(n12633) );
  INV_X1 U14943 ( .A(n12631), .ZN(n12632) );
  AND2_X1 U14944 ( .A1(n12633), .A2(n12632), .ZN(n12734) );
  AOI21_X1 U14945 ( .B1(n12733), .B2(n12634), .A(n12734), .ZN(n12635) );
  XNOR2_X1 U14946 ( .A(n13213), .B(n12673), .ZN(n12636) );
  NAND2_X1 U14947 ( .A1(n12835), .A2(n12664), .ZN(n12637) );
  NAND2_X1 U14948 ( .A1(n12636), .A2(n12637), .ZN(n12641) );
  INV_X1 U14949 ( .A(n12636), .ZN(n12639) );
  INV_X1 U14950 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U14951 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  AND2_X1 U14952 ( .A1(n12641), .A2(n12640), .ZN(n12747) );
  NAND2_X1 U14953 ( .A1(n12746), .A2(n12747), .ZN(n12745) );
  XNOR2_X1 U14954 ( .A(n13206), .B(n12673), .ZN(n12642) );
  NAND2_X1 U14955 ( .A1(n12834), .A2(n12664), .ZN(n12643) );
  XNOR2_X1 U14956 ( .A(n12642), .B(n12643), .ZN(n12785) );
  INV_X1 U14957 ( .A(n12642), .ZN(n12645) );
  INV_X1 U14958 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U14959 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  NAND2_X1 U14960 ( .A1(n12833), .A2(n12619), .ZN(n12692) );
  XOR2_X1 U14961 ( .A(n12649), .B(n12647), .Z(n12771) );
  XNOR2_X1 U14962 ( .A(n12651), .B(n12652), .ZN(n12715) );
  XNOR2_X1 U14963 ( .A(n13179), .B(n12663), .ZN(n12654) );
  AND2_X1 U14964 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  NOR2_X2 U14965 ( .A1(n12784), .A2(n12656), .ZN(n12660) );
  XNOR2_X1 U14966 ( .A(n13025), .B(n12663), .ZN(n12658) );
  AND2_X1 U14967 ( .A1(n12829), .A2(n12664), .ZN(n12657) );
  INV_X1 U14968 ( .A(n12658), .ZN(n12659) );
  XNOR2_X1 U14969 ( .A(n13168), .B(n12673), .ZN(n12725) );
  NAND2_X1 U14970 ( .A1(n12828), .A2(n12619), .ZN(n12661) );
  NOR2_X1 U14971 ( .A1(n12725), .A2(n12661), .ZN(n12662) );
  AOI21_X1 U14972 ( .B1(n12725), .B2(n12661), .A(n12662), .ZN(n12756) );
  XNOR2_X1 U14973 ( .A(n13002), .B(n6554), .ZN(n12665) );
  AND2_X1 U14974 ( .A1(n12827), .A2(n12664), .ZN(n12666) );
  NAND2_X1 U14975 ( .A1(n12665), .A2(n12666), .ZN(n12669) );
  INV_X1 U14976 ( .A(n12665), .ZN(n12796) );
  INV_X1 U14977 ( .A(n12666), .ZN(n12667) );
  NAND2_X1 U14978 ( .A1(n12796), .A2(n12667), .ZN(n12668) );
  NAND2_X1 U14979 ( .A1(n12669), .A2(n12668), .ZN(n12723) );
  INV_X1 U14980 ( .A(n12669), .ZN(n12670) );
  XNOR2_X1 U14981 ( .A(n12672), .B(n12671), .ZN(n12799) );
  XNOR2_X1 U14982 ( .A(n13149), .B(n12673), .ZN(n12675) );
  NAND2_X1 U14983 ( .A1(n12825), .A2(n12619), .ZN(n12674) );
  NOR2_X1 U14984 ( .A1(n12675), .A2(n12674), .ZN(n12701) );
  AOI21_X1 U14985 ( .B1(n12675), .B2(n12674), .A(n12701), .ZN(n12676) );
  NAND2_X1 U14986 ( .A1(n12677), .A2(n12676), .ZN(n12703) );
  OAI211_X1 U14987 ( .C1(n12677), .C2(n12676), .A(n12703), .B(n14688), .ZN(
        n12683) );
  NAND2_X1 U14988 ( .A1(n12824), .A2(n12801), .ZN(n12679) );
  NAND2_X1 U14989 ( .A1(n12826), .A2(n12800), .ZN(n12678) );
  NAND2_X1 U14990 ( .A1(n12679), .A2(n12678), .ZN(n12978) );
  OAI22_X1 U14991 ( .A1(n12972), .A2(n14694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12680), .ZN(n12681) );
  AOI21_X1 U14992 ( .B1(n12978), .B2(n14685), .A(n12681), .ZN(n12682) );
  OAI211_X1 U14993 ( .C1(n7131), .C2(n12821), .A(n12683), .B(n12682), .ZN(
        P2_U3186) );
  INV_X1 U14994 ( .A(n12684), .ZN(n12691) );
  AOI22_X1 U14995 ( .A1(n12685), .A2(n14688), .B1(n12813), .B2(n12829), .ZN(
        n12690) );
  AOI22_X1 U14996 ( .A1(n12828), .A2(n12801), .B1(n12800), .B2(n12830), .ZN(
        n13172) );
  INV_X1 U14997 ( .A(n12686), .ZN(n13022) );
  AOI22_X1 U14998 ( .A1(n13022), .A2(n12803), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12687) );
  OAI21_X1 U14999 ( .B1(n13172), .B2(n12806), .A(n12687), .ZN(n12688) );
  AOI21_X1 U15000 ( .B1(n13025), .B2(n14690), .A(n12688), .ZN(n12689) );
  OAI21_X1 U15001 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(P2_U3188) );
  XNOR2_X1 U15002 ( .A(n12764), .B(n12692), .ZN(n12693) );
  XNOR2_X1 U15003 ( .A(n12765), .B(n12693), .ZN(n12700) );
  NAND2_X1 U15004 ( .A1(n12832), .A2(n12801), .ZN(n12695) );
  NAND2_X1 U15005 ( .A1(n12834), .A2(n12800), .ZN(n12694) );
  AND2_X1 U15006 ( .A1(n12695), .A2(n12694), .ZN(n13198) );
  INV_X1 U15007 ( .A(n13198), .ZN(n13077) );
  NAND2_X1 U15008 ( .A1(n13077), .A2(n14685), .ZN(n12697) );
  OAI211_X1 U15009 ( .C1(n14694), .C2(n13074), .A(n12697), .B(n12696), .ZN(
        n12698) );
  AOI21_X1 U15010 ( .B1(n13078), .B2(n14690), .A(n12698), .ZN(n12699) );
  OAI21_X1 U15011 ( .B1(n12700), .B2(n12792), .A(n12699), .ZN(P2_U3191) );
  INV_X1 U15012 ( .A(n12701), .ZN(n12702) );
  NAND2_X1 U15013 ( .A1(n12703), .A2(n12702), .ZN(n12707) );
  NAND2_X1 U15014 ( .A1(n12824), .A2(n12619), .ZN(n12704) );
  XNOR2_X1 U15015 ( .A(n12704), .B(n6554), .ZN(n12705) );
  XNOR2_X1 U15016 ( .A(n13144), .B(n12705), .ZN(n12706) );
  XNOR2_X1 U15017 ( .A(n12707), .B(n12706), .ZN(n12713) );
  AOI22_X1 U15018 ( .A1(n12708), .A2(n12803), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12709) );
  OAI21_X1 U15019 ( .B1(n12710), .B2(n12806), .A(n12709), .ZN(n12711) );
  AOI21_X1 U15020 ( .B1(n13144), .B2(n14690), .A(n12711), .ZN(n12712) );
  OAI21_X1 U15021 ( .B1(n12713), .B2(n12792), .A(n12712), .ZN(P2_U3192) );
  OAI211_X1 U15022 ( .C1(n12716), .C2(n12715), .A(n12714), .B(n14688), .ZN(
        n12722) );
  NAND2_X1 U15023 ( .A1(n12830), .A2(n12801), .ZN(n12718) );
  NAND2_X1 U15024 ( .A1(n12832), .A2(n12800), .ZN(n12717) );
  AND2_X1 U15025 ( .A1(n12718), .A2(n12717), .ZN(n13183) );
  INV_X1 U15026 ( .A(n13183), .ZN(n13052) );
  OAI22_X1 U15027 ( .A1(n14694), .A2(n13049), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12719), .ZN(n12720) );
  AOI21_X1 U15028 ( .B1(n13052), .B2(n14685), .A(n12720), .ZN(n12721) );
  OAI211_X1 U15029 ( .C1(n13185), .C2(n12821), .A(n12722), .B(n12721), .ZN(
        P2_U3195) );
  AOI21_X1 U15030 ( .B1(n12755), .B2(n12723), .A(n12792), .ZN(n12727) );
  NOR3_X1 U15031 ( .A1(n12725), .A2(n12724), .A3(n12794), .ZN(n12726) );
  NOR2_X1 U15032 ( .A1(n12727), .A2(n12726), .ZN(n12731) );
  AOI22_X1 U15033 ( .A1(n12826), .A2(n12801), .B1(n12800), .B2(n12828), .ZN(
        n13160) );
  AOI22_X1 U15034 ( .A1(n12999), .A2(n12803), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12728) );
  OAI21_X1 U15035 ( .B1(n13160), .B2(n12806), .A(n12728), .ZN(n12729) );
  AOI21_X1 U15036 ( .B1(n13002), .B2(n14690), .A(n12729), .ZN(n12730) );
  OAI21_X1 U15037 ( .B1(n12731), .B2(n12798), .A(n12730), .ZN(P2_U3197) );
  XNOR2_X1 U15038 ( .A(n12732), .B(n12733), .ZN(n12814) );
  OAI22_X1 U15039 ( .A1(n12814), .A2(n12812), .B1(n12733), .B2(n12732), .ZN(
        n12737) );
  NOR2_X1 U15040 ( .A1(n12735), .A2(n12734), .ZN(n12736) );
  XNOR2_X1 U15041 ( .A(n12737), .B(n12736), .ZN(n12744) );
  NAND2_X1 U15042 ( .A1(n12835), .A2(n12801), .ZN(n12739) );
  NAND2_X1 U15043 ( .A1(n12837), .A2(n12800), .ZN(n12738) );
  NAND2_X1 U15044 ( .A1(n12739), .A2(n12738), .ZN(n13218) );
  NAND2_X1 U15045 ( .A1(n13218), .A2(n14685), .ZN(n12741) );
  OAI211_X1 U15046 ( .C1(n14694), .C2(n13121), .A(n12741), .B(n12740), .ZN(
        n12742) );
  AOI21_X1 U15047 ( .B1(n13219), .B2(n14690), .A(n12742), .ZN(n12743) );
  OAI21_X1 U15048 ( .B1(n12744), .B2(n12792), .A(n12743), .ZN(P2_U3198) );
  OAI21_X1 U15049 ( .B1(n12747), .B2(n12746), .A(n12745), .ZN(n12748) );
  NAND2_X1 U15050 ( .A1(n12748), .A2(n14688), .ZN(n12754) );
  OAI22_X1 U15051 ( .A1(n12750), .A2(n14754), .B1(n12749), .B2(n14378), .ZN(
        n13212) );
  OAI21_X1 U15052 ( .B1(n14694), .B2(n13106), .A(n12751), .ZN(n12752) );
  AOI21_X1 U15053 ( .B1(n13212), .B2(n14685), .A(n12752), .ZN(n12753) );
  OAI211_X1 U15054 ( .C1(n13110), .C2(n12821), .A(n12754), .B(n12753), .ZN(
        P2_U3200) );
  INV_X1 U15055 ( .A(n13168), .ZN(n13013) );
  OAI211_X1 U15056 ( .C1(n12757), .C2(n12756), .A(n12755), .B(n14688), .ZN(
        n12762) );
  OAI22_X1 U15057 ( .A1(n12795), .A2(n14754), .B1(n12778), .B2(n14378), .ZN(
        n13008) );
  INV_X1 U15058 ( .A(n13011), .ZN(n12759) );
  OAI22_X1 U15059 ( .A1(n12759), .A2(n14694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12758), .ZN(n12760) );
  AOI21_X1 U15060 ( .B1(n13008), .B2(n14685), .A(n12760), .ZN(n12761) );
  OAI211_X1 U15061 ( .C1(n13013), .C2(n12821), .A(n12762), .B(n12761), .ZN(
        P2_U3201) );
  INV_X1 U15062 ( .A(n12763), .ZN(n12774) );
  INV_X1 U15063 ( .A(n12765), .ZN(n12766) );
  OAI33_X1 U15064 ( .A1(n12794), .A2(n12767), .A3(n12788), .B1(n12792), .B2(
        n7342), .B3(n12766), .ZN(n12772) );
  INV_X1 U15065 ( .A(n13194), .ZN(n13066) );
  AOI22_X1 U15066 ( .A1(n12803), .A2(n13063), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12769) );
  OAI22_X1 U15067 ( .A1(n12777), .A2(n14754), .B1(n12788), .B2(n14378), .ZN(
        n13193) );
  NAND2_X1 U15068 ( .A1(n13193), .A2(n14685), .ZN(n12768) );
  OAI211_X1 U15069 ( .C1(n13066), .C2(n12821), .A(n12769), .B(n12768), .ZN(
        n12770) );
  AOI21_X1 U15070 ( .B1(n12772), .B2(n12771), .A(n12770), .ZN(n12773) );
  OAI21_X1 U15071 ( .B1(n12774), .B2(n12792), .A(n12773), .ZN(P2_U3205) );
  INV_X1 U15072 ( .A(n12775), .ZN(n12776) );
  AOI22_X1 U15073 ( .A1(n12776), .A2(n14688), .B1(n12813), .B2(n12830), .ZN(
        n12783) );
  OAI22_X1 U15074 ( .A1(n12778), .A2(n14754), .B1(n12777), .B2(n14378), .ZN(
        n13030) );
  OAI22_X1 U15075 ( .A1(n13032), .A2(n14694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12779), .ZN(n12781) );
  INV_X1 U15076 ( .A(n13179), .ZN(n13035) );
  NOR2_X1 U15077 ( .A1(n13035), .A2(n12821), .ZN(n12780) );
  AOI211_X1 U15078 ( .C1(n14685), .C2(n13030), .A(n12781), .B(n12780), .ZN(
        n12782) );
  OAI21_X1 U15079 ( .B1(n12784), .B2(n12783), .A(n12782), .ZN(P2_U3207) );
  XNOR2_X1 U15080 ( .A(n12786), .B(n12785), .ZN(n12793) );
  OAI22_X1 U15081 ( .A1(n12788), .A2(n14754), .B1(n12787), .B2(n14378), .ZN(
        n13085) );
  OAI22_X1 U15082 ( .A1(n14694), .A2(n13088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15268), .ZN(n12790) );
  NOR2_X1 U15083 ( .A1(n13091), .A2(n12821), .ZN(n12789) );
  AOI211_X1 U15084 ( .C1(n14685), .C2(n13085), .A(n12790), .B(n12789), .ZN(
        n12791) );
  OAI21_X1 U15085 ( .B1(n12793), .B2(n12792), .A(n12791), .ZN(P2_U3210) );
  NOR3_X1 U15086 ( .A1(n12796), .A2(n12795), .A3(n12794), .ZN(n12797) );
  AOI21_X1 U15087 ( .B1(n12798), .B2(n14688), .A(n12797), .ZN(n12811) );
  INV_X1 U15088 ( .A(n12799), .ZN(n12810) );
  AOI22_X1 U15089 ( .A1(n12825), .A2(n12801), .B1(n12800), .B2(n12827), .ZN(
        n13153) );
  NAND2_X1 U15090 ( .A1(n12991), .A2(n14690), .ZN(n12805) );
  INV_X1 U15091 ( .A(n12802), .ZN(n12988) );
  AOI22_X1 U15092 ( .A1(n12988), .A2(n12803), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12804) );
  OAI211_X1 U15093 ( .C1(n13153), .C2(n12806), .A(n12805), .B(n12804), .ZN(
        n12807) );
  AOI21_X1 U15094 ( .B1(n12808), .B2(n14688), .A(n12807), .ZN(n12809) );
  OAI21_X1 U15095 ( .B1(n12811), .B2(n12810), .A(n12809), .ZN(P2_U3212) );
  NAND2_X1 U15096 ( .A1(n14688), .A2(n12812), .ZN(n12816) );
  NAND2_X1 U15097 ( .A1(n12813), .A2(n12837), .ZN(n12815) );
  MUX2_X1 U15098 ( .A(n12816), .B(n12815), .S(n12814), .Z(n12820) );
  OAI22_X1 U15099 ( .A1(n14694), .A2(n12817), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7667), .ZN(n12818) );
  AOI21_X1 U15100 ( .B1(n13227), .B2(n14685), .A(n12818), .ZN(n12819) );
  OAI211_X1 U15101 ( .C1(n7146), .C2(n12821), .A(n12820), .B(n12819), .ZN(
        P2_U3213) );
  MUX2_X1 U15102 ( .A(n12960), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12850), .Z(
        P2_U3562) );
  MUX2_X1 U15103 ( .A(n12822), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12850), .Z(
        P2_U3561) );
  MUX2_X1 U15104 ( .A(n12823), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12850), .Z(
        P2_U3560) );
  MUX2_X1 U15105 ( .A(n12824), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12850), .Z(
        P2_U3559) );
  MUX2_X1 U15106 ( .A(n12825), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12850), .Z(
        P2_U3558) );
  MUX2_X1 U15107 ( .A(n12826), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12850), .Z(
        P2_U3557) );
  MUX2_X1 U15108 ( .A(n12827), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12850), .Z(
        P2_U3556) );
  MUX2_X1 U15109 ( .A(n12828), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12850), .Z(
        P2_U3555) );
  MUX2_X1 U15110 ( .A(n12829), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12850), .Z(
        P2_U3554) );
  MUX2_X1 U15111 ( .A(n12830), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12850), .Z(
        P2_U3553) );
  MUX2_X1 U15112 ( .A(n12831), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12850), .Z(
        P2_U3552) );
  MUX2_X1 U15113 ( .A(n12832), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12850), .Z(
        P2_U3551) );
  INV_X2 U15114 ( .A(P2_U3947), .ZN(n12850) );
  MUX2_X1 U15115 ( .A(n12833), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12850), .Z(
        P2_U3550) );
  MUX2_X1 U15116 ( .A(n12834), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12850), .Z(
        P2_U3549) );
  MUX2_X1 U15117 ( .A(n12835), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12850), .Z(
        P2_U3548) );
  MUX2_X1 U15118 ( .A(n12836), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12850), .Z(
        P2_U3547) );
  MUX2_X1 U15119 ( .A(n12837), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12850), .Z(
        P2_U3546) );
  MUX2_X1 U15120 ( .A(n12838), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12850), .Z(
        P2_U3545) );
  MUX2_X1 U15121 ( .A(n12839), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12850), .Z(
        P2_U3544) );
  MUX2_X1 U15122 ( .A(n12840), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12850), .Z(
        P2_U3543) );
  MUX2_X1 U15123 ( .A(n12841), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12850), .Z(
        P2_U3542) );
  MUX2_X1 U15124 ( .A(n12842), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12850), .Z(
        P2_U3541) );
  MUX2_X1 U15125 ( .A(n12843), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12850), .Z(
        P2_U3540) );
  MUX2_X1 U15126 ( .A(n12844), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12850), .Z(
        P2_U3539) );
  MUX2_X1 U15127 ( .A(n12845), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12850), .Z(
        P2_U3538) );
  MUX2_X1 U15128 ( .A(n12846), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12850), .Z(
        P2_U3537) );
  MUX2_X1 U15129 ( .A(n12847), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12850), .Z(
        P2_U3536) );
  MUX2_X1 U15130 ( .A(n12848), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12850), .Z(
        P2_U3535) );
  MUX2_X1 U15131 ( .A(n12849), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12850), .Z(
        P2_U3534) );
  MUX2_X1 U15132 ( .A(n8876), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12850), .Z(
        P2_U3533) );
  MUX2_X1 U15133 ( .A(n8178), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12850), .Z(
        P2_U3532) );
  MUX2_X1 U15134 ( .A(n8862), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12850), .Z(
        P2_U3531) );
  OAI22_X1 U15135 ( .A1(n12925), .A2(n12857), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12851), .ZN(n12852) );
  AOI21_X1 U15136 ( .B1(n14718), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n12852), .ZN(
        n12865) );
  INV_X1 U15137 ( .A(n12853), .ZN(n12856) );
  OAI21_X1 U15138 ( .B1(n9181), .B2(n12860), .A(n12854), .ZN(n12855) );
  NAND3_X1 U15139 ( .A1(n14725), .A2(n12856), .A3(n12855), .ZN(n12864) );
  MUX2_X1 U15140 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n12858), .S(n12857), .Z(
        n12859) );
  OAI21_X1 U15141 ( .B1(n9360), .B2(n12860), .A(n12859), .ZN(n12861) );
  NAND3_X1 U15142 ( .A1(n6547), .A2(n12862), .A3(n12861), .ZN(n12863) );
  NAND3_X1 U15143 ( .A1(n12865), .A2(n12864), .A3(n12863), .ZN(P2_U3215) );
  OAI21_X1 U15144 ( .B1(n12925), .B2(n12867), .A(n12866), .ZN(n12868) );
  AOI21_X1 U15145 ( .B1(n14718), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n12868), .ZN(
        n12881) );
  INV_X1 U15146 ( .A(n12869), .ZN(n12872) );
  MUX2_X1 U15147 ( .A(n9336), .B(P2_REG1_REG_5__SCAN_IN), .S(n12870), .Z(
        n12871) );
  NAND2_X1 U15148 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  OAI211_X1 U15149 ( .C1(n12874), .C2(n12873), .A(n14725), .B(n12884), .ZN(
        n12880) );
  OR3_X1 U15150 ( .A1(n12877), .A2(n12876), .A3(n12875), .ZN(n12878) );
  NAND3_X1 U15151 ( .A1(n6547), .A2(n12892), .A3(n12878), .ZN(n12879) );
  NAND3_X1 U15152 ( .A1(n12881), .A2(n12880), .A3(n12879), .ZN(P2_U3219) );
  INV_X1 U15153 ( .A(n12904), .ZN(n12886) );
  NAND3_X1 U15154 ( .A1(n12884), .A2(n12883), .A3(n12882), .ZN(n12885) );
  NAND3_X1 U15155 ( .A1(n12886), .A2(n14725), .A3(n12885), .ZN(n12897) );
  OAI21_X1 U15156 ( .B1(n12925), .B2(n12888), .A(n12887), .ZN(n12889) );
  AOI21_X1 U15157 ( .B1(n14718), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n12889), .ZN(
        n12896) );
  INV_X1 U15158 ( .A(n12910), .ZN(n12894) );
  NAND3_X1 U15159 ( .A1(n12892), .A2(n12891), .A3(n12890), .ZN(n12893) );
  NAND3_X1 U15160 ( .A1(n12894), .A2(n6547), .A3(n12893), .ZN(n12895) );
  NAND3_X1 U15161 ( .A1(n12897), .A2(n12896), .A3(n12895), .ZN(P2_U3220) );
  MUX2_X1 U15162 ( .A(n9338), .B(P2_REG1_REG_7__SCAN_IN), .S(n12898), .Z(
        n12901) );
  INV_X1 U15163 ( .A(n12899), .ZN(n12900) );
  NAND2_X1 U15164 ( .A1(n12901), .A2(n12900), .ZN(n12903) );
  OAI211_X1 U15165 ( .C1(n12904), .C2(n12903), .A(n12902), .B(n14725), .ZN(
        n12915) );
  OAI21_X1 U15166 ( .B1(n12925), .B2(n12906), .A(n12905), .ZN(n12907) );
  AOI21_X1 U15167 ( .B1(n14718), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n12907), .ZN(
        n12914) );
  OR3_X1 U15168 ( .A1(n12910), .A2(n12909), .A3(n12908), .ZN(n12911) );
  NAND3_X1 U15169 ( .A1(n12912), .A2(n6547), .A3(n12911), .ZN(n12913) );
  NAND3_X1 U15170 ( .A1(n12915), .A2(n12914), .A3(n12913), .ZN(P2_U3221) );
  INV_X1 U15171 ( .A(n12916), .ZN(n12919) );
  MUX2_X1 U15172 ( .A(n15047), .B(P2_REG1_REG_11__SCAN_IN), .S(n12917), .Z(
        n12918) );
  NAND2_X1 U15173 ( .A1(n12919), .A2(n12918), .ZN(n12921) );
  OAI211_X1 U15174 ( .C1(n12922), .C2(n12921), .A(n12920), .B(n14725), .ZN(
        n12933) );
  OAI21_X1 U15175 ( .B1(n12925), .B2(n12924), .A(n12923), .ZN(n12926) );
  AOI21_X1 U15176 ( .B1(n14718), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n12926), 
        .ZN(n12932) );
  OAI21_X1 U15177 ( .B1(n12929), .B2(n12928), .A(n12927), .ZN(n12930) );
  NAND2_X1 U15178 ( .A1(n12930), .A2(n6547), .ZN(n12931) );
  NAND3_X1 U15179 ( .A1(n12933), .A2(n12932), .A3(n12931), .ZN(P2_U3225) );
  NAND2_X1 U15180 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14386)
         );
  OAI211_X1 U15181 ( .C1(n12936), .C2(n12935), .A(n12934), .B(n14725), .ZN(
        n12937) );
  AND2_X1 U15182 ( .A1(n14386), .A2(n12937), .ZN(n12943) );
  AOI22_X1 U15183 ( .A1(n14718), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n14720), 
        .B2(n12938), .ZN(n12942) );
  OAI211_X1 U15184 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n12940), .A(n6547), .B(
        n12939), .ZN(n12941) );
  NAND3_X1 U15185 ( .A1(n12943), .A2(n12942), .A3(n12941), .ZN(P2_U3228) );
  AOI21_X1 U15186 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12945), .A(n12944), 
        .ZN(n12947) );
  OR2_X1 U15187 ( .A1(n12947), .A2(n15310), .ZN(n12955) );
  NOR2_X1 U15188 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15268), .ZN(n12948) );
  AOI21_X1 U15189 ( .B1(n14720), .B2(n12949), .A(n12948), .ZN(n12954) );
  OAI211_X1 U15190 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n12951), .A(n14725), 
        .B(n12950), .ZN(n12953) );
  NAND2_X1 U15191 ( .A1(n14718), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n12952) );
  NAND4_X1 U15192 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        P2_U3232) );
  NAND2_X1 U15193 ( .A1(n12964), .A2(n13137), .ZN(n12963) );
  XNOR2_X1 U15194 ( .A(n13134), .B(n12963), .ZN(n12957) );
  NAND2_X1 U15195 ( .A1(n12957), .A2(n10011), .ZN(n13133) );
  INV_X1 U15196 ( .A(n12958), .ZN(n12959) );
  NAND2_X1 U15197 ( .A1(n12960), .A2(n12959), .ZN(n13135) );
  NOR2_X1 U15198 ( .A1(n14736), .A2(n13135), .ZN(n12966) );
  NOR2_X1 U15199 ( .A1(n13134), .A2(n14739), .ZN(n12961) );
  AOI211_X1 U15200 ( .C1(n14736), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12966), 
        .B(n12961), .ZN(n12962) );
  OAI21_X1 U15201 ( .B1(n13133), .B2(n13129), .A(n12962), .ZN(P2_U3234) );
  OAI211_X1 U15202 ( .C1(n13137), .C2(n12964), .A(n10011), .B(n12963), .ZN(
        n13136) );
  NOR2_X1 U15203 ( .A1(n13137), .A2(n14739), .ZN(n12965) );
  AOI211_X1 U15204 ( .C1(n14736), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12966), 
        .B(n12965), .ZN(n12967) );
  OAI21_X1 U15205 ( .B1(n13129), .B2(n13136), .A(n12967), .ZN(P2_U3235) );
  XNOR2_X1 U15206 ( .A(n12969), .B(n12968), .ZN(n13152) );
  INV_X1 U15207 ( .A(n12970), .ZN(n12971) );
  AOI211_X1 U15208 ( .C1(n13149), .C2(n12986), .A(n13104), .B(n12971), .ZN(
        n13148) );
  INV_X1 U15209 ( .A(n12972), .ZN(n12973) );
  AOI22_X1 U15210 ( .A1(n12973), .A2(n14734), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14736), .ZN(n12974) );
  OAI21_X1 U15211 ( .B1(n7131), .B2(n14739), .A(n12974), .ZN(n12981) );
  OAI21_X1 U15212 ( .B1(n12977), .B2(n12976), .A(n12975), .ZN(n12979) );
  NOR2_X1 U15213 ( .A1(n13151), .A2(n14736), .ZN(n12980) );
  OAI21_X1 U15214 ( .B1(n13152), .B2(n13114), .A(n12982), .ZN(P2_U3238) );
  XNOR2_X1 U15215 ( .A(n12983), .B(n12985), .ZN(n13159) );
  XOR2_X1 U15216 ( .A(n12985), .B(n12984), .Z(n13157) );
  INV_X1 U15217 ( .A(n12998), .ZN(n12987) );
  OAI211_X1 U15218 ( .C1(n12987), .C2(n13155), .A(n10011), .B(n12986), .ZN(
        n13154) );
  AOI22_X1 U15219 ( .A1(n12988), .A2(n14734), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14736), .ZN(n12989) );
  OAI21_X1 U15220 ( .B1(n13153), .B2(n14736), .A(n12989), .ZN(n12990) );
  AOI21_X1 U15221 ( .B1(n12991), .B2(n14393), .A(n12990), .ZN(n12992) );
  OAI21_X1 U15222 ( .B1(n13154), .B2(n13129), .A(n12992), .ZN(n12993) );
  AOI21_X1 U15223 ( .B1(n13157), .B2(n13131), .A(n12993), .ZN(n12994) );
  OAI21_X1 U15224 ( .B1(n13159), .B2(n13114), .A(n12994), .ZN(P2_U3239) );
  XOR2_X1 U15225 ( .A(n12996), .B(n12995), .Z(n13166) );
  XNOR2_X1 U15226 ( .A(n12997), .B(n12996), .ZN(n13164) );
  OAI211_X1 U15227 ( .C1(n13010), .C2(n13162), .A(n12998), .B(n10011), .ZN(
        n13161) );
  AOI22_X1 U15228 ( .A1(n12999), .A2(n14734), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14736), .ZN(n13000) );
  OAI21_X1 U15229 ( .B1(n13160), .B2(n14736), .A(n13000), .ZN(n13001) );
  AOI21_X1 U15230 ( .B1(n13002), .B2(n14393), .A(n13001), .ZN(n13003) );
  OAI21_X1 U15231 ( .B1(n13161), .B2(n13129), .A(n13003), .ZN(n13004) );
  AOI21_X1 U15232 ( .B1(n13164), .B2(n13131), .A(n13004), .ZN(n13005) );
  OAI21_X1 U15233 ( .B1(n13166), .B2(n13114), .A(n13005), .ZN(P2_U3240) );
  XNOR2_X1 U15234 ( .A(n13007), .B(n13006), .ZN(n13009) );
  AOI21_X1 U15235 ( .B1(n13009), .B2(n14753), .A(n13008), .ZN(n13170) );
  AOI211_X1 U15236 ( .C1(n13168), .C2(n13021), .A(n13104), .B(n13010), .ZN(
        n13167) );
  AOI22_X1 U15237 ( .A1(n13011), .A2(n14734), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14736), .ZN(n13012) );
  OAI21_X1 U15238 ( .B1(n13013), .B2(n14739), .A(n13012), .ZN(n13017) );
  XNOR2_X1 U15239 ( .A(n13015), .B(n13014), .ZN(n13171) );
  NOR2_X1 U15240 ( .A1(n13171), .A2(n13114), .ZN(n13016) );
  OAI21_X1 U15241 ( .B1(n13170), .B2(n14736), .A(n13018), .ZN(P2_U3241) );
  XNOR2_X1 U15242 ( .A(n6618), .B(n13020), .ZN(n13177) );
  XOR2_X1 U15243 ( .A(n13020), .B(n13019), .Z(n13175) );
  OAI211_X1 U15244 ( .C1(n7138), .C2(n7139), .A(n10011), .B(n13021), .ZN(
        n13173) );
  AOI22_X1 U15245 ( .A1(n13022), .A2(n14734), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14736), .ZN(n13023) );
  OAI21_X1 U15246 ( .B1(n13172), .B2(n14736), .A(n13023), .ZN(n13024) );
  AOI21_X1 U15247 ( .B1(n13025), .B2(n14393), .A(n13024), .ZN(n13026) );
  OAI21_X1 U15248 ( .B1(n13173), .B2(n13129), .A(n13026), .ZN(n13027) );
  AOI21_X1 U15249 ( .B1(n13175), .B2(n13131), .A(n13027), .ZN(n13028) );
  OAI21_X1 U15250 ( .B1(n13177), .B2(n13114), .A(n13028), .ZN(P2_U3242) );
  XOR2_X1 U15251 ( .A(n13036), .B(n13029), .Z(n13031) );
  AOI21_X1 U15252 ( .B1(n13031), .B2(n14753), .A(n13030), .ZN(n13181) );
  AOI211_X1 U15253 ( .C1(n13179), .C2(n13047), .A(n12664), .B(n7139), .ZN(
        n13178) );
  INV_X1 U15254 ( .A(n13032), .ZN(n13033) );
  AOI22_X1 U15255 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(n14736), .B1(n13033), 
        .B2(n14734), .ZN(n13034) );
  OAI21_X1 U15256 ( .B1(n13035), .B2(n14739), .A(n13034), .ZN(n13041) );
  NOR2_X1 U15257 ( .A1(n13037), .A2(n13036), .ZN(n13038) );
  OR2_X1 U15258 ( .A1(n13039), .A2(n13038), .ZN(n13182) );
  NOR2_X1 U15259 ( .A1(n13182), .A2(n13114), .ZN(n13040) );
  AOI211_X1 U15260 ( .C1(n13178), .C2(n14731), .A(n13041), .B(n13040), .ZN(
        n13042) );
  OAI21_X1 U15261 ( .B1(n13181), .B2(n14736), .A(n13042), .ZN(P2_U3243) );
  XNOR2_X1 U15262 ( .A(n13044), .B(n13043), .ZN(n13190) );
  XNOR2_X1 U15263 ( .A(n13046), .B(n13045), .ZN(n13187) );
  AOI21_X1 U15264 ( .B1(n13053), .B2(n13062), .A(n13104), .ZN(n13048) );
  NAND2_X1 U15265 ( .A1(n13048), .A2(n13047), .ZN(n13184) );
  OAI22_X1 U15266 ( .A1(n6558), .A2(n13050), .B1(n13049), .B2(n14751), .ZN(
        n13051) );
  AOI21_X1 U15267 ( .B1(n13052), .B2(n6558), .A(n13051), .ZN(n13055) );
  NAND2_X1 U15268 ( .A1(n13053), .A2(n14393), .ZN(n13054) );
  OAI211_X1 U15269 ( .C1(n13184), .C2(n13129), .A(n13055), .B(n13054), .ZN(
        n13056) );
  AOI21_X1 U15270 ( .B1(n13187), .B2(n10037), .A(n13056), .ZN(n13057) );
  OAI21_X1 U15271 ( .B1(n13190), .B2(n13058), .A(n13057), .ZN(P2_U3244) );
  XOR2_X1 U15272 ( .A(n13060), .B(n13059), .Z(n13197) );
  XNOR2_X1 U15273 ( .A(n13061), .B(n13060), .ZN(n13191) );
  NAND2_X1 U15274 ( .A1(n13191), .A2(n13131), .ZN(n13069) );
  AOI211_X1 U15275 ( .C1(n13194), .C2(n13073), .A(n13104), .B(n7140), .ZN(
        n13192) );
  AOI22_X1 U15276 ( .A1(n14736), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13063), 
        .B2(n14734), .ZN(n13065) );
  NAND2_X1 U15277 ( .A1(n13193), .A2(n6558), .ZN(n13064) );
  OAI211_X1 U15278 ( .C1(n13066), .C2(n14739), .A(n13065), .B(n13064), .ZN(
        n13067) );
  AOI21_X1 U15279 ( .B1(n13192), .B2(n14731), .A(n13067), .ZN(n13068) );
  OAI211_X1 U15280 ( .C1(n13197), .C2(n13114), .A(n13069), .B(n13068), .ZN(
        P2_U3245) );
  XOR2_X1 U15281 ( .A(n13071), .B(n13070), .Z(n13204) );
  XNOR2_X1 U15282 ( .A(n13072), .B(n13071), .ZN(n13202) );
  OAI211_X1 U15283 ( .C1(n13087), .C2(n13200), .A(n10011), .B(n13073), .ZN(
        n13199) );
  INV_X1 U15284 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13075) );
  OAI22_X1 U15285 ( .A1(n6558), .A2(n13075), .B1(n13074), .B2(n14751), .ZN(
        n13076) );
  AOI21_X1 U15286 ( .B1(n13077), .B2(n6558), .A(n13076), .ZN(n13080) );
  NAND2_X1 U15287 ( .A1(n13078), .A2(n14393), .ZN(n13079) );
  OAI211_X1 U15288 ( .C1(n13199), .C2(n13129), .A(n13080), .B(n13079), .ZN(
        n13081) );
  AOI21_X1 U15289 ( .B1(n13202), .B2(n13131), .A(n13081), .ZN(n13082) );
  OAI21_X1 U15290 ( .B1(n13114), .B2(n13204), .A(n13082), .ZN(P2_U3246) );
  XNOR2_X1 U15291 ( .A(n13084), .B(n13083), .ZN(n13086) );
  AOI21_X1 U15292 ( .B1(n13086), .B2(n14753), .A(n13085), .ZN(n13208) );
  AOI211_X1 U15293 ( .C1(n13206), .C2(n7147), .A(n13104), .B(n13087), .ZN(
        n13205) );
  INV_X1 U15294 ( .A(n13088), .ZN(n13089) );
  AOI22_X1 U15295 ( .A1(n14736), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13089), 
        .B2(n14734), .ZN(n13090) );
  OAI21_X1 U15296 ( .B1(n13091), .B2(n14739), .A(n13090), .ZN(n13097) );
  INV_X1 U15297 ( .A(n13092), .ZN(n13093) );
  AOI21_X1 U15298 ( .B1(n13095), .B2(n13094), .A(n13093), .ZN(n13209) );
  NOR2_X1 U15299 ( .A1(n13209), .A2(n13114), .ZN(n13096) );
  AOI211_X1 U15300 ( .C1(n13205), .C2(n14731), .A(n13097), .B(n13096), .ZN(
        n13098) );
  OAI21_X1 U15301 ( .B1(n13208), .B2(n14736), .A(n13098), .ZN(P2_U3247) );
  OAI21_X1 U15302 ( .B1(n13100), .B2(n13102), .A(n13099), .ZN(n13216) );
  XOR2_X1 U15303 ( .A(n13102), .B(n13101), .Z(n13210) );
  NAND2_X1 U15304 ( .A1(n13210), .A2(n13131), .ZN(n13113) );
  INV_X1 U15305 ( .A(n6707), .ZN(n13105) );
  AOI211_X1 U15306 ( .C1(n13213), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        n13211) );
  OAI22_X1 U15307 ( .A1(n6558), .A2(n13107), .B1(n13106), .B2(n14751), .ZN(
        n13108) );
  AOI21_X1 U15308 ( .B1(n13212), .B2(n6558), .A(n13108), .ZN(n13109) );
  OAI21_X1 U15309 ( .B1(n13110), .B2(n14739), .A(n13109), .ZN(n13111) );
  AOI21_X1 U15310 ( .B1(n13211), .B2(n14731), .A(n13111), .ZN(n13112) );
  OAI211_X1 U15311 ( .C1(n13216), .C2(n13114), .A(n13113), .B(n13112), .ZN(
        P2_U3248) );
  AOI21_X1 U15312 ( .B1(n13116), .B2(n13119), .A(n13115), .ZN(n13217) );
  NAND2_X1 U15313 ( .A1(n6700), .A2(n13219), .ZN(n13117) );
  NAND2_X1 U15314 ( .A1(n13117), .A2(n10011), .ZN(n13118) );
  OR2_X1 U15315 ( .A1(n13118), .A2(n6707), .ZN(n13222) );
  OR2_X1 U15316 ( .A1(n13120), .A2(n13119), .ZN(n13220) );
  NAND3_X1 U15317 ( .A1(n13220), .A2(n13221), .A3(n10037), .ZN(n13128) );
  NAND2_X1 U15318 ( .A1(n13218), .A2(n6558), .ZN(n13124) );
  INV_X1 U15319 ( .A(n13121), .ZN(n13122) );
  NAND2_X1 U15320 ( .A1(n14734), .A2(n13122), .ZN(n13123) );
  OAI211_X1 U15321 ( .C1(n6558), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        n13126) );
  AOI21_X1 U15322 ( .B1(n13219), .B2(n14393), .A(n13126), .ZN(n13127) );
  OAI211_X1 U15323 ( .C1(n13222), .C2(n13129), .A(n13128), .B(n13127), .ZN(
        n13130) );
  AOI21_X1 U15324 ( .B1(n13217), .B2(n13131), .A(n13130), .ZN(n13132) );
  INV_X1 U15325 ( .A(n13132), .ZN(P2_U3249) );
  OAI211_X1 U15326 ( .C1(n13134), .C2(n14819), .A(n13133), .B(n13135), .ZN(
        n13233) );
  INV_X2 U15327 ( .A(n14834), .ZN(n14833) );
  MUX2_X1 U15328 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13233), .S(n14833), .Z(
        P2_U3530) );
  OAI211_X1 U15329 ( .C1(n13137), .C2(n14819), .A(n13136), .B(n13135), .ZN(
        n13234) );
  MUX2_X1 U15330 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13234), .S(n14833), .Z(
        P2_U3529) );
  AOI21_X1 U15331 ( .B1(n14795), .B2(n13139), .A(n13138), .ZN(n13140) );
  MUX2_X1 U15332 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13235), .S(n14833), .Z(
        P2_U3528) );
  AOI21_X1 U15333 ( .B1(n14795), .B2(n13144), .A(n13143), .ZN(n13145) );
  OAI211_X1 U15334 ( .C1(n14799), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        n13236) );
  MUX2_X1 U15335 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13236), .S(n14833), .Z(
        P2_U3527) );
  AOI21_X1 U15336 ( .B1(n14795), .B2(n13149), .A(n13148), .ZN(n13150) );
  OAI211_X1 U15337 ( .C1(n14799), .C2(n13152), .A(n13151), .B(n13150), .ZN(
        n13237) );
  MUX2_X1 U15338 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13237), .S(n14833), .Z(
        P2_U3526) );
  OAI211_X1 U15339 ( .C1(n13155), .C2(n14819), .A(n13154), .B(n13153), .ZN(
        n13156) );
  AOI21_X1 U15340 ( .B1(n13157), .B2(n14753), .A(n13156), .ZN(n13158) );
  OAI21_X1 U15341 ( .B1(n14799), .B2(n13159), .A(n13158), .ZN(n13238) );
  MUX2_X1 U15342 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13238), .S(n14833), .Z(
        P2_U3525) );
  OAI211_X1 U15343 ( .C1(n13162), .C2(n14819), .A(n13161), .B(n13160), .ZN(
        n13163) );
  AOI21_X1 U15344 ( .B1(n13164), .B2(n14753), .A(n13163), .ZN(n13165) );
  OAI21_X1 U15345 ( .B1(n14799), .B2(n13166), .A(n13165), .ZN(n13239) );
  MUX2_X1 U15346 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13239), .S(n14833), .Z(
        P2_U3524) );
  AOI21_X1 U15347 ( .B1(n14795), .B2(n13168), .A(n13167), .ZN(n13169) );
  OAI211_X1 U15348 ( .C1(n14799), .C2(n13171), .A(n13170), .B(n13169), .ZN(
        n13240) );
  MUX2_X1 U15349 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13240), .S(n14833), .Z(
        P2_U3523) );
  OAI211_X1 U15350 ( .C1(n7138), .C2(n14819), .A(n13173), .B(n13172), .ZN(
        n13174) );
  AOI21_X1 U15351 ( .B1(n13175), .B2(n14753), .A(n13174), .ZN(n13176) );
  OAI21_X1 U15352 ( .B1(n14799), .B2(n13177), .A(n13176), .ZN(n13241) );
  MUX2_X1 U15353 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13241), .S(n14833), .Z(
        P2_U3522) );
  AOI21_X1 U15354 ( .B1(n14795), .B2(n13179), .A(n13178), .ZN(n13180) );
  OAI211_X1 U15355 ( .C1(n14799), .C2(n13182), .A(n13181), .B(n13180), .ZN(
        n13242) );
  MUX2_X1 U15356 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13242), .S(n14833), .Z(
        P2_U3521) );
  OAI211_X1 U15357 ( .C1(n13185), .C2(n14819), .A(n13184), .B(n13183), .ZN(
        n13186) );
  AOI21_X1 U15358 ( .B1(n13187), .B2(n7116), .A(n13186), .ZN(n13188) );
  OAI21_X1 U15359 ( .B1(n13190), .B2(n13189), .A(n13188), .ZN(n13243) );
  MUX2_X1 U15360 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13243), .S(n14833), .Z(
        P2_U3520) );
  NAND2_X1 U15361 ( .A1(n13191), .A2(n14753), .ZN(n13196) );
  AOI211_X1 U15362 ( .C1(n14795), .C2(n13194), .A(n13193), .B(n13192), .ZN(
        n13195) );
  OAI211_X1 U15363 ( .C1(n14799), .C2(n13197), .A(n13196), .B(n13195), .ZN(
        n13244) );
  MUX2_X1 U15364 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13244), .S(n14833), .Z(
        P2_U3519) );
  OAI211_X1 U15365 ( .C1(n13200), .C2(n14819), .A(n13199), .B(n13198), .ZN(
        n13201) );
  AOI21_X1 U15366 ( .B1(n13202), .B2(n14753), .A(n13201), .ZN(n13203) );
  OAI21_X1 U15367 ( .B1(n14799), .B2(n13204), .A(n13203), .ZN(n13245) );
  MUX2_X1 U15368 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13245), .S(n14833), .Z(
        P2_U3518) );
  AOI21_X1 U15369 ( .B1(n14795), .B2(n13206), .A(n13205), .ZN(n13207) );
  OAI211_X1 U15370 ( .C1(n14799), .C2(n13209), .A(n13208), .B(n13207), .ZN(
        n13246) );
  MUX2_X1 U15371 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13246), .S(n14833), .Z(
        P2_U3517) );
  NAND2_X1 U15372 ( .A1(n13210), .A2(n14753), .ZN(n13215) );
  AOI211_X1 U15373 ( .C1(n14795), .C2(n13213), .A(n13212), .B(n13211), .ZN(
        n13214) );
  OAI211_X1 U15374 ( .C1(n14799), .C2(n13216), .A(n13215), .B(n13214), .ZN(
        n13247) );
  MUX2_X1 U15375 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13247), .S(n14833), .Z(
        P2_U3516) );
  NAND2_X1 U15376 ( .A1(n13217), .A2(n14753), .ZN(n13225) );
  AOI21_X1 U15377 ( .B1(n13219), .B2(n14795), .A(n13218), .ZN(n13224) );
  NAND3_X1 U15378 ( .A1(n13221), .A2(n13220), .A3(n7116), .ZN(n13223) );
  NAND4_X1 U15379 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13248) );
  MUX2_X1 U15380 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13248), .S(n14833), .Z(
        P2_U3515) );
  AOI211_X1 U15381 ( .C1(n14795), .C2(n13228), .A(n13227), .B(n13226), .ZN(
        n13231) );
  NAND3_X1 U15382 ( .A1(n6699), .A2(n14753), .A3(n13229), .ZN(n13230) );
  OAI211_X1 U15383 ( .C1(n13232), .C2(n14799), .A(n13231), .B(n13230), .ZN(
        n13249) );
  MUX2_X1 U15384 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13249), .S(n14833), .Z(
        P2_U3514) );
  INV_X2 U15385 ( .A(n14824), .ZN(n14814) );
  MUX2_X1 U15386 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13233), .S(n14814), .Z(
        P2_U3498) );
  MUX2_X1 U15387 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13234), .S(n14814), .Z(
        P2_U3497) );
  MUX2_X1 U15388 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13236), .S(n14814), .Z(
        P2_U3495) );
  MUX2_X1 U15389 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13237), .S(n14814), .Z(
        P2_U3494) );
  MUX2_X1 U15390 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13238), .S(n14814), .Z(
        P2_U3493) );
  MUX2_X1 U15391 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13239), .S(n14814), .Z(
        P2_U3492) );
  MUX2_X1 U15392 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13240), .S(n14814), .Z(
        P2_U3491) );
  MUX2_X1 U15393 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13241), .S(n14814), .Z(
        P2_U3490) );
  MUX2_X1 U15394 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13242), .S(n14814), .Z(
        P2_U3489) );
  MUX2_X1 U15395 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13243), .S(n14814), .Z(
        P2_U3488) );
  MUX2_X1 U15396 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13244), .S(n14814), .Z(
        P2_U3487) );
  MUX2_X1 U15397 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13245), .S(n14814), .Z(
        P2_U3486) );
  MUX2_X1 U15398 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13246), .S(n14814), .Z(
        P2_U3484) );
  MUX2_X1 U15399 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13247), .S(n14814), .Z(
        P2_U3481) );
  MUX2_X1 U15400 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13248), .S(n14814), .Z(
        P2_U3478) );
  MUX2_X1 U15401 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13249), .S(n14814), .Z(
        P2_U3475) );
  INV_X1 U15402 ( .A(n13445), .ZN(n14138) );
  INV_X1 U15403 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13251) );
  NAND3_X1 U15404 ( .A1(n13251), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13253) );
  OAI22_X1 U15405 ( .A1(n13250), .A2(n13253), .B1(n13252), .B2(n13269), .ZN(
        n13254) );
  INV_X1 U15406 ( .A(n13254), .ZN(n13255) );
  OAI21_X1 U15407 ( .B1(n14138), .B2(n13272), .A(n13255), .ZN(P2_U3296) );
  OAI222_X1 U15408 ( .A1(n13272), .A2(n13454), .B1(n13257), .B2(P2_U3088), 
        .C1(n13256), .C2(n13269), .ZN(P2_U3297) );
  INV_X1 U15409 ( .A(n13258), .ZN(n14140) );
  OAI222_X1 U15410 ( .A1(n13272), .A2(n14140), .B1(n13259), .B2(P2_U3088), 
        .C1(n15002), .C2(n13269), .ZN(P2_U3298) );
  NAND2_X1 U15411 ( .A1(n13261), .A2(n13260), .ZN(n13263) );
  OAI211_X1 U15412 ( .C1(n13269), .C2(n13264), .A(n13263), .B(n13262), .ZN(
        P2_U3299) );
  INV_X1 U15413 ( .A(n13265), .ZN(n14143) );
  OAI222_X1 U15414 ( .A1(n13272), .A2(n14143), .B1(n8140), .B2(P2_U3088), .C1(
        n13266), .C2(n13269), .ZN(P2_U3300) );
  INV_X1 U15415 ( .A(n13267), .ZN(n14147) );
  OAI222_X1 U15416 ( .A1(n13269), .A2(n15228), .B1(n13268), .B2(P2_U3088), 
        .C1(n13272), .C2(n14147), .ZN(P2_U3301) );
  OAI222_X1 U15417 ( .A1(n13269), .A2(n13273), .B1(n13272), .B2(n13271), .C1(
        P2_U3088), .C2(n13270), .ZN(P2_U3302) );
  INV_X1 U15418 ( .A(n13274), .ZN(n13275) );
  MUX2_X1 U15419 ( .A(n13275), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15420 ( .A1(n13669), .A2(n13398), .ZN(n13280) );
  NAND2_X1 U15421 ( .A1(n13671), .A2(n13662), .ZN(n13279) );
  NAND2_X1 U15422 ( .A1(n13280), .A2(n13279), .ZN(n13849) );
  AOI22_X1 U15423 ( .A1(n14433), .A2(n13849), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13281) );
  OAI21_X1 U15424 ( .B1(n13852), .B2(n14463), .A(n13281), .ZN(n13282) );
  AOI21_X1 U15425 ( .B1(n14040), .B2(n14447), .A(n13282), .ZN(n13283) );
  OAI21_X1 U15426 ( .B1(n13286), .B2(n13285), .A(n13284), .ZN(n13287) );
  NAND2_X1 U15427 ( .A1(n13287), .A2(n14440), .ZN(n13291) );
  AND2_X1 U15428 ( .A1(n13673), .A2(n13398), .ZN(n13288) );
  AOI21_X1 U15429 ( .B1(n13582), .B2(n13662), .A(n13288), .ZN(n14063) );
  OAI22_X1 U15430 ( .A1(n14063), .A2(n14456), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15150), .ZN(n13289) );
  AOI21_X1 U15431 ( .B1(n13916), .B2(n13410), .A(n13289), .ZN(n13290) );
  OAI211_X1 U15432 ( .C1(n14065), .C2(n13414), .A(n13291), .B(n13290), .ZN(
        P1_U3216) );
  OAI211_X1 U15433 ( .C1(n13294), .C2(n13293), .A(n13292), .B(n14440), .ZN(
        n13298) );
  AOI22_X1 U15434 ( .A1(n14447), .A2(n14596), .B1(n14433), .B2(n13295), .ZN(
        n13297) );
  MUX2_X1 U15435 ( .A(n14463), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n13296) );
  NAND3_X1 U15436 ( .A1(n13298), .A2(n13297), .A3(n13296), .ZN(P1_U3218) );
  OAI21_X1 U15437 ( .B1(n6599), .B2(n13300), .A(n13299), .ZN(n13302) );
  NAND3_X1 U15438 ( .A1(n13302), .A2(n14440), .A3(n13301), .ZN(n13305) );
  OAI22_X1 U15439 ( .A1(n13573), .A2(n13388), .B1(n13342), .B2(n13387), .ZN(
        n13975) );
  AND2_X1 U15440 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13821) );
  NOR2_X1 U15441 ( .A1(n14463), .A2(n13982), .ZN(n13303) );
  AOI211_X1 U15442 ( .C1(n13975), .C2(n14433), .A(n13821), .B(n13303), .ZN(
        n13304) );
  OAI211_X1 U15443 ( .C1(n7159), .C2(n13414), .A(n13305), .B(n13304), .ZN(
        P1_U3219) );
  INV_X1 U15444 ( .A(n13306), .ZN(n13307) );
  AOI21_X1 U15445 ( .B1(n13309), .B2(n13308), .A(n13307), .ZN(n13314) );
  INV_X1 U15446 ( .A(n13954), .ZN(n13310) );
  NOR2_X1 U15447 ( .A1(n13310), .A2(n14655), .ZN(n14077) );
  OAI22_X1 U15448 ( .A1(n15203), .A2(n13388), .B1(n13573), .B2(n13387), .ZN(
        n14076) );
  AOI22_X1 U15449 ( .A1(n14076), .A2(n14433), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13311) );
  OAI21_X1 U15450 ( .B1(n13948), .B2(n14463), .A(n13311), .ZN(n13312) );
  AOI21_X1 U15451 ( .B1(n14077), .B2(n14451), .A(n13312), .ZN(n13313) );
  OAI21_X1 U15452 ( .B1(n13314), .B2(n14458), .A(n13313), .ZN(P1_U3223) );
  NAND2_X1 U15453 ( .A1(n13673), .A2(n13662), .ZN(n13316) );
  NAND2_X1 U15454 ( .A1(n13671), .A2(n13398), .ZN(n13315) );
  NAND2_X1 U15455 ( .A1(n13316), .A2(n13315), .ZN(n14050) );
  AOI22_X1 U15456 ( .A1(n14433), .A2(n14050), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13317) );
  OAI21_X1 U15457 ( .B1(n13882), .B2(n14463), .A(n13317), .ZN(n13325) );
  INV_X1 U15458 ( .A(n13319), .ZN(n13320) );
  NAND3_X1 U15459 ( .A1(n13318), .A2(n13321), .A3(n13320), .ZN(n13322) );
  AOI21_X1 U15460 ( .B1(n13323), .B2(n13322), .A(n14458), .ZN(n13324) );
  AOI211_X1 U15461 ( .C1(n14447), .C2(n14051), .A(n13325), .B(n13324), .ZN(
        n13326) );
  INV_X1 U15462 ( .A(n13326), .ZN(P1_U3225) );
  INV_X1 U15463 ( .A(n13327), .ZN(n13328) );
  AOI21_X1 U15464 ( .B1(n13330), .B2(n13329), .A(n13328), .ZN(n13336) );
  NAND2_X1 U15465 ( .A1(n14433), .A2(n14105), .ZN(n13331) );
  OAI211_X1 U15466 ( .C1(n14463), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        n13334) );
  AOI21_X1 U15467 ( .B1(n14106), .B2(n14447), .A(n13334), .ZN(n13335) );
  OAI21_X1 U15468 ( .B1(n13336), .B2(n14458), .A(n13335), .ZN(P1_U3226) );
  XNOR2_X1 U15469 ( .A(n13338), .B(n13337), .ZN(n13339) );
  XNOR2_X1 U15470 ( .A(n13340), .B(n13339), .ZN(n13347) );
  OAI22_X1 U15471 ( .A1(n13342), .A2(n13388), .B1(n13341), .B2(n13387), .ZN(
        n14009) );
  NAND2_X1 U15472 ( .A1(n14009), .A2(n14433), .ZN(n13344) );
  OAI211_X1 U15473 ( .C1(n14463), .C2(n14011), .A(n13344), .B(n13343), .ZN(
        n13345) );
  AOI21_X1 U15474 ( .B1(n13435), .B2(n14447), .A(n13345), .ZN(n13346) );
  OAI21_X1 U15475 ( .B1(n13347), .B2(n14458), .A(n13346), .ZN(P1_U3228) );
  NOR2_X1 U15476 ( .A1(n13349), .A2(n13348), .ZN(n13351) );
  INV_X1 U15477 ( .A(n13318), .ZN(n13350) );
  AOI21_X1 U15478 ( .B1(n13351), .B2(n13284), .A(n13350), .ZN(n13357) );
  AND2_X1 U15479 ( .A1(n13900), .A2(n14636), .ZN(n14058) );
  NAND2_X1 U15480 ( .A1(n13674), .A2(n13662), .ZN(n13353) );
  NAND2_X1 U15481 ( .A1(n13672), .A2(n13398), .ZN(n13352) );
  NAND2_X1 U15482 ( .A1(n13353), .A2(n13352), .ZN(n14057) );
  AOI22_X1 U15483 ( .A1(n14433), .A2(n14057), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13354) );
  OAI21_X1 U15484 ( .B1(n13903), .B2(n14463), .A(n13354), .ZN(n13355) );
  AOI21_X1 U15485 ( .B1(n14058), .B2(n14451), .A(n13355), .ZN(n13356) );
  OAI21_X1 U15486 ( .B1(n13357), .B2(n14458), .A(n13356), .ZN(P1_U3229) );
  XNOR2_X1 U15487 ( .A(n13359), .B(n13358), .ZN(n13365) );
  NAND2_X1 U15488 ( .A1(n13675), .A2(n13398), .ZN(n13361) );
  NAND2_X1 U15489 ( .A1(n13677), .A2(n13662), .ZN(n13360) );
  NAND2_X1 U15490 ( .A1(n13361), .A2(n13360), .ZN(n13959) );
  AOI22_X1 U15491 ( .A1(n13959), .A2(n14433), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13362) );
  OAI21_X1 U15492 ( .B1(n13967), .B2(n14463), .A(n13362), .ZN(n13363) );
  AOI21_X1 U15493 ( .B1(n14083), .B2(n14447), .A(n13363), .ZN(n13364) );
  OAI21_X1 U15494 ( .B1(n13365), .B2(n14458), .A(n13364), .ZN(P1_U3233) );
  OAI211_X1 U15495 ( .C1(n13368), .C2(n13367), .A(n13366), .B(n14440), .ZN(
        n13374) );
  INV_X1 U15496 ( .A(n13369), .ZN(n13372) );
  OAI21_X1 U15497 ( .B1(n14456), .B2(n14474), .A(n13370), .ZN(n13371) );
  AOI21_X1 U15498 ( .B1(n13372), .B2(n13410), .A(n13371), .ZN(n13373) );
  OAI211_X1 U15499 ( .C1(n7091), .C2(n13414), .A(n13374), .B(n13373), .ZN(
        P1_U3234) );
  OAI21_X1 U15500 ( .B1(n13377), .B2(n13376), .A(n13375), .ZN(n13383) );
  NAND2_X1 U15501 ( .A1(n13675), .A2(n13662), .ZN(n13379) );
  NAND2_X1 U15502 ( .A1(n13674), .A2(n13398), .ZN(n13378) );
  NAND2_X1 U15503 ( .A1(n13379), .A2(n13378), .ZN(n14071) );
  AOI22_X1 U15504 ( .A1(n14071), .A2(n14433), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13381) );
  NAND2_X1 U15505 ( .A1(n13935), .A2(n13410), .ZN(n13380) );
  OAI211_X1 U15506 ( .C1(n13937), .C2(n13414), .A(n13381), .B(n13380), .ZN(
        n13382) );
  AOI21_X1 U15507 ( .B1(n13383), .B2(n14440), .A(n13382), .ZN(n13384) );
  INV_X1 U15508 ( .A(n13384), .ZN(P1_U3235) );
  AOI21_X1 U15509 ( .B1(n13386), .B2(n13385), .A(n6599), .ZN(n13393) );
  OAI22_X1 U15510 ( .A1(n13568), .A2(n13388), .B1(n13434), .B2(n13387), .ZN(
        n13992) );
  NAND2_X1 U15511 ( .A1(n13992), .A2(n14433), .ZN(n13390) );
  OAI211_X1 U15512 ( .C1(n14463), .C2(n13997), .A(n13390), .B(n13389), .ZN(
        n13391) );
  AOI21_X1 U15513 ( .B1(n14094), .B2(n14447), .A(n13391), .ZN(n13392) );
  OAI21_X1 U15514 ( .B1(n13393), .B2(n14458), .A(n13392), .ZN(P1_U3238) );
  OAI21_X1 U15515 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(n13397) );
  INV_X1 U15516 ( .A(n13397), .ZN(n13404) );
  NAND2_X1 U15517 ( .A1(n13670), .A2(n13398), .ZN(n13400) );
  NAND2_X1 U15518 ( .A1(n13672), .A2(n13662), .ZN(n13399) );
  NAND2_X1 U15519 ( .A1(n13400), .A2(n13399), .ZN(n13864) );
  AOI22_X1 U15520 ( .A1(n14433), .A2(n13864), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13401) );
  OAI21_X1 U15521 ( .B1(n13868), .B2(n14463), .A(n13401), .ZN(n13402) );
  AOI21_X1 U15522 ( .B1(n14045), .B2(n14447), .A(n13402), .ZN(n13403) );
  OAI21_X1 U15523 ( .B1(n13404), .B2(n14458), .A(n13403), .ZN(P1_U3240) );
  OAI211_X1 U15524 ( .C1(n13407), .C2(n13406), .A(n13405), .B(n14440), .ZN(
        n13413) );
  NAND2_X1 U15525 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14539)
         );
  OAI21_X1 U15526 ( .B1(n14456), .B2(n13408), .A(n14539), .ZN(n13409) );
  AOI21_X1 U15527 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13412) );
  OAI211_X1 U15528 ( .C1(n7089), .C2(n13414), .A(n13413), .B(n13412), .ZN(
        P1_U3241) );
  NOR2_X1 U15529 ( .A1(n13416), .A2(n13415), .ZN(n13420) );
  NAND4_X1 U15530 ( .A1(n13420), .A2(n13419), .A3(n13418), .A4(n13417), .ZN(
        n13421) );
  NOR3_X1 U15531 ( .A1(n14547), .A2(n13422), .A3(n13421), .ZN(n13424) );
  NAND4_X1 U15532 ( .A1(n13426), .A2(n13425), .A3(n13424), .A4(n13423), .ZN(
        n13427) );
  OR4_X1 U15533 ( .A1(n14266), .A2(n13429), .A3(n13428), .A4(n13427), .ZN(
        n13430) );
  XNOR2_X1 U15534 ( .A(n13435), .B(n13434), .ZN(n14006) );
  OR4_X1 U15535 ( .A1(n13437), .A2(n7224), .A3(n13436), .A4(n14006), .ZN(
        n13438) );
  NOR2_X1 U15536 ( .A1(n13930), .A2(n13440), .ZN(n13441) );
  NAND4_X1 U15537 ( .A1(n13890), .A2(n13441), .A3(n13895), .A4(n13909), .ZN(
        n13442) );
  NOR4_X1 U15538 ( .A1(n13443), .A2(n13857), .A3(n13871), .A4(n13442), .ZN(
        n13460) );
  NAND2_X1 U15539 ( .A1(n13445), .A2(n13444), .ZN(n13447) );
  NAND2_X1 U15540 ( .A1(n13455), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U15541 ( .A1(n10245), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U15542 ( .A1(n13448), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U15543 ( .A1(n11778), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n13450) );
  NAND3_X1 U15544 ( .A1(n13452), .A2(n13451), .A3(n13450), .ZN(n13828) );
  XNOR2_X1 U15545 ( .A(n13646), .B(n13828), .ZN(n13641) );
  NAND2_X1 U15546 ( .A1(n13455), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13456) );
  XNOR2_X1 U15547 ( .A(n13824), .B(n13667), .ZN(n13458) );
  NAND4_X1 U15548 ( .A1(n13460), .A2(n13459), .A3(n13641), .A4(n13458), .ZN(
        n13461) );
  XNOR2_X1 U15549 ( .A(n13461), .B(n13952), .ZN(n13659) );
  NAND2_X1 U15550 ( .A1(n13465), .A2(n13464), .ZN(n13613) );
  MUX2_X1 U15551 ( .A(n13669), .B(n14033), .S(n6825), .Z(n13622) );
  XNOR2_X1 U15552 ( .A(n13467), .B(n6620), .ZN(n13470) );
  NAND2_X1 U15553 ( .A1(n13470), .A2(n13469), .ZN(n13475) );
  MUX2_X1 U15554 ( .A(n13696), .B(n13473), .S(n6620), .Z(n13471) );
  NAND2_X1 U15555 ( .A1(n13696), .A2(n13473), .ZN(n13474) );
  NOR2_X1 U15556 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  OAI21_X1 U15557 ( .B1(n13477), .B2(n13476), .A(n14566), .ZN(n13485) );
  INV_X1 U15558 ( .A(n13478), .ZN(n13481) );
  INV_X1 U15559 ( .A(n13479), .ZN(n13480) );
  NAND2_X1 U15560 ( .A1(n13485), .A2(n13484), .ZN(n13489) );
  MUX2_X1 U15561 ( .A(n13487), .B(n13486), .S(n13596), .Z(n13488) );
  MUX2_X1 U15562 ( .A(n13490), .B(n14603), .S(n13596), .Z(n13493) );
  MUX2_X1 U15563 ( .A(n13491), .B(n13692), .S(n13596), .Z(n13492) );
  NAND2_X1 U15564 ( .A1(n13494), .A2(n13493), .ZN(n13495) );
  MUX2_X1 U15565 ( .A(n13497), .B(n13691), .S(n13596), .Z(n13499) );
  MUX2_X1 U15566 ( .A(n13691), .B(n13497), .S(n13596), .Z(n13498) );
  MUX2_X1 U15567 ( .A(n13690), .B(n14559), .S(n13596), .Z(n13502) );
  MUX2_X1 U15568 ( .A(n14559), .B(n13690), .S(n13596), .Z(n13500) );
  NAND2_X1 U15569 ( .A1(n13501), .A2(n13500), .ZN(n13505) );
  OR2_X1 U15570 ( .A1(n13503), .A2(n13502), .ZN(n13504) );
  MUX2_X1 U15571 ( .A(n13689), .B(n13506), .S(n6825), .Z(n13509) );
  NAND2_X1 U15572 ( .A1(n13510), .A2(n13509), .ZN(n13508) );
  NAND2_X1 U15573 ( .A1(n13508), .A2(n13507), .ZN(n13511) );
  MUX2_X1 U15574 ( .A(n13688), .B(n14635), .S(n13596), .Z(n13513) );
  MUX2_X1 U15575 ( .A(n13688), .B(n14635), .S(n6825), .Z(n13512) );
  MUX2_X1 U15576 ( .A(n13687), .B(n13514), .S(n6825), .Z(n13518) );
  NAND2_X1 U15577 ( .A1(n13517), .A2(n13518), .ZN(n13516) );
  MUX2_X1 U15578 ( .A(n13687), .B(n13514), .S(n13617), .Z(n13515) );
  MUX2_X1 U15579 ( .A(n13686), .B(n14653), .S(n13596), .Z(n13521) );
  MUX2_X1 U15580 ( .A(n13686), .B(n14653), .S(n6825), .Z(n13520) );
  MUX2_X1 U15581 ( .A(n13685), .B(n14450), .S(n6825), .Z(n13525) );
  NAND2_X1 U15582 ( .A1(n13524), .A2(n13525), .ZN(n13523) );
  MUX2_X1 U15583 ( .A(n13685), .B(n14450), .S(n13596), .Z(n13522) );
  NAND2_X1 U15584 ( .A1(n13523), .A2(n13522), .ZN(n13529) );
  INV_X1 U15585 ( .A(n13524), .ZN(n13527) );
  INV_X1 U15586 ( .A(n13525), .ZN(n13526) );
  NAND2_X1 U15587 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  MUX2_X1 U15588 ( .A(n13684), .B(n14274), .S(n13617), .Z(n13532) );
  MUX2_X1 U15589 ( .A(n13684), .B(n14274), .S(n6825), .Z(n13530) );
  MUX2_X1 U15590 ( .A(n13683), .B(n14476), .S(n6825), .Z(n13542) );
  NAND2_X1 U15591 ( .A1(n14476), .A2(n13617), .ZN(n13533) );
  OAI211_X1 U15592 ( .C1(n13534), .C2(n13617), .A(n13542), .B(n13533), .ZN(
        n13535) );
  AOI21_X1 U15593 ( .B1(n13549), .B2(n13537), .A(n13617), .ZN(n13541) );
  NAND2_X1 U15594 ( .A1(n14431), .A2(n13538), .ZN(n13539) );
  AOI21_X1 U15595 ( .B1(n13550), .B2(n13539), .A(n6825), .ZN(n13540) );
  NOR2_X1 U15596 ( .A1(n13541), .A2(n13540), .ZN(n13547) );
  INV_X1 U15597 ( .A(n13542), .ZN(n13544) );
  MUX2_X1 U15598 ( .A(n13683), .B(n14476), .S(n13617), .Z(n13543) );
  NAND3_X1 U15599 ( .A1(n13545), .A2(n13544), .A3(n13543), .ZN(n13546) );
  MUX2_X1 U15600 ( .A(n13550), .B(n13549), .S(n13596), .Z(n13551) );
  MUX2_X1 U15601 ( .A(n13680), .B(n14106), .S(n6825), .Z(n13555) );
  MUX2_X1 U15602 ( .A(n13680), .B(n14106), .S(n13617), .Z(n13553) );
  INV_X1 U15603 ( .A(n13553), .ZN(n13554) );
  NAND2_X1 U15604 ( .A1(n13556), .A2(n13555), .ZN(n13558) );
  MUX2_X1 U15605 ( .A(n13561), .B(n13560), .S(n13617), .Z(n13557) );
  MUX2_X1 U15606 ( .A(n13561), .B(n13560), .S(n6825), .Z(n13562) );
  MUX2_X1 U15607 ( .A(n13564), .B(n13563), .S(n6825), .Z(n13565) );
  NAND2_X1 U15608 ( .A1(n13567), .A2(n13566), .ZN(n13572) );
  OR2_X1 U15609 ( .A1(n14089), .A2(n13568), .ZN(n13570) );
  MUX2_X1 U15610 ( .A(n13570), .B(n13569), .S(n13617), .Z(n13571) );
  MUX2_X1 U15611 ( .A(n13573), .B(n13962), .S(n6825), .Z(n13576) );
  MUX2_X1 U15612 ( .A(n13573), .B(n13962), .S(n13617), .Z(n13574) );
  INV_X1 U15613 ( .A(n13574), .ZN(n13575) );
  NAND2_X1 U15614 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  MUX2_X1 U15615 ( .A(n13675), .B(n13954), .S(n13617), .Z(n13581) );
  MUX2_X1 U15616 ( .A(n13675), .B(n13954), .S(n6825), .Z(n13580) );
  MUX2_X1 U15617 ( .A(n13582), .B(n14072), .S(n6825), .Z(n13584) );
  MUX2_X1 U15618 ( .A(n15203), .B(n13937), .S(n13617), .Z(n13583) );
  AOI21_X1 U15619 ( .B1(n13585), .B2(n13584), .A(n13583), .ZN(n13587) );
  NOR2_X1 U15620 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  MUX2_X1 U15621 ( .A(n13674), .B(n13919), .S(n6825), .Z(n13588) );
  MUX2_X1 U15622 ( .A(n13673), .B(n13900), .S(n6825), .Z(n13592) );
  NAND2_X1 U15623 ( .A1(n13593), .A2(n13592), .ZN(n13591) );
  MUX2_X1 U15624 ( .A(n13673), .B(n13900), .S(n13617), .Z(n13590) );
  NAND2_X1 U15625 ( .A1(n13591), .A2(n13590), .ZN(n13595) );
  MUX2_X1 U15626 ( .A(n13672), .B(n14051), .S(n13596), .Z(n13599) );
  MUX2_X1 U15627 ( .A(n13672), .B(n14051), .S(n6825), .Z(n13597) );
  NAND2_X1 U15628 ( .A1(n13598), .A2(n13597), .ZN(n13601) );
  MUX2_X1 U15629 ( .A(n13671), .B(n14045), .S(n6825), .Z(n13603) );
  MUX2_X1 U15630 ( .A(n13671), .B(n14045), .S(n13617), .Z(n13602) );
  MUX2_X1 U15631 ( .A(n13670), .B(n14040), .S(n13596), .Z(n13607) );
  NAND2_X1 U15632 ( .A1(n13606), .A2(n13607), .ZN(n13605) );
  MUX2_X1 U15633 ( .A(n14040), .B(n13670), .S(n13617), .Z(n13604) );
  INV_X1 U15634 ( .A(n13606), .ZN(n13609) );
  INV_X1 U15635 ( .A(n13607), .ZN(n13608) );
  MUX2_X1 U15636 ( .A(n13669), .B(n14033), .S(n13617), .Z(n13610) );
  NAND2_X1 U15637 ( .A1(n13828), .A2(n13617), .ZN(n13612) );
  AOI21_X1 U15638 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13614) );
  AOI21_X1 U15639 ( .B1(n13824), .B2(n6825), .A(n13614), .ZN(n13629) );
  OAI21_X1 U15640 ( .B1(n13828), .B2(n13615), .A(n13667), .ZN(n13616) );
  INV_X1 U15641 ( .A(n13616), .ZN(n13618) );
  MUX2_X1 U15642 ( .A(n13618), .B(n13824), .S(n13617), .Z(n13627) );
  INV_X1 U15643 ( .A(n13668), .ZN(n13620) );
  MUX2_X1 U15644 ( .A(n13620), .B(n13619), .S(n6825), .Z(n13624) );
  MUX2_X1 U15645 ( .A(n13668), .B(n14029), .S(n13617), .Z(n13623) );
  AOI22_X1 U15646 ( .A1(n13629), .A2(n13627), .B1(n13624), .B2(n13623), .ZN(
        n13621) );
  INV_X1 U15647 ( .A(n13623), .ZN(n13626) );
  INV_X1 U15648 ( .A(n13624), .ZN(n13625) );
  NAND2_X1 U15649 ( .A1(n13626), .A2(n13625), .ZN(n13628) );
  NAND2_X1 U15650 ( .A1(n13629), .A2(n13628), .ZN(n13633) );
  INV_X1 U15651 ( .A(n13627), .ZN(n13632) );
  INV_X1 U15652 ( .A(n13628), .ZN(n13631) );
  INV_X1 U15653 ( .A(n13629), .ZN(n13630) );
  AOI22_X1 U15654 ( .A1(n13633), .A2(n13632), .B1(n13631), .B2(n13630), .ZN(
        n13634) );
  NAND2_X1 U15655 ( .A1(n9433), .A2(n13636), .ZN(n13637) );
  NAND2_X1 U15656 ( .A1(n13638), .A2(n13637), .ZN(n13640) );
  NAND2_X1 U15657 ( .A1(n13639), .A2(n13952), .ZN(n14275) );
  NAND2_X1 U15658 ( .A1(n13640), .A2(n14275), .ZN(n13645) );
  INV_X1 U15659 ( .A(n13645), .ZN(n13642) );
  OR2_X1 U15660 ( .A1(n13646), .A2(n13596), .ZN(n13653) );
  XNOR2_X1 U15661 ( .A(n13653), .B(n13645), .ZN(n13643) );
  NAND4_X1 U15662 ( .A1(n13643), .A2(n14022), .A3(n13828), .A4(n13644), .ZN(
        n13650) );
  AND2_X1 U15663 ( .A1(n13646), .A2(n13596), .ZN(n13656) );
  INV_X1 U15664 ( .A(n13656), .ZN(n13647) );
  OR3_X1 U15665 ( .A1(n13647), .A2(n13828), .A3(n13645), .ZN(n13649) );
  INV_X1 U15666 ( .A(n13828), .ZN(n13657) );
  AND2_X1 U15667 ( .A1(n13645), .A2(n13644), .ZN(n13652) );
  NAND4_X1 U15668 ( .A1(n13647), .A2(n13657), .A3(n13652), .A4(n13646), .ZN(
        n13648) );
  OAI21_X1 U15669 ( .B1(n13653), .B2(n13657), .A(n13652), .ZN(n13655) );
  AOI211_X1 U15670 ( .C1(n13657), .C2(n13656), .A(n13655), .B(n13654), .ZN(
        n13658) );
  NOR2_X1 U15671 ( .A1(n14142), .A2(P1_U3086), .ZN(n13661) );
  NAND3_X1 U15672 ( .A1(n13663), .A2(n13662), .A3(n13661), .ZN(n13664) );
  OAI211_X1 U15673 ( .C1(n6847), .C2(n13666), .A(n13664), .B(P1_B_REG_SCAN_IN), 
        .ZN(n13665) );
  MUX2_X1 U15674 ( .A(n13828), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13695), .Z(
        P1_U3591) );
  MUX2_X1 U15675 ( .A(n13667), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13695), .Z(
        P1_U3590) );
  MUX2_X1 U15676 ( .A(n13668), .B(P1_DATAO_REG_29__SCAN_IN), .S(n13695), .Z(
        P1_U3589) );
  MUX2_X1 U15677 ( .A(n13669), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13695), .Z(
        P1_U3588) );
  MUX2_X1 U15678 ( .A(n13670), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13695), .Z(
        P1_U3587) );
  MUX2_X1 U15679 ( .A(n13671), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13695), .Z(
        P1_U3586) );
  MUX2_X1 U15680 ( .A(n13672), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13695), .Z(
        P1_U3585) );
  MUX2_X1 U15681 ( .A(n13673), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13695), .Z(
        P1_U3584) );
  MUX2_X1 U15682 ( .A(n13674), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13695), .Z(
        P1_U3583) );
  MUX2_X1 U15683 ( .A(n13675), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13695), .Z(
        P1_U3581) );
  MUX2_X1 U15684 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13676), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15685 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13677), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15686 ( .A(n13678), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13695), .Z(
        P1_U3578) );
  MUX2_X1 U15687 ( .A(n13679), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13695), .Z(
        P1_U3577) );
  MUX2_X1 U15688 ( .A(n13680), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13695), .Z(
        P1_U3576) );
  MUX2_X1 U15689 ( .A(n13681), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13695), .Z(
        P1_U3575) );
  MUX2_X1 U15690 ( .A(n13682), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13695), .Z(
        P1_U3574) );
  MUX2_X1 U15691 ( .A(n13683), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13695), .Z(
        P1_U3573) );
  MUX2_X1 U15692 ( .A(n13684), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13695), .Z(
        P1_U3572) );
  MUX2_X1 U15693 ( .A(n13685), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13695), .Z(
        P1_U3571) );
  MUX2_X1 U15694 ( .A(n13686), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13695), .Z(
        P1_U3570) );
  MUX2_X1 U15695 ( .A(n13687), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13695), .Z(
        P1_U3569) );
  MUX2_X1 U15696 ( .A(n13688), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13695), .Z(
        P1_U3568) );
  MUX2_X1 U15697 ( .A(n13689), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13695), .Z(
        P1_U3567) );
  MUX2_X1 U15698 ( .A(n13690), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13695), .Z(
        P1_U3566) );
  MUX2_X1 U15699 ( .A(n13691), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13695), .Z(
        P1_U3565) );
  MUX2_X1 U15700 ( .A(n13692), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13695), .Z(
        P1_U3564) );
  MUX2_X1 U15701 ( .A(n13693), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13695), .Z(
        P1_U3563) );
  MUX2_X1 U15702 ( .A(n13694), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13695), .Z(
        P1_U3562) );
  MUX2_X1 U15703 ( .A(n13696), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13695), .Z(
        P1_U3561) );
  MUX2_X1 U15704 ( .A(n13698), .B(n13697), .S(n14142), .Z(n13702) );
  INV_X1 U15705 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U15706 ( .A1(n14517), .A2(n13699), .ZN(n13700) );
  NAND2_X1 U15707 ( .A1(n13701), .A2(n13700), .ZN(n14518) );
  INV_X1 U15708 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14520) );
  NAND2_X1 U15709 ( .A1(n14518), .A2(n14520), .ZN(n14523) );
  OAI211_X1 U15710 ( .C1(n13702), .C2(n9233), .A(P1_U4016), .B(n14523), .ZN(
        n13747) );
  AOI22_X1 U15711 ( .A1(n14525), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13715) );
  OAI21_X1 U15712 ( .B1(n13704), .B2(n13703), .A(n13718), .ZN(n13710) );
  MUX2_X1 U15713 ( .A(n9205), .B(P1_REG1_REG_2__SCAN_IN), .S(n13712), .Z(
        n13707) );
  INV_X1 U15714 ( .A(n13705), .ZN(n13706) );
  NAND2_X1 U15715 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  NAND3_X1 U15716 ( .A1(n13819), .A2(n13723), .A3(n13708), .ZN(n13709) );
  OAI21_X1 U15717 ( .B1(n14534), .B2(n13710), .A(n13709), .ZN(n13711) );
  INV_X1 U15718 ( .A(n13711), .ZN(n13714) );
  NAND2_X1 U15719 ( .A1(n13817), .A2(n13712), .ZN(n13713) );
  NAND4_X1 U15720 ( .A1(n13747), .A2(n13715), .A3(n13714), .A4(n13713), .ZN(
        P1_U3245) );
  MUX2_X1 U15721 ( .A(n15054), .B(P1_REG2_REG_3__SCAN_IN), .S(n13720), .Z(
        n13716) );
  NAND3_X1 U15722 ( .A1(n13718), .A2(n13717), .A3(n13716), .ZN(n13719) );
  NAND3_X1 U15723 ( .A1(n13813), .A2(n13742), .A3(n13719), .ZN(n13728) );
  AOI22_X1 U15724 ( .A1(n14525), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13727) );
  NAND2_X1 U15725 ( .A1(n13817), .A2(n13720), .ZN(n13726) );
  MUX2_X1 U15726 ( .A(n9212), .B(P1_REG1_REG_3__SCAN_IN), .S(n13720), .Z(
        n13721) );
  NAND3_X1 U15727 ( .A1(n13723), .A2(n13722), .A3(n13721), .ZN(n13724) );
  NAND3_X1 U15728 ( .A1(n13819), .A2(n13736), .A3(n13724), .ZN(n13725) );
  NAND4_X1 U15729 ( .A1(n13728), .A2(n13727), .A3(n13726), .A4(n13725), .ZN(
        P1_U3246) );
  NAND2_X1 U15730 ( .A1(n14525), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U15731 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  AOI21_X1 U15732 ( .B1(n13732), .B2(n13817), .A(n13731), .ZN(n13746) );
  INV_X1 U15733 ( .A(n13733), .ZN(n13738) );
  NAND3_X1 U15734 ( .A1(n13736), .A2(n13735), .A3(n13734), .ZN(n13737) );
  NAND3_X1 U15735 ( .A1(n13819), .A2(n13738), .A3(n13737), .ZN(n13745) );
  INV_X1 U15736 ( .A(n13739), .ZN(n13759) );
  NAND3_X1 U15737 ( .A1(n13742), .A2(n13741), .A3(n13740), .ZN(n13743) );
  NAND3_X1 U15738 ( .A1(n13813), .A2(n13759), .A3(n13743), .ZN(n13744) );
  NAND4_X1 U15739 ( .A1(n13747), .A2(n13746), .A3(n13745), .A4(n13744), .ZN(
        P1_U3247) );
  INV_X1 U15740 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U15741 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13748) );
  OAI21_X1 U15742 ( .B1(n14541), .B2(n14160), .A(n13748), .ZN(n13749) );
  AOI21_X1 U15743 ( .B1(n13750), .B2(n13817), .A(n13749), .ZN(n13764) );
  OAI21_X1 U15744 ( .B1(n13753), .B2(n13752), .A(n13751), .ZN(n13754) );
  NAND2_X1 U15745 ( .A1(n13819), .A2(n13754), .ZN(n13763) );
  INV_X1 U15746 ( .A(n13755), .ZN(n13758) );
  MUX2_X1 U15747 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10387), .S(n13756), .Z(
        n13757) );
  NAND3_X1 U15748 ( .A1(n13759), .A2(n13758), .A3(n13757), .ZN(n13760) );
  NAND3_X1 U15749 ( .A1(n13813), .A2(n13761), .A3(n13760), .ZN(n13762) );
  NAND3_X1 U15750 ( .A1(n13764), .A2(n13763), .A3(n13762), .ZN(P1_U3248) );
  INV_X1 U15751 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13766) );
  OAI21_X1 U15752 ( .B1(n14541), .B2(n13766), .A(n13765), .ZN(n13767) );
  AOI21_X1 U15753 ( .B1(n13775), .B2(n13817), .A(n13767), .ZN(n13783) );
  INV_X1 U15754 ( .A(n13768), .ZN(n13770) );
  MUX2_X1 U15755 ( .A(n14671), .B(P1_REG1_REG_7__SCAN_IN), .S(n13775), .Z(
        n13769) );
  NAND2_X1 U15756 ( .A1(n13770), .A2(n13769), .ZN(n13772) );
  OAI211_X1 U15757 ( .C1(n13773), .C2(n13772), .A(n13819), .B(n13771), .ZN(
        n13782) );
  INV_X1 U15758 ( .A(n13774), .ZN(n13777) );
  MUX2_X1 U15759 ( .A(n10537), .B(P1_REG2_REG_7__SCAN_IN), .S(n13775), .Z(
        n13776) );
  NAND2_X1 U15760 ( .A1(n13777), .A2(n13776), .ZN(n13779) );
  OAI211_X1 U15761 ( .C1(n13780), .C2(n13779), .A(n13813), .B(n13778), .ZN(
        n13781) );
  NAND3_X1 U15762 ( .A1(n13783), .A2(n13782), .A3(n13781), .ZN(P1_U3250) );
  INV_X1 U15763 ( .A(n13784), .ZN(n13789) );
  NOR3_X1 U15764 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(n13788) );
  OAI21_X1 U15765 ( .B1(n13789), .B2(n13788), .A(n13819), .ZN(n13801) );
  INV_X1 U15766 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14172) );
  NAND2_X1 U15767 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13790) );
  OAI21_X1 U15768 ( .B1(n14541), .B2(n14172), .A(n13790), .ZN(n13791) );
  AOI21_X1 U15769 ( .B1(n13792), .B2(n13817), .A(n13791), .ZN(n13800) );
  MUX2_X1 U15770 ( .A(n9493), .B(P1_REG2_REG_9__SCAN_IN), .S(n13792), .Z(
        n13795) );
  INV_X1 U15771 ( .A(n13793), .ZN(n13794) );
  NAND2_X1 U15772 ( .A1(n13795), .A2(n13794), .ZN(n13797) );
  OAI211_X1 U15773 ( .C1(n13798), .C2(n13797), .A(n13796), .B(n13813), .ZN(
        n13799) );
  NAND3_X1 U15774 ( .A1(n13801), .A2(n13800), .A3(n13799), .ZN(P1_U3252) );
  INV_X1 U15775 ( .A(n13802), .ZN(n13803) );
  NAND2_X1 U15776 ( .A1(n13808), .A2(n13803), .ZN(n13804) );
  NAND2_X1 U15777 ( .A1(n13805), .A2(n13804), .ZN(n13806) );
  XOR2_X1 U15778 ( .A(n13806), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13815) );
  NAND2_X1 U15779 ( .A1(n13808), .A2(n13807), .ZN(n13809) );
  NAND2_X1 U15780 ( .A1(n13810), .A2(n13809), .ZN(n13812) );
  XNOR2_X1 U15781 ( .A(n13812), .B(n13811), .ZN(n13814) );
  AOI22_X1 U15782 ( .A1(n13815), .A2(n13813), .B1(n13814), .B2(n13819), .ZN(
        n13820) );
  INV_X1 U15783 ( .A(n13814), .ZN(n13818) );
  NOR2_X1 U15784 ( .A1(n13815), .A2(n14534), .ZN(n13816) );
  INV_X1 U15785 ( .A(n13821), .ZN(n13822) );
  OAI211_X1 U15786 ( .C1(n7580), .C2(n14541), .A(n13823), .B(n13822), .ZN(
        P1_U3262) );
  NAND2_X1 U15787 ( .A1(n13832), .A2(n14025), .ZN(n13831) );
  XNOR2_X1 U15788 ( .A(n13831), .B(n14022), .ZN(n14021) );
  NAND2_X1 U15789 ( .A1(n14021), .A2(n13825), .ZN(n13830) );
  INV_X1 U15790 ( .A(n13826), .ZN(n13827) );
  NAND2_X1 U15791 ( .A1(n13828), .A2(n13827), .ZN(n14023) );
  NOR2_X1 U15792 ( .A1(n14276), .A2(n14023), .ZN(n13834) );
  AOI21_X1 U15793 ( .B1(n14276), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13834), 
        .ZN(n13829) );
  OAI211_X1 U15794 ( .C1(n14022), .C2(n14012), .A(n13830), .B(n13829), .ZN(
        P1_U3263) );
  OAI211_X1 U15795 ( .C1(n13832), .C2(n14025), .A(n14577), .B(n13831), .ZN(
        n14024) );
  NOR2_X1 U15796 ( .A1(n14025), .A2(n14012), .ZN(n13833) );
  AOI211_X1 U15797 ( .C1(n14276), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13834), 
        .B(n13833), .ZN(n13835) );
  OAI21_X1 U15798 ( .B1(n14016), .B2(n14024), .A(n13835), .ZN(P1_U3264) );
  XNOR2_X1 U15799 ( .A(n13836), .B(n13845), .ZN(n13838) );
  OAI22_X1 U15800 ( .A1(n14002), .A2(n15271), .B1(n13839), .B2(n14010), .ZN(
        n13843) );
  OAI211_X1 U15801 ( .C1(n13841), .C2(n13851), .A(n14577), .B(n13840), .ZN(
        n14035) );
  NOR2_X1 U15802 ( .A1(n14035), .A2(n14016), .ZN(n13842) );
  AOI211_X1 U15803 ( .C1(n14572), .C2(n14033), .A(n13843), .B(n13842), .ZN(
        n13847) );
  NAND2_X1 U15804 ( .A1(n13845), .A2(n13844), .ZN(n14034) );
  NAND3_X1 U15805 ( .A1(n6606), .A2(n13922), .A3(n14034), .ZN(n13846) );
  OAI211_X1 U15806 ( .C1(n14038), .C2(n14276), .A(n13847), .B(n13846), .ZN(
        P1_U3265) );
  XNOR2_X1 U15807 ( .A(n13848), .B(n13857), .ZN(n13850) );
  AOI211_X1 U15808 ( .C1(n14040), .C2(n13866), .A(n6570), .B(n13851), .ZN(
        n14039) );
  INV_X1 U15809 ( .A(n13852), .ZN(n13853) );
  AOI22_X1 U15810 ( .A1(n14276), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13853), 
        .B2(n14574), .ZN(n13854) );
  OAI21_X1 U15811 ( .B1(n13855), .B2(n14012), .A(n13854), .ZN(n13861) );
  OAI21_X1 U15812 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13859) );
  INV_X1 U15813 ( .A(n13859), .ZN(n14043) );
  NOR2_X1 U15814 ( .A1(n14043), .A2(n14020), .ZN(n13860) );
  AOI211_X1 U15815 ( .C1(n14039), .C2(n14581), .A(n13861), .B(n13860), .ZN(
        n13862) );
  OAI21_X1 U15816 ( .B1(n14042), .B2(n14575), .A(n13862), .ZN(P1_U3266) );
  XNOR2_X1 U15817 ( .A(n13863), .B(n7166), .ZN(n13865) );
  AOI21_X1 U15818 ( .B1(n13865), .B2(n14571), .A(n13864), .ZN(n14047) );
  INV_X1 U15819 ( .A(n13866), .ZN(n13867) );
  AOI211_X1 U15820 ( .C1(n14045), .C2(n13880), .A(n6570), .B(n13867), .ZN(
        n14044) );
  INV_X1 U15821 ( .A(n13868), .ZN(n13869) );
  AOI22_X1 U15822 ( .A1(n14276), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13869), 
        .B2(n14574), .ZN(n13870) );
  OAI21_X1 U15823 ( .B1(n7085), .B2(n14012), .A(n13870), .ZN(n13876) );
  NOR2_X1 U15824 ( .A1(n13872), .A2(n13871), .ZN(n13873) );
  NOR2_X1 U15825 ( .A1(n14048), .A2(n14020), .ZN(n13875) );
  AOI211_X1 U15826 ( .C1(n14044), .C2(n14581), .A(n13876), .B(n13875), .ZN(
        n13877) );
  OAI21_X1 U15827 ( .B1(n14047), .B2(n14575), .A(n13877), .ZN(P1_U3267) );
  OAI21_X1 U15828 ( .B1(n13879), .B2(n13890), .A(n13878), .ZN(n14049) );
  INV_X1 U15829 ( .A(n14049), .ZN(n13894) );
  AOI21_X1 U15830 ( .B1(n13901), .B2(n14051), .A(n6570), .ZN(n13881) );
  NAND2_X1 U15831 ( .A1(n13881), .A2(n13880), .ZN(n14053) );
  INV_X1 U15832 ( .A(n14053), .ZN(n13888) );
  INV_X1 U15833 ( .A(n14050), .ZN(n13883) );
  OAI22_X1 U15834 ( .A1(n14575), .A2(n13883), .B1(n13882), .B2(n14010), .ZN(
        n13884) );
  AOI21_X1 U15835 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14276), .A(n13884), 
        .ZN(n13885) );
  OAI21_X1 U15836 ( .B1(n13886), .B2(n14012), .A(n13885), .ZN(n13887) );
  AOI21_X1 U15837 ( .B1(n13888), .B2(n14581), .A(n13887), .ZN(n13893) );
  NAND2_X1 U15838 ( .A1(n13891), .A2(n13890), .ZN(n14052) );
  NAND3_X1 U15839 ( .A1(n13889), .A2(n14052), .A3(n13922), .ZN(n13892) );
  OAI211_X1 U15840 ( .C1(n13894), .C2(n13924), .A(n13893), .B(n13892), .ZN(
        P1_U3268) );
  XNOR2_X1 U15841 ( .A(n13896), .B(n13895), .ZN(n14062) );
  AOI211_X1 U15842 ( .C1(n13899), .C2(n13898), .A(n14550), .B(n13897), .ZN(
        n14060) );
  OAI21_X1 U15843 ( .B1(n14060), .B2(n14057), .A(n14002), .ZN(n13908) );
  AOI21_X1 U15844 ( .B1(n13914), .B2(n13900), .A(n6570), .ZN(n13902) );
  AND2_X1 U15845 ( .A1(n13902), .A2(n13901), .ZN(n14059) );
  INV_X1 U15846 ( .A(n13903), .ZN(n13904) );
  AOI22_X1 U15847 ( .A1(n14276), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13904), 
        .B2(n14574), .ZN(n13905) );
  OAI21_X1 U15848 ( .B1(n7087), .B2(n14012), .A(n13905), .ZN(n13906) );
  AOI21_X1 U15849 ( .B1(n14059), .B2(n14581), .A(n13906), .ZN(n13907) );
  OAI211_X1 U15850 ( .C1(n14020), .C2(n14062), .A(n13908), .B(n13907), .ZN(
        P1_U3269) );
  XNOR2_X1 U15851 ( .A(n13910), .B(n13909), .ZN(n14069) );
  XNOR2_X1 U15852 ( .A(n13912), .B(n13911), .ZN(n14067) );
  AOI21_X1 U15853 ( .B1(n13919), .B2(n13913), .A(n6570), .ZN(n13915) );
  NAND2_X1 U15854 ( .A1(n13915), .A2(n13914), .ZN(n14064) );
  AOI22_X1 U15855 ( .A1(n14276), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13916), 
        .B2(n14574), .ZN(n13917) );
  OAI21_X1 U15856 ( .B1(n14063), .B2(n14575), .A(n13917), .ZN(n13918) );
  AOI21_X1 U15857 ( .B1(n13919), .B2(n14572), .A(n13918), .ZN(n13920) );
  OAI21_X1 U15858 ( .B1(n14064), .B2(n14016), .A(n13920), .ZN(n13921) );
  AOI21_X1 U15859 ( .B1(n14067), .B2(n13922), .A(n13921), .ZN(n13923) );
  OAI21_X1 U15860 ( .B1(n14069), .B2(n13924), .A(n13923), .ZN(P1_U3270) );
  OAI21_X1 U15861 ( .B1(n13930), .B2(n13926), .A(n13925), .ZN(n13927) );
  INV_X1 U15862 ( .A(n13927), .ZN(n14075) );
  AOI21_X1 U15863 ( .B1(n13930), .B2(n13929), .A(n13928), .ZN(n13931) );
  INV_X1 U15864 ( .A(n14074), .ZN(n13932) );
  OAI21_X1 U15865 ( .B1(n13932), .B2(n14071), .A(n14002), .ZN(n13940) );
  XNOR2_X1 U15866 ( .A(n13937), .B(n13933), .ZN(n13934) );
  AND2_X1 U15867 ( .A1(n13934), .A2(n14577), .ZN(n14070) );
  AOI22_X1 U15868 ( .A1(n13935), .A2(n14574), .B1(n14575), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n13936) );
  OAI21_X1 U15869 ( .B1(n13937), .B2(n14012), .A(n13936), .ZN(n13938) );
  AOI21_X1 U15870 ( .B1(n14070), .B2(n14581), .A(n13938), .ZN(n13939) );
  OAI211_X1 U15871 ( .C1(n14075), .C2(n14020), .A(n13940), .B(n13939), .ZN(
        P1_U3271) );
  INV_X1 U15872 ( .A(n13941), .ZN(n13942) );
  AOI21_X1 U15873 ( .B1(n13946), .B2(n13943), .A(n13942), .ZN(n14081) );
  AOI211_X1 U15874 ( .C1(n13954), .C2(n13964), .A(n6570), .B(n13944), .ZN(
        n14078) );
  INV_X1 U15875 ( .A(n14078), .ZN(n13951) );
  OAI211_X1 U15876 ( .C1(n13947), .C2(n13946), .A(n14571), .B(n13945), .ZN(
        n14080) );
  INV_X1 U15877 ( .A(n13948), .ZN(n13949) );
  AOI21_X1 U15878 ( .B1(n13949), .B2(n14574), .A(n14076), .ZN(n13950) );
  OAI211_X1 U15879 ( .C1(n13952), .C2(n13951), .A(n14080), .B(n13950), .ZN(
        n13953) );
  NAND2_X1 U15880 ( .A1(n13953), .A2(n14002), .ZN(n13956) );
  AOI22_X1 U15881 ( .A1(n13954), .A2(n14572), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14575), .ZN(n13955) );
  OAI211_X1 U15882 ( .C1(n14081), .C2(n14020), .A(n13956), .B(n13955), .ZN(
        P1_U3272) );
  OAI21_X1 U15883 ( .B1(n6703), .B2(n13958), .A(n13957), .ZN(n14086) );
  AOI21_X1 U15884 ( .B1(n6704), .B2(n13958), .A(n14550), .ZN(n13961) );
  AOI21_X1 U15885 ( .B1(n13961), .B2(n13960), .A(n13959), .ZN(n14085) );
  OR2_X1 U15886 ( .A1(n13962), .A2(n13980), .ZN(n13963) );
  AND3_X1 U15887 ( .A1(n13964), .A2(n14577), .A3(n13963), .ZN(n14082) );
  NAND2_X1 U15888 ( .A1(n14082), .A2(n13965), .ZN(n13966) );
  OAI211_X1 U15889 ( .C1(n14010), .C2(n13967), .A(n14085), .B(n13966), .ZN(
        n13968) );
  NAND2_X1 U15890 ( .A1(n13968), .A2(n14002), .ZN(n13970) );
  AOI22_X1 U15891 ( .A1(n14083), .A2(n14572), .B1(n14575), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n13969) );
  OAI211_X1 U15892 ( .C1(n14086), .C2(n14020), .A(n13970), .B(n13969), .ZN(
        P1_U3273) );
  XNOR2_X1 U15893 ( .A(n13971), .B(n13974), .ZN(n14091) );
  AOI21_X1 U15894 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13977) );
  INV_X1 U15895 ( .A(n13975), .ZN(n13976) );
  OAI21_X1 U15896 ( .B1(n13977), .B2(n14550), .A(n13976), .ZN(n14087) );
  NAND2_X1 U15897 ( .A1(n6596), .A2(n14089), .ZN(n13978) );
  NAND2_X1 U15898 ( .A1(n13978), .A2(n14577), .ZN(n13979) );
  NOR2_X1 U15899 ( .A1(n13980), .A2(n13979), .ZN(n14088) );
  NAND2_X1 U15900 ( .A1(n14088), .A2(n14581), .ZN(n13985) );
  NAND2_X1 U15901 ( .A1(n14575), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n13981) );
  OAI21_X1 U15902 ( .B1(n14010), .B2(n13982), .A(n13981), .ZN(n13983) );
  AOI21_X1 U15903 ( .B1(n14089), .B2(n14572), .A(n13983), .ZN(n13984) );
  NAND2_X1 U15904 ( .A1(n13985), .A2(n13984), .ZN(n13986) );
  AOI21_X1 U15905 ( .B1(n14087), .B2(n14002), .A(n13986), .ZN(n13987) );
  OAI21_X1 U15906 ( .B1(n14091), .B2(n14020), .A(n13987), .ZN(P1_U3274) );
  XNOR2_X1 U15907 ( .A(n13988), .B(n13990), .ZN(n14096) );
  OAI211_X1 U15908 ( .C1(n13991), .C2(n13990), .A(n13989), .B(n14571), .ZN(
        n13994) );
  INV_X1 U15909 ( .A(n13992), .ZN(n13993) );
  NAND2_X1 U15910 ( .A1(n13994), .A2(n13993), .ZN(n14092) );
  AOI21_X1 U15911 ( .B1(n14007), .B2(n14094), .A(n6570), .ZN(n13995) );
  AND2_X1 U15912 ( .A1(n13995), .A2(n6596), .ZN(n14093) );
  NAND2_X1 U15913 ( .A1(n14093), .A2(n14581), .ZN(n14000) );
  NAND2_X1 U15914 ( .A1(n14575), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n13996) );
  OAI21_X1 U15915 ( .B1(n14010), .B2(n13997), .A(n13996), .ZN(n13998) );
  AOI21_X1 U15916 ( .B1(n14094), .B2(n14572), .A(n13998), .ZN(n13999) );
  NAND2_X1 U15917 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  AOI21_X1 U15918 ( .B1(n14092), .B2(n14002), .A(n14001), .ZN(n14003) );
  OAI21_X1 U15919 ( .B1(n14020), .B2(n14096), .A(n14003), .ZN(P1_U3275) );
  XNOR2_X1 U15920 ( .A(n14004), .B(n14006), .ZN(n14103) );
  XOR2_X1 U15921 ( .A(n14006), .B(n14005), .Z(n14101) );
  OAI211_X1 U15922 ( .C1(n14008), .C2(n14099), .A(n14577), .B(n14007), .ZN(
        n14098) );
  INV_X1 U15923 ( .A(n14009), .ZN(n14097) );
  OAI22_X1 U15924 ( .A1(n14097), .A2(n14276), .B1(n14011), .B2(n14010), .ZN(
        n14014) );
  NOR2_X1 U15925 ( .A1(n14099), .A2(n14012), .ZN(n14013) );
  AOI211_X1 U15926 ( .C1(n14575), .C2(P1_REG2_REG_17__SCAN_IN), .A(n14014), 
        .B(n14013), .ZN(n14015) );
  OAI21_X1 U15927 ( .B1(n14098), .B2(n14016), .A(n14015), .ZN(n14017) );
  AOI21_X1 U15928 ( .B1(n14101), .B2(n14018), .A(n14017), .ZN(n14019) );
  OAI21_X1 U15929 ( .B1(n14103), .B2(n14020), .A(n14019), .ZN(P1_U3276) );
  MUX2_X1 U15930 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14117), .S(n14679), .Z(
        P1_U3559) );
  OAI211_X1 U15931 ( .C1(n14025), .C2(n14655), .A(n14024), .B(n14023), .ZN(
        n14118) );
  MUX2_X1 U15932 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14118), .S(n14679), .Z(
        P1_U3558) );
  NAND3_X1 U15933 ( .A1(n14032), .A2(n14031), .A3(n14030), .ZN(n14119) );
  MUX2_X1 U15934 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14119), .S(n14679), .Z(
        P1_U3557) );
  NAND2_X1 U15935 ( .A1(n14033), .A2(n14636), .ZN(n14037) );
  NAND3_X1 U15936 ( .A1(n6606), .A2(n14660), .A3(n14034), .ZN(n14036) );
  NAND4_X1 U15937 ( .A1(n14038), .A2(n14037), .A3(n14036), .A4(n14035), .ZN(
        n14120) );
  MUX2_X1 U15938 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14120), .S(n14679), .Z(
        P1_U3556) );
  AOI21_X1 U15939 ( .B1(n14636), .B2(n14040), .A(n14039), .ZN(n14041) );
  OAI211_X1 U15940 ( .C1(n14639), .C2(n14043), .A(n14042), .B(n14041), .ZN(
        n14121) );
  MUX2_X1 U15941 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14121), .S(n14679), .Z(
        P1_U3555) );
  AOI21_X1 U15942 ( .B1(n14636), .B2(n14045), .A(n14044), .ZN(n14046) );
  OAI211_X1 U15943 ( .C1(n14639), .C2(n14048), .A(n14047), .B(n14046), .ZN(
        n14122) );
  MUX2_X1 U15944 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14122), .S(n14679), .Z(
        P1_U3554) );
  NAND2_X1 U15945 ( .A1(n14049), .A2(n14571), .ZN(n14056) );
  AOI21_X1 U15946 ( .B1(n14051), .B2(n14636), .A(n14050), .ZN(n14055) );
  NAND3_X1 U15947 ( .A1(n13889), .A2(n14660), .A3(n14052), .ZN(n14054) );
  NAND4_X1 U15948 ( .A1(n14056), .A2(n14055), .A3(n14054), .A4(n14053), .ZN(
        n14123) );
  MUX2_X1 U15949 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14123), .S(n14679), .Z(
        P1_U3553) );
  NOR4_X1 U15950 ( .A1(n14060), .A2(n14059), .A3(n14058), .A4(n14057), .ZN(
        n14061) );
  OAI21_X1 U15951 ( .B1(n14639), .B2(n14062), .A(n14061), .ZN(n14124) );
  MUX2_X1 U15952 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14124), .S(n14679), .Z(
        P1_U3552) );
  OAI211_X1 U15953 ( .C1(n14065), .C2(n14655), .A(n14064), .B(n14063), .ZN(
        n14066) );
  AOI21_X1 U15954 ( .B1(n14067), .B2(n14660), .A(n14066), .ZN(n14068) );
  OAI21_X1 U15955 ( .B1(n14069), .B2(n14550), .A(n14068), .ZN(n14125) );
  MUX2_X1 U15956 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14125), .S(n14679), .Z(
        P1_U3551) );
  AOI211_X1 U15957 ( .C1(n14636), .C2(n14072), .A(n14071), .B(n14070), .ZN(
        n14073) );
  OAI211_X1 U15958 ( .C1(n14639), .C2(n14075), .A(n14074), .B(n14073), .ZN(
        n14126) );
  MUX2_X1 U15959 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14126), .S(n14679), .Z(
        P1_U3550) );
  NOR3_X1 U15960 ( .A1(n14078), .A2(n14077), .A3(n14076), .ZN(n14079) );
  OAI211_X1 U15961 ( .C1(n14081), .C2(n14639), .A(n14080), .B(n14079), .ZN(
        n14127) );
  MUX2_X1 U15962 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14127), .S(n14679), .Z(
        P1_U3549) );
  AOI21_X1 U15963 ( .B1(n14636), .B2(n14083), .A(n14082), .ZN(n14084) );
  OAI211_X1 U15964 ( .C1(n14639), .C2(n14086), .A(n14085), .B(n14084), .ZN(
        n14128) );
  MUX2_X1 U15965 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14128), .S(n14679), .Z(
        P1_U3548) );
  AOI211_X1 U15966 ( .C1(n14636), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        n14090) );
  OAI21_X1 U15967 ( .B1(n14639), .B2(n14091), .A(n14090), .ZN(n14129) );
  MUX2_X1 U15968 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14129), .S(n14679), .Z(
        P1_U3547) );
  AOI211_X1 U15969 ( .C1(n14636), .C2(n14094), .A(n14093), .B(n14092), .ZN(
        n14095) );
  OAI21_X1 U15970 ( .B1(n14639), .B2(n14096), .A(n14095), .ZN(n14130) );
  MUX2_X1 U15971 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14130), .S(n14679), .Z(
        P1_U3546) );
  OAI211_X1 U15972 ( .C1(n14099), .C2(n14655), .A(n14098), .B(n14097), .ZN(
        n14100) );
  AOI21_X1 U15973 ( .B1(n14101), .B2(n14571), .A(n14100), .ZN(n14102) );
  OAI21_X1 U15974 ( .B1(n14639), .B2(n14103), .A(n14102), .ZN(n14131) );
  MUX2_X1 U15975 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14131), .S(n14679), .Z(
        P1_U3545) );
  AOI211_X1 U15976 ( .C1(n14636), .C2(n14106), .A(n14105), .B(n14104), .ZN(
        n14109) );
  NAND2_X1 U15977 ( .A1(n14107), .A2(n14660), .ZN(n14108) );
  OAI211_X1 U15978 ( .C1(n14110), .C2(n14550), .A(n14109), .B(n14108), .ZN(
        n14132) );
  MUX2_X1 U15979 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14132), .S(n14679), .Z(
        P1_U3544) );
  AND2_X1 U15980 ( .A1(n14111), .A2(n14660), .ZN(n14114) );
  OAI21_X1 U15981 ( .B1(n7089), .B2(n14655), .A(n14112), .ZN(n14113) );
  MUX2_X1 U15982 ( .A(n14133), .B(P1_REG1_REG_15__SCAN_IN), .S(n14676), .Z(
        P1_U3543) );
  MUX2_X1 U15983 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14116), .S(n14679), .Z(
        P1_U3528) );
  MUX2_X1 U15984 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14117), .S(n14663), .Z(
        P1_U3527) );
  MUX2_X1 U15985 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14118), .S(n14663), .Z(
        P1_U3526) );
  MUX2_X1 U15986 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14119), .S(n14663), .Z(
        P1_U3525) );
  MUX2_X1 U15987 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14120), .S(n14663), .Z(
        P1_U3524) );
  MUX2_X1 U15988 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14121), .S(n14663), .Z(
        P1_U3523) );
  MUX2_X1 U15989 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14122), .S(n14663), .Z(
        P1_U3522) );
  MUX2_X1 U15990 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14123), .S(n14663), .Z(
        P1_U3521) );
  MUX2_X1 U15991 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14124), .S(n14663), .Z(
        P1_U3520) );
  MUX2_X1 U15992 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14125), .S(n14663), .Z(
        P1_U3519) );
  MUX2_X1 U15993 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14126), .S(n14663), .Z(
        P1_U3518) );
  MUX2_X1 U15994 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14127), .S(n14663), .Z(
        P1_U3517) );
  MUX2_X1 U15995 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14128), .S(n14663), .Z(
        P1_U3516) );
  MUX2_X1 U15996 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14129), .S(n14663), .Z(
        P1_U3515) );
  MUX2_X1 U15997 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14130), .S(n14663), .Z(
        P1_U3513) );
  MUX2_X1 U15998 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14131), .S(n14663), .Z(
        P1_U3510) );
  MUX2_X1 U15999 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14132), .S(n14663), .Z(
        P1_U3507) );
  MUX2_X1 U16000 ( .A(n14133), .B(P1_REG0_REG_15__SCAN_IN), .S(n14661), .Z(
        P1_U3504) );
  NOR4_X1 U16001 ( .A1(n14134), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9479), .A4(
        P1_U3086), .ZN(n14135) );
  AOI21_X1 U16002 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14136), .A(n14135), 
        .ZN(n14137) );
  OAI21_X1 U16003 ( .B1(n14138), .B2(n14148), .A(n14137), .ZN(P1_U3324) );
  OAI222_X1 U16004 ( .A1(n14145), .A2(n14141), .B1(n14148), .B2(n14140), .C1(
        n14139), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16005 ( .A1(n14145), .A2(n14144), .B1(n14148), .B2(n14143), .C1(
        n14142), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U16006 ( .A1(P1_U3086), .A2(n14149), .B1(n14148), .B2(n14147), 
        .C1(n14146), .C2(n14145), .ZN(P1_U3329) );
  MUX2_X1 U16007 ( .A(n6847), .B(n14150), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16008 ( .A(n14152), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16009 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14183) );
  INV_X1 U16010 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15187) );
  NAND2_X1 U16011 ( .A1(n15187), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n14242) );
  INV_X1 U16012 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15261) );
  INV_X1 U16013 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14542) );
  XNOR2_X1 U16014 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14238) );
  INV_X1 U16015 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U16016 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n15115), .ZN(n15216) );
  INV_X1 U16017 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14879) );
  INV_X1 U16018 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14179) );
  XOR2_X1 U16019 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14187) );
  XNOR2_X1 U16020 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14225) );
  XNOR2_X1 U16021 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14172), .ZN(n14190) );
  XNOR2_X1 U16022 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14218) );
  NAND2_X1 U16023 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14154), .ZN(n14155) );
  NAND2_X1 U16024 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14156), .ZN(n14158) );
  NAND2_X1 U16025 ( .A1(n14191), .A2(n6734), .ZN(n14157) );
  NAND2_X1 U16026 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14159), .ZN(n14162) );
  NAND2_X1 U16027 ( .A1(n14205), .A2(n14160), .ZN(n14161) );
  OR2_X1 U16028 ( .A1(n14164), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14163) );
  INV_X1 U16029 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U16030 ( .A1(n14166), .A2(n14165), .ZN(n14168) );
  XNOR2_X1 U16031 ( .A(n14166), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14214) );
  NAND2_X1 U16032 ( .A1(n14214), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U16033 ( .A1(n14168), .A2(n14167), .ZN(n14219) );
  NAND2_X1 U16034 ( .A1(n14218), .A2(n14219), .ZN(n14169) );
  NAND2_X1 U16035 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14173), .ZN(n14175) );
  XOR2_X1 U16036 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14173), .Z(n14223) );
  INV_X1 U16037 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U16038 ( .A1(n14223), .A2(n14224), .ZN(n14174) );
  NAND2_X1 U16039 ( .A1(n14175), .A2(n14174), .ZN(n14226) );
  NAND2_X1 U16040 ( .A1(n14225), .A2(n14226), .ZN(n14176) );
  AND2_X1 U16041 ( .A1(n14879), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14180) );
  INV_X1 U16042 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15172) );
  OAI22_X1 U16043 ( .A1(n15216), .A2(n14236), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n15172), .ZN(n14237) );
  NAND2_X1 U16044 ( .A1(n14238), .A2(n14237), .ZN(n14181) );
  OAI21_X1 U16045 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n14542), .A(n14181), 
        .ZN(n14186) );
  XOR2_X1 U16046 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n14185) );
  OR2_X1 U16047 ( .A1(n14186), .A2(n14185), .ZN(n14182) );
  OAI21_X1 U16048 ( .B1(n15261), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14182), 
        .ZN(n14243) );
  AOI22_X1 U16049 ( .A1(n14183), .A2(P3_ADDR_REG_17__SCAN_IN), .B1(n14242), 
        .B2(n14243), .ZN(n14184) );
  INV_X1 U16050 ( .A(n14184), .ZN(n14298) );
  XOR2_X1 U16051 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14297) );
  XNOR2_X1 U16052 ( .A(n14298), .B(n14297), .ZN(n14301) );
  XOR2_X1 U16053 ( .A(n14186), .B(n14185), .Z(n14240) );
  XOR2_X1 U16054 ( .A(n14188), .B(n14187), .Z(n14500) );
  XOR2_X1 U16055 ( .A(n14190), .B(n14189), .Z(n14259) );
  AND2_X1 U16056 ( .A1(n14203), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14204) );
  XNOR2_X1 U16057 ( .A(n14192), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15301) );
  XOR2_X1 U16058 ( .A(n14194), .B(n14193), .Z(n14251) );
  INV_X1 U16059 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14199) );
  NOR2_X1 U16060 ( .A1(n14198), .A2(n14199), .ZN(n14200) );
  AOI21_X1 U16061 ( .B1(n15116), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14196), .ZN(
        n15295) );
  INV_X1 U16062 ( .A(n15295), .ZN(n14197) );
  NAND2_X1 U16063 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n14197), .ZN(n15305) );
  NOR2_X1 U16064 ( .A1(n15305), .A2(n15304), .ZN(n15303) );
  NOR2_X1 U16065 ( .A1(n14251), .A2(n14250), .ZN(n14201) );
  NAND2_X1 U16066 ( .A1(n14251), .A2(n14250), .ZN(n14249) );
  NAND2_X1 U16067 ( .A1(n15301), .A2(n15300), .ZN(n14202) );
  NOR2_X1 U16068 ( .A1(n15301), .A2(n15300), .ZN(n15299) );
  XNOR2_X1 U16069 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14205), .ZN(n14207) );
  NAND2_X1 U16070 ( .A1(n14206), .A2(n14207), .ZN(n14208) );
  INV_X1 U16071 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15293) );
  INV_X1 U16072 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14209) );
  NOR2_X1 U16073 ( .A1(n14210), .A2(n14209), .ZN(n14213) );
  XOR2_X1 U16074 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n14211) );
  XNOR2_X1 U16075 ( .A(n14212), .B(n14211), .ZN(n14254) );
  INV_X1 U16076 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14216) );
  NOR2_X1 U16077 ( .A1(n14215), .A2(n14216), .ZN(n14217) );
  XNOR2_X1 U16078 ( .A(n14214), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15298) );
  XNOR2_X1 U16079 ( .A(n14219), .B(n14218), .ZN(n14221) );
  NAND2_X1 U16080 ( .A1(n14220), .A2(n14221), .ZN(n14222) );
  INV_X1 U16081 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15241) );
  NAND2_X1 U16082 ( .A1(n14259), .A2(n14260), .ZN(n14258) );
  XNOR2_X1 U16083 ( .A(n14224), .B(n14223), .ZN(n14263) );
  XOR2_X1 U16084 ( .A(n14226), .B(n14225), .Z(n14228) );
  INV_X1 U16085 ( .A(n14494), .ZN(n14495) );
  INV_X1 U16086 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14497) );
  NAND2_X1 U16087 ( .A1(n14228), .A2(n14227), .ZN(n14496) );
  NAND2_X1 U16088 ( .A1(n14500), .A2(n14499), .ZN(n14229) );
  XNOR2_X1 U16089 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14231) );
  XNOR2_X1 U16090 ( .A(n14231), .B(n14230), .ZN(n14233) );
  NAND2_X1 U16091 ( .A1(n14232), .A2(n14233), .ZN(n14234) );
  INV_X1 U16092 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14503) );
  AOI21_X1 U16093 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15115), .A(n15216), 
        .ZN(n14235) );
  XOR2_X1 U16094 ( .A(n14236), .B(n14235), .Z(n14506) );
  NAND2_X1 U16095 ( .A1(n14507), .A2(n14506), .ZN(n14505) );
  XNOR2_X1 U16096 ( .A(n14238), .B(n14237), .ZN(n14510) );
  NOR2_X1 U16097 ( .A1(n14511), .A2(n14510), .ZN(n14239) );
  NAND2_X1 U16098 ( .A1(n14511), .A2(n14510), .ZN(n14509) );
  NAND2_X1 U16099 ( .A1(n14240), .A2(n14241), .ZN(n14515) );
  INV_X1 U16100 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15017) );
  OAI21_X1 U16101 ( .B1(n15187), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14242), 
        .ZN(n14244) );
  XOR2_X1 U16102 ( .A(n14244), .B(n14243), .Z(n14245) );
  INV_X1 U16103 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U16104 ( .A1(n14246), .A2(n14245), .ZN(n14295) );
  NAND2_X1 U16105 ( .A1(n14296), .A2(n14295), .ZN(n14292) );
  AOI21_X1 U16106 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14247) );
  OAI21_X1 U16107 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14247), 
        .ZN(U28) );
  AOI21_X1 U16108 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14248) );
  OAI21_X1 U16109 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14248), 
        .ZN(U29) );
  OAI21_X1 U16110 ( .B1(n14251), .B2(n14250), .A(n14249), .ZN(n14252) );
  XNOR2_X1 U16111 ( .A(n14252), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16112 ( .B1(n14255), .B2(n14254), .A(n14253), .ZN(SUB_1596_U57) );
  OAI21_X1 U16113 ( .B1(n14257), .B2(n15241), .A(n14256), .ZN(SUB_1596_U55) );
  OAI21_X1 U16114 ( .B1(n14260), .B2(n14259), .A(n14258), .ZN(n14261) );
  XNOR2_X1 U16115 ( .A(n14261), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  AOI21_X1 U16116 ( .B1(n14264), .B2(n14263), .A(n14262), .ZN(n14265) );
  XOR2_X1 U16117 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14265), .Z(SUB_1596_U70)
         );
  INV_X1 U16118 ( .A(n14628), .ZN(n14649) );
  XNOR2_X1 U16119 ( .A(n14267), .B(n14266), .ZN(n14288) );
  XNOR2_X1 U16120 ( .A(n14269), .B(n14268), .ZN(n14271) );
  OAI21_X1 U16121 ( .B1(n14271), .B2(n14550), .A(n14270), .ZN(n14272) );
  AOI21_X1 U16122 ( .B1(n14649), .B2(n14288), .A(n14272), .ZN(n14285) );
  AOI222_X1 U16123 ( .A1(n14274), .A2(n14572), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14575), .C1(n14574), .C2(n14273), .ZN(n14282) );
  NOR2_X1 U16124 ( .A1(n14276), .A2(n14275), .ZN(n14582) );
  INV_X1 U16125 ( .A(n14277), .ZN(n14279) );
  OAI211_X1 U16126 ( .C1(n14279), .C2(n14284), .A(n14577), .B(n14278), .ZN(
        n14283) );
  INV_X1 U16127 ( .A(n14283), .ZN(n14280) );
  AOI22_X1 U16128 ( .A1(n14288), .A2(n14582), .B1(n14581), .B2(n14280), .ZN(
        n14281) );
  OAI211_X1 U16129 ( .C1(n14276), .C2(n14285), .A(n14282), .B(n14281), .ZN(
        P1_U3281) );
  INV_X1 U16130 ( .A(n14642), .ZN(n14631) );
  OAI21_X1 U16131 ( .B1(n14284), .B2(n14655), .A(n14283), .ZN(n14287) );
  INV_X1 U16132 ( .A(n14285), .ZN(n14286) );
  AOI211_X1 U16133 ( .C1(n14631), .C2(n14288), .A(n14287), .B(n14286), .ZN(
        n14291) );
  INV_X1 U16134 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U16135 ( .A1(n14663), .A2(n14291), .B1(n14289), .B2(n14661), .ZN(
        P1_U3495) );
  AOI22_X1 U16136 ( .A1(n14679), .A2(n14291), .B1(n14290), .B2(n14676), .ZN(
        P1_U3540) );
  OAI222_X1 U16137 ( .A1(n14296), .A2(n14295), .B1(n14296), .B2(n14294), .C1(
        n14293), .C2(n14292), .ZN(SUB_1596_U63) );
  NOR2_X1 U16138 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  AOI21_X1 U16139 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n12191), .A(n14299), 
        .ZN(n14304) );
  XNOR2_X1 U16140 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14303) );
  AOI21_X1 U16141 ( .B1(n14308), .B2(n14307), .A(n14306), .ZN(n14325) );
  INV_X1 U16142 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U16143 ( .B1(n14310), .B2(P3_REG1_REG_15__SCAN_IN), .A(n14309), 
        .ZN(n14311) );
  INV_X1 U16144 ( .A(n14311), .ZN(n14312) );
  OR2_X1 U16145 ( .A1(n14313), .A2(n14312), .ZN(n14315) );
  OAI211_X1 U16146 ( .C1(n14878), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        n14322) );
  OAI211_X1 U16147 ( .C1(n14319), .C2(n14318), .A(n14317), .B(n14903), .ZN(
        n14320) );
  INV_X1 U16148 ( .A(n14320), .ZN(n14321) );
  AOI211_X1 U16149 ( .C1(n14906), .C2(n14323), .A(n14322), .B(n14321), .ZN(
        n14324) );
  OAI21_X1 U16150 ( .B1(n14325), .B2(n14912), .A(n14324), .ZN(P3_U3197) );
  AOI22_X1 U16151 ( .A1(n14906), .A2(n14326), .B1(n14899), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14343) );
  XNOR2_X1 U16152 ( .A(n14328), .B(n14327), .ZN(n14334) );
  NAND2_X1 U16153 ( .A1(n14330), .A2(n14329), .ZN(n14331) );
  AOI21_X1 U16154 ( .B1(n14332), .B2(n14331), .A(n14882), .ZN(n14333) );
  AOI21_X1 U16155 ( .B1(n14334), .B2(n14895), .A(n14333), .ZN(n14342) );
  INV_X1 U16156 ( .A(n14335), .ZN(n14341) );
  INV_X1 U16157 ( .A(n14336), .ZN(n14339) );
  OAI221_X1 U16158 ( .B1(n14339), .B2(n14338), .C1(n14339), .C2(n14337), .A(
        n14843), .ZN(n14340) );
  NAND4_X1 U16159 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n14340), .ZN(
        P3_U3198) );
  AOI21_X1 U16160 ( .B1(n14346), .B2(n14345), .A(n14344), .ZN(n14362) );
  OAI21_X1 U16161 ( .B1(n14348), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14347), 
        .ZN(n14360) );
  NAND2_X1 U16162 ( .A1(n14350), .A2(n14349), .ZN(n14351) );
  NAND2_X1 U16163 ( .A1(n14351), .A2(n14903), .ZN(n14352) );
  NOR2_X1 U16164 ( .A1(n14353), .A2(n14352), .ZN(n14359) );
  AOI21_X1 U16165 ( .B1(n14899), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n14354), 
        .ZN(n14355) );
  OAI21_X1 U16166 ( .B1(n14357), .B2(n14356), .A(n14355), .ZN(n14358) );
  AOI211_X1 U16167 ( .C1(n14360), .C2(n14895), .A(n14359), .B(n14358), .ZN(
        n14361) );
  OAI21_X1 U16168 ( .B1(n14362), .B2(n14912), .A(n14361), .ZN(P3_U3199) );
  OAI21_X1 U16169 ( .B1(n14364), .B2(n14971), .A(n14363), .ZN(n14373) );
  OAI22_X1 U16170 ( .A1(n14986), .A2(n14373), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n14989), .ZN(n14365) );
  INV_X1 U16171 ( .A(n14365), .ZN(P3_U3489) );
  AOI211_X1 U16172 ( .C1(n14368), .C2(n14963), .A(n14367), .B(n14366), .ZN(
        n14376) );
  AOI22_X1 U16173 ( .A1(n14989), .A2(n14376), .B1(n12193), .B2(n14986), .ZN(
        P3_U3471) );
  AOI211_X1 U16174 ( .C1(n14963), .C2(n14371), .A(n14370), .B(n14369), .ZN(
        n14377) );
  INV_X1 U16175 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U16176 ( .A1(n14989), .A2(n14377), .B1(n14372), .B2(n14986), .ZN(
        P3_U3470) );
  OAI22_X1 U16177 ( .A1(n14977), .A2(n14373), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n14979), .ZN(n14374) );
  INV_X1 U16178 ( .A(n14374), .ZN(P3_U3457) );
  INV_X1 U16179 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U16180 ( .A1(n14979), .A2(n14376), .B1(n14375), .B2(n14977), .ZN(
        P3_U3426) );
  INV_X1 U16181 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U16182 ( .A1(n14979), .A2(n14377), .B1(n15257), .B2(n14977), .ZN(
        P3_U3423) );
  OAI22_X1 U16183 ( .A1(n14380), .A2(n14754), .B1(n14379), .B2(n14378), .ZN(
        n14389) );
  NAND2_X1 U16184 ( .A1(n14382), .A2(n14381), .ZN(n14383) );
  NAND2_X1 U16185 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  AOI222_X1 U16186 ( .A1(n14690), .A2(n14396), .B1(n14389), .B2(n14685), .C1(
        n14385), .C2(n14688), .ZN(n14387) );
  OAI211_X1 U16187 ( .C1(n14694), .C2(n14391), .A(n14387), .B(n14386), .ZN(
        P2_U3187) );
  XNOR2_X1 U16188 ( .A(n14388), .B(n14395), .ZN(n14390) );
  AOI21_X1 U16189 ( .B1(n14390), .B2(n14753), .A(n14389), .ZN(n14405) );
  INV_X1 U16190 ( .A(n14391), .ZN(n14392) );
  AOI222_X1 U16191 ( .A1(n14396), .A2(n14393), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14736), .C1(n14734), .C2(n14392), .ZN(n14402) );
  XOR2_X1 U16192 ( .A(n14394), .B(n14395), .Z(n14408) );
  INV_X1 U16193 ( .A(n14396), .ZN(n14404) );
  INV_X1 U16194 ( .A(n14397), .ZN(n14399) );
  OAI211_X1 U16195 ( .C1(n14404), .C2(n14399), .A(n10011), .B(n14398), .ZN(
        n14403) );
  INV_X1 U16196 ( .A(n14403), .ZN(n14400) );
  AOI22_X1 U16197 ( .A1(n14408), .A2(n10037), .B1(n14731), .B2(n14400), .ZN(
        n14401) );
  OAI211_X1 U16198 ( .C1(n14736), .C2(n14405), .A(n14402), .B(n14401), .ZN(
        P2_U3251) );
  OAI21_X1 U16199 ( .B1(n14404), .B2(n14819), .A(n14403), .ZN(n14407) );
  INV_X1 U16200 ( .A(n14405), .ZN(n14406) );
  AOI211_X1 U16201 ( .C1(n7116), .C2(n14408), .A(n14407), .B(n14406), .ZN(
        n14424) );
  AOI22_X1 U16202 ( .A1(n14833), .A2(n14424), .B1(n7910), .B2(n14834), .ZN(
        P2_U3513) );
  AOI21_X1 U16203 ( .B1(n14410), .B2(n14795), .A(n14409), .ZN(n14412) );
  OAI211_X1 U16204 ( .C1(n14413), .C2(n14799), .A(n14412), .B(n14411), .ZN(
        n14414) );
  AOI21_X1 U16205 ( .B1(n14415), .B2(n14753), .A(n14414), .ZN(n14425) );
  AOI22_X1 U16206 ( .A1(n14833), .A2(n14425), .B1(n10987), .B2(n14834), .ZN(
        P2_U3512) );
  NOR2_X1 U16207 ( .A1(n14416), .A2(n6774), .ZN(n14421) );
  INV_X1 U16208 ( .A(n14689), .ZN(n14419) );
  OAI211_X1 U16209 ( .C1(n14419), .C2(n14819), .A(n14418), .B(n14417), .ZN(
        n14420) );
  AOI211_X1 U16210 ( .C1(n8861), .C2(n14422), .A(n14421), .B(n14420), .ZN(
        n14426) );
  AOI22_X1 U16211 ( .A1(n14833), .A2(n14426), .B1(n9891), .B2(n14834), .ZN(
        P2_U3511) );
  INV_X1 U16212 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U16213 ( .A1(n14814), .A2(n14424), .B1(n14423), .B2(n14824), .ZN(
        P2_U3472) );
  INV_X1 U16214 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U16215 ( .A1(n14814), .A2(n14425), .B1(n15243), .B2(n14824), .ZN(
        P2_U3469) );
  INV_X1 U16216 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15250) );
  AOI22_X1 U16217 ( .A1(n14814), .A2(n14426), .B1(n15250), .B2(n14824), .ZN(
        P2_U3466) );
  NAND2_X1 U16218 ( .A1(n14428), .A2(n14427), .ZN(n14429) );
  NAND2_X1 U16219 ( .A1(n14430), .A2(n14429), .ZN(n14432) );
  AOI222_X1 U16220 ( .A1(n14434), .A2(n14433), .B1(n14432), .B2(n14440), .C1(
        n14431), .C2(n14447), .ZN(n14436) );
  OAI211_X1 U16221 ( .C1(n14463), .C2(n14437), .A(n14436), .B(n14435), .ZN(
        P1_U3215) );
  OAI21_X1 U16222 ( .B1(n14456), .B2(n14439), .A(n14438), .ZN(n14446) );
  OAI211_X1 U16223 ( .C1(n14443), .C2(n14442), .A(n14441), .B(n14440), .ZN(
        n14444) );
  INV_X1 U16224 ( .A(n14444), .ZN(n14445) );
  AOI211_X1 U16225 ( .C1(n14447), .C2(n14653), .A(n14446), .B(n14445), .ZN(
        n14448) );
  OAI21_X1 U16226 ( .B1(n14449), .B2(n14463), .A(n14448), .ZN(P1_U3217) );
  NAND2_X1 U16227 ( .A1(n14450), .A2(n14636), .ZN(n14483) );
  INV_X1 U16228 ( .A(n14483), .ZN(n14452) );
  AOI22_X1 U16229 ( .A1(n14452), .A2(n14451), .B1(P1_REG3_REG_11__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14462) );
  AOI21_X1 U16230 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14459) );
  OAI22_X1 U16231 ( .A1(n14459), .A2(n14458), .B1(n14457), .B2(n14456), .ZN(
        n14460) );
  INV_X1 U16232 ( .A(n14460), .ZN(n14461) );
  OAI211_X1 U16233 ( .C1(n14464), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        P1_U3236) );
  OAI211_X1 U16234 ( .C1(n14467), .C2(n14655), .A(n14466), .B(n14465), .ZN(
        n14470) );
  AND3_X1 U16235 ( .A1(n11256), .A2(n14468), .A3(n14660), .ZN(n14469) );
  AOI211_X1 U16236 ( .C1(n14471), .C2(n14571), .A(n14470), .B(n14469), .ZN(
        n14488) );
  AOI22_X1 U16237 ( .A1(n14679), .A2(n14488), .B1(n14472), .B2(n14676), .ZN(
        P1_U3542) );
  NAND2_X1 U16238 ( .A1(n14473), .A2(n14571), .ZN(n14478) );
  INV_X1 U16239 ( .A(n14474), .ZN(n14475) );
  AOI21_X1 U16240 ( .B1(n14476), .B2(n14636), .A(n14475), .ZN(n14477) );
  OAI211_X1 U16241 ( .C1(n6570), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14480) );
  AOI21_X1 U16242 ( .B1(n14481), .B2(n14660), .A(n14480), .ZN(n14490) );
  AOI22_X1 U16243 ( .A1(n14679), .A2(n14490), .B1(n10153), .B2(n14676), .ZN(
        P1_U3541) );
  OAI211_X1 U16244 ( .C1(n14484), .C2(n14639), .A(n14483), .B(n14482), .ZN(
        n14485) );
  NOR2_X1 U16245 ( .A1(n14486), .A2(n14485), .ZN(n14492) );
  AOI22_X1 U16246 ( .A1(n14679), .A2(n14492), .B1(n9485), .B2(n14676), .ZN(
        P1_U3539) );
  INV_X1 U16247 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16248 ( .A1(n14663), .A2(n14488), .B1(n14487), .B2(n14661), .ZN(
        P1_U3501) );
  INV_X1 U16249 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U16250 ( .A1(n14663), .A2(n14490), .B1(n14489), .B2(n14661), .ZN(
        P1_U3498) );
  INV_X1 U16251 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U16252 ( .A1(n14663), .A2(n14492), .B1(n14491), .B2(n14661), .ZN(
        P1_U3492) );
  OAI222_X1 U16253 ( .A1(n14497), .A2(n14496), .B1(n14497), .B2(n14495), .C1(
        n14494), .C2(n14493), .ZN(SUB_1596_U69) );
  AOI21_X1 U16254 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n14501) );
  XOR2_X1 U16255 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14501), .Z(SUB_1596_U68)
         );
  OAI21_X1 U16256 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(SUB_1596_U67) );
  OAI21_X1 U16257 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n14508) );
  XNOR2_X1 U16258 ( .A(n14508), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI21_X1 U16259 ( .B1(n14511), .B2(n14510), .A(n14509), .ZN(n14512) );
  XNOR2_X1 U16260 ( .A(n14512), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U16261 ( .A(n14515), .ZN(n14514) );
  OAI222_X1 U16262 ( .A1(n15017), .A2(n14516), .B1(n15017), .B2(n14515), .C1(
        n14514), .C2(n14513), .ZN(SUB_1596_U64) );
  NOR2_X1 U16263 ( .A1(n14517), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n14519) );
  OR2_X1 U16264 ( .A1(n14518), .A2(n14519), .ZN(n14522) );
  INV_X1 U16265 ( .A(n14519), .ZN(n14521) );
  MUX2_X1 U16266 ( .A(n14522), .B(n14521), .S(n14520), .Z(n14524) );
  NAND2_X1 U16267 ( .A1(n14524), .A2(n14523), .ZN(n14527) );
  AOI22_X1 U16268 ( .A1(n14525), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14526) );
  OAI21_X1 U16269 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(P1_U3243) );
  AOI21_X1 U16270 ( .B1(n14530), .B2(P1_REG1_REG_15__SCAN_IN), .A(n14529), 
        .ZN(n14535) );
  AOI21_X1 U16271 ( .B1(n14532), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14531), 
        .ZN(n14533) );
  OAI222_X1 U16272 ( .A1(n6779), .A2(n14537), .B1(n14536), .B2(n14535), .C1(
        n14534), .C2(n14533), .ZN(n14538) );
  INV_X1 U16273 ( .A(n14538), .ZN(n14540) );
  OAI211_X1 U16274 ( .C1(n14542), .C2(n14541), .A(n14540), .B(n14539), .ZN(
        P1_U3258) );
  XOR2_X1 U16275 ( .A(n14547), .B(n14543), .Z(n14618) );
  INV_X1 U16276 ( .A(n14618), .ZN(n14560) );
  INV_X1 U16277 ( .A(n14544), .ZN(n14545) );
  AOI21_X1 U16278 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14551) );
  INV_X1 U16279 ( .A(n14548), .ZN(n14549) );
  OAI21_X1 U16280 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(n14622) );
  AOI21_X1 U16281 ( .B1(n14649), .B2(n14560), .A(n14622), .ZN(n14563) );
  INV_X1 U16282 ( .A(n14552), .ZN(n14553) );
  AOI222_X1 U16283 ( .A1(n14559), .A2(n14572), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14575), .C1(n14574), .C2(n14553), .ZN(n14562) );
  INV_X1 U16284 ( .A(n14554), .ZN(n14558) );
  INV_X1 U16285 ( .A(n14555), .ZN(n14556) );
  AOI211_X1 U16286 ( .C1(n14559), .C2(n14558), .A(n6570), .B(n14556), .ZN(
        n14619) );
  AOI22_X1 U16287 ( .A1(n14560), .A2(n14582), .B1(n14581), .B2(n14619), .ZN(
        n14561) );
  OAI211_X1 U16288 ( .C1(n14276), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        P1_U3287) );
  OAI21_X1 U16289 ( .B1(n14566), .B2(n14565), .A(n14564), .ZN(n14570) );
  XNOR2_X1 U16290 ( .A(n14567), .B(n14566), .ZN(n14576) );
  NOR2_X1 U16291 ( .A1(n14576), .A2(n14628), .ZN(n14568) );
  AOI211_X1 U16292 ( .C1(n14571), .C2(n14570), .A(n14569), .B(n14568), .ZN(
        n14591) );
  AOI222_X1 U16293 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n14575), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14574), .C1(n14573), .C2(n14572), .ZN(
        n14584) );
  INV_X1 U16294 ( .A(n14576), .ZN(n14594) );
  OAI211_X1 U16295 ( .C1(n14579), .C2(n14590), .A(n14578), .B(n14577), .ZN(
        n14589) );
  INV_X1 U16296 ( .A(n14589), .ZN(n14580) );
  AOI22_X1 U16297 ( .A1(n14582), .A2(n14594), .B1(n14581), .B2(n14580), .ZN(
        n14583) );
  OAI211_X1 U16298 ( .C1(n14276), .C2(n14591), .A(n14584), .B(n14583), .ZN(
        P1_U3291) );
  AND2_X1 U16299 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14586), .ZN(P1_U3294) );
  INV_X1 U16300 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15185) );
  NOR2_X1 U16301 ( .A1(n14585), .A2(n15185), .ZN(P1_U3295) );
  INV_X1 U16302 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15042) );
  NOR2_X1 U16303 ( .A1(n14585), .A2(n15042), .ZN(P1_U3296) );
  INV_X1 U16304 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15095) );
  NOR2_X1 U16305 ( .A1(n14585), .A2(n15095), .ZN(P1_U3297) );
  AND2_X1 U16306 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14586), .ZN(P1_U3298) );
  AND2_X1 U16307 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14586), .ZN(P1_U3299) );
  AND2_X1 U16308 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14586), .ZN(P1_U3300) );
  AND2_X1 U16309 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14586), .ZN(P1_U3301) );
  AND2_X1 U16310 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14586), .ZN(P1_U3302) );
  AND2_X1 U16311 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14586), .ZN(P1_U3303) );
  AND2_X1 U16312 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14586), .ZN(P1_U3304) );
  AND2_X1 U16313 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14586), .ZN(P1_U3305) );
  AND2_X1 U16314 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14586), .ZN(P1_U3306) );
  AND2_X1 U16315 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14586), .ZN(P1_U3307) );
  AND2_X1 U16316 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14586), .ZN(P1_U3308) );
  AND2_X1 U16317 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14586), .ZN(P1_U3309) );
  AND2_X1 U16318 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14586), .ZN(P1_U3310) );
  AND2_X1 U16319 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14586), .ZN(P1_U3311) );
  INV_X1 U16320 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15104) );
  NOR2_X1 U16321 ( .A1(n14585), .A2(n15104), .ZN(P1_U3312) );
  AND2_X1 U16322 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14586), .ZN(P1_U3313) );
  AND2_X1 U16323 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14586), .ZN(P1_U3314) );
  INV_X1 U16324 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15189) );
  NOR2_X1 U16325 ( .A1(n14585), .A2(n15189), .ZN(P1_U3315) );
  AND2_X1 U16326 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14586), .ZN(P1_U3316) );
  AND2_X1 U16327 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14586), .ZN(P1_U3317) );
  AND2_X1 U16328 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14586), .ZN(P1_U3318) );
  AND2_X1 U16329 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14586), .ZN(P1_U3319) );
  AND2_X1 U16330 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14586), .ZN(P1_U3320) );
  AND2_X1 U16331 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14586), .ZN(P1_U3321) );
  AND2_X1 U16332 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14586), .ZN(P1_U3322) );
  AND2_X1 U16333 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14586), .ZN(P1_U3323) );
  INV_X1 U16334 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U16335 ( .A1(n14663), .A2(n14588), .B1(n14587), .B2(n14661), .ZN(
        P1_U3462) );
  OAI21_X1 U16336 ( .B1(n14590), .B2(n14655), .A(n14589), .ZN(n14593) );
  INV_X1 U16337 ( .A(n14591), .ZN(n14592) );
  AOI211_X1 U16338 ( .C1(n14631), .C2(n14594), .A(n14593), .B(n14592), .ZN(
        n14664) );
  INV_X1 U16339 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15267) );
  AOI22_X1 U16340 ( .A1(n14663), .A2(n14664), .B1(n15267), .B2(n14661), .ZN(
        P1_U3465) );
  INV_X1 U16341 ( .A(n14599), .ZN(n14601) );
  AOI21_X1 U16342 ( .B1(n14636), .B2(n14596), .A(n14595), .ZN(n14598) );
  OAI211_X1 U16343 ( .C1(n14599), .C2(n14642), .A(n14598), .B(n14597), .ZN(
        n14600) );
  AOI21_X1 U16344 ( .B1(n14649), .B2(n14601), .A(n14600), .ZN(n14665) );
  INV_X1 U16345 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U16346 ( .A1(n14663), .A2(n14665), .B1(n14602), .B2(n14661), .ZN(
        P1_U3468) );
  NOR2_X1 U16347 ( .A1(n14603), .A2(n14655), .ZN(n14604) );
  NOR2_X1 U16348 ( .A1(n14605), .A2(n14604), .ZN(n14608) );
  OR2_X1 U16349 ( .A1(n14606), .A2(n14639), .ZN(n14607) );
  AND3_X1 U16350 ( .A1(n14609), .A2(n14608), .A3(n14607), .ZN(n14666) );
  AOI22_X1 U16351 ( .A1(n14663), .A2(n14666), .B1(n10246), .B2(n14661), .ZN(
        P1_U3471) );
  INV_X1 U16352 ( .A(n14610), .ZN(n14616) );
  OR4_X1 U16353 ( .A1(n14614), .A2(n14613), .A3(n14612), .A4(n14611), .ZN(
        n14615) );
  AOI21_X1 U16354 ( .B1(n14616), .B2(n14660), .A(n14615), .ZN(n14668) );
  INV_X1 U16355 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14617) );
  AOI22_X1 U16356 ( .A1(n14663), .A2(n14668), .B1(n14617), .B2(n14661), .ZN(
        P1_U3474) );
  NOR2_X1 U16357 ( .A1(n14618), .A2(n14639), .ZN(n14621) );
  NOR4_X1 U16358 ( .A1(n14622), .A2(n14621), .A3(n14620), .A4(n14619), .ZN(
        n14670) );
  INV_X1 U16359 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15206) );
  AOI22_X1 U16360 ( .A1(n14663), .A2(n14670), .B1(n15206), .B2(n14661), .ZN(
        P1_U3477) );
  INV_X1 U16361 ( .A(n14627), .ZN(n14630) );
  NOR2_X1 U16362 ( .A1(n14624), .A2(n14623), .ZN(n14625) );
  OAI211_X1 U16363 ( .C1(n14628), .C2(n14627), .A(n14626), .B(n14625), .ZN(
        n14629) );
  AOI21_X1 U16364 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14672) );
  INV_X1 U16365 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U16366 ( .A1(n14663), .A2(n14672), .B1(n14632), .B2(n14661), .ZN(
        P1_U3480) );
  AOI211_X1 U16367 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14637) );
  OAI21_X1 U16368 ( .B1(n14639), .B2(n14638), .A(n14637), .ZN(n14640) );
  INV_X1 U16369 ( .A(n14640), .ZN(n14673) );
  INV_X1 U16370 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14641) );
  AOI22_X1 U16371 ( .A1(n14663), .A2(n14673), .B1(n14641), .B2(n14661), .ZN(
        P1_U3483) );
  INV_X1 U16372 ( .A(n14643), .ZN(n14650) );
  NOR2_X1 U16373 ( .A1(n14643), .A2(n14642), .ZN(n14648) );
  OAI211_X1 U16374 ( .C1(n14646), .C2(n14655), .A(n14645), .B(n14644), .ZN(
        n14647) );
  AOI211_X1 U16375 ( .C1(n14650), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14675) );
  INV_X1 U16376 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14651) );
  AOI22_X1 U16377 ( .A1(n14663), .A2(n14675), .B1(n14651), .B2(n14661), .ZN(
        P1_U3486) );
  INV_X1 U16378 ( .A(n14652), .ZN(n14659) );
  INV_X1 U16379 ( .A(n14653), .ZN(n14656) );
  OAI21_X1 U16380 ( .B1(n14656), .B2(n14655), .A(n14654), .ZN(n14658) );
  AOI211_X1 U16381 ( .C1(n14660), .C2(n14659), .A(n14658), .B(n14657), .ZN(
        n14678) );
  INV_X1 U16382 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14662) );
  AOI22_X1 U16383 ( .A1(n14663), .A2(n14678), .B1(n14662), .B2(n14661), .ZN(
        P1_U3489) );
  AOI22_X1 U16384 ( .A1(n14679), .A2(n14664), .B1(n9205), .B2(n14676), .ZN(
        P1_U3530) );
  AOI22_X1 U16385 ( .A1(n14679), .A2(n14665), .B1(n9212), .B2(n14676), .ZN(
        P1_U3531) );
  AOI22_X1 U16386 ( .A1(n14679), .A2(n14666), .B1(n15086), .B2(n14676), .ZN(
        P1_U3532) );
  AOI22_X1 U16387 ( .A1(n14679), .A2(n14668), .B1(n14667), .B2(n14676), .ZN(
        P1_U3533) );
  AOI22_X1 U16388 ( .A1(n14679), .A2(n14670), .B1(n14669), .B2(n14676), .ZN(
        P1_U3534) );
  AOI22_X1 U16389 ( .A1(n14679), .A2(n14672), .B1(n14671), .B2(n14676), .ZN(
        P1_U3535) );
  AOI22_X1 U16390 ( .A1(n14679), .A2(n14673), .B1(n9488), .B2(n14676), .ZN(
        P1_U3536) );
  AOI22_X1 U16391 ( .A1(n14679), .A2(n14675), .B1(n14674), .B2(n14676), .ZN(
        P1_U3537) );
  AOI22_X1 U16392 ( .A1(n14679), .A2(n14678), .B1(n14677), .B2(n14676), .ZN(
        P1_U3538) );
  NOR2_X1 U16393 ( .A1(n14718), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16394 ( .A(n14680), .ZN(n14682) );
  NOR2_X1 U16395 ( .A1(n14682), .A2(n14681), .ZN(n14683) );
  XNOR2_X1 U16396 ( .A(n14684), .B(n14683), .ZN(n14687) );
  AOI222_X1 U16397 ( .A1(n14690), .A2(n14689), .B1(n14688), .B2(n14687), .C1(
        n14686), .C2(n14685), .ZN(n14692) );
  OAI211_X1 U16398 ( .C1(n14694), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        P2_U3196) );
  OAI21_X1 U16399 ( .B1(n14697), .B2(n14696), .A(n14695), .ZN(n14703) );
  OAI21_X1 U16400 ( .B1(n14700), .B2(n14699), .A(n14698), .ZN(n14701) );
  AOI222_X1 U16401 ( .A1(n14703), .A2(n14725), .B1(n14702), .B2(n14720), .C1(
        n14701), .C2(n6547), .ZN(n14705) );
  OAI211_X1 U16402 ( .C1(n6827), .C2(n14706), .A(n14705), .B(n14704), .ZN(
        P2_U3223) );
  AOI22_X1 U16403 ( .A1(n14718), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14717) );
  OAI211_X1 U16404 ( .C1(n14709), .C2(n14708), .A(n14707), .B(n6547), .ZN(
        n14716) );
  NAND2_X1 U16405 ( .A1(n14720), .A2(n14710), .ZN(n14715) );
  OAI211_X1 U16406 ( .C1(n14713), .C2(n14712), .A(n14711), .B(n14725), .ZN(
        n14714) );
  NAND4_X1 U16407 ( .A1(n14717), .A2(n14716), .A3(n14715), .A4(n14714), .ZN(
        P2_U3227) );
  AOI22_X1 U16408 ( .A1(n14718), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14730) );
  NAND2_X1 U16409 ( .A1(n14720), .A2(n14719), .ZN(n14729) );
  XNOR2_X1 U16410 ( .A(n14721), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U16411 ( .A1(n14723), .A2(n6547), .ZN(n14728) );
  XNOR2_X1 U16412 ( .A(n14724), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U16413 ( .A1(n14726), .A2(n14725), .ZN(n14727) );
  NAND4_X1 U16414 ( .A1(n14730), .A2(n14729), .A3(n14728), .A4(n14727), .ZN(
        P2_U3229) );
  NAND2_X1 U16415 ( .A1(n14732), .A2(n14731), .ZN(n14738) );
  INV_X1 U16416 ( .A(n14733), .ZN(n14735) );
  AOI22_X1 U16417 ( .A1(n14736), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14735), 
        .B2(n14734), .ZN(n14737) );
  OAI211_X1 U16418 ( .C1(n14740), .C2(n14739), .A(n14738), .B(n14737), .ZN(
        n14741) );
  AOI21_X1 U16419 ( .B1(n10037), .B2(n14742), .A(n14741), .ZN(n14743) );
  OAI21_X1 U16420 ( .B1(n14736), .B2(n14744), .A(n14743), .ZN(P2_U3258) );
  INV_X1 U16421 ( .A(n14756), .ZN(n14770) );
  INV_X1 U16422 ( .A(n14745), .ZN(n14746) );
  NOR2_X1 U16423 ( .A1(n14747), .A2(n14746), .ZN(n14769) );
  OAI21_X1 U16424 ( .B1(n14749), .B2(n14748), .A(n14769), .ZN(n14750) );
  OAI21_X1 U16425 ( .B1(n14752), .B2(n14751), .A(n14750), .ZN(n14757) );
  NOR2_X1 U16426 ( .A1(n14816), .A2(n14753), .ZN(n14755) );
  OAI22_X1 U16427 ( .A1(n14756), .A2(n14755), .B1(n7686), .B2(n14754), .ZN(
        n14768) );
  AOI211_X1 U16428 ( .C1(n6720), .C2(n14770), .A(n14757), .B(n14768), .ZN(
        n14758) );
  AOI22_X1 U16429 ( .A1(n14736), .A2(n9360), .B1(n14758), .B2(n6558), .ZN(
        P2_U3265) );
  NAND2_X1 U16430 ( .A1(n14767), .A2(n14759), .ZN(n14760) );
  AND2_X1 U16431 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14760), .ZN(P2_U3266) );
  INV_X1 U16432 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15077) );
  NOR2_X1 U16433 ( .A1(n14761), .A2(n15077), .ZN(P2_U3267) );
  AND2_X1 U16434 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14760), .ZN(P2_U3268) );
  INV_X1 U16435 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15079) );
  NOR2_X1 U16436 ( .A1(n14761), .A2(n15079), .ZN(P2_U3269) );
  AND2_X1 U16437 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14760), .ZN(P2_U3270) );
  AND2_X1 U16438 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14760), .ZN(P2_U3271) );
  AND2_X1 U16439 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14760), .ZN(P2_U3272) );
  NOR2_X1 U16440 ( .A1(n14761), .A2(n15109), .ZN(P2_U3273) );
  AND2_X1 U16441 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14760), .ZN(P2_U3274) );
  AND2_X1 U16442 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14760), .ZN(P2_U3275) );
  NOR2_X1 U16443 ( .A1(n14761), .A2(n15048), .ZN(P2_U3276) );
  NOR2_X1 U16444 ( .A1(n14761), .A2(n15065), .ZN(P2_U3277) );
  AND2_X1 U16445 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14760), .ZN(P2_U3278) );
  AND2_X1 U16446 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14760), .ZN(P2_U3279) );
  AND2_X1 U16447 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14760), .ZN(P2_U3280) );
  AND2_X1 U16448 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14760), .ZN(P2_U3281) );
  AND2_X1 U16449 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14760), .ZN(P2_U3282) );
  NOR2_X1 U16450 ( .A1(n14761), .A2(n15045), .ZN(P2_U3283) );
  AND2_X1 U16451 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14760), .ZN(P2_U3284) );
  NOR2_X1 U16452 ( .A1(n14761), .A2(n14992), .ZN(P2_U3285) );
  AND2_X1 U16453 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14760), .ZN(P2_U3286) );
  AND2_X1 U16454 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14760), .ZN(P2_U3287) );
  AND2_X1 U16455 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14760), .ZN(P2_U3288) );
  INV_X1 U16456 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U16457 ( .A1(n14761), .A2(n15124), .ZN(P2_U3289) );
  AND2_X1 U16458 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14760), .ZN(P2_U3290) );
  AND2_X1 U16459 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14760), .ZN(P2_U3291) );
  AND2_X1 U16460 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14760), .ZN(P2_U3292) );
  AND2_X1 U16461 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14760), .ZN(P2_U3293) );
  NOR2_X1 U16462 ( .A1(n14761), .A2(n15084), .ZN(P2_U3294) );
  AND2_X1 U16463 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14760), .ZN(P2_U3295) );
  OAI22_X1 U16464 ( .A1(n14764), .A2(n14762), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n14761), .ZN(n14763) );
  INV_X1 U16465 ( .A(n14763), .ZN(P2_U3416) );
  INV_X1 U16466 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U16467 ( .A1(n14767), .A2(n14766), .B1(n14765), .B2(n14764), .ZN(
        P2_U3417) );
  AOI211_X1 U16468 ( .C1(n14770), .C2(n8861), .A(n14769), .B(n14768), .ZN(
        n14825) );
  AOI22_X1 U16469 ( .A1(n14814), .A2(n14825), .B1(n7688), .B2(n14824), .ZN(
        P2_U3430) );
  OAI21_X1 U16470 ( .B1(n14772), .B2(n14819), .A(n14771), .ZN(n14774) );
  AOI211_X1 U16471 ( .C1(n8861), .C2(n14775), .A(n14774), .B(n14773), .ZN(
        n14826) );
  INV_X1 U16472 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14776) );
  AOI22_X1 U16473 ( .A1(n14814), .A2(n14826), .B1(n14776), .B2(n14824), .ZN(
        P2_U3433) );
  INV_X1 U16474 ( .A(n14777), .ZN(n14783) );
  NOR2_X1 U16475 ( .A1(n14777), .A2(n6774), .ZN(n14782) );
  OAI211_X1 U16476 ( .C1(n14780), .C2(n14819), .A(n14779), .B(n14778), .ZN(
        n14781) );
  AOI211_X1 U16477 ( .C1(n8861), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14827) );
  INV_X1 U16478 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U16479 ( .A1(n14814), .A2(n14827), .B1(n14784), .B2(n14824), .ZN(
        P2_U3436) );
  INV_X1 U16480 ( .A(n14785), .ZN(n14791) );
  INV_X1 U16481 ( .A(n14786), .ZN(n14787) );
  OAI211_X1 U16482 ( .C1(n14789), .C2(n14819), .A(n14788), .B(n14787), .ZN(
        n14790) );
  AOI21_X1 U16483 ( .B1(n7116), .B2(n14791), .A(n14790), .ZN(n14828) );
  INV_X1 U16484 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14792) );
  AOI22_X1 U16485 ( .A1(n14814), .A2(n14828), .B1(n14792), .B2(n14824), .ZN(
        P2_U3439) );
  AOI21_X1 U16486 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14797) );
  OAI211_X1 U16487 ( .C1(n14799), .C2(n14798), .A(n14797), .B(n14796), .ZN(
        n14800) );
  INV_X1 U16488 ( .A(n14800), .ZN(n14829) );
  INV_X1 U16489 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16490 ( .A1(n14814), .A2(n14829), .B1(n14801), .B2(n14824), .ZN(
        P2_U3442) );
  OAI21_X1 U16491 ( .B1(n14803), .B2(n14819), .A(n14802), .ZN(n14805) );
  AOI211_X1 U16492 ( .C1(n14806), .C2(n7116), .A(n14805), .B(n14804), .ZN(
        n14830) );
  INV_X1 U16493 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U16494 ( .A1(n14814), .A2(n14830), .B1(n15230), .B2(n14824), .ZN(
        P2_U3454) );
  AOI21_X1 U16495 ( .B1(n14809), .B2(n6774), .A(n14807), .ZN(n14812) );
  NOR2_X1 U16496 ( .A1(n7148), .A2(n14819), .ZN(n14810) );
  NOR4_X1 U16497 ( .A1(n14813), .A2(n14812), .A3(n14811), .A4(n14810), .ZN(
        n14832) );
  AOI22_X1 U16498 ( .A1(n14814), .A2(n14832), .B1(n7853), .B2(n14824), .ZN(
        P2_U3460) );
  OAI21_X1 U16499 ( .B1(n8861), .B2(n14816), .A(n14815), .ZN(n14817) );
  INV_X1 U16500 ( .A(n14817), .ZN(n14822) );
  OAI21_X1 U16501 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14821) );
  NOR3_X1 U16502 ( .A1(n14823), .A2(n14822), .A3(n14821), .ZN(n14835) );
  AOI22_X1 U16503 ( .A1(n14814), .A2(n14835), .B1(n7865), .B2(n14824), .ZN(
        P2_U3463) );
  AOI22_X1 U16504 ( .A1(n14833), .A2(n14825), .B1(n9181), .B2(n14834), .ZN(
        P2_U3499) );
  AOI22_X1 U16505 ( .A1(n14833), .A2(n14826), .B1(n7680), .B2(n14834), .ZN(
        P2_U3500) );
  AOI22_X1 U16506 ( .A1(n14833), .A2(n14827), .B1(n7699), .B2(n14834), .ZN(
        P2_U3501) );
  AOI22_X1 U16507 ( .A1(n14833), .A2(n14828), .B1(n7716), .B2(n14834), .ZN(
        P2_U3502) );
  AOI22_X1 U16508 ( .A1(n14833), .A2(n14829), .B1(n9335), .B2(n14834), .ZN(
        P2_U3503) );
  AOI22_X1 U16509 ( .A1(n14833), .A2(n14830), .B1(n7815), .B2(n14834), .ZN(
        P2_U3507) );
  AOI22_X1 U16510 ( .A1(n14833), .A2(n14832), .B1(n14831), .B2(n14834), .ZN(
        P2_U3509) );
  AOI22_X1 U16511 ( .A1(n14833), .A2(n14835), .B1(n15047), .B2(n14834), .ZN(
        P2_U3510) );
  NOR2_X1 U16512 ( .A1(P3_U3897), .A2(n14899), .ZN(P3_U3150) );
  AOI22_X1 U16513 ( .A1(n14906), .A2(n14836), .B1(n14899), .B2(
        P3_ADDR_REG_11__SCAN_IN), .ZN(n14849) );
  XNOR2_X1 U16514 ( .A(n14838), .B(n14837), .ZN(n14842) );
  OAI21_X1 U16515 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n14840), .A(n14839), 
        .ZN(n14841) );
  AOI22_X1 U16516 ( .A1(n14842), .A2(n14903), .B1(n14841), .B2(n14895), .ZN(
        n14848) );
  OAI221_X1 U16517 ( .B1(n14845), .B2(n11322), .C1(n14845), .C2(n14844), .A(
        n14843), .ZN(n14846) );
  NAND4_X1 U16518 ( .A1(n14849), .A2(n14848), .A3(n14847), .A4(n14846), .ZN(
        P3_U3193) );
  AOI21_X1 U16519 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14869) );
  OAI21_X1 U16520 ( .B1(n14855), .B2(n14854), .A(n14853), .ZN(n14867) );
  INV_X1 U16521 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14861) );
  INV_X1 U16522 ( .A(n14856), .ZN(n14857) );
  NAND2_X1 U16523 ( .A1(n14906), .A2(n14857), .ZN(n14860) );
  INV_X1 U16524 ( .A(n14858), .ZN(n14859) );
  OAI211_X1 U16525 ( .C1(n14861), .C2(n14878), .A(n14860), .B(n14859), .ZN(
        n14866) );
  XNOR2_X1 U16526 ( .A(n14863), .B(n14862), .ZN(n14864) );
  NOR2_X1 U16527 ( .A1(n14864), .A2(n14882), .ZN(n14865) );
  AOI211_X1 U16528 ( .C1(n14895), .C2(n14867), .A(n14866), .B(n14865), .ZN(
        n14868) );
  OAI21_X1 U16529 ( .B1(n14869), .B2(n14912), .A(n14868), .ZN(P3_U3194) );
  AOI21_X1 U16530 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n14889) );
  OAI21_X1 U16531 ( .B1(n14874), .B2(P3_REG1_REG_13__SCAN_IN), .A(n14873), 
        .ZN(n14887) );
  NAND2_X1 U16532 ( .A1(n14906), .A2(n14875), .ZN(n14877) );
  OAI211_X1 U16533 ( .C1(n14879), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        n14886) );
  NAND2_X1 U16534 ( .A1(n14881), .A2(n14880), .ZN(n14883) );
  AOI21_X1 U16535 ( .B1(n14884), .B2(n14883), .A(n14882), .ZN(n14885) );
  AOI211_X1 U16536 ( .C1(n14887), .C2(n14895), .A(n14886), .B(n14885), .ZN(
        n14888) );
  OAI21_X1 U16537 ( .B1(n14889), .B2(n14912), .A(n14888), .ZN(P3_U3195) );
  AOI21_X1 U16538 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n14913) );
  XNOR2_X1 U16539 ( .A(n14894), .B(n14893), .ZN(n14896) );
  NAND2_X1 U16540 ( .A1(n14896), .A2(n14895), .ZN(n14910) );
  INV_X1 U16541 ( .A(n14897), .ZN(n14898) );
  AOI21_X1 U16542 ( .B1(n14899), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n14898), 
        .ZN(n14909) );
  NAND2_X1 U16543 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  NAND3_X1 U16544 ( .A1(n14904), .A2(n14903), .A3(n14902), .ZN(n14908) );
  NAND2_X1 U16545 ( .A1(n14906), .A2(n14905), .ZN(n14907) );
  AND4_X1 U16546 ( .A1(n14910), .A2(n14909), .A3(n14908), .A4(n14907), .ZN(
        n14911) );
  OAI21_X1 U16547 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(P3_U3196) );
  OAI21_X1 U16548 ( .B1(n14915), .B2(n14919), .A(n14914), .ZN(n14957) );
  NAND2_X1 U16549 ( .A1(n14916), .A2(n14966), .ZN(n14954) );
  OAI22_X1 U16550 ( .A1(n14954), .A2(n14935), .B1(n14934), .B2(n14917), .ZN(
        n14927) );
  XNOR2_X1 U16551 ( .A(n14919), .B(n14918), .ZN(n14926) );
  INV_X1 U16552 ( .A(n14920), .ZN(n14924) );
  OAI22_X1 U16553 ( .A1(n14922), .A2(n14941), .B1(n14921), .B2(n14943), .ZN(
        n14923) );
  AOI21_X1 U16554 ( .B1(n14957), .B2(n14924), .A(n14923), .ZN(n14925) );
  OAI21_X1 U16555 ( .B1(n14939), .B2(n14926), .A(n14925), .ZN(n14955) );
  AOI211_X1 U16556 ( .C1(n14928), .C2(n14957), .A(n14927), .B(n14955), .ZN(
        n14929) );
  AOI22_X1 U16557 ( .A1(n14949), .A2(n15262), .B1(n14929), .B2(n14946), .ZN(
        P3_U3231) );
  XOR2_X1 U16558 ( .A(n14930), .B(n14937), .Z(n14953) );
  NAND2_X1 U16559 ( .A1(n14932), .A2(n14966), .ZN(n14950) );
  OAI22_X1 U16560 ( .A1(n14950), .A2(n14935), .B1(n14934), .B2(n14933), .ZN(
        n14944) );
  XNOR2_X1 U16561 ( .A(n14937), .B(n14936), .ZN(n14938) );
  OAI222_X1 U16562 ( .A1(n14943), .A2(n14942), .B1(n14941), .B2(n14940), .C1(
        n14939), .C2(n14938), .ZN(n14951) );
  AOI211_X1 U16563 ( .C1(n14945), .C2(n14953), .A(n14944), .B(n14951), .ZN(
        n14947) );
  AOI22_X1 U16564 ( .A1(n14949), .A2(n14948), .B1(n14947), .B2(n14946), .ZN(
        P3_U3232) );
  INV_X1 U16565 ( .A(n14950), .ZN(n14952) );
  AOI211_X1 U16566 ( .C1(n14963), .C2(n14953), .A(n14952), .B(n14951), .ZN(
        n14980) );
  AOI22_X1 U16567 ( .A1(n14979), .A2(n14980), .B1(n8258), .B2(n14977), .ZN(
        P3_U3393) );
  INV_X1 U16568 ( .A(n14954), .ZN(n14956) );
  AOI211_X1 U16569 ( .C1(n14958), .C2(n14957), .A(n14956), .B(n14955), .ZN(
        n14981) );
  INV_X1 U16570 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15231) );
  AOI22_X1 U16571 ( .A1(n14979), .A2(n14981), .B1(n15231), .B2(n14977), .ZN(
        P3_U3396) );
  NOR2_X1 U16572 ( .A1(n14959), .A2(n14971), .ZN(n14961) );
  AOI211_X1 U16573 ( .C1(n14963), .C2(n14962), .A(n14961), .B(n14960), .ZN(
        n14983) );
  INV_X1 U16574 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U16575 ( .A1(n14979), .A2(n14983), .B1(n14964), .B2(n14977), .ZN(
        P3_U3414) );
  AOI21_X1 U16576 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(n14968) );
  OAI21_X1 U16577 ( .B1(n14973), .B2(n14969), .A(n14968), .ZN(n14984) );
  OAI22_X1 U16578 ( .A1(n14977), .A2(n14984), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n14979), .ZN(n14970) );
  INV_X1 U16579 ( .A(n14970), .ZN(P3_U3417) );
  OAI22_X1 U16580 ( .A1(n14974), .A2(n14973), .B1(n14972), .B2(n14971), .ZN(
        n14976) );
  NOR2_X1 U16581 ( .A1(n14976), .A2(n14975), .ZN(n14988) );
  INV_X1 U16582 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16583 ( .A1(n14979), .A2(n14988), .B1(n14978), .B2(n14977), .ZN(
        P3_U3420) );
  AOI22_X1 U16584 ( .A1(n14989), .A2(n14980), .B1(n8259), .B2(n14986), .ZN(
        P3_U3460) );
  AOI22_X1 U16585 ( .A1(n14989), .A2(n14981), .B1(n9581), .B2(n14986), .ZN(
        P3_U3461) );
  AOI22_X1 U16586 ( .A1(n14989), .A2(n14983), .B1(n14982), .B2(n14986), .ZN(
        P3_U3467) );
  OAI22_X1 U16587 ( .A1(n14986), .A2(n14984), .B1(P3_REG1_REG_9__SCAN_IN), 
        .B2(n14989), .ZN(n14985) );
  INV_X1 U16588 ( .A(n14985), .ZN(P3_U3468) );
  AOI22_X1 U16589 ( .A1(n14989), .A2(n14988), .B1(n14987), .B2(n14986), .ZN(
        P3_U3469) );
  AOI22_X1 U16590 ( .A1(n15207), .A2(keyinput43), .B1(keyinput111), .B2(n15206), .ZN(n14990) );
  OAI221_X1 U16591 ( .B1(n15207), .B2(keyinput43), .C1(n15206), .C2(
        keyinput111), .A(n14990), .ZN(n14999) );
  AOI22_X1 U16592 ( .A1(n14992), .A2(keyinput50), .B1(n15208), .B2(keyinput89), 
        .ZN(n14991) );
  OAI221_X1 U16593 ( .B1(n14992), .B2(keyinput50), .C1(n15208), .C2(keyinput89), .A(n14991), .ZN(n14998) );
  XNOR2_X1 U16594 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput39), .ZN(n14996)
         );
  XNOR2_X1 U16595 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput74), .ZN(n14995) );
  XNOR2_X1 U16596 ( .A(P3_REG0_REG_28__SCAN_IN), .B(keyinput6), .ZN(n14994) );
  XNOR2_X1 U16597 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput13), .ZN(n14993) );
  NAND4_X1 U16598 ( .A1(n14996), .A2(n14995), .A3(n14994), .A4(n14993), .ZN(
        n14997) );
  NOR3_X1 U16599 ( .A1(n14999), .A2(n14998), .A3(n14997), .ZN(n15040) );
  INV_X1 U16600 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n15210) );
  AOI22_X1 U16601 ( .A1(n15210), .A2(keyinput27), .B1(keyinput0), .B2(n15209), 
        .ZN(n15000) );
  OAI221_X1 U16602 ( .B1(n15210), .B2(keyinput27), .C1(n15209), .C2(keyinput0), 
        .A(n15000), .ZN(n15007) );
  INV_X1 U16603 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15003) );
  AOI22_X1 U16604 ( .A1(n15003), .A2(keyinput84), .B1(n15002), .B2(keyinput116), .ZN(n15001) );
  OAI221_X1 U16605 ( .B1(n15003), .B2(keyinput84), .C1(n15002), .C2(
        keyinput116), .A(n15001), .ZN(n15006) );
  XNOR2_X1 U16606 ( .A(n15004), .B(keyinput54), .ZN(n15005) );
  OR3_X1 U16607 ( .A1(n15007), .A2(n15006), .A3(n15005), .ZN(n15013) );
  AOI22_X1 U16608 ( .A1(n15009), .A2(keyinput105), .B1(keyinput7), .B2(n7896), 
        .ZN(n15008) );
  OAI221_X1 U16609 ( .B1(n15009), .B2(keyinput105), .C1(n7896), .C2(keyinput7), 
        .A(n15008), .ZN(n15012) );
  XNOR2_X1 U16610 ( .A(n15010), .B(keyinput21), .ZN(n15011) );
  NOR3_X1 U16611 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(n15039) );
  AOI22_X1 U16612 ( .A1(n15015), .A2(keyinput87), .B1(keyinput40), .B2(n9181), 
        .ZN(n15014) );
  OAI221_X1 U16613 ( .B1(n15015), .B2(keyinput87), .C1(n9181), .C2(keyinput40), 
        .A(n15014), .ZN(n15024) );
  AOI22_X1 U16614 ( .A1(n15250), .A2(keyinput82), .B1(keyinput67), .B2(n15017), 
        .ZN(n15016) );
  OAI221_X1 U16615 ( .B1(n15250), .B2(keyinput82), .C1(n15017), .C2(keyinput67), .A(n15016), .ZN(n15023) );
  AOI22_X1 U16616 ( .A1(n6729), .A2(keyinput5), .B1(keyinput76), .B2(n15019), 
        .ZN(n15018) );
  OAI221_X1 U16617 ( .B1(n6729), .B2(keyinput5), .C1(n15019), .C2(keyinput76), 
        .A(n15018), .ZN(n15022) );
  AOI22_X1 U16618 ( .A1(n15249), .A2(keyinput65), .B1(n7865), .B2(keyinput88), 
        .ZN(n15020) );
  OAI221_X1 U16619 ( .B1(n15249), .B2(keyinput65), .C1(n7865), .C2(keyinput88), 
        .A(n15020), .ZN(n15021) );
  NOR4_X1 U16620 ( .A1(n15024), .A2(n15023), .A3(n15022), .A4(n15021), .ZN(
        n15038) );
  AOI22_X1 U16621 ( .A1(n15026), .A2(keyinput37), .B1(n15251), .B2(keyinput102), .ZN(n15025) );
  OAI221_X1 U16622 ( .B1(n15026), .B2(keyinput37), .C1(n15251), .C2(
        keyinput102), .A(n15025), .ZN(n15036) );
  INV_X1 U16623 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n15029) );
  INV_X1 U16624 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15028) );
  AOI22_X1 U16625 ( .A1(n15029), .A2(keyinput19), .B1(n15028), .B2(keyinput10), 
        .ZN(n15027) );
  OAI221_X1 U16626 ( .B1(n15029), .B2(keyinput19), .C1(n15028), .C2(keyinput10), .A(n15027), .ZN(n15035) );
  XOR2_X1 U16627 ( .A(n8053), .B(keyinput123), .Z(n15033) );
  XNOR2_X1 U16628 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput110), .ZN(n15032)
         );
  XNOR2_X1 U16629 ( .A(P2_REG0_REG_17__SCAN_IN), .B(keyinput122), .ZN(n15031)
         );
  XNOR2_X1 U16630 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput97), .ZN(n15030) );
  NAND4_X1 U16631 ( .A1(n15033), .A2(n15032), .A3(n15031), .A4(n15030), .ZN(
        n15034) );
  NOR3_X1 U16632 ( .A1(n15036), .A2(n15035), .A3(n15034), .ZN(n15037) );
  NAND4_X1 U16633 ( .A1(n15040), .A2(n15039), .A3(n15038), .A4(n15037), .ZN(
        n15201) );
  AOI22_X1 U16634 ( .A1(n15241), .A2(keyinput56), .B1(n15042), .B2(keyinput23), 
        .ZN(n15041) );
  OAI221_X1 U16635 ( .B1(n15241), .B2(keyinput56), .C1(n15042), .C2(keyinput23), .A(n15041), .ZN(n15052) );
  AOI22_X1 U16636 ( .A1(n12599), .A2(keyinput4), .B1(n15242), .B2(keyinput28), 
        .ZN(n15043) );
  OAI221_X1 U16637 ( .B1(n12599), .B2(keyinput4), .C1(n15242), .C2(keyinput28), 
        .A(n15043), .ZN(n15051) );
  AOI22_X1 U16638 ( .A1(n7832), .A2(keyinput51), .B1(n15045), .B2(keyinput2), 
        .ZN(n15044) );
  OAI221_X1 U16639 ( .B1(n7832), .B2(keyinput51), .C1(n15045), .C2(keyinput2), 
        .A(n15044), .ZN(n15050) );
  AOI22_X1 U16640 ( .A1(n15048), .A2(keyinput41), .B1(keyinput3), .B2(n15047), 
        .ZN(n15046) );
  OAI221_X1 U16641 ( .B1(n15048), .B2(keyinput41), .C1(n15047), .C2(keyinput3), 
        .A(n15046), .ZN(n15049) );
  NOR4_X1 U16642 ( .A1(n15052), .A2(n15051), .A3(n15050), .A4(n15049), .ZN(
        n15093) );
  AOI22_X1 U16643 ( .A1(n15054), .A2(keyinput103), .B1(n9336), .B2(keyinput62), 
        .ZN(n15053) );
  OAI221_X1 U16644 ( .B1(n15054), .B2(keyinput103), .C1(n9336), .C2(keyinput62), .A(n15053), .ZN(n15063) );
  AOI22_X1 U16645 ( .A1(n15243), .A2(keyinput78), .B1(keyinput73), .B2(n9310), 
        .ZN(n15055) );
  OAI221_X1 U16646 ( .B1(n15243), .B2(keyinput78), .C1(n9310), .C2(keyinput73), 
        .A(n15055), .ZN(n15062) );
  AOI22_X1 U16647 ( .A1(n15244), .A2(keyinput8), .B1(keyinput99), .B2(n9756), 
        .ZN(n15056) );
  OAI221_X1 U16648 ( .B1(n15244), .B2(keyinput8), .C1(n9756), .C2(keyinput99), 
        .A(n15056), .ZN(n15061) );
  INV_X1 U16649 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16650 ( .A1(n15059), .A2(keyinput114), .B1(keyinput22), .B2(n15058), .ZN(n15057) );
  OAI221_X1 U16651 ( .B1(n15059), .B2(keyinput114), .C1(n15058), .C2(
        keyinput22), .A(n15057), .ZN(n15060) );
  NOR4_X1 U16652 ( .A1(n15063), .A2(n15062), .A3(n15061), .A4(n15060), .ZN(
        n15092) );
  AOI22_X1 U16653 ( .A1(n15066), .A2(keyinput69), .B1(keyinput72), .B2(n15065), 
        .ZN(n15064) );
  OAI221_X1 U16654 ( .B1(n15066), .B2(keyinput69), .C1(n15065), .C2(keyinput72), .A(n15064), .ZN(n15074) );
  XOR2_X1 U16655 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput119), .Z(n15073) );
  XNOR2_X1 U16656 ( .A(keyinput94), .B(n9493), .ZN(n15072) );
  XNOR2_X1 U16657 ( .A(P2_B_REG_SCAN_IN), .B(keyinput71), .ZN(n15070) );
  XNOR2_X1 U16658 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput29), .ZN(n15069)
         );
  XNOR2_X1 U16659 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput81), .ZN(n15068) );
  XNOR2_X1 U16660 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput100), .ZN(n15067) );
  NAND4_X1 U16661 ( .A1(n15070), .A2(n15069), .A3(n15068), .A4(n15067), .ZN(
        n15071) );
  NOR4_X1 U16662 ( .A1(n15074), .A2(n15073), .A3(n15072), .A4(n15071), .ZN(
        n15091) );
  AOI22_X1 U16663 ( .A1(n15077), .A2(keyinput18), .B1(keyinput46), .B2(n15076), 
        .ZN(n15075) );
  OAI221_X1 U16664 ( .B1(n15077), .B2(keyinput18), .C1(n15076), .C2(keyinput46), .A(n15075), .ZN(n15082) );
  XNOR2_X1 U16665 ( .A(n15078), .B(keyinput109), .ZN(n15081) );
  XNOR2_X1 U16666 ( .A(n15079), .B(keyinput1), .ZN(n15080) );
  OR3_X1 U16667 ( .A1(n15082), .A2(n15081), .A3(n15080), .ZN(n15089) );
  AOI22_X1 U16668 ( .A1(n15084), .A2(keyinput127), .B1(keyinput59), .B2(n7716), 
        .ZN(n15083) );
  OAI221_X1 U16669 ( .B1(n15084), .B2(keyinput127), .C1(n7716), .C2(keyinput59), .A(n15083), .ZN(n15088) );
  AOI22_X1 U16670 ( .A1(n8000), .A2(keyinput112), .B1(keyinput49), .B2(n15086), 
        .ZN(n15085) );
  OAI221_X1 U16671 ( .B1(n8000), .B2(keyinput112), .C1(n15086), .C2(keyinput49), .A(n15085), .ZN(n15087) );
  NOR3_X1 U16672 ( .A1(n15089), .A2(n15088), .A3(n15087), .ZN(n15090) );
  NAND4_X1 U16673 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15200) );
  AOI22_X1 U16674 ( .A1(n15095), .A2(keyinput95), .B1(n15223), .B2(keyinput55), 
        .ZN(n15094) );
  OAI221_X1 U16675 ( .B1(n15095), .B2(keyinput95), .C1(n15223), .C2(keyinput55), .A(n15094), .ZN(n15101) );
  AOI22_X1 U16676 ( .A1(n15097), .A2(keyinput70), .B1(n15224), .B2(keyinput126), .ZN(n15096) );
  OAI221_X1 U16677 ( .B1(n15097), .B2(keyinput70), .C1(n15224), .C2(
        keyinput126), .A(n15096), .ZN(n15100) );
  XNOR2_X1 U16678 ( .A(n15098), .B(keyinput11), .ZN(n15099) );
  OR3_X1 U16679 ( .A1(n15101), .A2(n15100), .A3(n15099), .ZN(n15107) );
  AOI22_X1 U16680 ( .A1(n15103), .A2(keyinput33), .B1(keyinput124), .B2(n7853), 
        .ZN(n15102) );
  OAI221_X1 U16681 ( .B1(n15103), .B2(keyinput33), .C1(n7853), .C2(keyinput124), .A(n15102), .ZN(n15106) );
  XNOR2_X1 U16682 ( .A(n15104), .B(keyinput92), .ZN(n15105) );
  NOR3_X1 U16683 ( .A1(n15107), .A2(n15106), .A3(n15105), .ZN(n15148) );
  AOI22_X1 U16684 ( .A1(n15110), .A2(keyinput53), .B1(keyinput31), .B2(n15109), 
        .ZN(n15108) );
  OAI221_X1 U16685 ( .B1(n15110), .B2(keyinput53), .C1(n15109), .C2(keyinput31), .A(n15108), .ZN(n15122) );
  AOI22_X1 U16686 ( .A1(n15113), .A2(keyinput68), .B1(keyinput24), .B2(n15112), 
        .ZN(n15111) );
  OAI221_X1 U16687 ( .B1(n15113), .B2(keyinput68), .C1(n15112), .C2(keyinput24), .A(n15111), .ZN(n15121) );
  AOI22_X1 U16688 ( .A1(n15116), .A2(keyinput121), .B1(n15115), .B2(keyinput32), .ZN(n15114) );
  OAI221_X1 U16689 ( .B1(n15116), .B2(keyinput121), .C1(n15115), .C2(
        keyinput32), .A(n15114), .ZN(n15120) );
  AOI22_X1 U16690 ( .A1(n15118), .A2(keyinput75), .B1(n15228), .B2(keyinput125), .ZN(n15117) );
  OAI221_X1 U16691 ( .B1(n15118), .B2(keyinput75), .C1(n15228), .C2(
        keyinput125), .A(n15117), .ZN(n15119) );
  NOR4_X1 U16692 ( .A1(n15122), .A2(n15121), .A3(n15120), .A4(n15119), .ZN(
        n15147) );
  INV_X1 U16693 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15229) );
  AOI22_X1 U16694 ( .A1(n15229), .A2(keyinput106), .B1(keyinput30), .B2(n15124), .ZN(n15123) );
  OAI221_X1 U16695 ( .B1(n15229), .B2(keyinput106), .C1(n15124), .C2(
        keyinput30), .A(n15123), .ZN(n15133) );
  AOI22_X1 U16696 ( .A1(n12191), .A2(keyinput107), .B1(n7562), .B2(keyinput64), 
        .ZN(n15125) );
  OAI221_X1 U16697 ( .B1(n12191), .B2(keyinput107), .C1(n7562), .C2(keyinput64), .A(n15125), .ZN(n15132) );
  INV_X1 U16698 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n15232) );
  INV_X1 U16699 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n15127) );
  AOI22_X1 U16700 ( .A1(n15232), .A2(keyinput86), .B1(keyinput93), .B2(n15127), 
        .ZN(n15126) );
  OAI221_X1 U16701 ( .B1(n15232), .B2(keyinput86), .C1(n15127), .C2(keyinput93), .A(n15126), .ZN(n15131) );
  AOI22_X1 U16702 ( .A1(n15129), .A2(keyinput20), .B1(n9951), .B2(keyinput108), 
        .ZN(n15128) );
  OAI221_X1 U16703 ( .B1(n15129), .B2(keyinput20), .C1(n9951), .C2(keyinput108), .A(n15128), .ZN(n15130) );
  NOR4_X1 U16704 ( .A1(n15133), .A2(n15132), .A3(n15131), .A4(n15130), .ZN(
        n15146) );
  AOI22_X1 U16705 ( .A1(n15135), .A2(keyinput26), .B1(keyinput79), .B2(n15231), 
        .ZN(n15134) );
  OAI221_X1 U16706 ( .B1(n15135), .B2(keyinput26), .C1(n15231), .C2(keyinput79), .A(n15134), .ZN(n15144) );
  AOI22_X1 U16707 ( .A1(n15270), .A2(keyinput42), .B1(keyinput12), .B2(n15137), 
        .ZN(n15136) );
  OAI221_X1 U16708 ( .B1(n15270), .B2(keyinput42), .C1(n15137), .C2(keyinput12), .A(n15136), .ZN(n15143) );
  INV_X1 U16709 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U16710 ( .A1(n15268), .A2(keyinput44), .B1(n15269), .B2(keyinput66), 
        .ZN(n15138) );
  OAI221_X1 U16711 ( .B1(n15268), .B2(keyinput44), .C1(n15269), .C2(keyinput66), .A(n15138), .ZN(n15142) );
  XOR2_X1 U16712 ( .A(n15230), .B(keyinput57), .Z(n15140) );
  XNOR2_X1 U16713 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput115), .ZN(n15139) );
  NAND2_X1 U16714 ( .A1(n15140), .A2(n15139), .ZN(n15141) );
  NOR4_X1 U16715 ( .A1(n15144), .A2(n15143), .A3(n15142), .A4(n15141), .ZN(
        n15145) );
  NAND4_X1 U16716 ( .A1(n15148), .A2(n15147), .A3(n15146), .A4(n15145), .ZN(
        n15199) );
  AOI22_X1 U16717 ( .A1(n15267), .A2(keyinput117), .B1(n15150), .B2(keyinput58), .ZN(n15149) );
  OAI221_X1 U16718 ( .B1(n15267), .B2(keyinput117), .C1(n15150), .C2(
        keyinput58), .A(n15149), .ZN(n15159) );
  INV_X1 U16719 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U16720 ( .A1(n15271), .A2(keyinput45), .B1(n14917), .B2(keyinput96), 
        .ZN(n15151) );
  OAI221_X1 U16721 ( .B1(n15271), .B2(keyinput45), .C1(n14917), .C2(keyinput96), .A(n15151), .ZN(n15158) );
  AOI22_X1 U16722 ( .A1(n15154), .A2(keyinput63), .B1(n15153), .B2(keyinput48), 
        .ZN(n15152) );
  OAI221_X1 U16723 ( .B1(n15154), .B2(keyinput63), .C1(n15153), .C2(keyinput48), .A(n15152), .ZN(n15157) );
  AOI22_X1 U16724 ( .A1(n15293), .A2(keyinput77), .B1(n8032), .B2(keyinput9), 
        .ZN(n15155) );
  OAI221_X1 U16725 ( .B1(n15293), .B2(keyinput77), .C1(n8032), .C2(keyinput9), 
        .A(n15155), .ZN(n15156) );
  NOR4_X1 U16726 ( .A1(n15159), .A2(n15158), .A3(n15157), .A4(n15156), .ZN(
        n15197) );
  AOI22_X1 U16727 ( .A1(n7815), .A2(keyinput16), .B1(n15161), .B2(keyinput52), 
        .ZN(n15160) );
  OAI221_X1 U16728 ( .B1(n7815), .B2(keyinput16), .C1(n15161), .C2(keyinput52), 
        .A(n15160), .ZN(n15170) );
  XNOR2_X1 U16729 ( .A(n15273), .B(keyinput120), .ZN(n15169) );
  XNOR2_X1 U16730 ( .A(n15162), .B(keyinput15), .ZN(n15168) );
  XNOR2_X1 U16731 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput98), .ZN(n15166) );
  XNOR2_X1 U16732 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput85), .ZN(n15165) );
  XNOR2_X1 U16733 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput101), .ZN(n15164) );
  XNOR2_X1 U16734 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput91), .ZN(n15163)
         );
  NAND4_X1 U16735 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        n15167) );
  NOR4_X1 U16736 ( .A1(n15170), .A2(n15169), .A3(n15168), .A4(n15167), .ZN(
        n15196) );
  AOI22_X1 U16737 ( .A1(n15172), .A2(keyinput90), .B1(n8011), .B2(keyinput113), 
        .ZN(n15171) );
  OAI221_X1 U16738 ( .B1(n15172), .B2(keyinput90), .C1(n8011), .C2(keyinput113), .A(n15171), .ZN(n15181) );
  AOI22_X1 U16739 ( .A1(n13251), .A2(keyinput80), .B1(keyinput83), .B2(n15174), 
        .ZN(n15173) );
  OAI221_X1 U16740 ( .B1(n13251), .B2(keyinput80), .C1(n15174), .C2(keyinput83), .A(n15173), .ZN(n15180) );
  AOI22_X1 U16741 ( .A1(n15176), .A2(keyinput118), .B1(n15256), .B2(keyinput61), .ZN(n15175) );
  OAI221_X1 U16742 ( .B1(n15176), .B2(keyinput118), .C1(n15256), .C2(
        keyinput61), .A(n15175), .ZN(n15179) );
  AOI22_X1 U16743 ( .A1(n15257), .A2(keyinput60), .B1(keyinput17), .B2(n15258), 
        .ZN(n15177) );
  OAI221_X1 U16744 ( .B1(n15257), .B2(keyinput60), .C1(n15258), .C2(keyinput17), .A(n15177), .ZN(n15178) );
  NOR4_X1 U16745 ( .A1(n15181), .A2(n15180), .A3(n15179), .A4(n15178), .ZN(
        n15195) );
  AOI22_X1 U16746 ( .A1(n15183), .A2(keyinput35), .B1(n15262), .B2(keyinput25), 
        .ZN(n15182) );
  OAI221_X1 U16747 ( .B1(n15183), .B2(keyinput35), .C1(n15262), .C2(keyinput25), .A(n15182), .ZN(n15193) );
  AOI22_X1 U16748 ( .A1(n15185), .A2(keyinput36), .B1(keyinput38), .B2(n15261), 
        .ZN(n15184) );
  OAI221_X1 U16749 ( .B1(n15185), .B2(keyinput36), .C1(n15261), .C2(keyinput38), .A(n15184), .ZN(n15192) );
  AOI22_X1 U16750 ( .A1(n15187), .A2(keyinput14), .B1(n15259), .B2(keyinput47), 
        .ZN(n15186) );
  OAI221_X1 U16751 ( .B1(n15187), .B2(keyinput14), .C1(n15259), .C2(keyinput47), .A(n15186), .ZN(n15191) );
  AOI22_X1 U16752 ( .A1(n15260), .A2(keyinput34), .B1(n15189), .B2(keyinput104), .ZN(n15188) );
  OAI221_X1 U16753 ( .B1(n15260), .B2(keyinput34), .C1(n15189), .C2(
        keyinput104), .A(n15188), .ZN(n15190) );
  NOR4_X1 U16754 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15194) );
  NAND4_X1 U16755 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15198) );
  NOR4_X1 U16756 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15205) );
  MUX2_X1 U16757 ( .A(n15203), .B(n15202), .S(n13695), .Z(n15204) );
  XNOR2_X1 U16758 ( .A(n15205), .B(n15204), .ZN(n15288) );
  NAND4_X1 U16759 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n15208), .A3(n15207), 
        .A4(n15206), .ZN(n15215) );
  NAND4_X1 U16760 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG3_REG_12__SCAN_IN), .A4(P1_REG3_REG_16__SCAN_IN), .ZN(n15214) );
  NAND4_X1 U16761 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(P1_REG0_REG_30__SCAN_IN), .A3(n15210), .A4(n15209), .ZN(n15213) );
  NAND4_X1 U16762 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), 
        .A3(P1_ADDR_REG_10__SCAN_IN), .A4(n15211), .ZN(n15212) );
  NOR4_X1 U16763 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15286) );
  INV_X1 U16764 ( .A(n15216), .ZN(n15220) );
  NOR4_X1 U16765 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .A3(P3_ADDR_REG_0__SCAN_IN), .A4(P2_ADDR_REG_2__SCAN_IN), .ZN(n15217)
         );
  NAND4_X1 U16766 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n15218), .A3(n15217), 
        .A4(n15293), .ZN(n15219) );
  NOR4_X1 U16767 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15285) );
  NOR4_X1 U16768 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), 
        .A3(n15223), .A4(n7716), .ZN(n15225) );
  NAND3_X1 U16769 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15225), .A3(n15224), .ZN(
        n15240) );
  NAND4_X1 U16770 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P1_REG2_REG_8__SCAN_IN), .A4(n15226), .ZN(n15227) );
  NOR3_X1 U16771 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(P1_REG1_REG_4__SCAN_IN), 
        .A3(n15227), .ZN(n15238) );
  NAND4_X1 U16772 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P3_ADDR_REG_18__SCAN_IN), 
        .A3(n15229), .A4(n15228), .ZN(n15236) );
  NAND4_X1 U16773 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(P2_REG0_REG_10__SCAN_IN), 
        .A3(P1_REG2_REG_6__SCAN_IN), .A4(P3_DATAO_REG_18__SCAN_IN), .ZN(n15235) );
  NAND4_X1 U16774 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_REG2_REG_4__SCAN_IN), 
        .A3(n15231), .A4(n15230), .ZN(n15234) );
  NAND4_X1 U16775 ( .A1(P3_REG2_REG_19__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .A3(P1_REG0_REG_27__SCAN_IN), .A4(n15232), .ZN(n15233) );
  NOR4_X1 U16776 ( .A1(n15236), .A2(n15235), .A3(n15234), .A4(n15233), .ZN(
        n15237) );
  NAND4_X1 U16777 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(n15238), .A3(n15237), .A4(
        n9493), .ZN(n15239) );
  NOR4_X1 U16778 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), 
        .A3(n15240), .A4(n15239), .ZN(n15284) );
  NOR4_X1 U16779 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(P2_REG1_REG_5__SCAN_IN), 
        .A3(P1_REG2_REG_3__SCAN_IN), .A4(n7832), .ZN(n15248) );
  NOR4_X1 U16780 ( .A1(P1_D_REG_29__SCAN_IN), .A2(SI_31_), .A3(n15242), .A4(
        n15241), .ZN(n15247) );
  NOR4_X1 U16781 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(P3_REG2_REG_3__SCAN_IN), 
        .A3(P3_REG1_REG_20__SCAN_IN), .A4(P2_B_REG_SCAN_IN), .ZN(n15246) );
  NOR4_X1 U16782 ( .A1(SI_27_), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n15244), .A4(
        n15243), .ZN(n15245) );
  NAND4_X1 U16783 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        n15282) );
  NOR4_X1 U16784 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .A3(n6729), .A4(n15249), .ZN(n15255) );
  NOR4_X1 U16785 ( .A1(P3_REG1_REG_19__SCAN_IN), .A2(n7896), .A3(n15250), .A4(
        n9181), .ZN(n15254) );
  NOR4_X1 U16786 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .A3(
        P2_REG0_REG_17__SCAN_IN), .A4(n15251), .ZN(n15253) );
  NOR4_X1 U16787 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_11__SCAN_IN), .A4(n8053), .ZN(n15252) );
  NAND4_X1 U16788 ( .A1(n15255), .A2(n15254), .A3(n15253), .A4(n15252), .ZN(
        n15281) );
  NOR4_X1 U16789 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(n15258), .A3(n15257), 
        .A4(n15256), .ZN(n15266) );
  NOR4_X1 U16790 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P2_REG2_REG_23__SCAN_IN), .A4(P3_DATAO_REG_5__SCAN_IN), .ZN(n15265) );
  NOR4_X1 U16791 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P3_ADDR_REG_17__SCAN_IN), 
        .A3(n15260), .A4(n15259), .ZN(n15264) );
  NOR4_X1 U16792 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P3_REG1_REG_31__SCAN_IN), 
        .A3(n15262), .A4(n15261), .ZN(n15263) );
  NAND4_X1 U16793 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15280) );
  NOR4_X1 U16794 ( .A1(n15270), .A2(n15269), .A3(n15268), .A4(n15267), .ZN(
        n15278) );
  NOR4_X1 U16795 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .A3(P1_REG2_REG_12__SCAN_IN), .A4(n15271), .ZN(n15277) );
  NOR4_X1 U16796 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(n15273), .A3(n15272), .A4(
        n7815), .ZN(n15274) );
  AND4_X1 U16797 ( .A1(n15275), .A2(P3_IR_REG_14__SCAN_IN), .A3(n15274), .A4(
        P2_REG2_REG_24__SCAN_IN), .ZN(n15276) );
  NAND4_X1 U16798 ( .A1(n15278), .A2(n15277), .A3(n15276), .A4(
        P3_D_REG_15__SCAN_IN), .ZN(n15279) );
  NOR4_X1 U16799 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        n15283) );
  NAND4_X1 U16800 ( .A1(n15286), .A2(n15285), .A3(n15284), .A4(n15283), .ZN(
        n15287) );
  XNOR2_X1 U16801 ( .A(n15288), .B(n15287), .ZN(P1_U3582) );
  AOI21_X1 U16802 ( .B1(n15291), .B2(n15290), .A(n15289), .ZN(SUB_1596_U59) );
  OAI21_X1 U16803 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(SUB_1596_U58) );
  XNOR2_X1 U16804 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15295), .ZN(SUB_1596_U53)
         );
  AOI21_X1 U16805 ( .B1(n15298), .B2(n15297), .A(n15296), .ZN(SUB_1596_U56) );
  AOI21_X1 U16806 ( .B1(n15301), .B2(n15300), .A(n15299), .ZN(n15302) );
  XOR2_X1 U16807 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15302), .Z(SUB_1596_U60) );
  AOI21_X1 U16808 ( .B1(n15305), .B2(n15304), .A(n15303), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7567 ( .A(n8213), .Z(n11044) );
  INV_X1 U7300 ( .A(n6825), .ZN(n13617) );
  BUF_X2 U7301 ( .A(n8135), .Z(n8101) );
  OR2_X1 U7306 ( .A1(n8281), .A2(n10050), .ZN(n11438) );
  CLKBUF_X1 U7320 ( .A(n8311), .Z(n11401) );
  INV_X1 U7336 ( .A(n10011), .ZN(n13104) );
  INV_X2 U7346 ( .A(n10011), .ZN(n12664) );
  NAND2_X2 U7357 ( .A1(n9233), .A2(n14142), .ZN(n11671) );
  CLKBUF_X1 U7364 ( .A(n9926), .Z(n6555) );
  NAND2_X1 U7371 ( .A1(n12716), .A2(n12715), .ZN(n12714) );
  OR2_X1 U7402 ( .A1(n9179), .A2(n8140), .ZN(n15310) );
endmodule

