

module b21_C_gen_AntiSAT_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086;

  OR2_X1 U4815 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  INV_X2 U4816 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR2_X1 U4817 ( .A1(n5515), .A2(n8500), .ZN(n6059) );
  CLKBUF_X2 U4818 ( .A(n4960), .Z(n5328) );
  CLKBUF_X2 U4819 ( .A(n4333), .Z(n5330) );
  XNOR2_X1 U4820 ( .A(n5019), .B(n5018), .ZN(n6080) );
  INV_X1 U4821 ( .A(n5346), .ZN(n5377) );
  CLKBUF_X2 U4822 ( .A(n5481), .Z(n8888) );
  INV_X1 U4823 ( .A(n5967), .ZN(n8388) );
  INV_X1 U4824 ( .A(n5481), .ZN(n8623) );
  INV_X1 U4825 ( .A(n5523), .ZN(n8204) );
  INV_X1 U4826 ( .A(n8509), .ZN(n6762) );
  CLKBUF_X2 U4827 ( .A(n8409), .Z(n4311) );
  AND2_X1 U4828 ( .A1(n6027), .A2(n6284), .ZN(n8409) );
  NOR2_X1 U4829 ( .A1(n4753), .A2(n4965), .ZN(n7866) );
  INV_X4 U4830 ( .A(n5894), .ZN(n5644) );
  INV_X1 U4831 ( .A(n5540), .ZN(n6216) );
  NAND2_X1 U4832 ( .A1(n7730), .A2(n4686), .ZN(n4684) );
  INV_X2 U4834 ( .A(n8409), .ZN(n6381) );
  INV_X1 U4835 ( .A(n9912), .ZN(n4400) );
  NAND2_X1 U4836 ( .A1(n8054), .A2(n7783), .ZN(n7865) );
  AND4_X1 U4837 ( .A1(n5459), .A2(n5458), .A3(n5457), .A4(n5456), .ZN(n8505)
         );
  NAND2_X2 U4839 ( .A1(n5378), .A2(n5382), .ZN(n6039) );
  AOI21_X2 U4840 ( .B1(n8141), .B2(n8140), .A(n9211), .ZN(n9194) );
  OAI22_X1 U4841 ( .A1(n9194), .A2(n9195), .B1(n8147), .B2(n8146), .ZN(n9266)
         );
  INV_X1 U4842 ( .A(n5330), .ZN(n5275) );
  INV_X1 U4843 ( .A(n5039), .ZN(n7859) );
  NAND4_X1 U4844 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n8552)
         );
  INV_X2 U4845 ( .A(n8946), .ZN(n9019) );
  NAND2_X1 U4846 ( .A1(n9266), .A2(n4346), .ZN(n4661) );
  INV_X2 U4847 ( .A(n8213), .ZN(n5970) );
  INV_X2 U4848 ( .A(n6751), .ZN(n10001) );
  OAI21_X2 U4849 ( .B1(n7545), .B2(n7544), .A(n7543), .ZN(n7658) );
  OAI22_X2 U4850 ( .A1(n9543), .A2(n5141), .B1(n9283), .B2(n9556), .ZN(n9521)
         );
  OAI211_X2 U4851 ( .C1(n6075), .C2(n5523), .A(n5522), .B(n5521), .ZN(n6990)
         );
  INV_X2 U4852 ( .A(n5796), .ZN(n5544) );
  OAI211_X1 U4853 ( .C1(n6080), .C2(n5523), .A(n5498), .B(n5497), .ZN(n8509)
         );
  XNOR2_X2 U4854 ( .A(n5038), .B(n5037), .ZN(n6082) );
  NAND2_X1 U4855 ( .A1(n4599), .A2(n4833), .ZN(n5038) );
  XNOR2_X2 U4856 ( .A(n5340), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5342) );
  NAND2_X2 U4857 ( .A1(n5337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5340) );
  AND2_X4 U4858 ( .A1(n6285), .A2(n6291), .ZN(n8411) );
  OAI21_X1 U4859 ( .B1(n9487), .B2(n5259), .A(n5269), .ZN(n9375) );
  NAND2_X1 U4860 ( .A1(n4393), .A2(n4371), .ZN(n4392) );
  NAND2_X1 U4861 ( .A1(n9230), .A2(n9231), .ZN(n9229) );
  NOR2_X1 U4862 ( .A1(n4390), .A2(n8304), .ZN(n8795) );
  OR2_X1 U4863 ( .A1(n4338), .A2(n5267), .ZN(n9390) );
  NAND2_X1 U4864 ( .A1(n7664), .A2(n7663), .ZN(n7730) );
  OR2_X1 U4865 ( .A1(n8864), .A2(n8856), .ZN(n8865) );
  NAND2_X1 U4866 ( .A1(n5233), .A2(n5232), .ZN(n9601) );
  OR2_X1 U4867 ( .A1(n9687), .A2(n4510), .ZN(n4654) );
  NAND2_X1 U4868 ( .A1(n5215), .A2(n5214), .ZN(n9611) );
  NAND2_X1 U4869 ( .A1(n7286), .A2(n8261), .ZN(n7562) );
  OR2_X1 U4870 ( .A1(n6970), .A2(n4408), .ZN(n7286) );
  OR2_X1 U4871 ( .A1(n9851), .A2(n9842), .ZN(n9852) );
  NAND2_X1 U4872 ( .A1(n5092), .A2(n5091), .ZN(n7641) );
  INV_X2 U4873 ( .A(n9884), .ZN(n9856) );
  NAND2_X2 U4874 ( .A1(n6820), .A2(n8943), .ZN(n8946) );
  NAND2_X1 U4875 ( .A1(n8057), .A2(n9840), .ZN(n7864) );
  NAND2_X2 U4876 ( .A1(n6721), .A2(n9880), .ZN(n9884) );
  NAND4_X2 U4877 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n4970), .ZN(n9290)
         );
  INV_X1 U4878 ( .A(n9874), .ZN(n4444) );
  INV_X1 U4879 ( .A(n6658), .ZN(n7017) );
  NAND4_X1 U4880 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n9291)
         );
  OAI211_X1 U4881 ( .C1(n6039), .C2(n6148), .A(n4981), .B(n4980), .ZN(n9905)
         );
  OAI22_X1 U4882 ( .A1(n6985), .A2(n5970), .B1(n9979), .B2(n5644), .ZN(n6459)
         );
  NAND2_X1 U4883 ( .A1(n8554), .A2(n8213), .ZN(n5569) );
  OAI211_X1 U4884 ( .C1(n6086), .C2(n5523), .A(n5555), .B(n5554), .ZN(n6958)
         );
  AND3_X1 U4885 ( .A1(n5518), .A2(n5519), .A3(n4559), .ZN(n6472) );
  AND4_X1 U4886 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n6826)
         );
  INV_X1 U4887 ( .A(n5562), .ZN(n5816) );
  NAND2_X2 U4888 ( .A1(n6039), .A2(n5475), .ZN(n7857) );
  CLKBUF_X1 U4889 ( .A(n5382), .Z(n9755) );
  NAND2_X1 U4890 ( .A1(n4812), .A2(n4811), .ZN(n4990) );
  AND2_X1 U4892 ( .A1(n5448), .A2(n9158), .ZN(n7751) );
  NAND2_X2 U4893 ( .A1(n8388), .A2(n8193), .ZN(n5976) );
  OR2_X1 U4894 ( .A1(n5447), .A2(n5468), .ZN(n5445) );
  XNOR2_X1 U4895 ( .A(n4828), .B(n4827), .ZN(n5010) );
  MUX2_X1 U4896 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5470), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5472) );
  NOR2_X1 U4897 ( .A1(n4675), .A2(n4523), .ZN(n4522) );
  XNOR2_X1 U4898 ( .A(n4831), .B(SI_6_), .ZN(n5018) );
  OR2_X2 U4899 ( .A1(n7852), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9165) );
  OAI21_X1 U4900 ( .B1(n5769), .B2(n4719), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5947) );
  AND2_X1 U4901 ( .A1(n5753), .A2(n5443), .ZN(n4565) );
  INV_X1 U4902 ( .A(n4987), .ZN(n4766) );
  INV_X2 U4903 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AND2_X1 U4904 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7535) );
  NOR2_X1 U4905 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4412) );
  NOR2_X1 U4906 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4413) );
  INV_X1 U4907 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5460) );
  NOR2_X1 U4908 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5434) );
  INV_X1 U4909 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5950) );
  INV_X1 U4910 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5463) );
  OAI21_X1 U4911 ( .B1(n6034), .B2(n9922), .A(n4321), .ZN(n6021) );
  NAND2_X1 U4912 ( .A1(n9219), .A2(n9221), .ZN(n9220) );
  XNOR2_X1 U4913 ( .A(n4926), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5378) );
  XNOR2_X2 U4914 ( .A(n5864), .B(n5862), .ZN(n8481) );
  AOI211_X1 U4915 ( .C1(n4310), .C2(n8508), .A(n8507), .B(n8506), .ZN(n8514)
         );
  XNOR2_X2 U4916 ( .A(n5445), .B(n5444), .ZN(n5454) );
  INV_X1 U4917 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U4918 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  INV_X1 U4919 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U4920 ( .A1(n7839), .A2(n7838), .ZN(n7846) );
  NAND2_X1 U4921 ( .A1(n7834), .A2(n7833), .ZN(n7839) );
  OAI21_X1 U4922 ( .B1(n5205), .B2(n5204), .A(n4885), .ZN(n5221) );
  AND2_X1 U4923 ( .A1(n4889), .A2(n4888), .ZN(n5220) );
  NAND2_X1 U4924 ( .A1(n4454), .A2(n4456), .ZN(n4453) );
  NAND2_X1 U4925 ( .A1(n7915), .A2(n5352), .ZN(n7782) );
  AND2_X1 U4926 ( .A1(n7904), .A2(n7915), .ZN(n8058) );
  NAND2_X1 U4927 ( .A1(n8392), .A2(n8193), .ZN(n5483) );
  INV_X1 U4928 ( .A(n7751), .ZN(n4556) );
  OR2_X1 U4929 ( .A1(n9029), .A2(n8192), .ZN(n8347) );
  INV_X1 U4930 ( .A(n4544), .ZN(n4543) );
  NAND2_X1 U4931 ( .A1(n8806), .A2(n8693), .ZN(n4550) );
  AND2_X1 U4932 ( .A1(n8771), .A2(n8757), .ZN(n8762) );
  NOR2_X1 U4933 ( .A1(n6821), .A2(n6658), .ZN(n6904) );
  AND2_X1 U4934 ( .A1(n6284), .A2(n6442), .ZN(n6291) );
  NAND2_X1 U4935 ( .A1(n6585), .A2(n4383), .ZN(n6587) );
  INV_X1 U4936 ( .A(n6586), .ZN(n4383) );
  OR2_X1 U4937 ( .A1(n7862), .A2(n7861), .ZN(n8040) );
  AND2_X1 U4938 ( .A1(n5372), .A2(n9362), .ZN(n8066) );
  OR2_X1 U4939 ( .A1(n9591), .A2(n9380), .ZN(n7991) );
  INV_X1 U4940 ( .A(n4434), .ZN(n4433) );
  OAI21_X1 U4941 ( .B1(n5264), .B2(n4435), .A(n9420), .ZN(n4434) );
  INV_X1 U4942 ( .A(n7979), .ZN(n4435) );
  INV_X1 U4943 ( .A(n9827), .ZN(n4515) );
  NAND2_X1 U4944 ( .A1(n6394), .A2(n4444), .ZN(n8050) );
  NAND2_X1 U4946 ( .A1(n4919), .A2(n4918), .ZN(n5306) );
  OAI21_X1 U4947 ( .B1(n5143), .B2(n5142), .A(n4867), .ZN(n5159) );
  AND2_X1 U4948 ( .A1(n4843), .A2(n4842), .ZN(n5057) );
  AND2_X1 U4949 ( .A1(n5883), .A2(n6001), .ZN(n5884) );
  OR2_X1 U4950 ( .A1(n5889), .A2(n8796), .ZN(n5883) );
  NAND2_X1 U4951 ( .A1(n8434), .A2(n5822), .ZN(n8439) );
  AND2_X1 U4952 ( .A1(n5656), .A2(n5640), .ZN(n4711) );
  OR2_X1 U4953 ( .A1(n5574), .A2(n6910), .ZN(n5514) );
  XNOR2_X1 U4954 ( .A(n4566), .B(n8609), .ZN(n8595) );
  OR2_X1 U4955 ( .A1(n9042), .A2(n8545), .ZN(n8187) );
  OR2_X1 U4956 ( .A1(n9053), .A2(n8695), .ZN(n8696) );
  AOI21_X1 U4957 ( .B1(n4544), .B2(n4542), .A(n4541), .ZN(n4540) );
  INV_X1 U4958 ( .A(n4545), .ZN(n4542) );
  NAND2_X1 U4959 ( .A1(n4342), .A2(n4565), .ZN(n5471) );
  INV_X2 U4960 ( .A(n4824), .ZN(n5475) );
  OAI211_X1 U4961 ( .C1(n4522), .C2(n5164), .A(n4405), .B(n4777), .ZN(n4926)
         );
  NAND2_X1 U4962 ( .A1(n5132), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U4963 ( .A1(n4781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4928) );
  AND2_X1 U4964 ( .A1(n8170), .A2(n9669), .ZN(n4960) );
  AND2_X1 U4965 ( .A1(n8170), .A2(n4785), .ZN(n4958) );
  OR2_X1 U4966 ( .A1(n9577), .A2(n9282), .ZN(n8015) );
  NAND2_X1 U4967 ( .A1(n9438), .A2(n4369), .ZN(n9382) );
  INV_X1 U4968 ( .A(n9588), .ZN(n4526) );
  NOR2_X1 U4969 ( .A1(n9382), .A2(n5293), .ZN(n9356) );
  OAI21_X1 U4970 ( .B1(n9375), .B2(n5281), .A(n5280), .ZN(n7756) );
  OR2_X1 U4971 ( .A1(n9588), .A2(n9403), .ZN(n5280) );
  XNOR2_X1 U4972 ( .A(n9588), .B(n9198), .ZN(n9378) );
  INV_X1 U4973 ( .A(n7304), .ZN(n4447) );
  INV_X1 U4974 ( .A(n7857), .ZN(n5213) );
  OAI21_X1 U4975 ( .B1(n6890), .B2(n7911), .A(n5027), .ZN(n6720) );
  INV_X1 U4976 ( .A(n9529), .ZN(n9875) );
  XNOR2_X1 U4977 ( .A(n7856), .B(n7855), .ZN(n9157) );
  NAND2_X1 U4978 ( .A1(n7851), .A2(n7850), .ZN(n7856) );
  NAND2_X1 U4979 ( .A1(n4580), .A2(n4579), .ZN(n5250) );
  AOI21_X1 U4980 ( .B1(n4581), .B2(n4328), .A(n5248), .ZN(n4579) );
  OAI21_X1 U4981 ( .B1(n4314), .B2(n7561), .A(n4370), .ZN(n4458) );
  NOR2_X1 U4982 ( .A1(n4408), .A2(n7561), .ZN(n4459) );
  NAND2_X1 U4983 ( .A1(n8314), .A2(n8310), .ZN(n4466) );
  NOR2_X1 U4984 ( .A1(n4468), .A2(n8180), .ZN(n4467) );
  OAI21_X1 U4985 ( .B1(n7996), .B2(n7995), .A(n7997), .ZN(n4615) );
  NAND2_X1 U4986 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  INV_X1 U4987 ( .A(n4454), .ZN(n4450) );
  OR2_X1 U4988 ( .A1(n8671), .A2(n8904), .ZN(n8674) );
  AND2_X1 U4989 ( .A1(n6762), .A2(n10001), .ZN(n4734) );
  NAND2_X1 U4990 ( .A1(n8010), .A2(n7993), .ZN(n4616) );
  NAND2_X1 U4991 ( .A1(n4679), .A2(n4678), .ZN(n4677) );
  INV_X1 U4992 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4678) );
  INV_X1 U4993 ( .A(n4680), .ZN(n4679) );
  NAND2_X1 U4994 ( .A1(n4343), .A2(n4319), .ZN(n4523) );
  NOR2_X1 U4995 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4430) );
  NOR2_X1 U4996 ( .A1(n5051), .A2(n4490), .ZN(n4486) );
  INV_X1 U4997 ( .A(n5057), .ZN(n4490) );
  INV_X1 U4998 ( .A(n4843), .ZN(n4488) );
  NAND2_X1 U4999 ( .A1(n4840), .A2(n7449), .ZN(n4843) );
  INV_X1 U5000 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4799) );
  INV_X1 U5001 ( .A(n8519), .ZN(n4697) );
  AOI21_X1 U5002 ( .B1(n4558), .B2(n4557), .A(n7751), .ZN(n4560) );
  INV_X1 U5003 ( .A(n8187), .ZN(n4627) );
  INV_X1 U5004 ( .A(n4629), .ZN(n4628) );
  OR2_X1 U5005 ( .A1(n5922), .A2(n7371), .ZN(n5986) );
  NOR2_X1 U5006 ( .A1(n9072), .A2(n9077), .ZN(n4743) );
  OR2_X1 U5007 ( .A1(n9077), .A2(n8690), .ZN(n8310) );
  NOR2_X1 U5008 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  OR2_X1 U5009 ( .A1(n9106), .A2(n8908), .ZN(n8289) );
  NAND2_X1 U5010 ( .A1(n5718), .A2(n4644), .ZN(n8283) );
  NOR2_X1 U5011 ( .A1(n8977), .A2(n4645), .ZN(n4644) );
  INV_X1 U5012 ( .A(n5717), .ZN(n4645) );
  NAND2_X1 U5013 ( .A1(n9111), .A2(n8977), .ZN(n8284) );
  OR2_X1 U5014 ( .A1(n9121), .A2(n8978), .ZN(n8921) );
  NOR2_X1 U5015 ( .A1(n4731), .A2(n9121), .ZN(n4730) );
  INV_X1 U5016 ( .A(n4732), .ZN(n4731) );
  OR2_X1 U5017 ( .A1(n9127), .A2(n7600), .ZN(n8267) );
  AND2_X1 U5018 ( .A1(n6756), .A2(n8219), .ZN(n4402) );
  NAND2_X1 U5019 ( .A1(n4404), .A2(n8221), .ZN(n4403) );
  AND2_X1 U5020 ( .A1(n5621), .A2(n5620), .ZN(n5659) );
  INV_X1 U5021 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4416) );
  INV_X1 U5022 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U5023 ( .A1(n7205), .A2(n7270), .ZN(n4651) );
  INV_X1 U5024 ( .A(n8136), .ZN(n4499) );
  NAND2_X1 U5025 ( .A1(n9186), .A2(n9185), .ZN(n8131) );
  NOR2_X1 U5026 ( .A1(n7742), .A2(n4683), .ZN(n4682) );
  INV_X1 U5027 ( .A(n4685), .ZN(n4683) );
  INV_X1 U5028 ( .A(n8089), .ZN(n4504) );
  OAI21_X1 U5029 ( .B1(n4593), .B2(n8033), .A(n8037), .ZN(n4589) );
  OAI21_X1 U5030 ( .B1(n4593), .B2(n8034), .A(n4592), .ZN(n4591) );
  NAND2_X1 U5031 ( .A1(n8074), .A2(n8030), .ZN(n4592) );
  OR2_X1 U5032 ( .A1(n9572), .A2(n9272), .ZN(n8020) );
  OR2_X1 U5033 ( .A1(n9330), .A2(n9347), .ZN(n8023) );
  INV_X1 U5034 ( .A(n9378), .ZN(n4443) );
  INV_X1 U5035 ( .A(n4616), .ZN(n9361) );
  AND2_X1 U5036 ( .A1(n7899), .A2(n4422), .ZN(n4421) );
  NAND2_X1 U5037 ( .A1(n4425), .A2(n4423), .ZN(n4422) );
  INV_X1 U5038 ( .A(n7965), .ZN(n4423) );
  INV_X1 U5039 ( .A(n7818), .ZN(n4418) );
  NAND2_X1 U5040 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U5041 ( .A1(n5014), .A2(n5015), .ZN(n7904) );
  NAND2_X1 U5042 ( .A1(n4399), .A2(n9912), .ZN(n8057) );
  INV_X1 U5043 ( .A(n9845), .ZN(n4399) );
  INV_X1 U5044 ( .A(n5132), .ZN(n4774) );
  NAND2_X1 U5045 ( .A1(n4578), .A2(n5271), .ZN(n5283) );
  NAND2_X1 U5046 ( .A1(n4617), .A2(n4880), .ZN(n5205) );
  NAND2_X1 U5047 ( .A1(n5193), .A2(n4878), .ZN(n4617) );
  NOR2_X1 U5048 ( .A1(n5163), .A2(n5162), .ZN(n5179) );
  AND2_X1 U5049 ( .A1(n4605), .A2(n4862), .ZN(n4604) );
  NAND2_X1 U5050 ( .A1(n4852), .A2(n7471), .ZN(n4855) );
  AND4_X1 U5051 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4771)
         );
  INV_X1 U5052 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4768) );
  INV_X1 U5053 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4767) );
  OAI21_X1 U5054 ( .B1(n5088), .B2(n4851), .A(n4850), .ZN(n5103) );
  NAND2_X1 U5055 ( .A1(n4848), .A2(n4847), .ZN(n5088) );
  NAND2_X1 U5056 ( .A1(n4836), .A2(n4835), .ZN(n4839) );
  AOI21_X1 U5057 ( .B1(n4598), .B2(n5037), .A(n4355), .ZN(n4595) );
  INV_X1 U5058 ( .A(n4833), .ZN(n4598) );
  AND2_X1 U5059 ( .A1(n5037), .A2(n5018), .ZN(n4597) );
  OAI21_X1 U5060 ( .B1(n4824), .B2(n4813), .A(n4618), .ZN(n4814) );
  NAND2_X1 U5061 ( .A1(n4824), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4618) );
  NOR2_X1 U5062 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4952) );
  NAND2_X1 U5063 ( .A1(n5539), .A2(n4947), .ZN(n4594) );
  NOR2_X1 U5064 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NOR2_X1 U5065 ( .A1(n5556), .A2(n5557), .ZN(n4702) );
  NAND2_X1 U5066 ( .A1(n8466), .A2(n8467), .ZN(n4710) );
  AND2_X1 U5067 ( .A1(n5839), .A2(n5826), .ZN(n4712) );
  INV_X1 U5068 ( .A(n8475), .ZN(n5839) );
  OR2_X1 U5069 ( .A1(n5829), .A2(n7478), .ZN(n5856) );
  NAND2_X1 U5070 ( .A1(n5664), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5685) );
  INV_X1 U5071 ( .A(n5666), .ZN(n5664) );
  OR2_X1 U5072 ( .A1(n5645), .A2(n7463), .ZN(n5666) );
  NOR2_X1 U5073 ( .A1(n6042), .A2(n4709), .ZN(n4708) );
  INV_X1 U5074 ( .A(n5768), .ZN(n4709) );
  INV_X1 U5075 ( .A(n8467), .ZN(n4706) );
  INV_X1 U5076 ( .A(n5788), .ZN(n4705) );
  AND2_X1 U5077 ( .A1(n5821), .A2(n5805), .ZN(n8488) );
  NAND2_X1 U5078 ( .A1(n4697), .A2(n5904), .ZN(n4696) );
  NAND2_X1 U5079 ( .A1(n4471), .A2(n8358), .ZN(n4470) );
  OAI21_X1 U5080 ( .B1(n8345), .B2(n4475), .A(n4472), .ZN(n4471) );
  INV_X1 U5081 ( .A(n8357), .ZN(n4469) );
  AND2_X1 U5082 ( .A1(n5993), .A2(n5992), .ZN(n8188) );
  OR2_X1 U5083 ( .A1(n7131), .A2(n7130), .ZN(n4571) );
  OR2_X1 U5084 ( .A1(n8592), .A2(n4380), .ZN(n4566) );
  NAND2_X1 U5085 ( .A1(n8196), .A2(n8195), .ZN(n8639) );
  NAND2_X1 U5086 ( .A1(n8347), .A2(n8348), .ZN(n8700) );
  AND2_X1 U5087 ( .A1(n8762), .A2(n4322), .ZN(n8702) );
  NAND2_X1 U5088 ( .A1(n4552), .A2(n4554), .ZN(n8715) );
  AOI21_X1 U5089 ( .B1(n8728), .B2(n4555), .A(n4352), .ZN(n4554) );
  INV_X1 U5090 ( .A(n8697), .ZN(n4555) );
  NAND2_X1 U5091 ( .A1(n8343), .A2(n8341), .ZN(n8714) );
  OR2_X1 U5092 ( .A1(n8728), .A2(n4455), .ZN(n4629) );
  NAND2_X1 U5093 ( .A1(n8630), .A2(n8546), .ZN(n8697) );
  AND2_X1 U5094 ( .A1(n8185), .A2(n8328), .ZN(n8744) );
  NAND2_X1 U5095 ( .A1(n8795), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5096 ( .A1(n8744), .A2(n8186), .ZN(n8743) );
  NAND2_X1 U5097 ( .A1(n8738), .A2(n8742), .ZN(n8737) );
  AND2_X1 U5098 ( .A1(n5902), .A2(n5901), .ZN(n8781) );
  NAND2_X1 U5099 ( .A1(n8794), .A2(n8184), .ZN(n8775) );
  NAND2_X1 U5100 ( .A1(n8795), .A2(n4541), .ZN(n8794) );
  AND2_X1 U5101 ( .A1(n4550), .A2(n8692), .ZN(n4545) );
  NAND2_X1 U5102 ( .A1(n4362), .A2(n4550), .ZN(n4544) );
  OR2_X1 U5103 ( .A1(n8858), .A2(n9083), .ZN(n4754) );
  NOR2_X1 U5104 ( .A1(n4754), .A2(n9077), .ZN(n8830) );
  OR2_X1 U5105 ( .A1(n5793), .A2(n8493), .ZN(n5813) );
  OR2_X1 U5106 ( .A1(n8876), .A2(n4564), .ZN(n4563) );
  NOR2_X1 U5107 ( .A1(n9093), .A2(n8906), .ZN(n4564) );
  NAND2_X1 U5108 ( .A1(n5450), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5491) );
  INV_X1 U5109 ( .A(n5508), .ZN(n5450) );
  NOR2_X1 U5110 ( .A1(n4535), .A2(n6754), .ZN(n4534) );
  INV_X1 U5111 ( .A(n6749), .ZN(n4535) );
  INV_X1 U5112 ( .A(n9014), .ZN(n8968) );
  AND2_X1 U5113 ( .A1(n6217), .A2(n6662), .ZN(n8965) );
  NAND2_X1 U5114 ( .A1(n6656), .A2(n6837), .ZN(n6821) );
  XNOR2_X1 U5115 ( .A(n8554), .B(n6837), .ZN(n8363) );
  INV_X1 U5116 ( .A(n6958), .ZN(n6648) );
  NAND2_X1 U5118 ( .A1(n5921), .A2(n5920), .ZN(n9042) );
  NAND2_X1 U5119 ( .A1(n5893), .A2(n5892), .ZN(n9053) );
  NAND2_X1 U5120 ( .A1(n5869), .A2(n5868), .ZN(n9057) );
  AND2_X1 U5121 ( .A1(n5625), .A2(n5624), .ZN(n10011) );
  OR2_X1 U5122 ( .A1(n9973), .A2(n5961), .ZN(n6496) );
  XNOR2_X1 U5123 ( .A(n5474), .B(n5473), .ZN(n8398) );
  NAND2_X1 U5124 ( .A1(n5954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  AND2_X1 U5125 ( .A1(n5462), .A2(n5461), .ZN(n4721) );
  NOR2_X1 U5126 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5436) );
  NOR2_X1 U5127 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5435) );
  AND2_X1 U5128 ( .A1(n6598), .A2(n6587), .ZN(n4671) );
  NAND2_X1 U5129 ( .A1(n9176), .A2(n9177), .ZN(n9175) );
  XNOR2_X1 U5130 ( .A(n6382), .B(n6381), .ZN(n6383) );
  OR2_X1 U5131 ( .A1(n7063), .A2(n7064), .ZN(n4649) );
  NOR2_X1 U5132 ( .A1(n6290), .A2(n6289), .ZN(n6296) );
  NAND2_X1 U5133 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  OR2_X1 U5134 ( .A1(n7728), .A2(n7729), .ZN(n4686) );
  INV_X1 U5135 ( .A(n7891), .ZN(n5373) );
  XNOR2_X1 U5136 ( .A(n8029), .B(n9325), .ZN(n7891) );
  OAI21_X1 U5137 ( .B1(n9355), .B2(n4389), .A(n4385), .ZN(n9319) );
  INV_X1 U5138 ( .A(n4386), .ZN(n4385) );
  NAND2_X1 U5139 ( .A1(n9345), .A2(n7888), .ZN(n4389) );
  OAI21_X1 U5140 ( .B1(n8067), .B2(n4387), .A(n5318), .ZN(n4386) );
  NAND2_X1 U5141 ( .A1(n9362), .A2(n8010), .ZN(n7887) );
  AOI21_X1 U5142 ( .B1(n4433), .B2(n4435), .A(n4359), .ZN(n4431) );
  OR2_X1 U5143 ( .A1(n9377), .A2(n9378), .ZN(n9376) );
  AND2_X1 U5144 ( .A1(n7822), .A2(n9400), .ZN(n9420) );
  NAND2_X1 U5145 ( .A1(n5369), .A2(n5264), .ZN(n9434) );
  NAND2_X1 U5146 ( .A1(n9467), .A2(n4519), .ZN(n4518) );
  NOR2_X1 U5147 ( .A1(n4520), .A2(n9606), .ZN(n4519) );
  AND2_X1 U5148 ( .A1(n7897), .A2(n7818), .ZN(n9486) );
  AOI21_X1 U5149 ( .B1(n5367), .B2(n7965), .A(n4426), .ZN(n4425) );
  INV_X1 U5150 ( .A(n7863), .ZN(n4426) );
  NAND2_X1 U5151 ( .A1(n9515), .A2(n7965), .ZN(n4420) );
  OR2_X1 U5152 ( .A1(n9630), .A2(n9530), .ZN(n7965) );
  OR2_X1 U5153 ( .A1(n9533), .A2(n9630), .ZN(n9507) );
  OAI21_X1 U5154 ( .B1(n9521), .B2(n5157), .A(n5156), .ZN(n9506) );
  NAND2_X1 U5155 ( .A1(n4438), .A2(n4436), .ZN(n9522) );
  NOR2_X1 U5156 ( .A1(n9525), .A2(n4437), .ZN(n4436) );
  INV_X1 U5157 ( .A(n7930), .ZN(n4437) );
  NAND2_X1 U5158 ( .A1(n7693), .A2(n4439), .ZN(n4438) );
  NOR2_X1 U5159 ( .A1(n4440), .A2(n9544), .ZN(n4439) );
  INV_X1 U5160 ( .A(n7794), .ZN(n4440) );
  NAND2_X1 U5161 ( .A1(n5134), .A2(n5133), .ZN(n9556) );
  NAND2_X1 U5162 ( .A1(n5119), .A2(n5118), .ZN(n7702) );
  OR2_X1 U5163 ( .A1(n7583), .A2(n7187), .ZN(n4756) );
  OAI21_X1 U5164 ( .B1(n6938), .B2(n5359), .A(n7923), .ZN(n7304) );
  NOR2_X1 U5165 ( .A1(n7872), .A2(n4410), .ZN(n4409) );
  INV_X1 U5166 ( .A(n5042), .ZN(n4410) );
  OR2_X1 U5167 ( .A1(n5039), .A2(n6080), .ZN(n5020) );
  NAND2_X1 U5168 ( .A1(n5351), .A2(n8054), .ZN(n6556) );
  NAND2_X1 U5169 ( .A1(n4967), .A2(n4966), .ZN(n6635) );
  INV_X1 U5170 ( .A(n7866), .ZN(n4966) );
  NOR2_X1 U5171 ( .A1(n9862), .A2(n6394), .ZN(n6639) );
  OR2_X1 U5172 ( .A1(n6378), .A2(n9860), .ZN(n9862) );
  INV_X1 U5173 ( .A(n9531), .ZN(n9873) );
  NAND2_X1 U5174 ( .A1(n5184), .A2(n5183), .ZN(n9623) );
  XNOR2_X1 U5175 ( .A(n4784), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4785) );
  XNOR2_X1 U5176 ( .A(n7846), .B(n7845), .ZN(n9161) );
  XNOR2_X1 U5177 ( .A(n4780), .B(n4779), .ZN(n4786) );
  INV_X1 U5178 ( .A(n4893), .ZN(n4583) );
  INV_X1 U5179 ( .A(n4582), .ZN(n4581) );
  OAI21_X1 U5180 ( .B1(n4585), .B2(n4328), .A(n4899), .ZN(n4582) );
  NAND2_X1 U5181 ( .A1(n4584), .A2(n4893), .ZN(n5240) );
  NAND2_X1 U5182 ( .A1(n4890), .A2(n4585), .ZN(n4584) );
  INV_X1 U5183 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5209) );
  XNOR2_X1 U5184 ( .A(n5103), .B(n5102), .ZN(n6111) );
  XNOR2_X1 U5185 ( .A(n4834), .B(n7460), .ZN(n5037) );
  INV_X1 U5186 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U5187 ( .A1(n6618), .A2(n5636), .ZN(n6622) );
  AND2_X1 U5188 ( .A1(n6518), .A2(n6517), .ZN(n8192) );
  AND2_X1 U5189 ( .A1(n8193), .A2(n8888), .ZN(n4716) );
  NAND2_X1 U5190 ( .A1(n5983), .A2(n5968), .ZN(n8518) );
  INV_X1 U5191 ( .A(n8508), .ZN(n8544) );
  INV_X1 U5192 ( .A(n8188), .ZN(n8725) );
  NOR2_X1 U5193 ( .A1(n5553), .A2(n4573), .ZN(n8561) );
  OAI21_X1 U5194 ( .B1(n4576), .B2(n5551), .A(n4574), .ZN(n4573) );
  NAND2_X1 U5195 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4576) );
  NOR2_X1 U5196 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5551) );
  NOR2_X1 U5197 ( .A1(n7712), .A2(n7711), .ZN(n8592) );
  NAND2_X1 U5198 ( .A1(n8207), .A2(n8206), .ZN(n9025) );
  NAND2_X1 U5199 ( .A1(n5253), .A2(n5252), .ZN(n9591) );
  INV_X1 U5200 ( .A(n9403), .ZN(n9198) );
  NAND2_X1 U5201 ( .A1(n7651), .A2(n7859), .ZN(n5286) );
  NAND2_X1 U5202 ( .A1(n5065), .A2(n5064), .ZN(n9827) );
  OR2_X1 U5203 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  NAND2_X1 U5204 ( .A1(n6039), .A2(n4323), .ZN(n4957) );
  OR2_X1 U5205 ( .A1(n4955), .A2(n6086), .ZN(n4956) );
  NAND2_X1 U5206 ( .A1(n5298), .A2(n5297), .ZN(n9577) );
  NAND2_X1 U5207 ( .A1(n7676), .A2(n7859), .ZN(n5298) );
  MUX2_X1 U5208 ( .A(n8044), .B(n8043), .S(n9867), .Z(n8081) );
  NAND2_X1 U5209 ( .A1(n8048), .A2(n8047), .ZN(n8080) );
  NAND4_X1 U5210 ( .A1(n5098), .A2(n5097), .A3(n5096), .A4(n5095), .ZN(n9684)
         );
  AOI21_X1 U5211 ( .B1(n9157), .B2(n7859), .A(n7858), .ZN(n9701) );
  XNOR2_X1 U5212 ( .A(n9563), .B(n9701), .ZN(n9703) );
  NAND2_X1 U5213 ( .A1(n9313), .A2(n9566), .ZN(n9563) );
  NAND2_X1 U5214 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U5215 ( .A1(n5273), .A2(n5272), .ZN(n9588) );
  OR2_X1 U5216 ( .A1(n9946), .A2(n6025), .ZN(n9880) );
  INV_X1 U5217 ( .A(n9440), .ZN(n9504) );
  AOI21_X1 U5218 ( .B1(n5340), .B2(n5339), .A(n5164), .ZN(n4382) );
  NAND2_X1 U5219 ( .A1(n4461), .A2(n8371), .ZN(n4460) );
  INV_X1 U5220 ( .A(n8257), .ZN(n4461) );
  OR2_X1 U5221 ( .A1(n8273), .A2(n8272), .ZN(n8277) );
  AND2_X1 U5222 ( .A1(n8377), .A2(n8290), .ZN(n4476) );
  INV_X1 U5223 ( .A(n8330), .ZN(n4456) );
  AOI21_X1 U5224 ( .B1(n8330), .B2(n4353), .A(n4455), .ZN(n4454) );
  NOR2_X1 U5225 ( .A1(n8304), .A2(n8346), .ZN(n4464) );
  AOI21_X1 U5226 ( .B1(n8303), .B2(n4467), .A(n4466), .ZN(n4465) );
  NAND2_X1 U5227 ( .A1(n8305), .A2(n8346), .ZN(n4462) );
  OAI21_X1 U5228 ( .B1(n4616), .B2(n4615), .A(n4613), .ZN(n8000) );
  INV_X1 U5229 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U5230 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4429) );
  OAI21_X1 U5231 ( .B1(n8326), .B2(n4452), .A(n4324), .ZN(n8338) );
  INV_X1 U5232 ( .A(n8217), .ZN(n4643) );
  NAND2_X1 U5233 ( .A1(n6479), .A2(n6478), .ZN(n8229) );
  INV_X1 U5234 ( .A(n5106), .ZN(n4509) );
  AOI21_X1 U5235 ( .B1(n5106), .B2(n5039), .A(n7186), .ZN(n4508) );
  INV_X1 U5236 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5160) );
  NOR2_X1 U5237 ( .A1(n4607), .A2(n4602), .ZN(n4601) );
  INV_X1 U5238 ( .A(n4847), .ZN(n4602) );
  NAND2_X1 U5239 ( .A1(n4608), .A2(n5130), .ZN(n4607) );
  INV_X1 U5240 ( .A(n4611), .ZN(n4606) );
  INV_X1 U5241 ( .A(n4859), .ZN(n4621) );
  INV_X1 U5242 ( .A(n4855), .ZN(n4622) );
  NAND2_X1 U5243 ( .A1(n5115), .A2(n4623), .ZN(n4619) );
  INV_X1 U5244 ( .A(n6502), .ZN(n5585) );
  NAND2_X1 U5245 ( .A1(n8449), .A2(n5851), .ZN(n5864) );
  NOR2_X1 U5246 ( .A1(n4474), .A2(n4473), .ZN(n4472) );
  NAND2_X1 U5247 ( .A1(n8351), .A2(n8350), .ZN(n4473) );
  INV_X1 U5248 ( .A(n8349), .ZN(n4474) );
  OR2_X1 U5249 ( .A1(n8700), .A2(n8344), .ZN(n4475) );
  OR2_X1 U5250 ( .A1(n9025), .A2(n8209), .ZN(n8353) );
  NOR2_X1 U5251 ( .A1(n8724), .A2(n8186), .ZN(n4553) );
  AND2_X1 U5252 ( .A1(n4737), .A2(n4738), .ZN(n4736) );
  NOR2_X1 U5253 ( .A1(n9042), .A2(n9048), .ZN(n4738) );
  NOR2_X1 U5254 ( .A1(n4643), .A2(n8788), .ZN(n4642) );
  OR2_X1 U5255 ( .A1(n9048), .A2(n8546), .ZN(n8334) );
  AND2_X1 U5256 ( .A1(n8217), .A2(n8319), .ZN(n8776) );
  NAND2_X1 U5257 ( .A1(n8806), .A2(n4743), .ZN(n4742) );
  OR2_X1 U5258 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  OR2_X1 U5259 ( .A1(n8179), .A2(n8178), .ZN(n8902) );
  NAND2_X1 U5260 ( .A1(n8176), .A2(n4313), .ZN(n8903) );
  NOR2_X1 U5261 ( .A1(n8652), .A2(n9127), .ZN(n4732) );
  NAND2_X1 U5262 ( .A1(n8555), .A2(n6648), .ZN(n8230) );
  NAND2_X1 U5263 ( .A1(n6483), .A2(n9986), .ZN(n6478) );
  INV_X1 U5264 ( .A(n6496), .ZN(n6816) );
  NAND2_X1 U5265 ( .A1(n6904), .A2(n4318), .ZN(n4760) );
  NAND2_X1 U5266 ( .A1(n6904), .A2(n4734), .ZN(n6880) );
  NAND2_X1 U5267 ( .A1(n6654), .A2(n8232), .ZN(n6824) );
  AND2_X1 U5268 ( .A1(n5442), .A2(n4725), .ZN(n4724) );
  NOR2_X1 U5269 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4725) );
  NAND2_X1 U5270 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U5271 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4720) );
  NOR2_X1 U5272 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5433) );
  INV_X1 U5273 ( .A(n5609), .ZN(n5617) );
  AND2_X1 U5274 ( .A1(n9244), .A2(n4499), .ZN(n4497) );
  OR2_X1 U5275 ( .A1(n4498), .A2(n9244), .ZN(n4496) );
  XNOR2_X1 U5276 ( .A(n7188), .B(n6381), .ZN(n7192) );
  NAND2_X1 U5277 ( .A1(n4506), .A2(n4505), .ZN(n7188) );
  NAND2_X1 U5278 ( .A1(n6111), .A2(n4508), .ZN(n4506) );
  AOI21_X1 U5279 ( .B1(n4508), .B2(n4509), .A(n4351), .ZN(n4505) );
  INV_X1 U5280 ( .A(n7202), .ZN(n4510) );
  INV_X1 U5281 ( .A(n7269), .ZN(n4653) );
  AND2_X1 U5282 ( .A1(n8130), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5283 ( .A1(n4388), .A2(n7888), .ZN(n4387) );
  INV_X1 U5284 ( .A(n8015), .ZN(n4388) );
  NAND2_X1 U5285 ( .A1(n5293), .A2(n9381), .ZN(n8010) );
  NAND2_X1 U5286 ( .A1(n4614), .A2(n9367), .ZN(n9362) );
  NOR2_X1 U5287 ( .A1(n9597), .A2(n9591), .ZN(n4527) );
  INV_X1 U5288 ( .A(n9491), .ZN(n4393) );
  OR2_X1 U5289 ( .A1(n9618), .A2(n9623), .ZN(n4520) );
  AND2_X1 U5290 ( .A1(n9553), .A2(n9714), .ZN(n9532) );
  OR2_X1 U5291 ( .A1(n5067), .A2(n5066), .ZN(n5079) );
  AND2_X1 U5292 ( .A1(n7782), .A2(n7781), .ZN(n5354) );
  NAND2_X1 U5293 ( .A1(n6930), .A2(n5026), .ZN(n7915) );
  NAND2_X1 U5294 ( .A1(n4400), .A2(n9845), .ZN(n9840) );
  INV_X1 U5295 ( .A(n8050), .ZN(n4965) );
  NOR2_X1 U5296 ( .A1(n6394), .A2(n4444), .ZN(n4753) );
  NAND2_X1 U5297 ( .A1(n4676), .A2(n4776), .ZN(n4675) );
  INV_X1 U5298 ( .A(n4677), .ZN(n4676) );
  NAND2_X1 U5299 ( .A1(n5325), .A2(n5324), .ZN(n7834) );
  NAND2_X1 U5300 ( .A1(n5320), .A2(n5319), .ZN(n5325) );
  NAND2_X1 U5301 ( .A1(n4914), .A2(n4913), .ZN(n5296) );
  NAND2_X1 U5302 ( .A1(n4775), .A2(n4681), .ZN(n4680) );
  INV_X1 U5303 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4681) );
  INV_X1 U5304 ( .A(n4523), .ZN(n4773) );
  NAND2_X1 U5305 ( .A1(n5250), .A2(n4905), .ZN(n5270) );
  NOR2_X1 U5306 ( .A1(n4894), .A2(n4586), .ZN(n4585) );
  INV_X1 U5307 ( .A(n4889), .ZN(n4586) );
  NOR2_X1 U5308 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4381) );
  NOR2_X1 U5309 ( .A1(n4619), .A2(n4612), .ZN(n4611) );
  INV_X1 U5310 ( .A(n4850), .ZN(n4612) );
  INV_X1 U5311 ( .A(n4609), .ZN(n4608) );
  OAI21_X1 U5312 ( .B1(n4619), .B2(n4610), .A(n4620), .ZN(n4609) );
  NAND2_X1 U5313 ( .A1(n4851), .A2(n4850), .ZN(n4610) );
  AOI21_X1 U5314 ( .B1(n5115), .B2(n4622), .A(n4621), .ZN(n4620) );
  XNOR2_X1 U5315 ( .A(n4849), .B(n7375), .ZN(n5087) );
  AOI21_X1 U5316 ( .B1(n5057), .B2(n4489), .A(n4488), .ZN(n4487) );
  INV_X1 U5317 ( .A(n4839), .ZN(n4489) );
  OR2_X1 U5318 ( .A1(n5049), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5059) );
  OAI21_X1 U5319 ( .B1(n7852), .B2(n4826), .A(n4825), .ZN(n4828) );
  NAND2_X1 U5320 ( .A1(n7852), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U5321 ( .A1(n7535), .A2(n4800), .ZN(n4801) );
  INV_X1 U5322 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4800) );
  NAND2_X1 U5323 ( .A1(n4696), .A2(n5972), .ZN(n4695) );
  AND2_X1 U5324 ( .A1(n5890), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5325 ( .A1(n4695), .A2(n4691), .ZN(n4690) );
  INV_X1 U5326 ( .A(n4758), .ZN(n4691) );
  NAND2_X1 U5327 ( .A1(n5590), .A2(n5589), .ZN(n6052) );
  INV_X1 U5328 ( .A(n6459), .ZN(n5541) );
  AND3_X1 U5329 ( .A1(n5834), .A2(n5833), .A3(n5832), .ZN(n8690) );
  NAND2_X1 U5330 ( .A1(n5468), .A2(n4575), .ZN(n4574) );
  INV_X1 U5331 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4575) );
  NOR2_X1 U5332 ( .A1(n7241), .A2(n4569), .ZN(n6741) );
  AND2_X1 U5333 ( .A1(n7246), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5334 ( .A1(n6741), .A2(n6740), .ZN(n6783) );
  NAND2_X1 U5335 ( .A1(n6783), .A2(n4568), .ZN(n6785) );
  OR2_X1 U5336 ( .A1(n6784), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4568) );
  NAND2_X1 U5337 ( .A1(n6785), .A2(n6786), .ZN(n7161) );
  AOI21_X1 U5338 ( .B1(n8743), .B2(n4345), .A(n4625), .ZN(n8643) );
  NAND2_X1 U5339 ( .A1(n4626), .A2(n8343), .ZN(n4625) );
  NAND2_X1 U5340 ( .A1(n8383), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U5341 ( .A1(n8762), .A2(n4736), .ZN(n8716) );
  AND2_X1 U5342 ( .A1(n5986), .A2(n5923), .ZN(n8732) );
  NAND2_X1 U5343 ( .A1(n8762), .A2(n4738), .ZN(n8730) );
  NAND2_X1 U5344 ( .A1(n8743), .A2(n8331), .ZN(n4398) );
  NAND2_X1 U5345 ( .A1(n8725), .A2(n8968), .ZN(n4396) );
  NOR2_X1 U5346 ( .A1(n8790), .A2(n9057), .ZN(n8771) );
  NAND2_X1 U5347 ( .A1(n4538), .A2(n4537), .ZN(n8770) );
  AOI21_X1 U5348 ( .B1(n4540), .B2(n4543), .A(n4372), .ZN(n4537) );
  AOI21_X1 U5349 ( .B1(n8846), .B2(n4633), .A(n4391), .ZN(n4390) );
  OAI21_X1 U5350 ( .B1(n4634), .B2(n8181), .A(n8183), .ZN(n4391) );
  AOI21_X1 U5351 ( .B1(n8181), .B2(n8844), .A(n4637), .ZN(n4636) );
  INV_X1 U5352 ( .A(n8310), .ZN(n4637) );
  NAND2_X1 U5353 ( .A1(n4358), .A2(n4633), .ZN(n8820) );
  NOR2_X1 U5354 ( .A1(n4754), .A2(n4741), .ZN(n8815) );
  INV_X1 U5355 ( .A(n4743), .ZN(n4741) );
  NAND2_X1 U5356 ( .A1(n5811), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5829) );
  INV_X1 U5357 ( .A(n5813), .ZN(n5811) );
  AOI21_X1 U5358 ( .B1(n4563), .B2(n4562), .A(n4561), .ZN(n8845) );
  NAND2_X1 U5359 ( .A1(n9087), .A2(n8879), .ZN(n4562) );
  NOR2_X1 U5360 ( .A1(n9087), .A2(n8879), .ZN(n4561) );
  NOR2_X1 U5361 ( .A1(n8914), .A2(n9093), .ZN(n8887) );
  NAND2_X1 U5362 ( .A1(n8887), .A2(n8863), .ZN(n8858) );
  NAND2_X1 U5363 ( .A1(n4406), .A2(n8291), .ZN(n8878) );
  NAND2_X1 U5364 ( .A1(n8903), .A2(n4407), .ZN(n4406) );
  AND2_X1 U5365 ( .A1(n8902), .A2(n8292), .ZN(n4407) );
  INV_X1 U5366 ( .A(n5776), .ZN(n5775) );
  OR2_X1 U5367 ( .A1(n5759), .A2(n7440), .ZN(n5776) );
  NAND2_X1 U5368 ( .A1(n4727), .A2(n4726), .ZN(n8914) );
  NAND2_X1 U5369 ( .A1(n5740), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5759) );
  INV_X1 U5370 ( .A(n5742), .ZN(n5740) );
  NAND2_X1 U5371 ( .A1(n8933), .A2(n8938), .ZN(n8934) );
  AND2_X1 U5372 ( .A1(n8284), .A2(n4364), .ZN(n8961) );
  AND2_X1 U5373 ( .A1(n8284), .A2(n8283), .ZN(n8963) );
  AND2_X1 U5374 ( .A1(n8896), .A2(n8895), .ZN(n8981) );
  AND2_X1 U5375 ( .A1(n7572), .A2(n4728), .ZN(n8987) );
  NOR2_X1 U5376 ( .A1(n9116), .A2(n4729), .ZN(n4728) );
  INV_X1 U5377 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5378 ( .B1(n8173), .B2(n8664), .A(n8274), .ZN(n9011) );
  OR2_X1 U5379 ( .A1(n9011), .A2(n8654), .ZN(n9017) );
  NAND2_X1 U5380 ( .A1(n7572), .A2(n4732), .ZN(n9003) );
  NAND2_X1 U5381 ( .A1(n7598), .A2(n8267), .ZN(n8173) );
  NAND2_X1 U5382 ( .A1(n7572), .A2(n7571), .ZN(n7601) );
  AND2_X1 U5383 ( .A1(n8267), .A2(n8266), .ZN(n8658) );
  OR2_X1 U5384 ( .A1(n8656), .A2(n8655), .ZN(n7558) );
  AND2_X1 U5385 ( .A1(n6904), .A2(n4374), .ZN(n7293) );
  AND2_X1 U5386 ( .A1(n7293), .A2(n10011), .ZN(n7572) );
  NAND2_X1 U5387 ( .A1(n6969), .A2(n8256), .ZN(n6970) );
  INV_X1 U5388 ( .A(n8965), .ZN(n9012) );
  NOR2_X1 U5389 ( .A1(n4533), .A2(n6758), .ZN(n4531) );
  INV_X1 U5390 ( .A(n4534), .ZN(n4533) );
  INV_X1 U5391 ( .A(n4530), .ZN(n4529) );
  OAI21_X1 U5392 ( .B1(n6753), .B2(n6758), .A(n4357), .ZN(n4530) );
  AND2_X1 U5393 ( .A1(n4401), .A2(n4403), .ZN(n6757) );
  NAND2_X1 U5394 ( .A1(n5449), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U5395 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5573) );
  NAND2_X1 U5396 ( .A1(n5828), .A2(n5827), .ZN(n9077) );
  NAND2_X1 U5397 ( .A1(n5738), .A2(n5737), .ZN(n9106) );
  NAND2_X1 U5398 ( .A1(n5718), .A2(n5717), .ZN(n9111) );
  INV_X1 U5399 ( .A(n10024), .ZN(n9125) );
  AND2_X1 U5400 ( .A1(n7656), .A2(n5952), .ZN(n5956) );
  NAND2_X1 U5401 ( .A1(n5753), .A2(n4724), .ZN(n5954) );
  AND2_X1 U5402 ( .A1(n5442), .A2(n4723), .ZN(n4722) );
  INV_X1 U5403 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5404 ( .A1(n5465), .A2(n5468), .ZN(n4715) );
  AOI21_X1 U5405 ( .B1(n5464), .B2(P2_IR_REG_31__SCAN_IN), .A(
        P2_IR_REG_20__SCAN_IN), .ZN(n4714) );
  AND2_X1 U5406 ( .A1(n5659), .A2(n5658), .ZN(n5679) );
  NOR2_X1 U5407 ( .A1(n5552), .A2(n4703), .ZN(n5502) );
  NAND2_X1 U5408 ( .A1(n5429), .A2(n4416), .ZN(n4703) );
  AND2_X1 U5409 ( .A1(n4493), .A2(n4494), .ZN(n8139) );
  AND2_X1 U5410 ( .A1(n4496), .A2(n4495), .ZN(n4494) );
  OR2_X1 U5411 ( .A1(n8131), .A2(n4497), .ZN(n4493) );
  OR2_X1 U5412 ( .A1(n8130), .A2(n4499), .ZN(n4495) );
  AND2_X1 U5413 ( .A1(n6377), .A2(n6376), .ZN(n6384) );
  XNOR2_X1 U5414 ( .A(n7192), .B(n7191), .ZN(n9691) );
  AND2_X1 U5415 ( .A1(n9691), .A2(n9686), .ZN(n9687) );
  NAND2_X1 U5416 ( .A1(n7728), .A2(n7729), .ZN(n4685) );
  AND2_X1 U5417 ( .A1(n5185), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5198) );
  AOI21_X1 U5418 ( .B1(n9241), .B2(n4670), .A(n9168), .ZN(n4669) );
  NAND2_X1 U5419 ( .A1(n9246), .A2(n4670), .ZN(n4666) );
  NAND2_X1 U5420 ( .A1(n8139), .A2(n8138), .ZN(n9167) );
  NAND2_X1 U5421 ( .A1(n7063), .A2(n7064), .ZN(n4648) );
  NAND2_X1 U5422 ( .A1(n9175), .A2(n8113), .ZN(n9230) );
  AND2_X1 U5423 ( .A1(n5243), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5254) );
  AOI21_X1 U5424 ( .B1(n8131), .B2(n8130), .A(n4499), .ZN(n9241) );
  NOR2_X1 U5425 ( .A1(n7273), .A2(n7201), .ZN(n7275) );
  XNOR2_X1 U5426 ( .A(n7200), .B(n7199), .ZN(n7273) );
  NAND2_X1 U5427 ( .A1(n4502), .A2(n4504), .ZN(n4501) );
  AOI21_X1 U5428 ( .B1(n9618), .B2(n8412), .A(n8103), .ZN(n9255) );
  INV_X1 U5429 ( .A(n8040), .ZN(n8071) );
  AND2_X1 U5430 ( .A1(n8039), .A2(n8040), .ZN(n4587) );
  NAND2_X1 U5431 ( .A1(n4589), .A2(n7997), .ZN(n4588) );
  AND2_X1 U5432 ( .A1(n9356), .A2(n4365), .ZN(n9313) );
  AND2_X1 U5433 ( .A1(n8023), .A2(n8024), .ZN(n9323) );
  OAI21_X1 U5434 ( .B1(n9377), .B2(n4442), .A(n4441), .ZN(n9346) );
  NAND2_X1 U5435 ( .A1(n4315), .A2(n4349), .ZN(n4441) );
  NAND2_X1 U5436 ( .A1(n4315), .A2(n4443), .ZN(n4442) );
  OR2_X1 U5437 ( .A1(n9346), .A2(n9345), .ZN(n9350) );
  NAND2_X1 U5438 ( .A1(n9356), .A2(n4316), .ZN(n9339) );
  NAND2_X1 U5439 ( .A1(n9438), .A2(n4527), .ZN(n9393) );
  NOR2_X1 U5440 ( .A1(n9449), .A2(n9601), .ZN(n9438) );
  NAND2_X1 U5441 ( .A1(n9438), .A2(n9418), .ZN(n9412) );
  NOR2_X1 U5442 ( .A1(n5234), .A2(n9187), .ZN(n5243) );
  AOI21_X1 U5443 ( .B1(n4421), .B2(n4424), .A(n4418), .ZN(n4417) );
  INV_X1 U5444 ( .A(n4425), .ZN(n4424) );
  NOR2_X1 U5445 ( .A1(n9507), .A2(n9623), .ZN(n9492) );
  NOR2_X1 U5446 ( .A1(n5150), .A2(n5149), .ZN(n5168) );
  NAND2_X1 U5447 ( .A1(n7693), .A2(n7794), .ZN(n9546) );
  OR2_X1 U5448 ( .A1(n5121), .A2(n5120), .ZN(n5135) );
  NOR2_X1 U5449 ( .A1(n4756), .A2(n7702), .ZN(n9553) );
  NAND2_X1 U5450 ( .A1(n5101), .A2(n5100), .ZN(n7581) );
  NAND2_X1 U5451 ( .A1(n4507), .A2(n5106), .ZN(n7187) );
  NOR2_X1 U5452 ( .A1(n5079), .A2(n6256), .ZN(n5093) );
  OAI21_X1 U5453 ( .B1(n7304), .B2(n4360), .A(n7952), .ZN(n7589) );
  INV_X1 U5454 ( .A(n7927), .ZN(n4446) );
  NOR2_X1 U5455 ( .A1(n4513), .A2(n7641), .ZN(n4511) );
  NAND2_X1 U5456 ( .A1(n5389), .A2(n4329), .ZN(n7301) );
  AOI21_X1 U5457 ( .B1(n7300), .B2(n5073), .A(n4761), .ZN(n7262) );
  NAND2_X1 U5458 ( .A1(n4448), .A2(n7916), .ZN(n6938) );
  NAND2_X1 U5459 ( .A1(n5389), .A2(n5055), .ZN(n7303) );
  NOR2_X1 U5460 ( .A1(n6562), .A2(n4525), .ZN(n6893) );
  NOR2_X1 U5461 ( .A1(n6562), .A2(n4524), .ZN(n9836) );
  NAND2_X1 U5462 ( .A1(n9839), .A2(n4400), .ZN(n4524) );
  NAND2_X1 U5463 ( .A1(n5388), .A2(n4400), .ZN(n9837) );
  INV_X1 U5464 ( .A(n6562), .ZN(n5388) );
  AND2_X1 U5465 ( .A1(n6440), .A2(n9889), .ZN(n6300) );
  NAND2_X1 U5466 ( .A1(n5309), .A2(n5308), .ZN(n9572) );
  NAND2_X1 U5467 ( .A1(n5148), .A2(n5147), .ZN(n9635) );
  OR2_X1 U5468 ( .A1(n7857), .A2(n6088), .ZN(n4981) );
  NAND3_X1 U5469 ( .A1(n5417), .A2(n5416), .A3(n5421), .ZN(n6442) );
  NAND2_X1 U5470 ( .A1(n4774), .A2(n4522), .ZN(n4781) );
  XNOR2_X1 U5471 ( .A(n7834), .B(n7833), .ZN(n8189) );
  NAND2_X1 U5472 ( .A1(n4925), .A2(n4924), .ZN(n5320) );
  NAND2_X1 U5473 ( .A1(n5306), .A2(n5305), .ZN(n4925) );
  XNOR2_X1 U5474 ( .A(n5306), .B(n5305), .ZN(n7679) );
  XNOR2_X1 U5475 ( .A(n5296), .B(n5295), .ZN(n7676) );
  XNOR2_X1 U5476 ( .A(n4577), .B(n5284), .ZN(n7651) );
  NAND2_X1 U5477 ( .A1(n5336), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5341) );
  INV_X1 U5478 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5161) );
  XNOR2_X1 U5479 ( .A(n5131), .B(n5130), .ZN(n6277) );
  NAND2_X1 U5480 ( .A1(n4603), .A2(n4608), .ZN(n5131) );
  NAND2_X1 U5481 ( .A1(n5088), .A2(n4611), .ZN(n4603) );
  OAI21_X1 U5482 ( .B1(n5103), .B2(n5102), .A(n4855), .ZN(n5116) );
  NOR2_X1 U5483 ( .A1(n4672), .A2(n4674), .ZN(n5104) );
  INV_X1 U5484 ( .A(n4771), .ZN(n4672) );
  NAND2_X1 U5485 ( .A1(n4491), .A2(n4839), .ZN(n5058) );
  NAND2_X1 U5486 ( .A1(n4354), .A2(n4596), .ZN(n4491) );
  NAND2_X1 U5487 ( .A1(n4823), .A2(n4822), .ZN(n5011) );
  XNOR2_X1 U5488 ( .A(n4814), .B(n7385), .ZN(n4993) );
  NAND2_X1 U5489 ( .A1(n4688), .A2(n4693), .ZN(n7767) );
  AND2_X1 U5490 ( .A1(n4694), .A2(n5973), .ZN(n4693) );
  NAND2_X1 U5491 ( .A1(n5891), .A2(n4689), .ZN(n4688) );
  OR2_X1 U5492 ( .A1(n4340), .A2(n4695), .ZN(n4694) );
  AND4_X1 U5493 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n9015)
         );
  OAI21_X1 U5494 ( .B1(n6531), .B2(n6530), .A(n4701), .ZN(n6525) );
  INV_X1 U5495 ( .A(n4702), .ZN(n4701) );
  AND4_X1 U5496 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n9013)
         );
  NAND2_X1 U5497 ( .A1(n5683), .A2(n5682), .ZN(n9121) );
  NAND2_X1 U5498 ( .A1(n8458), .A2(n8457), .ZN(n8456) );
  AND4_X1 U5499 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n8908)
         );
  INV_X1 U5500 ( .A(n8551), .ZN(n6878) );
  NAND2_X1 U5501 ( .A1(n4710), .A2(n5768), .ZN(n6043) );
  NAND2_X1 U5502 ( .A1(n8439), .A2(n5826), .ZN(n8474) );
  AND4_X1 U5503 ( .A1(n5690), .A2(n5689), .A3(n5688), .A4(n5687), .ZN(n8978)
         );
  NAND2_X1 U5504 ( .A1(n5853), .A2(n5852), .ZN(n9067) );
  AND4_X1 U5505 ( .A1(n5651), .A2(n5650), .A3(n5649), .A4(n5648), .ZN(n7600)
         );
  AOI21_X1 U5506 ( .B1(n4708), .B2(n4706), .A(n4705), .ZN(n4704) );
  INV_X1 U5507 ( .A(n4708), .ZN(n4707) );
  NAND2_X1 U5508 ( .A1(n8458), .A2(n4340), .ZN(n4692) );
  AOI21_X1 U5509 ( .B1(n4470), .B2(n4469), .A(n4717), .ZN(n8396) );
  OR2_X1 U5510 ( .A1(n5796), .A2(n5530), .ZN(n5533) );
  OR2_X1 U5511 ( .A1(n5574), .A2(n5529), .ZN(n5534) );
  NAND2_X1 U5512 ( .A1(n6811), .A2(n6812), .ZN(n6810) );
  NOR2_X1 U5513 ( .A1(n7120), .A2(n7119), .ZN(n7118) );
  AND2_X1 U5514 ( .A1(n6810), .A2(n4572), .ZN(n7120) );
  NAND2_X1 U5515 ( .A1(n6702), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4572) );
  NOR2_X1 U5516 ( .A1(n7106), .A2(n4368), .ZN(n7131) );
  INV_X1 U5517 ( .A(n4571), .ZN(n7129) );
  NOR2_X1 U5518 ( .A1(n7096), .A2(n7095), .ZN(n7094) );
  AND2_X1 U5519 ( .A1(n4571), .A2(n4570), .ZN(n7096) );
  NAND2_X1 U5520 ( .A1(n6688), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4570) );
  NOR2_X1 U5521 ( .A1(n7708), .A2(n4567), .ZN(n7712) );
  AND2_X1 U5522 ( .A1(n7715), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4567) );
  INV_X1 U5523 ( .A(n4566), .ZN(n8603) );
  XNOR2_X1 U5524 ( .A(n8631), .B(n9025), .ZN(n9027) );
  INV_X1 U5525 ( .A(n8639), .ZN(n9708) );
  OR2_X1 U5526 ( .A1(n9036), .A2(n8725), .ZN(n8699) );
  OAI21_X1 U5527 ( .B1(n4624), .B2(n4629), .A(n8187), .ZN(n8709) );
  NAND2_X1 U5528 ( .A1(n8729), .A2(n8728), .ZN(n8727) );
  NAND2_X1 U5529 ( .A1(n8737), .A2(n8697), .ZN(n8729) );
  AOI21_X1 U5530 ( .B1(n4397), .B2(n8986), .A(n4394), .ZN(n9045) );
  NAND2_X1 U5531 ( .A1(n4396), .A2(n4395), .ZN(n4394) );
  XNOR2_X1 U5532 ( .A(n4398), .B(n8724), .ZN(n4397) );
  NAND2_X1 U5533 ( .A1(n8726), .A2(n8965), .ZN(n4395) );
  NAND2_X1 U5534 ( .A1(n8775), .A2(n8217), .ZN(n8759) );
  NAND2_X1 U5535 ( .A1(n4539), .A2(n4544), .ZN(n8789) );
  NAND2_X1 U5536 ( .A1(n8814), .A2(n4545), .ZN(n4539) );
  AND2_X1 U5537 ( .A1(n4547), .A2(n4551), .ZN(n8801) );
  NAND2_X1 U5538 ( .A1(n8814), .A2(n8692), .ZN(n4547) );
  NAND2_X1 U5539 ( .A1(n5810), .A2(n5809), .ZN(n9083) );
  INV_X1 U5540 ( .A(n4563), .ZN(n8857) );
  NAND2_X1 U5541 ( .A1(n6750), .A2(n4534), .ZN(n4532) );
  NAND2_X1 U5542 ( .A1(n6750), .A2(n6749), .ZN(n6903) );
  OR2_X1 U5543 ( .A1(n5523), .A2(n4332), .ZN(n5561) );
  CLKBUF_X1 U5544 ( .A(n9022), .Z(n8995) );
  NAND2_X1 U5545 ( .A1(n8946), .A2(n6819), .ZN(n9008) );
  NAND2_X1 U5546 ( .A1(n5540), .A2(n4344), .ZN(n5555) );
  AND2_X1 U5547 ( .A1(n8946), .A2(n6832), .ZN(n8940) );
  NAND2_X1 U5548 ( .A1(n8194), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5522) );
  INV_X1 U5549 ( .A(n9008), .ZN(n8892) );
  INV_X1 U5550 ( .A(n8940), .ZN(n9024) );
  INV_X1 U5551 ( .A(n10017), .ZN(n10026) );
  AND2_X1 U5552 ( .A1(n6215), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9978) );
  MUX2_X1 U5553 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5446), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5448) );
  OAI21_X1 U5554 ( .B1(n5769), .B2(n4361), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4484) );
  INV_X1 U5555 ( .A(n4721), .ZN(n4718) );
  INV_X1 U5556 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5557 ( .A1(n9220), .A2(n4671), .ZN(n6604) );
  NOR2_X1 U5558 ( .A1(n8425), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U5559 ( .A1(n4664), .A2(n4659), .ZN(n4656) );
  AND2_X1 U5560 ( .A1(n8417), .A2(n9694), .ZN(n4664) );
  NAND2_X1 U5561 ( .A1(n5167), .A2(n5166), .ZN(n9630) );
  NAND2_X1 U5562 ( .A1(n8090), .A2(n8089), .ZN(n9205) );
  NOR2_X1 U5563 ( .A1(n9224), .A2(n4400), .ZN(n9225) );
  NAND2_X1 U5564 ( .A1(n5223), .A2(n5222), .ZN(n9606) );
  INV_X1 U5565 ( .A(n9224), .ZN(n9276) );
  AND2_X1 U5566 ( .A1(n6297), .A2(n6439), .ZN(n9694) );
  NAND4_X1 U5567 ( .A1(n5112), .A2(n5111), .A3(n5110), .A4(n5109), .ZN(n9284)
         );
  NAND4_X1 U5568 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n9289)
         );
  OR2_X1 U5569 ( .A1(n5275), .A2(n9838), .ZN(n5005) );
  NAND2_X1 U5570 ( .A1(n4960), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U5571 ( .A1(n4960), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4944) );
  AND2_X1 U5572 ( .A1(n7841), .A2(n7840), .ZN(n9566) );
  INV_X1 U5573 ( .A(n5385), .ZN(n5386) );
  AOI21_X1 U5574 ( .B1(n9281), .B2(n9875), .A(n5384), .ZN(n5385) );
  NAND2_X1 U5575 ( .A1(n4384), .A2(n7888), .ZN(n9337) );
  NAND2_X1 U5576 ( .A1(n9355), .A2(n8015), .ZN(n4384) );
  INV_X1 U5577 ( .A(n9376), .ZN(n5371) );
  NAND2_X1 U5578 ( .A1(n9434), .A2(n7979), .ZN(n9419) );
  NAND2_X1 U5579 ( .A1(n4420), .A2(n4425), .ZN(n9476) );
  NAND2_X1 U5580 ( .A1(n4438), .A2(n7930), .ZN(n9524) );
  NAND2_X1 U5581 ( .A1(n4447), .A2(n7927), .ZN(n7258) );
  OAI211_X1 U5582 ( .C1(n6039), .C2(n6180), .A(n5054), .B(n5053), .ZN(n6947)
         );
  NAND2_X1 U5583 ( .A1(n4411), .A2(n5042), .ZN(n6942) );
  OAI21_X1 U5584 ( .B1(n6556), .B2(n5357), .A(n5356), .ZN(n6726) );
  OAI21_X1 U5585 ( .B1(n6039), .B2(n4950), .A(n4949), .ZN(n9860) );
  NAND2_X1 U5586 ( .A1(n6039), .A2(n6069), .ZN(n4949) );
  AOI21_X1 U5587 ( .B1(n9703), .B2(n9914), .A(n9702), .ZN(n9706) );
  OAI22_X1 U5588 ( .A1(n9899), .A2(n9946), .B1(n9898), .B2(n4445), .ZN(n9901)
         );
  INV_X1 U5589 ( .A(n6394), .ZN(n4445) );
  XNOR2_X1 U5590 ( .A(n5320), .B(n5319), .ZN(n7768) );
  OAI21_X1 U5591 ( .B1(n4890), .B2(n4328), .A(n4581), .ZN(n5247) );
  NAND2_X1 U5592 ( .A1(n5211), .A2(n5336), .ZN(n9850) );
  MUX2_X1 U5593 ( .A(n5208), .B(P1_IR_REG_31__SCAN_IN), .S(n5209), .Z(n5211)
         );
  NAND2_X1 U5594 ( .A1(n6622), .A2(n5640), .ZN(n6918) );
  NAND2_X1 U5595 ( .A1(n6008), .A2(n6007), .ZN(n6015) );
  OAI21_X1 U5596 ( .B1(n4632), .B2(n4631), .A(n4630), .ZN(P2_U3244) );
  NAND2_X1 U5597 ( .A1(n4330), .A2(n7028), .ZN(n4631) );
  XNOR2_X1 U5598 ( .A(n8211), .B(n8888), .ZN(n4632) );
  AOI21_X1 U5599 ( .B1(n8397), .B2(n7028), .A(n4331), .ZN(n4630) );
  OAI211_X1 U5600 ( .C1(n4661), .C2(n4657), .A(n4665), .B(n4655), .ZN(P1_U3218) );
  INV_X1 U5601 ( .A(n4664), .ZN(n4657) );
  AND2_X1 U5602 ( .A1(n8424), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U5603 ( .A1(n4661), .A2(n4658), .ZN(n4665) );
  OAI21_X1 U5604 ( .B1(n8081), .B2(n8080), .A(n8079), .ZN(n8087) );
  NOR2_X1 U5605 ( .A1(n9580), .A2(n9856), .ZN(n9372) );
  NOR2_X1 U5606 ( .A1(n9584), .A2(n9856), .ZN(n7763) );
  OAI22_X1 U5607 ( .A1(n9539), .A2(n4400), .B1(n6563), .B2(n9880), .ZN(n6564)
         );
  NAND2_X1 U5608 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NOR2_X1 U5609 ( .A1(n8179), .A2(n8654), .ZN(n4313) );
  AND2_X1 U5610 ( .A1(n8262), .A2(n4460), .ZN(n4314) );
  OR2_X1 U5611 ( .A1(n7830), .A2(n8066), .ZN(n4315) );
  INV_X2 U5612 ( .A(n4969), .ZN(n5236) );
  INV_X1 U5613 ( .A(n8788), .ZN(n4541) );
  INV_X1 U5614 ( .A(n4634), .ZN(n4633) );
  XNOR2_X1 U5615 ( .A(n9042), .B(n8545), .ZN(n8728) );
  AND2_X1 U5616 ( .A1(n9344), .A2(n9360), .ZN(n4316) );
  AND2_X1 U5617 ( .A1(n4765), .A2(n4673), .ZN(n4317) );
  INV_X1 U5618 ( .A(n8331), .ZN(n4455) );
  AND2_X1 U5619 ( .A1(n4734), .A2(n10004), .ZN(n4318) );
  AND4_X1 U5620 ( .A1(n5338), .A2(n4428), .A3(n5178), .A4(n4427), .ZN(n4319)
         );
  INV_X1 U5621 ( .A(n8813), .ZN(n4635) );
  OR3_X1 U5622 ( .A1(n5769), .A2(P2_IR_REG_18__SCAN_IN), .A3(
        P2_IR_REG_17__SCAN_IN), .ZN(n4320) );
  AND2_X1 U5623 ( .A1(n6026), .A2(n5390), .ZN(n4321) );
  NAND2_X1 U5624 ( .A1(n5553), .A2(n5429), .ZN(n5580) );
  AND2_X1 U5625 ( .A1(n4736), .A2(n4735), .ZN(n4322) );
  AND2_X1 U5626 ( .A1(n5475), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4323) );
  AND2_X1 U5627 ( .A1(n8921), .A2(n8279), .ZN(n8666) );
  AND2_X1 U5628 ( .A1(n4747), .A2(n4449), .ZN(n4324) );
  AND2_X1 U5629 ( .A1(n4316), .A2(n4516), .ZN(n4325) );
  AND2_X1 U5630 ( .A1(n5475), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4326) );
  AND2_X1 U5631 ( .A1(n4501), .A2(n8098), .ZN(n4327) );
  OR2_X1 U5632 ( .A1(n5239), .A2(n4583), .ZN(n4328) );
  XNOR2_X1 U5633 ( .A(n4484), .B(n5437), .ZN(n8193) );
  AND2_X1 U5634 ( .A1(n5055), .A2(n4515), .ZN(n4329) );
  NAND2_X1 U5635 ( .A1(n4684), .A2(n4682), .ZN(n8090) );
  AND2_X1 U5636 ( .A1(n5882), .A2(n5881), .ZN(n8780) );
  INV_X1 U5637 ( .A(n8780), .ZN(n4549) );
  NAND2_X1 U5638 ( .A1(n8213), .A2(n8212), .ZN(n4330) );
  NOR2_X1 U5639 ( .A1(n8401), .A2(n8400), .ZN(n4331) );
  NAND2_X2 U5640 ( .A1(n4556), .A2(n5454), .ZN(n5564) );
  XOR2_X1 U5641 ( .A(n4990), .B(n4979), .Z(n4332) );
  INV_X1 U5642 ( .A(n8138), .ZN(n4670) );
  AND2_X1 U5643 ( .A1(n4786), .A2(n4785), .ZN(n4333) );
  OR2_X1 U5644 ( .A1(n5398), .A2(n4680), .ZN(n5394) );
  AND2_X1 U5645 ( .A1(n4692), .A2(n4696), .ZN(n4334) );
  OR2_X1 U5646 ( .A1(n5398), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4335) );
  NAND2_X2 U5647 ( .A1(n4556), .A2(n9163), .ZN(n5796) );
  OR2_X1 U5648 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4336) );
  AND2_X1 U5649 ( .A1(n4698), .A2(n5572), .ZN(n4337) );
  NOR2_X1 U5650 ( .A1(n9597), .A2(n9435), .ZN(n4338) );
  INV_X1 U5651 ( .A(n6930), .ZN(n6891) );
  OAI211_X1 U5652 ( .C1(n6039), .C2(n6274), .A(n5021), .B(n5020), .ZN(n6930)
         );
  OR2_X1 U5653 ( .A1(n5398), .A2(n4677), .ZN(n4339) );
  AND2_X1 U5654 ( .A1(n4697), .A2(n8457), .ZN(n4340) );
  XNOR2_X1 U5655 ( .A(n4860), .B(SI_14_), .ZN(n5130) );
  NAND2_X1 U5656 ( .A1(n5342), .A2(n6029), .ZN(n6284) );
  OR2_X1 U5657 ( .A1(n8139), .A2(n8138), .ZN(n4341) );
  AND2_X1 U5658 ( .A1(n4724), .A2(n5473), .ZN(n4342) );
  AND4_X1 U5659 ( .A1(n4430), .A2(n4429), .A3(n5209), .A4(n5160), .ZN(n4343)
         );
  NAND2_X1 U5660 ( .A1(n8334), .A2(n8331), .ZN(n8742) );
  NAND2_X1 U5661 ( .A1(n5327), .A2(n5326), .ZN(n8029) );
  INV_X1 U5662 ( .A(n8694), .ZN(n4546) );
  AND2_X1 U5663 ( .A1(n7852), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4344) );
  AND2_X1 U5664 ( .A1(n8383), .A2(n4628), .ZN(n4345) );
  NOR2_X1 U5665 ( .A1(n8162), .A2(n4663), .ZN(n4346) );
  NAND2_X1 U5666 ( .A1(n4766), .A2(n4765), .ZN(n5006) );
  AND2_X1 U5667 ( .A1(n4358), .A2(n4636), .ZN(n4347) );
  NAND2_X1 U5668 ( .A1(n5906), .A2(n5905), .ZN(n9048) );
  AND2_X1 U5669 ( .A1(n5842), .A2(n5841), .ZN(n8819) );
  INV_X1 U5670 ( .A(n8819), .ZN(n9072) );
  NAND2_X1 U5671 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4348) );
  NAND2_X1 U5672 ( .A1(n9361), .A2(n8009), .ZN(n4349) );
  AND2_X1 U5673 ( .A1(n8102), .A2(n8098), .ZN(n4350) );
  AND2_X1 U5674 ( .A1(n9284), .A2(n8412), .ZN(n4351) );
  AND2_X1 U5675 ( .A1(n8698), .A2(n8545), .ZN(n4352) );
  AND4_X1 U5676 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n8977)
         );
  INV_X1 U5677 ( .A(n8977), .ZN(n4646) );
  NAND2_X1 U5678 ( .A1(n8381), .A2(n8327), .ZN(n4353) );
  NAND2_X1 U5679 ( .A1(n4839), .A2(n4838), .ZN(n5051) );
  OR2_X1 U5680 ( .A1(n9036), .A2(n8188), .ZN(n8343) );
  AND2_X1 U5681 ( .A1(n4595), .A2(n4492), .ZN(n4354) );
  AND2_X1 U5682 ( .A1(n4834), .A2(SI_7_), .ZN(n4355) );
  NAND2_X1 U5683 ( .A1(n4414), .A2(n4415), .ZN(n5552) );
  NAND2_X1 U5684 ( .A1(n9840), .A2(n5354), .ZN(n4356) );
  NAND2_X1 U5685 ( .A1(n8551), .A2(n4310), .ZN(n4357) );
  INV_X1 U5686 ( .A(n5102), .ZN(n4623) );
  NAND2_X1 U5687 ( .A1(n4855), .A2(n4854), .ZN(n5102) );
  OR2_X1 U5688 ( .A1(n8846), .A2(n4638), .ZN(n4358) );
  INV_X1 U5689 ( .A(n4452), .ZN(n4451) );
  NAND2_X1 U5690 ( .A1(n8333), .A2(n4453), .ZN(n4452) );
  OR2_X1 U5691 ( .A1(n7990), .A2(n7981), .ZN(n4359) );
  AND2_X1 U5692 ( .A1(n8020), .A2(n8019), .ZN(n8067) );
  OR2_X1 U5693 ( .A1(n5361), .A2(n4446), .ZN(n4360) );
  OR2_X1 U5694 ( .A1(n4718), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4361) );
  INV_X1 U5695 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5465) );
  AND2_X1 U5696 ( .A1(n4859), .A2(n4858), .ZN(n5115) );
  OR2_X1 U5697 ( .A1(n4546), .A2(n4548), .ZN(n4362) );
  NAND2_X1 U5698 ( .A1(n4766), .A2(n4317), .ZN(n4674) );
  AND2_X1 U5699 ( .A1(n6906), .A2(n8242), .ZN(n8243) );
  INV_X1 U5700 ( .A(n8243), .ZN(n4404) );
  NAND2_X1 U5701 ( .A1(n9597), .A2(n9435), .ZN(n4363) );
  AND2_X1 U5702 ( .A1(n8283), .A2(n8960), .ZN(n4364) );
  INV_X1 U5703 ( .A(n4503), .ZN(n4502) );
  OAI21_X1 U5704 ( .B1(n4682), .B2(n4504), .A(n9206), .ZN(n4503) );
  AND2_X1 U5705 ( .A1(n4325), .A2(n8034), .ZN(n4365) );
  AND2_X1 U5706 ( .A1(n4648), .A2(n4653), .ZN(n4366) );
  INV_X1 U5707 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4428) );
  INV_X1 U5708 ( .A(n8371), .ZN(n4408) );
  NAND2_X1 U5709 ( .A1(n4647), .A2(n4648), .ZN(n7206) );
  NAND2_X1 U5710 ( .A1(n4710), .A2(n4708), .ZN(n6040) );
  NAND2_X1 U5711 ( .A1(n4930), .A2(n4929), .ZN(n9330) );
  INV_X1 U5712 ( .A(n9330), .ZN(n4516) );
  INV_X1 U5713 ( .A(n6837), .ZN(n9991) );
  AND3_X1 U5714 ( .A1(n5561), .A2(n5560), .A3(n5559), .ZN(n6837) );
  OR2_X1 U5715 ( .A1(n5769), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4367) );
  INV_X1 U5716 ( .A(n9267), .ZN(n4662) );
  NAND2_X1 U5717 ( .A1(n4419), .A2(n4417), .ZN(n9468) );
  AND2_X1 U5718 ( .A1(n6689), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4368) );
  INV_X1 U5719 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5720 ( .A1(n7770), .A2(n7769), .ZN(n9036) );
  INV_X1 U5721 ( .A(n9036), .ZN(n4737) );
  NAND2_X1 U5722 ( .A1(n5613), .A2(n5612), .ZN(n7285) );
  NAND2_X1 U5723 ( .A1(n5286), .A2(n5285), .ZN(n5293) );
  INV_X1 U5724 ( .A(n5293), .ZN(n4614) );
  NAND2_X1 U5725 ( .A1(n9204), .A2(n4350), .ZN(n9254) );
  NAND2_X1 U5726 ( .A1(n4684), .A2(n4685), .ZN(n7740) );
  NAND2_X1 U5727 ( .A1(n8191), .A2(n8190), .ZN(n9029) );
  INV_X1 U5728 ( .A(n9029), .ZN(n4735) );
  NAND2_X1 U5729 ( .A1(n5242), .A2(n5241), .ZN(n9597) );
  NAND2_X1 U5730 ( .A1(n5792), .A2(n5791), .ZN(n9087) );
  NOR3_X1 U5731 ( .A1(n4754), .A2(n9062), .A3(n4742), .ZN(n4739) );
  NAND2_X1 U5732 ( .A1(n5774), .A2(n5773), .ZN(n9093) );
  AND2_X1 U5733 ( .A1(n4527), .A2(n4526), .ZN(n4369) );
  NOR2_X1 U5734 ( .A1(n9507), .A2(n4518), .ZN(n4521) );
  NAND2_X1 U5735 ( .A1(n5701), .A2(n5700), .ZN(n9116) );
  OR2_X1 U5736 ( .A1(n8162), .A2(n4662), .ZN(n4660) );
  INV_X1 U5737 ( .A(n4660), .ZN(n4659) );
  AND3_X1 U5738 ( .A1(n8264), .A2(n8267), .A3(n8268), .ZN(n4370) );
  INV_X1 U5739 ( .A(n4517), .ZN(n9463) );
  NOR3_X1 U5740 ( .A1(n9507), .A2(n9611), .A3(n4520), .ZN(n4517) );
  INV_X1 U5741 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U5742 ( .A1(n9623), .A2(n9478), .ZN(n4371) );
  INV_X1 U5743 ( .A(n4740), .ZN(n8802) );
  NOR2_X1 U5744 ( .A1(n4754), .A2(n4742), .ZN(n4740) );
  INV_X1 U5745 ( .A(n4513), .ZN(n4512) );
  NAND2_X1 U5746 ( .A1(n4329), .A2(n4514), .ZN(n4513) );
  NAND2_X1 U5747 ( .A1(n5867), .A2(n5866), .ZN(n9062) );
  NOR2_X1 U5748 ( .A1(n9507), .A2(n4520), .ZN(n9462) );
  AND2_X1 U5749 ( .A1(n9062), .A2(n4549), .ZN(n4372) );
  NAND2_X1 U5750 ( .A1(n5197), .A2(n5196), .ZN(n9618) );
  AND2_X1 U5751 ( .A1(n8963), .A2(n8975), .ZN(n4373) );
  AND2_X1 U5752 ( .A1(n4318), .A2(n8259), .ZN(n4374) );
  INV_X1 U5753 ( .A(n4551), .ZN(n4548) );
  NAND2_X1 U5754 ( .A1(n9072), .A2(n8838), .ZN(n4551) );
  NAND2_X1 U5755 ( .A1(n8305), .A2(n8807), .ZN(n4375) );
  INV_X1 U5756 ( .A(n4713), .ZN(n8361) );
  AOI21_X1 U5757 ( .B1(n5464), .B2(n4715), .A(n4714), .ZN(n4713) );
  AND2_X1 U5758 ( .A1(n9220), .A2(n6587), .ZN(n6768) );
  NAND2_X1 U5759 ( .A1(n6825), .A2(n8219), .ZN(n6755) );
  NAND2_X1 U5760 ( .A1(n6904), .A2(n10001), .ZN(n4376) );
  NAND2_X1 U5761 ( .A1(n5389), .A2(n4512), .ZN(n4377) );
  NAND2_X1 U5762 ( .A1(n4532), .A2(n6753), .ZN(n6875) );
  NAND2_X1 U5763 ( .A1(n4411), .A2(n4409), .ZN(n6940) );
  OAI21_X1 U5764 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(n9219) );
  NAND2_X1 U5765 ( .A1(n4774), .A2(n4773), .ZN(n5398) );
  NAND2_X1 U5766 ( .A1(n5753), .A2(n5442), .ZN(n5944) );
  NAND2_X1 U5767 ( .A1(n5753), .A2(n4722), .ZN(n4378) );
  NAND2_X1 U5768 ( .A1(n7572), .A2(n4730), .ZN(n4733) );
  INV_X1 U5769 ( .A(n4727), .ZN(n8941) );
  NOR2_X1 U5770 ( .A1(n8953), .A2(n9106), .ZN(n4727) );
  INV_X1 U5771 ( .A(n5976), .ZN(n5965) );
  AND2_X1 U5772 ( .A1(n4529), .A2(n4528), .ZN(n4379) );
  OAI21_X1 U5773 ( .B1(n6531), .B2(n4699), .A(n4337), .ZN(n6502) );
  NAND4_X1 U5774 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n9874)
         );
  NAND2_X1 U5775 ( .A1(n5758), .A2(n5757), .ZN(n9097) );
  INV_X1 U5776 ( .A(n9097), .ZN(n4726) );
  NAND2_X1 U5777 ( .A1(n5078), .A2(n5077), .ZN(n9672) );
  INV_X1 U5778 ( .A(n9672), .ZN(n4514) );
  AND2_X1 U5779 ( .A1(n8593), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4380) );
  XNOR2_X1 U5780 ( .A(n5341), .B(n4428), .ZN(n6029) );
  NOR2_X1 U5781 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7534) );
  INV_X1 U5782 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5783 ( .A1(n4591), .A2(n8032), .ZN(n4590) );
  AOI21_X1 U5784 ( .B1(n5387), .B2(n9871), .A(n5386), .ZN(n6026) );
  AOI21_X1 U5785 ( .B1(n9371), .B2(n9871), .A(n9370), .ZN(n9580) );
  AOI21_X1 U5786 ( .B1(n7762), .B2(n9871), .A(n7761), .ZN(n9584) );
  NAND2_X2 U5787 ( .A1(n6481), .A2(n8212), .ZN(n8986) );
  NAND2_X1 U5788 ( .A1(n4713), .A2(n5482), .ZN(n8212) );
  NOR2_X4 U5789 ( .A1(n5976), .A2(n4717), .ZN(n9993) );
  INV_X1 U5790 ( .A(n8361), .ZN(n4717) );
  NAND4_X1 U5791 ( .A1(n4771), .A2(n4766), .A3(n4317), .A4(n4772), .ZN(n5132)
         );
  NAND4_X1 U5792 ( .A1(n4771), .A2(n4766), .A3(n4317), .A4(n4381), .ZN(n5163)
         );
  XNOR2_X2 U5793 ( .A(n4382), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U5794 ( .A1(n9253), .A2(n9257), .ZN(n9176) );
  OAI21_X2 U5795 ( .B1(n4684), .B2(n4504), .A(n4502), .ZN(n9204) );
  NOR2_X1 U5796 ( .A1(n9242), .A2(n9244), .ZN(n9246) );
  AND2_X2 U5797 ( .A1(n8131), .A2(n4498), .ZN(n9242) );
  NAND2_X1 U5798 ( .A1(n6039), .A2(n4326), .ZN(n4936) );
  NOR2_X1 U5799 ( .A1(n9319), .A2(n9323), .ZN(n9320) );
  NAND2_X2 U5800 ( .A1(n4392), .A2(n5191), .ZN(n9487) );
  INV_X2 U5801 ( .A(n5807), .ZN(n8194) );
  NAND2_X2 U5802 ( .A1(n5540), .A2(n7852), .ZN(n5807) );
  NAND2_X2 U5803 ( .A1(n5984), .A2(n8398), .ZN(n5540) );
  NAND3_X1 U5804 ( .A1(n9839), .A2(n6891), .A3(n4400), .ZN(n4525) );
  NAND3_X1 U5805 ( .A1(n4401), .A2(n6758), .A3(n4403), .ZN(n6968) );
  NAND2_X1 U5806 ( .A1(n4402), .A2(n6825), .ZN(n4401) );
  NAND2_X1 U5807 ( .A1(n6720), .A2(n7869), .ZN(n4411) );
  XNOR2_X1 U5808 ( .A(n5335), .B(n7891), .ZN(n6034) );
  OR2_X1 U5809 ( .A1(n8229), .A2(n8362), .ZN(n6654) );
  NAND2_X1 U5810 ( .A1(n8230), .A2(n8232), .ZN(n8362) );
  AND2_X2 U5811 ( .A1(n5609), .A2(n4751), .ZN(n5753) );
  NAND3_X1 U5812 ( .A1(n4414), .A2(n4413), .A3(n4412), .ZN(n5476) );
  NOR2_X2 U5813 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4414) );
  NAND2_X1 U5814 ( .A1(n9515), .A2(n4421), .ZN(n4419) );
  OAI21_X1 U5815 ( .B1(n9515), .B2(n5367), .A(n7965), .ZN(n9497) );
  OAI21_X1 U5816 ( .B1(n5369), .B2(n4435), .A(n4433), .ZN(n9399) );
  NAND2_X1 U5817 ( .A1(n4432), .A2(n4431), .ZN(n5370) );
  NAND2_X1 U5818 ( .A1(n5369), .A2(n4433), .ZN(n4432) );
  INV_X1 U5819 ( .A(n7589), .ZN(n5363) );
  OAI211_X1 U5820 ( .C1(n6556), .C2(n5357), .A(n5358), .B(n5356), .ZN(n4448)
         );
  INV_X1 U5821 ( .A(n8258), .ZN(n4457) );
  AOI21_X1 U5822 ( .B1(n4457), .B2(n4459), .A(n4458), .ZN(n8273) );
  NAND2_X1 U5823 ( .A1(n4463), .A2(n4462), .ZN(n8318) );
  OAI21_X1 U5824 ( .B1(n4465), .B2(n4375), .A(n4464), .ZN(n4463) );
  INV_X1 U5825 ( .A(n8312), .ZN(n4468) );
  NAND2_X1 U5826 ( .A1(n4477), .A2(n4476), .ZN(n8294) );
  NAND2_X1 U5827 ( .A1(n4478), .A2(n8287), .ZN(n4477) );
  NAND3_X1 U5828 ( .A1(n4482), .A2(n4479), .A3(n4373), .ZN(n4478) );
  NAND2_X1 U5829 ( .A1(n4481), .A2(n4480), .ZN(n4479) );
  NOR2_X1 U5830 ( .A1(n8278), .A2(n8354), .ZN(n4480) );
  NAND2_X1 U5831 ( .A1(n8280), .A2(n8279), .ZN(n4481) );
  NAND2_X1 U5832 ( .A1(n4483), .A2(n8354), .ZN(n4482) );
  NAND2_X1 U5833 ( .A1(n8275), .A2(n8921), .ZN(n4483) );
  NAND2_X1 U5834 ( .A1(n4485), .A2(n4487), .ZN(n5074) );
  NAND3_X1 U5835 ( .A1(n4596), .A2(n4595), .A3(n4486), .ZN(n4485) );
  NAND2_X1 U5836 ( .A1(n4596), .A2(n4595), .ZN(n5052) );
  INV_X1 U5837 ( .A(n5051), .ZN(n4492) );
  INV_X1 U5838 ( .A(n4684), .ZN(n4500) );
  OAI21_X1 U5839 ( .B1(n4500), .B2(n4503), .A(n4327), .ZN(n8105) );
  NAND2_X1 U5840 ( .A1(n6111), .A2(n7859), .ZN(n4507) );
  NAND3_X1 U5841 ( .A1(n4647), .A2(n4366), .A3(n4654), .ZN(n4652) );
  NAND2_X1 U5842 ( .A1(n8105), .A2(n8104), .ZN(n9257) );
  NAND2_X1 U5843 ( .A1(n9229), .A2(n9233), .ZN(n9186) );
  NAND2_X1 U5844 ( .A1(n5074), .A2(n5075), .ZN(n4848) );
  NAND2_X1 U5845 ( .A1(n4652), .A2(n4650), .ZN(n7545) );
  NAND2_X1 U5846 ( .A1(n4808), .A2(n4807), .ZN(n4954) );
  NAND2_X1 U5847 ( .A1(n9350), .A2(n8020), .ZN(n9324) );
  NAND2_X1 U5848 ( .A1(n5368), .A2(n7970), .ZN(n9453) );
  NAND2_X1 U5849 ( .A1(n4666), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5850 ( .A1(n4356), .A2(n5355), .ZN(n5356) );
  NAND2_X1 U5851 ( .A1(n5389), .A2(n4511), .ZN(n7583) );
  NAND2_X1 U5852 ( .A1(n9356), .A2(n4325), .ZN(n9329) );
  AND2_X1 U5853 ( .A1(n9356), .A2(n9360), .ZN(n9338) );
  INV_X1 U5854 ( .A(n4521), .ZN(n9449) );
  NAND2_X1 U5855 ( .A1(n6750), .A2(n4531), .ZN(n4528) );
  NAND3_X1 U5856 ( .A1(n4529), .A2(n8369), .A3(n4528), .ZN(n6962) );
  NAND2_X1 U5857 ( .A1(n8814), .A2(n4540), .ZN(n4538) );
  NAND2_X1 U5858 ( .A1(n4536), .A2(n4540), .ZN(n8787) );
  OR2_X1 U5859 ( .A1(n8814), .A2(n4543), .ZN(n4536) );
  NAND2_X1 U5860 ( .A1(n8738), .A2(n4553), .ZN(n4552) );
  NAND2_X1 U5861 ( .A1(n5454), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4557) );
  OR2_X1 U5862 ( .A1(n5454), .A2(n6993), .ZN(n4558) );
  INV_X1 U5863 ( .A(n5454), .ZN(n9163) );
  INV_X1 U5864 ( .A(n4560), .ZN(n4559) );
  AND2_X1 U5865 ( .A1(n4342), .A2(n5753), .ZN(n5469) );
  NAND2_X1 U5866 ( .A1(n5471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U5867 ( .A1(n5283), .A2(n5282), .ZN(n4577) );
  INV_X1 U5868 ( .A(n5270), .ZN(n4578) );
  NAND2_X1 U5869 ( .A1(n4890), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U5870 ( .A1(n4890), .A2(n4889), .ZN(n5231) );
  NAND3_X1 U5871 ( .A1(n4590), .A2(n4588), .A3(n4587), .ZN(n8046) );
  NAND3_X1 U5872 ( .A1(n8027), .A2(n8037), .A3(n7842), .ZN(n4593) );
  NAND2_X1 U5873 ( .A1(n4594), .A2(SI_1_), .ZN(n4807) );
  XNOR2_X2 U5874 ( .A(n4594), .B(n4806), .ZN(n4934) );
  NAND2_X1 U5875 ( .A1(n5019), .A2(n5018), .ZN(n4599) );
  NAND2_X1 U5876 ( .A1(n5019), .A2(n4597), .ZN(n4596) );
  NAND2_X1 U5877 ( .A1(n4848), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U5878 ( .A1(n4600), .A2(n4604), .ZN(n5143) );
  NAND3_X1 U5879 ( .A1(n4606), .A2(n4608), .A3(n5130), .ZN(n4605) );
  NAND3_X1 U5880 ( .A1(n7994), .A2(n9362), .A3(n8032), .ZN(n4613) );
  OR2_X1 U5881 ( .A1(n4815), .A2(n4993), .ZN(n4817) );
  INV_X1 U5882 ( .A(n8743), .ZN(n4624) );
  NAND2_X1 U5883 ( .A1(n8846), .A2(n8847), .ZN(n8834) );
  INV_X1 U5884 ( .A(n8181), .ZN(n4638) );
  NAND2_X1 U5885 ( .A1(n4641), .A2(n4639), .ZN(n8185) );
  INV_X1 U5886 ( .A(n4640), .ZN(n4639) );
  OAI21_X1 U5887 ( .B1(n8184), .B2(n4643), .A(n8381), .ZN(n4640) );
  NAND2_X1 U5888 ( .A1(n7065), .A2(n4649), .ZN(n4647) );
  NAND2_X1 U5889 ( .A1(n4654), .A2(n4651), .ZN(n4650) );
  NAND2_X1 U5890 ( .A1(n4661), .A2(n4660), .ZN(n8426) );
  AOI21_X1 U5891 ( .B1(n9266), .B2(n9268), .A(n9267), .ZN(n8163) );
  INV_X1 U5892 ( .A(n9268), .ZN(n4663) );
  AND3_X2 U5893 ( .A1(n9167), .A2(n4667), .A3(n4668), .ZN(n9211) );
  NAND2_X1 U5894 ( .A1(n9167), .A2(n4668), .ZN(n9212) );
  INV_X1 U5895 ( .A(n9213), .ZN(n4667) );
  INV_X1 U5896 ( .A(n4674), .ZN(n5008) );
  AND2_X1 U5897 ( .A1(n5890), .A2(n4758), .ZN(n4687) );
  NAND2_X2 U5898 ( .A1(n5891), .A2(n4687), .ZN(n8458) );
  NAND2_X1 U5899 ( .A1(n6524), .A2(n4702), .ZN(n4698) );
  NAND2_X1 U5900 ( .A1(n6524), .A2(n4700), .ZN(n4699) );
  INV_X1 U5901 ( .A(n6530), .ZN(n4700) );
  OAI21_X1 U5902 ( .B1(n8466), .B2(n4707), .A(n4704), .ZN(n5806) );
  NAND2_X1 U5903 ( .A1(n6622), .A2(n4711), .ZN(n6916) );
  NAND2_X1 U5904 ( .A1(n8439), .A2(n4712), .ZN(n8445) );
  NAND3_X4 U5905 ( .A1(n4716), .A2(n8388), .A3(n8361), .ZN(n8213) );
  INV_X1 U5906 ( .A(n4733), .ZN(n9002) );
  NAND2_X1 U5907 ( .A1(n8762), .A2(n8630), .ZN(n8747) );
  INV_X1 U5908 ( .A(n4739), .ZN(n8790) );
  NOR2_X1 U5909 ( .A1(n6026), .A2(n9856), .ZN(n6036) );
  NAND4_X1 U5910 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n8557)
         );
  NAND2_X1 U5911 ( .A1(n6893), .A2(n6723), .ZN(n6943) );
  NAND2_X1 U5912 ( .A1(n5999), .A2(n5998), .ZN(P2_U3216) );
  INV_X1 U5913 ( .A(n6943), .ZN(n5389) );
  OAI21_X1 U5914 ( .B1(n6034), .B2(n9855), .A(n6033), .ZN(n6035) );
  CLKBUF_X1 U5915 ( .A(n6048), .Z(n6058) );
  NOR2_X1 U5916 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4764) );
  NAND4_X1 U5917 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), .ZN(n6292)
         );
  AND2_X1 U5918 ( .A1(n6292), .A2(n8411), .ZN(n6290) );
  XNOR2_X1 U5919 ( .A(n5947), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U5920 ( .A1(n5967), .A2(n8623), .ZN(n6481) );
  NAND2_X1 U5921 ( .A1(n5472), .A2(n5471), .ZN(n5984) );
  AOI21_X1 U5922 ( .B1(n9913), .B2(n8029), .A(n6028), .ZN(n5390) );
  AOI21_X1 U5923 ( .B1(n6028), .B2(n9535), .A(n6032), .ZN(n6033) );
  INV_X1 U5924 ( .A(n6472), .ZN(n6483) );
  NAND2_X1 U5925 ( .A1(n8987), .A2(n8959), .ZN(n8953) );
  NAND2_X1 U5926 ( .A1(n6477), .A2(n9979), .ZN(n7023) );
  INV_X1 U5927 ( .A(n6823), .ZN(n6656) );
  AND2_X1 U5928 ( .A1(n5887), .A2(n5886), .ZN(n6002) );
  AND2_X1 U5929 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  NAND2_X1 U5930 ( .A1(n5454), .A2(n7751), .ZN(n5546) );
  NOR2_X1 U5931 ( .A1(n9606), .A2(n9470), .ZN(n4744) );
  INV_X1 U5932 ( .A(n6291), .ZN(n7186) );
  OR2_X1 U5933 ( .A1(n9952), .A2(n6022), .ZN(n4745) );
  INV_X1 U5934 ( .A(n7874), .ZN(n5085) );
  INV_X1 U5935 ( .A(n8742), .ZN(n8186) );
  AND2_X1 U5936 ( .A1(n6429), .A2(n6401), .ZN(n4746) );
  AND2_X1 U5937 ( .A1(n8724), .A2(n8336), .ZN(n4747) );
  OR2_X1 U5938 ( .A1(n8833), .A2(n8690), .ZN(n4748) );
  OR2_X1 U5939 ( .A1(n8689), .A2(n8688), .ZN(n4749) );
  OR2_X1 U5940 ( .A1(n8777), .A2(n8346), .ZN(n4750) );
  AND4_X1 U5941 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n4751)
         );
  INV_X1 U5942 ( .A(n9042), .ZN(n8698) );
  AND2_X1 U5943 ( .A1(n9323), .A2(n8021), .ZN(n4752) );
  NOR2_X1 U5944 ( .A1(n9611), .A2(n9479), .ZN(n4755) );
  INV_X1 U5945 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4826) );
  AND3_X1 U5946 ( .A1(n5494), .A2(n5493), .A3(n5492), .ZN(n4757) );
  AND2_X1 U5947 ( .A1(n5930), .A2(n5929), .ZN(n8545) );
  OR2_X1 U5948 ( .A1(n6003), .A2(n6005), .ZN(n4758) );
  AND2_X1 U5949 ( .A1(n5915), .A2(n5914), .ZN(n8546) );
  NAND2_X1 U5950 ( .A1(n8668), .A2(n8667), .ZN(n4759) );
  AND2_X1 U5951 ( .A1(n9827), .A2(n9286), .ZN(n4761) );
  AND2_X1 U5952 ( .A1(n9591), .A2(n9421), .ZN(n4762) );
  NOR2_X1 U5953 ( .A1(n5268), .A2(n9390), .ZN(n4763) );
  AND2_X1 U5954 ( .A1(n8323), .A2(n4750), .ZN(n8324) );
  NAND2_X1 U5955 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  NAND2_X1 U5956 ( .A1(n8335), .A2(n8354), .ZN(n8336) );
  NOR4_X1 U5957 ( .A1(n8386), .A2(n8385), .A3(n8700), .A4(n8384), .ZN(n8387)
         );
  INV_X1 U5958 ( .A(n7796), .ZN(n5362) );
  INV_X1 U5959 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4772) );
  INV_X1 U5960 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5461) );
  INV_X1 U5961 ( .A(n7186), .ZN(n8406) );
  NOR2_X1 U5962 ( .A1(n4998), .A2(n7864), .ZN(n4999) );
  INV_X1 U5963 ( .A(n5721), .ZN(n5720) );
  NAND2_X1 U5964 ( .A1(n6481), .A2(n5976), .ZN(n8392) );
  NAND2_X1 U5965 ( .A1(n8551), .A2(n8213), .ZN(n5501) );
  INV_X1 U5966 ( .A(n5875), .ZN(n5870) );
  OR2_X1 U5967 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  INV_X1 U5968 ( .A(n5628), .ZN(n5626) );
  INV_X1 U5969 ( .A(n7186), .ZN(n8155) );
  AND2_X1 U5970 ( .A1(n9280), .A2(n9310), .ZN(n5384) );
  AND2_X1 U5971 ( .A1(n5360), .A2(n7932), .ZN(n7952) );
  INV_X1 U5972 ( .A(n9846), .ZN(n5026) );
  AND2_X1 U5973 ( .A1(n7904), .A2(n7905), .ZN(n9842) );
  XNOR2_X1 U5974 ( .A(n9893), .B(n9291), .ZN(n9865) );
  INV_X1 U5975 ( .A(n5491), .ZN(n5451) );
  NAND2_X1 U5976 ( .A1(n5720), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5742) );
  AND2_X1 U5977 ( .A1(n7766), .A2(n5935), .ZN(n5973) );
  OR2_X1 U5978 ( .A1(n5685), .A2(n7237), .ZN(n5703) );
  OR2_X1 U5979 ( .A1(n5703), .A2(n6743), .ZN(n5721) );
  NAND2_X1 U5980 ( .A1(n6483), .A2(n8213), .ZN(n5527) );
  NAND2_X1 U5981 ( .A1(n5870), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5895) );
  OR2_X1 U5982 ( .A1(n5600), .A2(n7434), .ZN(n5628) );
  NAND2_X1 U5983 ( .A1(n5626), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5645) );
  INV_X1 U5984 ( .A(n8193), .ZN(n5482) );
  NOR2_X1 U5985 ( .A1(n8669), .A2(n4759), .ZN(n8896) );
  NAND2_X1 U5986 ( .A1(n6478), .A2(n8225), .ZN(n6983) );
  NAND2_X1 U5987 ( .A1(n6604), .A2(n6603), .ZN(n6861) );
  INV_X1 U5988 ( .A(n7272), .ZN(n7201) );
  INV_X1 U5989 ( .A(n6039), .ZN(n5212) );
  OR2_X1 U5990 ( .A1(n5224), .A2(n4788), .ZN(n5234) );
  OR2_X1 U5991 ( .A1(n5135), .A2(n6421), .ZN(n5150) );
  NAND2_X1 U5992 ( .A1(n4959), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4941) );
  OR2_X1 U5993 ( .A1(n9623), .A2(n9478), .ZN(n5191) );
  AND2_X1 U5994 ( .A1(n5168), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5185) );
  OR2_X1 U5995 ( .A1(n9672), .A2(n7307), .ZN(n7928) );
  NAND2_X1 U5996 ( .A1(n9366), .A2(n9873), .ZN(n9369) );
  NAND2_X1 U5997 ( .A1(n6940), .A2(n5056), .ZN(n7300) );
  OR2_X1 U5998 ( .A1(n6930), .A2(n9846), .ZN(n5027) );
  NAND2_X1 U5999 ( .A1(n7846), .A2(n7845), .ZN(n7851) );
  INV_X1 U6000 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6001 ( .A1(n4864), .A2(n7458), .ZN(n4867) );
  INV_X1 U6002 ( .A(n5087), .ZN(n4851) );
  NAND2_X1 U6003 ( .A1(n5451), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U6004 ( .A1(n7177), .A2(n5728), .ZN(n7613) );
  INV_X1 U6005 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7434) );
  OR3_X1 U6006 ( .A1(n5895), .A2(n8461), .A3(n6009), .ZN(n5908) );
  NAND2_X1 U6007 ( .A1(n5775), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5793) );
  OR2_X1 U6008 ( .A1(n5856), .A2(n5854), .ZN(n5875) );
  AND2_X1 U6009 ( .A1(n6499), .A2(n5960), .ZN(n6818) );
  INV_X1 U6010 ( .A(n5574), .ZN(n5924) );
  OR2_X1 U6011 ( .A1(n5546), .A2(n6694), .ZN(n5547) );
  NAND2_X1 U6012 ( .A1(n8934), .A2(n8679), .ZN(n8898) );
  NAND2_X1 U6013 ( .A1(n9971), .A2(n5977), .ZN(n8943) );
  NOR2_X1 U6014 ( .A1(n5956), .A2(n7687), .ZN(n9969) );
  INV_X1 U6015 ( .A(n9288), .ZN(n6870) );
  AND2_X1 U6016 ( .A1(n5093), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5107) );
  AND2_X1 U6017 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5001) );
  OR2_X1 U6018 ( .A1(n6388), .A2(n6299), .ZN(n9682) );
  AND2_X1 U6019 ( .A1(n5313), .A2(n5312), .ZN(n9342) );
  OR2_X1 U6020 ( .A1(n9299), .A2(n6299), .ZN(n9808) );
  NOR2_X1 U6021 ( .A1(n4763), .A2(n4762), .ZN(n5269) );
  AND2_X1 U6022 ( .A1(n7808), .A2(n7794), .ZN(n7880) );
  AND2_X1 U6023 ( .A1(n7928), .A2(n7932), .ZN(n7874) );
  AND2_X1 U6024 ( .A1(n7915), .A2(n7781), .ZN(n7911) );
  INV_X1 U6025 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U6026 ( .A1(n7760), .A2(n7759), .ZN(n7761) );
  AND2_X1 U6027 ( .A1(n7924), .A2(n7923), .ZN(n7872) );
  OR2_X1 U6028 ( .A1(n6366), .A2(n8047), .ZN(n9946) );
  INV_X1 U6029 ( .A(n6378), .ZN(n9893) );
  AND2_X1 U6030 ( .A1(n4872), .A2(n4871), .ZN(n5158) );
  AND2_X1 U6031 ( .A1(n4847), .A2(n4846), .ZN(n5075) );
  OR3_X1 U6032 ( .A1(n7580), .A2(n7656), .A3(n7687), .ZN(n6663) );
  OAI21_X1 U6033 ( .B1(n8698), .B2(n8544), .A(n5996), .ZN(n5997) );
  AND2_X1 U6034 ( .A1(n5983), .A2(n5982), .ZN(n8460) );
  OAI21_X1 U6035 ( .B1(n8774), .B2(n8544), .A(n6012), .ZN(n6013) );
  AND2_X1 U6036 ( .A1(n6818), .A2(n5964), .ZN(n5983) );
  INV_X1 U6037 ( .A(n8518), .ZN(n8532) );
  NAND2_X1 U6038 ( .A1(n5978), .A2(n8943), .ZN(n8508) );
  AND4_X1 U6039 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n8538)
         );
  INV_X1 U6040 ( .A(n8613), .ZN(n7710) );
  INV_X1 U6041 ( .A(n8776), .ZN(n8769) );
  AND2_X1 U6042 ( .A1(n8268), .A2(n8265), .ZN(n8655) );
  AND2_X1 U6043 ( .A1(n8970), .A2(n8969), .ZN(n9114) );
  AND2_X1 U6044 ( .A1(n6663), .A2(n9978), .ZN(n9971) );
  AND2_X1 U6045 ( .A1(n5623), .A2(n5622), .ZN(n6688) );
  AND2_X1 U6046 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  INV_X1 U6047 ( .A(n9682), .ZN(n9222) );
  INV_X1 U6048 ( .A(n9898), .ZN(n9913) );
  AND4_X1 U6049 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n9347)
         );
  AND2_X1 U6050 ( .A1(n6171), .A2(n6172), .ZN(n6244) );
  AND2_X1 U6051 ( .A1(n6126), .A2(n6299), .ZN(n9817) );
  AND2_X1 U6052 ( .A1(n6120), .A2(n6119), .ZN(n9813) );
  INV_X1 U6053 ( .A(n8067), .ZN(n9345) );
  AND2_X1 U6054 ( .A1(n7898), .A2(n7970), .ZN(n9469) );
  AND2_X1 U6055 ( .A1(n7587), .A2(n7586), .ZN(n7955) );
  INV_X1 U6056 ( .A(n9946), .ZN(n9914) );
  OR2_X1 U6057 ( .A1(n6366), .A2(n5391), .ZN(n9898) );
  AND2_X1 U6058 ( .A1(n9878), .A2(n9918), .ZN(n9922) );
  AND2_X1 U6059 ( .A1(n5424), .A2(n6282), .ZN(n6020) );
  INV_X8 U6060 ( .A(n5475), .ZN(n7852) );
  INV_X1 U6061 ( .A(n8629), .ZN(n8599) );
  INV_X1 U6062 ( .A(n6013), .ZN(n6014) );
  OR2_X1 U6063 ( .A1(n8518), .A2(n5970), .ZN(n8516) );
  INV_X1 U6064 ( .A(n9087), .ZN(n8863) );
  OR3_X1 U6065 ( .A1(n5820), .A2(n5819), .A3(n5818), .ZN(n8868) );
  INV_X1 U6066 ( .A(n8538), .ZN(n8929) );
  INV_X1 U6067 ( .A(n6827), .ZN(n8555) );
  AND2_X1 U6068 ( .A1(n6219), .A2(n6218), .ZN(n8629) );
  AND2_X1 U6069 ( .A1(n8931), .A2(n8930), .ZN(n9109) );
  INV_X1 U6070 ( .A(n10039), .ZN(n10037) );
  NAND2_X1 U6071 ( .A1(n9971), .A2(n9970), .ZN(n9975) );
  XNOR2_X1 U6072 ( .A(n5951), .B(n5950), .ZN(n7580) );
  INV_X1 U6073 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6092) );
  INV_X1 U6074 ( .A(n9572), .ZN(n9344) );
  INV_X1 U6075 ( .A(n9611), .ZN(n9467) );
  AND2_X1 U6076 ( .A1(n6446), .A2(n6445), .ZN(n9699) );
  INV_X1 U6077 ( .A(n9694), .ZN(n9278) );
  INV_X1 U6078 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9765) );
  OR2_X1 U6079 ( .A1(n9321), .A2(n9320), .ZN(n9571) );
  INV_X1 U6080 ( .A(n9968), .ZN(n9965) );
  INV_X1 U6081 ( .A(n9952), .ZN(n9950) );
  AND2_X1 U6082 ( .A1(n6442), .A2(n5401), .ZN(n9889) );
  INV_X1 U6083 ( .A(n4785), .ZN(n9669) );
  INV_X1 U6084 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6090) );
  AND2_X1 U6085 ( .A1(n6037), .A2(n9978), .ZN(P2_U3966) );
  NAND2_X1 U6086 ( .A1(n4952), .A2(n4764), .ZN(n4987) );
  NOR2_X1 U6087 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4770) );
  NOR2_X1 U6088 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4769) );
  INV_X1 U6089 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4775) );
  INV_X1 U6090 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U6091 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4777) );
  INV_X1 U6092 ( .A(n4926), .ZN(n4778) );
  NAND2_X1 U6093 ( .A1(n4778), .A2(n4348), .ZN(n4780) );
  INV_X1 U6094 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4779) );
  INV_X1 U6095 ( .A(n4786), .ZN(n8170) );
  INV_X1 U6096 ( .A(n4781), .ZN(n4783) );
  NOR3_X1 U6097 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U6098 ( .A1(n4783), .A2(n4782), .ZN(n9662) );
  NAND2_X1 U6099 ( .A1(n9662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4784) );
  INV_X1 U6100 ( .A(n4958), .ZN(n4969) );
  NAND2_X1 U6101 ( .A1(n5236), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n4798) );
  AND2_X2 U6102 ( .A1(n4786), .A2(n9669), .ZN(n4959) );
  NAND2_X1 U6103 ( .A1(n6325), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U6104 ( .A1(n5328), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U6105 ( .A1(n5001), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6106 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n4787) );
  NOR2_X1 U6107 ( .A1(n5028), .A2(n4787), .ZN(n5043) );
  NAND2_X1 U6108 ( .A1(n5043), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5067) );
  INV_X1 U6109 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5066) );
  INV_X1 U6110 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U6111 ( .A1(n5107), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5121) );
  INV_X1 U6112 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5120) );
  INV_X1 U6113 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6421) );
  INV_X1 U6114 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6115 ( .A1(n5198), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6116 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n4788) );
  INV_X1 U6117 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U6118 ( .A1(n5254), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5255) );
  INV_X1 U6119 ( .A(n5255), .ZN(n5274) );
  NAND2_X1 U6120 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5274), .ZN(n5287) );
  INV_X1 U6121 ( .A(n5287), .ZN(n4789) );
  NAND2_X1 U6122 ( .A1(n4789), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5299) );
  INV_X1 U6123 ( .A(n5299), .ZN(n4790) );
  NAND2_X1 U6124 ( .A1(n4790), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5311) );
  INV_X1 U6125 ( .A(n5311), .ZN(n4791) );
  NAND2_X1 U6126 ( .A1(n4791), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5313) );
  INV_X1 U6127 ( .A(n5313), .ZN(n4792) );
  NAND2_X1 U6128 ( .A1(n4792), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5329) );
  INV_X1 U6129 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U6130 ( .A1(n5313), .A2(n4793), .ZN(n4794) );
  NAND2_X1 U6131 ( .A1(n5329), .A2(n4794), .ZN(n9331) );
  OR2_X1 U6132 ( .A1(n5275), .A2(n9331), .ZN(n4795) );
  INV_X1 U6133 ( .A(n9347), .ZN(n9281) );
  NAND2_X1 U6134 ( .A1(n7534), .A2(n4799), .ZN(n4802) );
  NAND2_X4 U6135 ( .A1(n4802), .A2(n4801), .ZN(n4824) );
  INV_X1 U6136 ( .A(n4824), .ZN(n4804) );
  AND2_X1 U6137 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U6138 ( .A1(n4804), .A2(n4803), .ZN(n5539) );
  AND2_X1 U6139 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U6140 ( .A1(n4824), .A2(n4805), .ZN(n4947) );
  INV_X1 U6141 ( .A(SI_1_), .ZN(n4806) );
  MUX2_X1 U6142 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4824), .Z(n4933) );
  NAND2_X1 U6143 ( .A1(n4934), .A2(n4933), .ZN(n4808) );
  MUX2_X1 U6144 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4824), .Z(n4810) );
  INV_X1 U6145 ( .A(SI_2_), .ZN(n4809) );
  XNOR2_X1 U6146 ( .A(n4810), .B(n4809), .ZN(n4953) );
  NAND2_X1 U6147 ( .A1(n4954), .A2(n4953), .ZN(n4812) );
  NAND2_X1 U6148 ( .A1(n4810), .A2(SI_2_), .ZN(n4811) );
  MUX2_X1 U6149 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4824), .Z(n4818) );
  XNOR2_X1 U6150 ( .A(n4818), .B(SI_3_), .ZN(n4979) );
  INV_X1 U6151 ( .A(n4979), .ZN(n4989) );
  NAND2_X1 U6152 ( .A1(n4814), .A2(SI_4_), .ZN(n4819) );
  INV_X1 U6153 ( .A(n4819), .ZN(n4815) );
  INV_X1 U6154 ( .A(SI_4_), .ZN(n7385) );
  AND2_X1 U6155 ( .A1(n4989), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U6156 ( .A1(n4990), .A2(n4816), .ZN(n4823) );
  INV_X1 U6157 ( .A(n4817), .ZN(n4821) );
  NAND2_X1 U6158 ( .A1(n4818), .A2(SI_3_), .ZN(n4991) );
  AND2_X1 U6159 ( .A1(n4991), .A2(n4819), .ZN(n4820) );
  OR2_X1 U6160 ( .A1(n4821), .A2(n4820), .ZN(n4822) );
  INV_X1 U6161 ( .A(SI_5_), .ZN(n4827) );
  NAND2_X1 U6162 ( .A1(n5011), .A2(n5010), .ZN(n4830) );
  NAND2_X1 U6163 ( .A1(n4828), .A2(SI_5_), .ZN(n4829) );
  NAND2_X2 U6164 ( .A1(n4830), .A2(n4829), .ZN(n5019) );
  INV_X1 U6165 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6074) );
  INV_X1 U6166 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6081) );
  MUX2_X1 U6167 ( .A(n6074), .B(n6081), .S(n7852), .Z(n4831) );
  INV_X1 U6168 ( .A(n4831), .ZN(n4832) );
  NAND2_X1 U6169 ( .A1(n4832), .A2(SI_6_), .ZN(n4833) );
  MUX2_X1 U6170 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7852), .Z(n4834) );
  INV_X1 U6171 ( .A(SI_7_), .ZN(n7460) );
  MUX2_X1 U6172 ( .A(n6092), .B(n6090), .S(n7852), .Z(n4836) );
  INV_X1 U6173 ( .A(SI_8_), .ZN(n4835) );
  INV_X1 U6174 ( .A(n4836), .ZN(n4837) );
  NAND2_X1 U6175 ( .A1(n4837), .A2(SI_8_), .ZN(n4838) );
  INV_X1 U6176 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6094) );
  INV_X1 U6177 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6095) );
  MUX2_X1 U6178 ( .A(n6094), .B(n6095), .S(n7852), .Z(n4840) );
  INV_X1 U6179 ( .A(SI_9_), .ZN(n7449) );
  INV_X1 U6180 ( .A(n4840), .ZN(n4841) );
  NAND2_X1 U6181 ( .A1(n4841), .A2(SI_9_), .ZN(n4842) );
  INV_X1 U6182 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6100) );
  INV_X1 U6183 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6098) );
  MUX2_X1 U6184 ( .A(n6100), .B(n6098), .S(n7852), .Z(n4844) );
  INV_X1 U6185 ( .A(SI_10_), .ZN(n7436) );
  NAND2_X1 U6186 ( .A1(n4844), .A2(n7436), .ZN(n4847) );
  INV_X1 U6187 ( .A(n4844), .ZN(n4845) );
  NAND2_X1 U6188 ( .A1(n4845), .A2(SI_10_), .ZN(n4846) );
  MUX2_X1 U6189 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7852), .Z(n4849) );
  INV_X1 U6190 ( .A(SI_11_), .ZN(n7375) );
  NAND2_X1 U6191 ( .A1(n4849), .A2(SI_11_), .ZN(n4850) );
  INV_X1 U6192 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6114) );
  INV_X1 U6193 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6112) );
  MUX2_X1 U6194 ( .A(n6114), .B(n6112), .S(n7852), .Z(n4852) );
  INV_X1 U6195 ( .A(n4852), .ZN(n4853) );
  NAND2_X1 U6196 ( .A1(n4853), .A2(SI_12_), .ZN(n4854) );
  INV_X1 U6197 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6185) );
  INV_X1 U6198 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6186) );
  MUX2_X1 U6199 ( .A(n6185), .B(n6186), .S(n7852), .Z(n4856) );
  INV_X1 U6200 ( .A(SI_13_), .ZN(n7475) );
  NAND2_X1 U6201 ( .A1(n4856), .A2(n7475), .ZN(n4859) );
  INV_X1 U6202 ( .A(n4856), .ZN(n4857) );
  NAND2_X1 U6203 ( .A1(n4857), .A2(SI_13_), .ZN(n4858) );
  INV_X1 U6204 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6278) );
  INV_X1 U6205 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6279) );
  MUX2_X1 U6206 ( .A(n6278), .B(n6279), .S(n7852), .Z(n4860) );
  INV_X1 U6207 ( .A(n4860), .ZN(n4861) );
  NAND2_X1 U6208 ( .A1(n4861), .A2(SI_14_), .ZN(n4862) );
  INV_X1 U6209 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6362) );
  INV_X1 U6210 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4863) );
  MUX2_X1 U6211 ( .A(n6362), .B(n4863), .S(n7852), .Z(n4864) );
  INV_X1 U6212 ( .A(n4864), .ZN(n4865) );
  NAND2_X1 U6213 ( .A1(n4865), .A2(SI_15_), .ZN(n4866) );
  NAND2_X1 U6214 ( .A1(n4867), .A2(n4866), .ZN(n5142) );
  INV_X1 U6215 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n4868) );
  INV_X1 U6216 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6415) );
  MUX2_X1 U6217 ( .A(n4868), .B(n6415), .S(n7852), .Z(n4869) );
  INV_X1 U6218 ( .A(SI_16_), .ZN(n7438) );
  NAND2_X1 U6219 ( .A1(n4869), .A2(n7438), .ZN(n4872) );
  INV_X1 U6220 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6221 ( .A1(n4870), .A2(SI_16_), .ZN(n4871) );
  NAND2_X1 U6222 ( .A1(n5159), .A2(n5158), .ZN(n4873) );
  NAND2_X1 U6223 ( .A1(n4873), .A2(n4872), .ZN(n5177) );
  INV_X1 U6224 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6454) );
  INV_X1 U6225 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6455) );
  MUX2_X1 U6226 ( .A(n6454), .B(n6455), .S(n7852), .Z(n4874) );
  XNOR2_X1 U6227 ( .A(n4874), .B(SI_17_), .ZN(n5176) );
  INV_X1 U6228 ( .A(n5176), .ZN(n4877) );
  INV_X1 U6229 ( .A(n4874), .ZN(n4875) );
  NAND2_X1 U6230 ( .A1(n4875), .A2(SI_17_), .ZN(n4876) );
  OAI21_X1 U6231 ( .B1(n5177), .B2(n4877), .A(n4876), .ZN(n5193) );
  MUX2_X1 U6232 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7852), .Z(n4879) );
  XNOR2_X1 U6233 ( .A(n4879), .B(SI_18_), .ZN(n5192) );
  INV_X1 U6234 ( .A(n5192), .ZN(n4878) );
  NAND2_X1 U6235 ( .A1(n4879), .A2(SI_18_), .ZN(n4880) );
  INV_X1 U6236 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8404) );
  INV_X1 U6237 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U6238 ( .A(n8404), .B(n6549), .S(n7852), .Z(n4882) );
  INV_X1 U6239 ( .A(SI_19_), .ZN(n4881) );
  NAND2_X1 U6240 ( .A1(n4882), .A2(n4881), .ZN(n4885) );
  INV_X1 U6241 ( .A(n4882), .ZN(n4883) );
  NAND2_X1 U6242 ( .A1(n4883), .A2(SI_19_), .ZN(n4884) );
  NAND2_X1 U6243 ( .A1(n4885), .A2(n4884), .ZN(n5204) );
  INV_X1 U6244 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6632) );
  INV_X1 U6245 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6716) );
  MUX2_X1 U6246 ( .A(n6632), .B(n6716), .S(n7852), .Z(n4886) );
  INV_X1 U6247 ( .A(SI_20_), .ZN(n7373) );
  NAND2_X1 U6248 ( .A1(n4886), .A2(n7373), .ZN(n4889) );
  INV_X1 U6249 ( .A(n4886), .ZN(n4887) );
  NAND2_X1 U6250 ( .A1(n4887), .A2(SI_20_), .ZN(n4888) );
  NAND2_X1 U6251 ( .A1(n5221), .A2(n5220), .ZN(n4890) );
  MUX2_X1 U6252 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7852), .Z(n4892) );
  INV_X1 U6253 ( .A(SI_21_), .ZN(n4891) );
  XNOR2_X1 U6254 ( .A(n4892), .B(n4891), .ZN(n5230) );
  INV_X1 U6255 ( .A(n5230), .ZN(n4894) );
  NAND2_X1 U6256 ( .A1(n4892), .A2(SI_21_), .ZN(n4893) );
  INV_X1 U6257 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6889) );
  INV_X1 U6258 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7061) );
  MUX2_X1 U6259 ( .A(n6889), .B(n7061), .S(n7852), .Z(n4896) );
  INV_X1 U6260 ( .A(SI_22_), .ZN(n4895) );
  NAND2_X1 U6261 ( .A1(n4896), .A2(n4895), .ZN(n4899) );
  INV_X1 U6262 ( .A(n4896), .ZN(n4897) );
  NAND2_X1 U6263 ( .A1(n4897), .A2(SI_22_), .ZN(n4898) );
  NAND2_X1 U6264 ( .A1(n4899), .A2(n4898), .ZN(n5239) );
  INV_X1 U6265 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4900) );
  INV_X1 U6266 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7093) );
  MUX2_X1 U6267 ( .A(n4900), .B(n7093), .S(n7852), .Z(n4902) );
  INV_X1 U6268 ( .A(SI_23_), .ZN(n4901) );
  NAND2_X1 U6269 ( .A1(n4902), .A2(n4901), .ZN(n4905) );
  INV_X1 U6270 ( .A(n4902), .ZN(n4903) );
  NAND2_X1 U6271 ( .A1(n4903), .A2(SI_23_), .ZN(n4904) );
  NAND2_X1 U6272 ( .A1(n4905), .A2(n4904), .ZN(n5248) );
  MUX2_X1 U6273 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7852), .Z(n4910) );
  INV_X1 U6274 ( .A(SI_24_), .ZN(n4906) );
  XNOR2_X1 U6275 ( .A(n4910), .B(n4906), .ZN(n5271) );
  INV_X1 U6276 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7654) );
  INV_X1 U6277 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7652) );
  MUX2_X1 U6278 ( .A(n7654), .B(n7652), .S(n7852), .Z(n4907) );
  INV_X1 U6279 ( .A(SI_25_), .ZN(n7356) );
  NAND2_X1 U6280 ( .A1(n4907), .A2(n7356), .ZN(n4913) );
  INV_X1 U6281 ( .A(n4907), .ZN(n4908) );
  NAND2_X1 U6282 ( .A1(n4908), .A2(SI_25_), .ZN(n4909) );
  NAND2_X1 U6283 ( .A1(n4913), .A2(n4909), .ZN(n5284) );
  INV_X1 U6284 ( .A(n5284), .ZN(n4911) );
  NAND2_X1 U6285 ( .A1(n4910), .A2(SI_24_), .ZN(n5282) );
  AND2_X1 U6286 ( .A1(n4911), .A2(n5282), .ZN(n4912) );
  NAND2_X1 U6287 ( .A1(n5283), .A2(n4912), .ZN(n4914) );
  INV_X1 U6288 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7686) );
  INV_X1 U6289 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7677) );
  MUX2_X1 U6290 ( .A(n7686), .B(n7677), .S(n7852), .Z(n4915) );
  INV_X1 U6291 ( .A(SI_26_), .ZN(n7353) );
  NAND2_X1 U6292 ( .A1(n4915), .A2(n7353), .ZN(n4918) );
  INV_X1 U6293 ( .A(n4915), .ZN(n4916) );
  NAND2_X1 U6294 ( .A1(n4916), .A2(SI_26_), .ZN(n4917) );
  AND2_X1 U6295 ( .A1(n4918), .A2(n4917), .ZN(n5295) );
  NAND2_X1 U6296 ( .A1(n5296), .A2(n5295), .ZN(n4919) );
  INV_X1 U6297 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n4920) );
  INV_X1 U6298 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5307) );
  MUX2_X1 U6299 ( .A(n4920), .B(n5307), .S(n7852), .Z(n4921) );
  INV_X1 U6300 ( .A(SI_27_), .ZN(n7477) );
  NAND2_X1 U6301 ( .A1(n4921), .A2(n7477), .ZN(n4924) );
  INV_X1 U6302 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6303 ( .A1(n4922), .A2(SI_27_), .ZN(n4923) );
  AND2_X1 U6304 ( .A1(n4924), .A2(n4923), .ZN(n5305) );
  MUX2_X1 U6305 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7852), .Z(n5321) );
  INV_X1 U6306 ( .A(SI_28_), .ZN(n5322) );
  XNOR2_X1 U6307 ( .A(n5321), .B(n5322), .ZN(n5319) );
  INV_X1 U6308 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4927) );
  XNOR2_X1 U6309 ( .A(n4928), .B(n4927), .ZN(n5382) );
  NAND2_X1 U6310 ( .A1(n6039), .A2(n7852), .ZN(n4955) );
  NAND2_X1 U6311 ( .A1(n7768), .A2(n7859), .ZN(n4930) );
  INV_X1 U6312 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7750) );
  OR2_X1 U6313 ( .A1(n7857), .A2(n7750), .ZN(n4929) );
  INV_X1 U6314 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4932) );
  NAND2_X1 U6315 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4931) );
  XNOR2_X1 U6316 ( .A(n4932), .B(n4931), .ZN(n6312) );
  INV_X1 U6317 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U6318 ( .A(n4934), .B(n4933), .ZN(n6075) );
  OR2_X1 U6319 ( .A1(n4955), .A2(n6075), .ZN(n4935) );
  OAI211_X1 U6320 ( .C1(n6039), .C2(n6312), .A(n4936), .B(n4935), .ZN(n6378)
         );
  NAND2_X1 U6321 ( .A1(n4958), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U6322 ( .A1(n4960), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U6323 ( .A1(n4333), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U6324 ( .A1(n4959), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6325 ( .A1(n4958), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6326 ( .A1(n4333), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4942) );
  INV_X1 U6327 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6328 ( .A1(n7852), .A2(SI_0_), .ZN(n4946) );
  INV_X1 U6329 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U6330 ( .A1(n4946), .A2(n4945), .ZN(n4948) );
  AND2_X1 U6331 ( .A1(n4948), .A2(n4947), .ZN(n6069) );
  AND2_X1 U6332 ( .A1(n6292), .A2(n9860), .ZN(n9864) );
  NAND2_X1 U6333 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  NAND2_X1 U6334 ( .A1(n9291), .A2(n6378), .ZN(n4951) );
  NAND2_X1 U6335 ( .A1(n9863), .A2(n4951), .ZN(n6633) );
  INV_X1 U6336 ( .A(n6633), .ZN(n4967) );
  INV_X1 U6337 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5164) );
  OR2_X1 U6338 ( .A1(n4952), .A2(n5164), .ZN(n4975) );
  INV_X1 U6339 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4974) );
  XNOR2_X1 U6340 ( .A(n4975), .B(n4974), .ZN(n9754) );
  INV_X1 U6341 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U6342 ( .A(n4954), .B(n4953), .ZN(n6086) );
  OAI211_X1 U6343 ( .C1(n6039), .C2(n9754), .A(n4957), .B(n4956), .ZN(n6394)
         );
  NAND2_X1 U6344 ( .A1(n4333), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6345 ( .A1(n4958), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6346 ( .A1(n4959), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4962) );
  OR2_X1 U6347 ( .A1(n9874), .A2(n6394), .ZN(n4968) );
  NAND2_X1 U6348 ( .A1(n6635), .A2(n4968), .ZN(n6536) );
  INV_X1 U6349 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U6350 ( .A1(n5330), .A2(n6447), .ZN(n4973) );
  NAND2_X1 U6351 ( .A1(n5236), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6352 ( .A1(n4959), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6353 ( .A1(n5328), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6354 ( .A1(n4975), .A2(n4974), .ZN(n4976) );
  NAND2_X1 U6355 ( .A1(n4976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4978) );
  INV_X1 U6356 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U6357 ( .A(n4978), .B(n4977), .ZN(n6148) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6088) );
  OR2_X1 U6359 ( .A1(n5039), .A2(n4332), .ZN(n4980) );
  INV_X1 U6360 ( .A(n9905), .ZN(n6544) );
  OR2_X1 U6361 ( .A1(n9290), .A2(n6544), .ZN(n8054) );
  NAND2_X1 U6362 ( .A1(n6544), .A2(n9290), .ZN(n7783) );
  NAND2_X1 U6363 ( .A1(n6536), .A2(n7865), .ZN(n6554) );
  OR2_X1 U6364 ( .A1(n9290), .A2(n9905), .ZN(n6553) );
  NAND2_X1 U6365 ( .A1(n5328), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6366 ( .A1(n5236), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U6367 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n4982) );
  NOR2_X1 U6368 ( .A1(n5001), .A2(n4982), .ZN(n9223) );
  NAND2_X1 U6369 ( .A1(n5330), .A2(n9223), .ZN(n4984) );
  NAND2_X1 U6370 ( .A1(n4959), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4983) );
  NAND4_X2 U6371 ( .A1(n4986), .A2(n4985), .A3(n4984), .A4(n4983), .ZN(n9845)
         );
  NAND2_X1 U6372 ( .A1(n4987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4988) );
  XNOR2_X1 U6373 ( .A(n4988), .B(n4765), .ZN(n9778) );
  INV_X1 U6374 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6085) );
  OR2_X1 U6375 ( .A1(n7857), .A2(n6085), .ZN(n4996) );
  NAND2_X1 U6376 ( .A1(n4990), .A2(n4989), .ZN(n4992) );
  NAND2_X1 U6377 ( .A1(n4992), .A2(n4991), .ZN(n4994) );
  XNOR2_X1 U6378 ( .A(n4994), .B(n4993), .ZN(n6084) );
  OR2_X1 U6379 ( .A1(n5039), .A2(n6084), .ZN(n4995) );
  OAI211_X1 U6380 ( .C1(n6039), .C2(n9778), .A(n4996), .B(n4995), .ZN(n9912)
         );
  OR2_X1 U6381 ( .A1(n9845), .A2(n9912), .ZN(n4997) );
  AND2_X1 U6382 ( .A1(n6553), .A2(n4997), .ZN(n5000) );
  INV_X1 U6383 ( .A(n4997), .ZN(n4998) );
  AOI21_X1 U6384 ( .B1(n6554), .B2(n5000), .A(n4999), .ZN(n9851) );
  OAI21_X1 U6385 ( .B1(n5001), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5028), .ZN(
        n9838) );
  NAND2_X1 U6386 ( .A1(n5328), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U6387 ( .A1(n5236), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6388 ( .A1(n4959), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5002) );
  INV_X1 U6389 ( .A(n9289), .ZN(n5014) );
  NAND2_X1 U6390 ( .A1(n5006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5007) );
  MUX2_X1 U6391 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5007), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5009) );
  AND2_X1 U6392 ( .A1(n5009), .A2(n4674), .ZN(n6167) );
  INV_X1 U6393 ( .A(n6167), .ZN(n6194) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6079) );
  OR2_X1 U6395 ( .A1(n7857), .A2(n6079), .ZN(n5013) );
  XNOR2_X1 U6396 ( .A(n5011), .B(n5010), .ZN(n6078) );
  OR2_X1 U6397 ( .A1(n5039), .A2(n6078), .ZN(n5012) );
  OAI211_X1 U6398 ( .C1(n6039), .C2(n6194), .A(n5013), .B(n5012), .ZN(n5015)
         );
  INV_X1 U6399 ( .A(n5015), .ZN(n9839) );
  NAND2_X1 U6400 ( .A1(n9839), .A2(n9289), .ZN(n7905) );
  NAND2_X1 U6401 ( .A1(n9289), .A2(n5015), .ZN(n5016) );
  NAND2_X1 U6402 ( .A1(n9852), .A2(n5016), .ZN(n6890) );
  OR2_X1 U6403 ( .A1(n5008), .A2(n5164), .ZN(n5017) );
  INV_X1 U6404 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U6405 ( .A(n5017), .B(n5035), .ZN(n6274) );
  OR2_X1 U6406 ( .A1(n7857), .A2(n6081), .ZN(n5021) );
  NAND2_X1 U6407 ( .A1(n5328), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6408 ( .A1(n5236), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5024) );
  XNOR2_X1 U6409 ( .A(n5028), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U6410 ( .A1(n5330), .A2(n6934), .ZN(n5023) );
  NAND2_X1 U6411 ( .A1(n4959), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5022) );
  NAND4_X1 U6412 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n9846)
         );
  NAND2_X1 U6413 ( .A1(n6891), .A2(n9846), .ZN(n7781) );
  INV_X1 U6414 ( .A(n5028), .ZN(n5029) );
  AOI21_X1 U6415 ( .B1(n5029), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n5030) );
  OR2_X1 U6416 ( .A1(n5030), .A2(n5043), .ZN(n6722) );
  OR2_X1 U6417 ( .A1(n5275), .A2(n6722), .ZN(n5034) );
  NAND2_X1 U6418 ( .A1(n5236), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6419 ( .A1(n5328), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6420 ( .A1(n4959), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5031) );
  NAND4_X1 U6421 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n9288)
         );
  NAND2_X1 U6422 ( .A1(n5008), .A2(n5035), .ZN(n5049) );
  NAND2_X1 U6423 ( .A1(n5049), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5036) );
  XNOR2_X1 U6424 ( .A(n5036), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6160) );
  INV_X1 U6425 ( .A(n6160), .ZN(n6207) );
  INV_X1 U6426 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6083) );
  OR2_X1 U6427 ( .A1(n7857), .A2(n6083), .ZN(n5041) );
  OR2_X1 U6428 ( .A1(n5039), .A2(n6082), .ZN(n5040) );
  OAI211_X1 U6429 ( .C1(n6039), .C2(n6207), .A(n5041), .B(n5040), .ZN(n6612)
         );
  NAND2_X1 U6430 ( .A1(n6870), .A2(n6612), .ZN(n7916) );
  INV_X1 U6431 ( .A(n6612), .ZN(n6723) );
  NAND2_X1 U6432 ( .A1(n6723), .A2(n9288), .ZN(n7917) );
  NAND2_X1 U6433 ( .A1(n7916), .A2(n7917), .ZN(n7869) );
  NAND2_X1 U6434 ( .A1(n6870), .A2(n6723), .ZN(n5042) );
  NAND2_X1 U6435 ( .A1(n5236), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6436 ( .A1(n5328), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5047) );
  OR2_X1 U6437 ( .A1(n5043), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5044) );
  AND2_X1 U6438 ( .A1(n5067), .A2(n5044), .ZN(n6869) );
  NAND2_X1 U6439 ( .A1(n5330), .A2(n6869), .ZN(n5046) );
  NAND2_X1 U6440 ( .A1(n4959), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5045) );
  NAND4_X1 U6441 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n9287)
         );
  INV_X1 U6442 ( .A(n9287), .ZN(n7306) );
  NAND2_X1 U6443 ( .A1(n5059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5050) );
  XNOR2_X1 U6444 ( .A(n5050), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6228) );
  INV_X1 U6445 ( .A(n6228), .ZN(n6180) );
  XNOR2_X1 U6446 ( .A(n5052), .B(n5051), .ZN(n6089) );
  NAND2_X1 U6447 ( .A1(n7859), .A2(n6089), .ZN(n5054) );
  OR2_X1 U6448 ( .A1(n7857), .A2(n6090), .ZN(n5053) );
  NAND2_X1 U6449 ( .A1(n7306), .A2(n6947), .ZN(n7924) );
  INV_X1 U6450 ( .A(n6947), .ZN(n5055) );
  NAND2_X1 U6451 ( .A1(n5055), .A2(n9287), .ZN(n7923) );
  NAND2_X1 U6452 ( .A1(n9287), .A2(n6947), .ZN(n5056) );
  XNOR2_X1 U6453 ( .A(n5058), .B(n5057), .ZN(n6093) );
  NAND2_X1 U6454 ( .A1(n6093), .A2(n7859), .ZN(n5065) );
  NOR2_X1 U6455 ( .A1(n5059), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5062) );
  OR2_X1 U6456 ( .A1(n5062), .A2(n5164), .ZN(n5060) );
  INV_X1 U6457 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5061) );
  MUX2_X1 U6458 ( .A(n5060), .B(P1_IR_REG_31__SCAN_IN), .S(n5061), .Z(n5063)
         );
  NAND2_X1 U6459 ( .A1(n5062), .A2(n5061), .ZN(n5089) );
  NAND2_X1 U6460 ( .A1(n5063), .A2(n5089), .ZN(n6245) );
  INV_X1 U6461 ( .A(n6245), .ZN(n6227) );
  AOI22_X1 U6462 ( .A1(n5213), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5212), .B2(
        n6227), .ZN(n5064) );
  NAND2_X1 U6463 ( .A1(n5328), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6464 ( .A1(n5236), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6465 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  AND2_X1 U6466 ( .A1(n5079), .A2(n5068), .ZN(n9825) );
  NAND2_X1 U6467 ( .A1(n5330), .A2(n9825), .ZN(n5070) );
  NAND2_X1 U6468 ( .A1(n6325), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5069) );
  NAND4_X1 U6469 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9286)
         );
  OR2_X1 U6470 ( .A1(n9827), .A2(n9286), .ZN(n5073) );
  XNOR2_X1 U6471 ( .A(n5074), .B(n5075), .ZN(n6097) );
  NAND2_X1 U6472 ( .A1(n6097), .A2(n7859), .ZN(n5078) );
  NAND2_X1 U6473 ( .A1(n5089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U6474 ( .A(n5076), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6224) );
  AOI22_X1 U6475 ( .A1(n5213), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5212), .B2(
        n6224), .ZN(n5077) );
  AND2_X1 U6476 ( .A1(n5079), .A2(n6256), .ZN(n5080) );
  NOR2_X1 U6477 ( .A1(n5093), .A2(n5080), .ZN(n7083) );
  NAND2_X1 U6478 ( .A1(n5330), .A2(n7083), .ZN(n5084) );
  NAND2_X1 U6479 ( .A1(n5236), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6480 ( .A1(n6325), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6481 ( .A1(n5328), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5081) );
  NAND4_X1 U6482 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n9285)
         );
  INV_X1 U6483 ( .A(n9285), .ZN(n7307) );
  NAND2_X1 U6484 ( .A1(n9672), .A2(n7307), .ZN(n7932) );
  NAND2_X1 U6485 ( .A1(n7262), .A2(n5085), .ZN(n7261) );
  OR2_X1 U6486 ( .A1(n9672), .A2(n9285), .ZN(n5086) );
  NAND2_X1 U6487 ( .A1(n7261), .A2(n5086), .ZN(n7314) );
  XNOR2_X1 U6488 ( .A(n5088), .B(n5087), .ZN(n6101) );
  NAND2_X1 U6489 ( .A1(n6101), .A2(n7859), .ZN(n5092) );
  OAI21_X1 U6490 ( .B1(n5089), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U6491 ( .A(n5090), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6234) );
  AOI22_X1 U6492 ( .A1(n5213), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5212), .B2(
        n6234), .ZN(n5091) );
  NOR2_X1 U6493 ( .A1(n5093), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5094) );
  OR2_X1 U6494 ( .A1(n5107), .A2(n5094), .ZN(n7318) );
  OR2_X1 U6495 ( .A1(n5275), .A2(n7318), .ZN(n5098) );
  NAND2_X1 U6496 ( .A1(n5328), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6497 ( .A1(n5236), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6498 ( .A1(n6325), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6499 ( .A1(n7641), .A2(n9684), .ZN(n5099) );
  NAND2_X1 U6500 ( .A1(n7314), .A2(n5099), .ZN(n5101) );
  OR2_X1 U6501 ( .A1(n7641), .A2(n9684), .ZN(n5100) );
  OR2_X1 U6502 ( .A1(n5104), .A2(n5164), .ZN(n5105) );
  XNOR2_X1 U6503 ( .A(n5105), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6335) );
  AOI22_X1 U6504 ( .A1(n5213), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5212), .B2(
        n6335), .ZN(n5106) );
  OR2_X1 U6505 ( .A1(n5107), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6506 ( .A1(n5121), .A2(n5108), .ZN(n9698) );
  OR2_X1 U6507 ( .A1(n5275), .A2(n9698), .ZN(n5112) );
  NAND2_X1 U6508 ( .A1(n5236), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6509 ( .A1(n6325), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6510 ( .A1(n5328), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6511 ( .A1(n7187), .A2(n9284), .ZN(n5114) );
  OR2_X1 U6512 ( .A1(n7187), .A2(n9284), .ZN(n5113) );
  NAND2_X1 U6513 ( .A1(n5114), .A2(n5113), .ZN(n7878) );
  OAI21_X1 U6514 ( .B1(n7581), .B2(n7878), .A(n5114), .ZN(n7689) );
  XNOR2_X1 U6515 ( .A(n5116), .B(n5115), .ZN(n6184) );
  NAND2_X1 U6516 ( .A1(n6184), .A2(n7859), .ZN(n5119) );
  NAND2_X1 U6517 ( .A1(n5132), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5117) );
  XNOR2_X1 U6518 ( .A(n5117), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6341) );
  AOI22_X1 U6519 ( .A1(n5213), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5212), .B2(
        n6341), .ZN(n5118) );
  NAND2_X1 U6520 ( .A1(n5236), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6521 ( .A1(n6325), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6522 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  AND2_X1 U6523 ( .A1(n5135), .A2(n5122), .ZN(n7701) );
  NAND2_X1 U6524 ( .A1(n5330), .A2(n7701), .ZN(n5124) );
  NAND2_X1 U6525 ( .A1(n5328), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5123) );
  NAND4_X1 U6526 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n9549)
         );
  OR2_X1 U6527 ( .A1(n7702), .A2(n9549), .ZN(n5127) );
  NAND2_X1 U6528 ( .A1(n7689), .A2(n5127), .ZN(n5129) );
  NAND2_X1 U6529 ( .A1(n7702), .A2(n9549), .ZN(n5128) );
  NAND2_X1 U6530 ( .A1(n5129), .A2(n5128), .ZN(n9543) );
  NAND2_X1 U6531 ( .A1(n6277), .A2(n7859), .ZN(n5134) );
  NAND2_X1 U6532 ( .A1(n5163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5144) );
  XNOR2_X1 U6533 ( .A(n5144), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7048) );
  AOI22_X1 U6534 ( .A1(n5213), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5212), .B2(
        n7048), .ZN(n5133) );
  NAND2_X1 U6535 ( .A1(n5328), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6536 ( .A1(n5236), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6537 ( .A1(n5135), .A2(n6421), .ZN(n5136) );
  AND2_X1 U6538 ( .A1(n5150), .A2(n5136), .ZN(n9554) );
  NAND2_X1 U6539 ( .A1(n5330), .A2(n9554), .ZN(n5138) );
  NAND2_X1 U6540 ( .A1(n6325), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5137) );
  NAND4_X1 U6541 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n9283)
         );
  AND2_X1 U6542 ( .A1(n9556), .A2(n9283), .ZN(n5141) );
  XNOR2_X1 U6543 ( .A(n5143), .B(n5142), .ZN(n6323) );
  NAND2_X1 U6544 ( .A1(n6323), .A2(n7859), .ZN(n5148) );
  NAND2_X1 U6545 ( .A1(n5144), .A2(n5161), .ZN(n5145) );
  NAND2_X1 U6546 ( .A1(n5145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5146) );
  XNOR2_X1 U6547 ( .A(n5146), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U6548 ( .A1(n5213), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5212), .B2(
        n9784), .ZN(n5147) );
  NAND2_X1 U6549 ( .A1(n5328), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6550 ( .A1(n5236), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5154) );
  AND2_X1 U6551 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  NOR2_X1 U6552 ( .A1(n5168), .A2(n5151), .ZN(n9536) );
  NAND2_X1 U6553 ( .A1(n5330), .A2(n9536), .ZN(n5153) );
  NAND2_X1 U6554 ( .A1(n6325), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6555 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n9548)
         );
  NOR2_X1 U6556 ( .A1(n9635), .A2(n9548), .ZN(n5157) );
  NAND2_X1 U6557 ( .A1(n9635), .A2(n9548), .ZN(n5156) );
  XNOR2_X1 U6558 ( .A(n5159), .B(n5158), .ZN(n6372) );
  NAND2_X1 U6559 ( .A1(n6372), .A2(n7859), .ZN(n5167) );
  NAND2_X1 U6560 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  OR2_X1 U6561 ( .A1(n5179), .A2(n5164), .ZN(n5165) );
  XNOR2_X1 U6562 ( .A(n5165), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7044) );
  AOI22_X1 U6563 ( .A1(n5213), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5212), .B2(
        n7044), .ZN(n5166) );
  NOR2_X1 U6564 ( .A1(n5168), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5169) );
  OR2_X1 U6565 ( .A1(n5185), .A2(n5169), .ZN(n9510) );
  OR2_X1 U6566 ( .A1(n5275), .A2(n9510), .ZN(n5173) );
  NAND2_X1 U6567 ( .A1(n5236), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6568 ( .A1(n6325), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6569 ( .A1(n5328), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5170) );
  NAND4_X1 U6570 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n9499)
         );
  INV_X1 U6571 ( .A(n9499), .ZN(n9530) );
  NAND2_X1 U6572 ( .A1(n9630), .A2(n9530), .ZN(n7964) );
  NAND2_X1 U6573 ( .A1(n7965), .A2(n7964), .ZN(n9514) );
  NAND2_X1 U6574 ( .A1(n9506), .A2(n9514), .ZN(n5175) );
  NAND2_X1 U6575 ( .A1(n9630), .A2(n9499), .ZN(n5174) );
  NAND2_X1 U6576 ( .A1(n5175), .A2(n5174), .ZN(n9491) );
  XNOR2_X1 U6577 ( .A(n5177), .B(n5176), .ZN(n6453) );
  NAND2_X1 U6578 ( .A1(n6453), .A2(n7859), .ZN(n5184) );
  INV_X1 U6579 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6580 ( .A1(n5179), .A2(n5178), .ZN(n5206) );
  NAND2_X1 U6581 ( .A1(n5206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5181) );
  INV_X1 U6582 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6583 ( .A1(n5181), .A2(n5180), .ZN(n5194) );
  OR2_X1 U6584 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  AND2_X1 U6585 ( .A1(n5194), .A2(n5182), .ZN(n7041) );
  AOI22_X1 U6586 ( .A1(n5213), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5212), .B2(
        n7041), .ZN(n5183) );
  NOR2_X1 U6587 ( .A1(n5185), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6588 ( .A1(n5198), .A2(n5186), .ZN(n9493) );
  OR2_X1 U6589 ( .A1(n5275), .A2(n9493), .ZN(n5190) );
  NAND2_X1 U6590 ( .A1(n5236), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6591 ( .A1(n6325), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6592 ( .A1(n5328), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5187) );
  NAND4_X1 U6593 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n9478)
         );
  XNOR2_X1 U6594 ( .A(n5193), .B(n5192), .ZN(n6491) );
  NAND2_X1 U6595 ( .A1(n6491), .A2(n7859), .ZN(n5197) );
  NAND2_X1 U6596 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6597 ( .A(n5195), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7031) );
  AOI22_X1 U6598 ( .A1(n5213), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5212), .B2(
        n7031), .ZN(n5196) );
  NAND2_X1 U6599 ( .A1(n5328), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6600 ( .A1(n5236), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5202) );
  OR2_X1 U6601 ( .A1(n5198), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5199) );
  AND2_X1 U6602 ( .A1(n5199), .A2(n5224), .ZN(n9482) );
  NAND2_X1 U6603 ( .A1(n5330), .A2(n9482), .ZN(n5201) );
  NAND2_X1 U6604 ( .A1(n6325), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5200) );
  NAND4_X1 U6605 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n9500)
         );
  INV_X1 U6606 ( .A(n9500), .ZN(n9180) );
  OR2_X1 U6607 ( .A1(n9618), .A2(n9180), .ZN(n7897) );
  NAND2_X1 U6608 ( .A1(n9618), .A2(n9180), .ZN(n7818) );
  XNOR2_X1 U6609 ( .A(n5205), .B(n5204), .ZN(n6548) );
  NAND2_X1 U6610 ( .A1(n6548), .A2(n7859), .ZN(n5215) );
  NOR2_X2 U6611 ( .A1(n5206), .A2(n4336), .ZN(n5210) );
  INV_X1 U6612 ( .A(n5210), .ZN(n5207) );
  NAND2_X1 U6613 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6614 ( .A1(n5210), .A2(n5209), .ZN(n5336) );
  INV_X1 U6615 ( .A(n9850), .ZN(n9867) );
  AOI22_X1 U6616 ( .A1(n5213), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9867), .B2(
        n5212), .ZN(n5214) );
  NAND2_X1 U6617 ( .A1(n5236), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6618 ( .A1(n6325), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6619 ( .A(n5224), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U6620 ( .A1(n5330), .A2(n9465), .ZN(n5217) );
  NAND2_X1 U6621 ( .A1(n5328), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5216) );
  NAND4_X1 U6622 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9479)
         );
  OR2_X1 U6623 ( .A1(n9486), .A2(n4755), .ZN(n9445) );
  XNOR2_X1 U6624 ( .A(n5221), .B(n5220), .ZN(n6631) );
  NAND2_X1 U6625 ( .A1(n6631), .A2(n7859), .ZN(n5223) );
  OR2_X1 U6626 ( .A1(n7857), .A2(n6716), .ZN(n5222) );
  NAND2_X1 U6627 ( .A1(n5236), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5229) );
  INV_X1 U6628 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9179) );
  INV_X1 U6629 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9235) );
  OAI21_X1 U6630 ( .B1(n5224), .B2(n9179), .A(n9235), .ZN(n5225) );
  AND2_X1 U6631 ( .A1(n5225), .A2(n5234), .ZN(n9450) );
  NAND2_X1 U6632 ( .A1(n9450), .A2(n5330), .ZN(n5228) );
  NAND2_X1 U6633 ( .A1(n6325), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6634 ( .A1(n5328), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5226) );
  NAND4_X1 U6635 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9470)
         );
  OR2_X1 U6636 ( .A1(n9445), .A2(n4744), .ZN(n9426) );
  XNOR2_X1 U6637 ( .A(n5231), .B(n5230), .ZN(n6718) );
  NAND2_X1 U6638 ( .A1(n6718), .A2(n7859), .ZN(n5233) );
  INV_X1 U6639 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7754) );
  OR2_X1 U6640 ( .A1(n7857), .A2(n7754), .ZN(n5232) );
  AND2_X1 U6641 ( .A1(n5234), .A2(n9187), .ZN(n5235) );
  OR2_X1 U6642 ( .A1(n5235), .A2(n5243), .ZN(n9437) );
  AOI22_X1 U6643 ( .A1(n5236), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5328), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6644 ( .A1(n6325), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5237) );
  OAI211_X1 U6645 ( .C1(n9437), .C2(n5275), .A(n5238), .B(n5237), .ZN(n9455)
         );
  INV_X1 U6646 ( .A(n9455), .ZN(n9248) );
  OR2_X1 U6647 ( .A1(n9601), .A2(n9248), .ZN(n7819) );
  NAND2_X1 U6648 ( .A1(n9601), .A2(n9248), .ZN(n7979) );
  NAND2_X1 U6649 ( .A1(n7819), .A2(n7979), .ZN(n9430) );
  INV_X1 U6650 ( .A(n9430), .ZN(n5264) );
  OR2_X1 U6651 ( .A1(n9426), .A2(n5264), .ZN(n9408) );
  XNOR2_X1 U6652 ( .A(n5240), .B(n5239), .ZN(n6888) );
  NAND2_X1 U6653 ( .A1(n6888), .A2(n7859), .ZN(n5242) );
  OR2_X1 U6654 ( .A1(n7857), .A2(n7061), .ZN(n5241) );
  NOR2_X1 U6655 ( .A1(n5243), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5244) );
  OR2_X1 U6656 ( .A1(n5254), .A2(n5244), .ZN(n9415) );
  AOI22_X1 U6657 ( .A1(n5236), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n5328), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6658 ( .A1(n6325), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5245) );
  OAI211_X1 U6659 ( .C1(n9415), .C2(n5275), .A(n5246), .B(n5245), .ZN(n9435)
         );
  OR2_X1 U6660 ( .A1(n9408), .A2(n4338), .ZN(n9389) );
  INV_X1 U6661 ( .A(n5247), .ZN(n5249) );
  NAND2_X1 U6662 ( .A1(n5249), .A2(n5248), .ZN(n5251) );
  NAND2_X1 U6663 ( .A1(n5251), .A2(n5250), .ZN(n7090) );
  NAND2_X1 U6664 ( .A1(n7090), .A2(n7859), .ZN(n5253) );
  OR2_X1 U6665 ( .A1(n7857), .A2(n7093), .ZN(n5252) );
  OR2_X1 U6666 ( .A1(n5254), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6667 ( .A1(n5256), .A2(n5255), .ZN(n9395) );
  AOI22_X1 U6668 ( .A1(n6325), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5236), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6669 ( .A1(n5328), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5257) );
  OAI211_X1 U6670 ( .C1(n9395), .C2(n5275), .A(n5258), .B(n5257), .ZN(n9421)
         );
  NOR2_X1 U6671 ( .A1(n9591), .A2(n9421), .ZN(n5268) );
  OR2_X1 U6672 ( .A1(n9389), .A2(n5268), .ZN(n5259) );
  NAND2_X1 U6673 ( .A1(n9618), .A2(n9500), .ZN(n9460) );
  NAND2_X1 U6674 ( .A1(n9611), .A2(n9479), .ZN(n5260) );
  AND2_X1 U6675 ( .A1(n9460), .A2(n5260), .ZN(n5261) );
  OR2_X1 U6676 ( .A1(n4755), .A2(n5261), .ZN(n9446) );
  OR2_X1 U6677 ( .A1(n4744), .A2(n9446), .ZN(n5263) );
  NAND2_X1 U6678 ( .A1(n9606), .A2(n9470), .ZN(n5262) );
  AND2_X1 U6679 ( .A1(n5263), .A2(n5262), .ZN(n9427) );
  OR2_X1 U6680 ( .A1(n5264), .A2(n9427), .ZN(n5266) );
  NAND2_X1 U6681 ( .A1(n9601), .A2(n9455), .ZN(n5265) );
  AND2_X1 U6682 ( .A1(n5266), .A2(n5265), .ZN(n9409) );
  AND2_X1 U6683 ( .A1(n4363), .A2(n9409), .ZN(n5267) );
  XNOR2_X1 U6684 ( .A(n5270), .B(n5271), .ZN(n7538) );
  NAND2_X1 U6685 ( .A1(n7538), .A2(n7859), .ZN(n5273) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7539) );
  OR2_X1 U6687 ( .A1(n7857), .A2(n7539), .ZN(n5272) );
  OAI21_X1 U6688 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5274), .A(n5287), .ZN(
        n9384) );
  OR2_X1 U6689 ( .A1(n5275), .A2(n9384), .ZN(n5279) );
  NAND2_X1 U6690 ( .A1(n5236), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6691 ( .A1(n5328), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6692 ( .A1(n6325), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5276) );
  NAND4_X1 U6693 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n9403)
         );
  AND2_X1 U6694 ( .A1(n9588), .A2(n9403), .ZN(n5281) );
  OR2_X1 U6695 ( .A1(n7857), .A2(n7652), .ZN(n5285) );
  NAND2_X1 U6696 ( .A1(n5328), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6697 ( .A1(n5236), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5291) );
  INV_X1 U6698 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U6699 ( .A1(n5287), .A2(n9196), .ZN(n5288) );
  AND2_X1 U6700 ( .A1(n5299), .A2(n5288), .ZN(n9197) );
  NAND2_X1 U6701 ( .A1(n5330), .A2(n9197), .ZN(n5290) );
  NAND2_X1 U6702 ( .A1(n6325), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5289) );
  NAND4_X1 U6703 ( .A1(n5292), .A2(n5291), .A3(n5290), .A4(n5289), .ZN(n9367)
         );
  INV_X1 U6704 ( .A(n9367), .ZN(n9381) );
  NOR2_X1 U6705 ( .A1(n5293), .A2(n9367), .ZN(n5294) );
  AOI21_X1 U6706 ( .B1(n7756), .B2(n7887), .A(n5294), .ZN(n9355) );
  OR2_X1 U6707 ( .A1(n7857), .A2(n7677), .ZN(n5297) );
  NAND2_X1 U6708 ( .A1(n5328), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6709 ( .A1(n5236), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5303) );
  INV_X1 U6710 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U6711 ( .A1(n5299), .A2(n9270), .ZN(n5300) );
  AND2_X1 U6712 ( .A1(n5311), .A2(n5300), .ZN(n9358) );
  NAND2_X1 U6713 ( .A1(n5330), .A2(n9358), .ZN(n5302) );
  NAND2_X1 U6714 ( .A1(n6325), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5301) );
  NAND4_X1 U6715 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9282)
         );
  NAND2_X1 U6716 ( .A1(n9577), .A2(n9282), .ZN(n7888) );
  NAND2_X1 U6717 ( .A1(n7679), .A2(n7859), .ZN(n5309) );
  OR2_X1 U6718 ( .A1(n7857), .A2(n5307), .ZN(n5308) );
  NAND2_X1 U6719 ( .A1(n5236), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6720 ( .A1(n5328), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5316) );
  INV_X1 U6721 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6722 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6723 ( .A1(n5330), .A2(n9342), .ZN(n5315) );
  NAND2_X1 U6724 ( .A1(n6325), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5314) );
  NAND4_X1 U6725 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n9366)
         );
  INV_X1 U6726 ( .A(n9366), .ZN(n9272) );
  NAND2_X1 U6727 ( .A1(n9572), .A2(n9272), .ZN(n8019) );
  OR2_X1 U6728 ( .A1(n9572), .A2(n9366), .ZN(n5318) );
  NAND2_X1 U6729 ( .A1(n9330), .A2(n9347), .ZN(n8024) );
  AOI21_X1 U6730 ( .B1(n9281), .B2(n9330), .A(n9320), .ZN(n5335) );
  INV_X1 U6731 ( .A(n5321), .ZN(n5323) );
  NAND2_X1 U6732 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  MUX2_X1 U6733 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7852), .Z(n7835) );
  INV_X1 U6734 ( .A(SI_29_), .ZN(n7836) );
  XNOR2_X1 U6735 ( .A(n7835), .B(n7836), .ZN(n7833) );
  NAND2_X1 U6736 ( .A1(n8189), .A2(n7859), .ZN(n5327) );
  OR2_X1 U6737 ( .A1(n7857), .A2(n8171), .ZN(n5326) );
  NAND2_X1 U6738 ( .A1(n5328), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6739 ( .A1(n5236), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5333) );
  INV_X1 U6740 ( .A(n5329), .ZN(n6030) );
  NAND2_X1 U6741 ( .A1(n5330), .A2(n6030), .ZN(n5332) );
  NAND2_X1 U6742 ( .A1(n6325), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5331) );
  NAND4_X1 U6743 ( .A1(n5334), .A2(n5333), .A3(n5332), .A4(n5331), .ZN(n9325)
         );
  NAND2_X1 U6744 ( .A1(n5341), .A2(n4428), .ZN(n5337) );
  INV_X1 U6745 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6746 ( .A1(n5377), .A2(n9850), .ZN(n6027) );
  INV_X1 U6747 ( .A(n6284), .ZN(n6286) );
  OR2_X1 U6748 ( .A1(n6027), .A2(n6286), .ZN(n5345) );
  AND2_X1 U6749 ( .A1(n6029), .A2(n9850), .ZN(n5391) );
  NAND2_X1 U6750 ( .A1(n5391), .A2(n5346), .ZN(n6285) );
  OR2_X1 U6751 ( .A1(n6285), .A2(n5343), .ZN(n5344) );
  AND2_X1 U6752 ( .A1(n5345), .A2(n5344), .ZN(n9878) );
  NAND2_X1 U6753 ( .A1(n5346), .A2(n9867), .ZN(n8032) );
  INV_X1 U6754 ( .A(n6029), .ZN(n8047) );
  OR2_X1 U6755 ( .A1(n8032), .A2(n8047), .ZN(n9918) );
  INV_X1 U6756 ( .A(n9865), .ZN(n9870) );
  INV_X1 U6757 ( .A(n9860), .ZN(n6367) );
  NOR2_X1 U6758 ( .A1(n6367), .A2(n6292), .ZN(n9869) );
  NAND2_X1 U6759 ( .A1(n9870), .A2(n9869), .ZN(n5348) );
  OR2_X1 U6760 ( .A1(n9291), .A2(n9893), .ZN(n5347) );
  NAND2_X1 U6761 ( .A1(n5348), .A2(n5347), .ZN(n8051) );
  NAND2_X1 U6762 ( .A1(n8051), .A2(n7866), .ZN(n5349) );
  NAND2_X1 U6763 ( .A1(n5349), .A2(n8050), .ZN(n7803) );
  INV_X1 U6764 ( .A(n7865), .ZN(n5350) );
  NAND2_X1 U6765 ( .A1(n7803), .A2(n5350), .ZN(n5351) );
  INV_X1 U6766 ( .A(n7905), .ZN(n5352) );
  INV_X1 U6767 ( .A(n8058), .ZN(n5353) );
  NAND2_X1 U6768 ( .A1(n8057), .A2(n5355), .ZN(n5357) );
  INV_X1 U6769 ( .A(n7869), .ZN(n5358) );
  INV_X1 U6770 ( .A(n7924), .ZN(n5359) );
  INV_X1 U6771 ( .A(n9286), .ZN(n7084) );
  OR2_X1 U6772 ( .A1(n7084), .A2(n9827), .ZN(n7927) );
  INV_X1 U6773 ( .A(n7928), .ZN(n5361) );
  AND2_X1 U6774 ( .A1(n9827), .A2(n7084), .ZN(n7257) );
  NAND2_X1 U6775 ( .A1(n7928), .A2(n7257), .ZN(n5360) );
  INV_X1 U6776 ( .A(n9284), .ZN(n7213) );
  NAND2_X1 U6777 ( .A1(n7187), .A2(n7213), .ZN(n7933) );
  INV_X1 U6778 ( .A(n9684), .ZN(n5364) );
  NAND2_X1 U6779 ( .A1(n7641), .A2(n5364), .ZN(n7586) );
  NAND2_X1 U6780 ( .A1(n7933), .A2(n7586), .ZN(n7796) );
  NAND2_X1 U6781 ( .A1(n5363), .A2(n5362), .ZN(n7690) );
  INV_X1 U6782 ( .A(n9549), .ZN(n9681) );
  OR2_X1 U6783 ( .A1(n7702), .A2(n9681), .ZN(n7808) );
  NAND2_X1 U6784 ( .A1(n7702), .A2(n9681), .ZN(n7794) );
  OR2_X1 U6785 ( .A1(n7187), .A2(n7213), .ZN(n7956) );
  NAND2_X1 U6786 ( .A1(n7796), .A2(n7956), .ZN(n7938) );
  OR2_X1 U6787 ( .A1(n7641), .A2(n5364), .ZN(n7587) );
  NAND2_X1 U6788 ( .A1(n7878), .A2(n7955), .ZN(n5365) );
  NAND2_X1 U6789 ( .A1(n7938), .A2(n5365), .ZN(n7943) );
  AND2_X1 U6790 ( .A1(n7880), .A2(n7943), .ZN(n5366) );
  NAND2_X1 U6791 ( .A1(n7690), .A2(n5366), .ZN(n7693) );
  INV_X1 U6792 ( .A(n9283), .ZN(n9528) );
  XNOR2_X1 U6793 ( .A(n9556), .B(n9528), .ZN(n9544) );
  OR2_X1 U6794 ( .A1(n9556), .A2(n9528), .ZN(n7930) );
  INV_X1 U6795 ( .A(n9548), .ZN(n9517) );
  OR2_X1 U6796 ( .A1(n9635), .A2(n9517), .ZN(n7941) );
  NAND2_X1 U6797 ( .A1(n9635), .A2(n9517), .ZN(n7942) );
  NAND2_X1 U6798 ( .A1(n7941), .A2(n7942), .ZN(n9525) );
  NAND2_X1 U6799 ( .A1(n9522), .A2(n7942), .ZN(n9515) );
  INV_X1 U6800 ( .A(n7964), .ZN(n5367) );
  INV_X1 U6801 ( .A(n9478), .ZN(n9518) );
  NAND2_X1 U6802 ( .A1(n9623), .A2(n9518), .ZN(n7863) );
  OR2_X1 U6803 ( .A1(n9623), .A2(n9518), .ZN(n9475) );
  AND2_X1 U6804 ( .A1(n7897), .A2(n9475), .ZN(n7899) );
  INV_X1 U6805 ( .A(n9479), .ZN(n9262) );
  OR2_X1 U6806 ( .A1(n9611), .A2(n9262), .ZN(n7898) );
  NAND2_X1 U6807 ( .A1(n9611), .A2(n9262), .ZN(n7970) );
  NAND2_X1 U6808 ( .A1(n9468), .A2(n9469), .ZN(n5368) );
  INV_X1 U6809 ( .A(n9470), .ZN(n9189) );
  OR2_X1 U6810 ( .A1(n9606), .A2(n9189), .ZN(n7978) );
  NAND2_X1 U6811 ( .A1(n9453), .A2(n7978), .ZN(n9432) );
  NAND2_X1 U6812 ( .A1(n9606), .A2(n9189), .ZN(n9431) );
  NAND2_X1 U6813 ( .A1(n9432), .A2(n9431), .ZN(n5369) );
  INV_X1 U6814 ( .A(n9435), .ZN(n9188) );
  OR2_X1 U6815 ( .A1(n9597), .A2(n9188), .ZN(n7822) );
  NAND2_X1 U6816 ( .A1(n9597), .A2(n9188), .ZN(n9400) );
  INV_X1 U6817 ( .A(n9421), .ZN(n9380) );
  NAND2_X1 U6818 ( .A1(n9591), .A2(n9380), .ZN(n7995) );
  NAND2_X1 U6819 ( .A1(n7991), .A2(n7995), .ZN(n7990) );
  INV_X1 U6820 ( .A(n9400), .ZN(n7981) );
  NAND2_X1 U6821 ( .A1(n5370), .A2(n7991), .ZN(n9377) );
  NAND2_X1 U6822 ( .A1(n9588), .A2(n9198), .ZN(n7993) );
  INV_X1 U6823 ( .A(n9282), .ZN(n9348) );
  NAND2_X1 U6824 ( .A1(n9577), .A2(n9348), .ZN(n8009) );
  INV_X1 U6825 ( .A(n8009), .ZN(n7830) );
  OR2_X1 U6826 ( .A1(n9577), .A2(n9348), .ZN(n5372) );
  NAND2_X1 U6827 ( .A1(n9324), .A2(n9323), .ZN(n9322) );
  NAND2_X1 U6828 ( .A1(n9322), .A2(n8023), .ZN(n5374) );
  XNOR2_X1 U6829 ( .A(n5374), .B(n5373), .ZN(n5387) );
  OR2_X1 U6830 ( .A1(n5346), .A2(n9850), .ZN(n5376) );
  OR2_X1 U6831 ( .A1(n5343), .A2(n6029), .ZN(n5375) );
  NAND2_X1 U6832 ( .A1(n5376), .A2(n5375), .ZN(n9871) );
  NAND2_X1 U6833 ( .A1(n5377), .A2(n5342), .ZN(n8042) );
  OR2_X1 U6834 ( .A1(n8042), .A2(n4312), .ZN(n9529) );
  NAND2_X1 U6835 ( .A1(n6325), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6836 ( .A1(n5236), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6837 ( .A1(n5328), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5379) );
  NAND3_X1 U6838 ( .A1(n5381), .A2(n5380), .A3(n5379), .ZN(n9280) );
  INV_X1 U6839 ( .A(n4312), .ZN(n6299) );
  OR2_X1 U6840 ( .A1(n8042), .A2(n6299), .ZN(n9531) );
  INV_X1 U6841 ( .A(P1_B_REG_SCAN_IN), .ZN(n5402) );
  NOR2_X1 U6842 ( .A1(n9755), .A2(n5402), .ZN(n5383) );
  NOR2_X1 U6843 ( .A1(n9531), .A2(n5383), .ZN(n9310) );
  NAND2_X1 U6844 ( .A1(n5346), .A2(n5343), .ZN(n6366) );
  NAND2_X1 U6845 ( .A1(n6639), .A2(n6544), .ZN(n6562) );
  INV_X1 U6846 ( .A(n7641), .ZN(n7317) );
  INV_X1 U6847 ( .A(n9556), .ZN(n9714) );
  INV_X1 U6848 ( .A(n9635), .ZN(n9540) );
  NAND2_X1 U6849 ( .A1(n9532), .A2(n9540), .ZN(n9533) );
  INV_X1 U6850 ( .A(n9618), .ZN(n9484) );
  INV_X1 U6851 ( .A(n9597), .ZN(n9418) );
  INV_X1 U6852 ( .A(n9577), .ZN(n9360) );
  AOI211_X1 U6853 ( .C1(n8029), .C2(n9329), .A(n9946), .B(n9313), .ZN(n6028)
         );
  OR2_X1 U6854 ( .A1(n8042), .A2(n5391), .ZN(n6440) );
  NAND2_X1 U6855 ( .A1(n4339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6856 ( .A(n5392), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6857 ( .A1(n4335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5393) );
  MUX2_X1 U6858 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5393), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5395) );
  NAND2_X1 U6859 ( .A1(n5395), .A2(n5394), .ZN(n7540) );
  INV_X1 U6860 ( .A(n7540), .ZN(n5416) );
  NAND2_X1 U6861 ( .A1(n5394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5396) );
  MUX2_X1 U6862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5396), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5397) );
  AND2_X1 U6863 ( .A1(n5397), .A2(n4339), .ZN(n5421) );
  NAND2_X1 U6864 ( .A1(n5398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5399) );
  MUX2_X1 U6865 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5399), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5400) );
  NAND2_X1 U6866 ( .A1(n5400), .A2(n4335), .ZN(n6441) );
  AND2_X1 U6867 ( .A1(n6441), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5401) );
  NOR2_X1 U6868 ( .A1(n5421), .A2(n5402), .ZN(n5403) );
  MUX2_X1 U6869 ( .A(n5403), .B(n5402), .S(n5416), .Z(n5404) );
  INV_X1 U6870 ( .A(n5417), .ZN(n7678) );
  NOR2_X1 U6871 ( .A1(n5404), .A2(n7678), .ZN(n6105) );
  NOR4_X1 U6872 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5408) );
  NOR4_X1 U6873 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5407) );
  NOR4_X1 U6874 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5406) );
  NOR4_X1 U6875 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5405) );
  NAND4_X1 U6876 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n5414)
         );
  NOR2_X1 U6877 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5412) );
  NOR4_X1 U6878 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5411) );
  NOR4_X1 U6879 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5410) );
  NOR4_X1 U6880 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5409) );
  NAND4_X1 U6881 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n5413)
         );
  NOR2_X1 U6882 ( .A1(n5414), .A2(n5413), .ZN(n6016) );
  NAND2_X1 U6883 ( .A1(n6016), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6884 ( .A1(n6105), .A2(n5415), .ZN(n5418) );
  OR2_X1 U6885 ( .A1(n5417), .A2(n5416), .ZN(n6107) );
  NAND2_X1 U6886 ( .A1(n5418), .A2(n6107), .ZN(n6281) );
  INV_X1 U6887 ( .A(n6281), .ZN(n5419) );
  AND2_X1 U6888 ( .A1(n6300), .A2(n5419), .ZN(n5425) );
  OR2_X1 U6889 ( .A1(n9946), .A2(n9850), .ZN(n5424) );
  INV_X1 U6890 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6891 ( .A1(n6105), .A2(n5420), .ZN(n5423) );
  INV_X1 U6892 ( .A(n5421), .ZN(n7653) );
  NAND2_X1 U6893 ( .A1(n7678), .A2(n7653), .ZN(n5422) );
  NAND2_X1 U6894 ( .A1(n5423), .A2(n5422), .ZN(n6282) );
  AND2_X2 U6895 ( .A1(n5425), .A2(n6020), .ZN(n9968) );
  NAND2_X1 U6896 ( .A1(n6021), .A2(n9968), .ZN(n5428) );
  INV_X1 U6897 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5426) );
  OR2_X1 U6898 ( .A1(n9968), .A2(n5426), .ZN(n5427) );
  NAND2_X1 U6899 ( .A1(n5428), .A2(n5427), .ZN(P1_U3552) );
  NOR2_X2 U6900 ( .A1(n5476), .A2(n5432), .ZN(n5609) );
  NOR2_X1 U6901 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5438) );
  INV_X1 U6902 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5466) );
  INV_X1 U6903 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5437) );
  NAND4_X1 U6904 ( .A1(n5438), .A2(n5466), .A3(n5437), .A4(n5463), .ZN(n5441)
         );
  INV_X1 U6905 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5439) );
  NAND4_X1 U6906 ( .A1(n5465), .A2(n5439), .A3(n5460), .A4(n5950), .ZN(n5440)
         );
  NOR2_X1 U6907 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  INV_X1 U6908 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5443) );
  NOR2_X2 U6909 ( .A1(n5471), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5447) );
  INV_X1 U6910 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5444) );
  INV_X1 U6911 ( .A(n5447), .ZN(n9158) );
  NAND2_X1 U6912 ( .A1(n5544), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5459) );
  INV_X4 U6913 ( .A(n5546), .ZN(n5562) );
  INV_X1 U6914 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6691) );
  OR2_X1 U6915 ( .A1(n5816), .A2(n6691), .ZN(n5458) );
  NAND2_X2 U6916 ( .A1(n7751), .A2(n9163), .ZN(n5574) );
  INV_X1 U6917 ( .A(n5573), .ZN(n5449) );
  INV_X1 U6918 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6919 ( .A1(n5491), .A2(n5452), .ZN(n5453) );
  NAND2_X1 U6920 ( .A1(n5600), .A2(n5453), .ZN(n6882) );
  OR2_X1 U6921 ( .A1(n5574), .A2(n6882), .ZN(n5457) );
  INV_X1 U6922 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5455) );
  OR2_X1 U6923 ( .A1(n5564), .A2(n5455), .ZN(n5456) );
  NAND2_X1 U6924 ( .A1(n5753), .A2(n5460), .ZN(n5769) );
  NOR2_X1 U6925 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5462) );
  NAND2_X1 U6926 ( .A1(n4320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6927 ( .A1(n5467), .A2(n5466), .ZN(n5464) );
  XNOR2_X1 U6928 ( .A(n5467), .B(n5466), .ZN(n5481) );
  NOR2_X1 U6929 ( .A1(n8505), .A2(n5970), .ZN(n5484) );
  INV_X1 U6930 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5468) );
  INV_X1 U6931 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6932 ( .A1(n5540), .A2(n5475), .ZN(n5523) );
  INV_X2 U6934 ( .A(n5807), .ZN(n8205) );
  NAND2_X1 U6935 ( .A1(n8205), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6936 ( .A1(n5476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6937 ( .A1(n5496), .A2(n5430), .ZN(n5477) );
  NAND2_X1 U6938 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U6939 ( .A(n5478), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U6940 ( .A1(n6216), .A2(n6690), .ZN(n5479) );
  OAI211_X1 U6941 ( .C1(n6082), .C2(n5523), .A(n5480), .B(n5479), .ZN(n6879)
         );
  INV_X1 U6942 ( .A(n6879), .ZN(n10004) );
  NAND2_X4 U6943 ( .A1(n5483), .A2(n8212), .ZN(n5894) );
  XNOR2_X1 U6944 ( .A(n10004), .B(n5894), .ZN(n5485) );
  NAND2_X1 U6945 ( .A1(n5484), .A2(n5485), .ZN(n5516) );
  INV_X1 U6946 ( .A(n5484), .ZN(n5486) );
  INV_X1 U6947 ( .A(n5485), .ZN(n6571) );
  NAND2_X1 U6948 ( .A1(n5486), .A2(n6571), .ZN(n5487) );
  NAND2_X1 U6949 ( .A1(n5516), .A2(n5487), .ZN(n6063) );
  INV_X1 U6950 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6693) );
  OR2_X1 U6951 ( .A1(n5816), .A2(n6693), .ZN(n5495) );
  INV_X1 U6952 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5488) );
  OR2_X1 U6953 ( .A1(n5564), .A2(n5488), .ZN(n5494) );
  INV_X1 U6954 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U6955 ( .A1(n5508), .A2(n5489), .ZN(n5490) );
  NAND2_X1 U6956 ( .A1(n5491), .A2(n5490), .ZN(n8504) );
  OR2_X1 U6957 ( .A1(n5574), .A2(n8504), .ZN(n5493) );
  NAND2_X1 U6958 ( .A1(n5544), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5492) );
  NAND2_X2 U6959 ( .A1(n5495), .A2(n4757), .ZN(n8551) );
  NAND2_X1 U6960 ( .A1(n8205), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5498) );
  XNOR2_X1 U6961 ( .A(n5496), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U6962 ( .A1(n6216), .A2(n6692), .ZN(n5497) );
  XNOR2_X1 U6963 ( .A(n6762), .B(n5894), .ZN(n5500) );
  INV_X1 U6964 ( .A(n5500), .ZN(n5499) );
  NAND2_X1 U6965 ( .A1(n5501), .A2(n5499), .ZN(n5596) );
  INV_X1 U6966 ( .A(n5596), .ZN(n5515) );
  XNOR2_X1 U6967 ( .A(n5501), .B(n5500), .ZN(n8499) );
  NAND2_X1 U6968 ( .A1(n8205), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5505) );
  OR2_X1 U6969 ( .A1(n5502), .A2(n5468), .ZN(n5503) );
  XNOR2_X1 U6970 ( .A(n5503), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U6971 ( .A1(n6216), .A2(n6702), .ZN(n5504) );
  OAI211_X1 U6972 ( .C1(n6078), .C2(n5523), .A(n5505), .B(n5504), .ZN(n6751)
         );
  XNOR2_X1 U6973 ( .A(n10001), .B(n5894), .ZN(n5587) );
  INV_X1 U6974 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U6975 ( .A1(n5573), .A2(n5506), .ZN(n5507) );
  NAND2_X1 U6976 ( .A1(n5508), .A2(n5507), .ZN(n6910) );
  NAND2_X1 U6977 ( .A1(n5562), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5513) );
  INV_X1 U6978 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5509) );
  OR2_X1 U6979 ( .A1(n5796), .A2(n5509), .ZN(n5512) );
  INV_X1 U6980 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5510) );
  OR2_X1 U6981 ( .A1(n5564), .A2(n5510), .ZN(n5511) );
  AND2_X1 U6982 ( .A1(n8552), .A2(n8213), .ZN(n5586) );
  NAND2_X1 U6983 ( .A1(n5587), .A2(n5586), .ZN(n5589) );
  AND2_X1 U6984 ( .A1(n8499), .A2(n5589), .ZN(n8500) );
  OR2_X2 U6985 ( .A1(n6063), .A2(n6059), .ZN(n6061) );
  AND2_X1 U6986 ( .A1(n5516), .A2(n6061), .ZN(n5599) );
  NAND2_X1 U6987 ( .A1(n5562), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5519) );
  INV_X1 U6988 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6993) );
  INV_X1 U6989 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6988) );
  OR2_X1 U6990 ( .A1(n5574), .A2(n6988), .ZN(n5518) );
  INV_X1 U6991 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5517) );
  INV_X1 U6992 ( .A(n5527), .ZN(n5525) );
  NAND2_X1 U6993 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5520) );
  XNOR2_X1 U6994 ( .A(n5520), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7232) );
  NAND2_X1 U6995 ( .A1(n6216), .A2(n7232), .ZN(n5521) );
  XNOR2_X1 U6996 ( .A(n5894), .B(n6990), .ZN(n5526) );
  INV_X1 U6997 ( .A(n5526), .ZN(n5524) );
  NAND2_X1 U6998 ( .A1(n5525), .A2(n5524), .ZN(n5528) );
  NAND2_X1 U6999 ( .A1(n5527), .A2(n5526), .ZN(n5543) );
  NAND2_X1 U7000 ( .A1(n5528), .A2(n5543), .ZN(n6460) );
  INV_X1 U7001 ( .A(n6460), .ZN(n5542) );
  NAND2_X1 U7002 ( .A1(n5562), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5535) );
  INV_X1 U7003 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5529) );
  INV_X1 U7004 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5530) );
  INV_X1 U7005 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5531) );
  OR2_X1 U7006 ( .A1(n5564), .A2(n5531), .ZN(n5532) );
  INV_X1 U7007 ( .A(SI_0_), .ZN(n5537) );
  INV_X1 U7008 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5536) );
  OAI21_X1 U7009 ( .B1(n7852), .B2(n5537), .A(n5536), .ZN(n5538) );
  AND2_X1 U7010 ( .A1(n5539), .A2(n5538), .ZN(n9166) );
  MUX2_X1 U7011 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9166), .S(n6667), .Z(n9979) );
  NAND2_X1 U7012 ( .A1(n8557), .A2(n9979), .ZN(n6985) );
  NAND2_X1 U7013 ( .A1(n5542), .A2(n5541), .ZN(n6457) );
  NAND2_X1 U7014 ( .A1(n6457), .A2(n5543), .ZN(n6531) );
  NAND2_X1 U7015 ( .A1(n5544), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5550) );
  INV_X1 U7016 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5545) );
  OR2_X1 U7017 ( .A1(n5564), .A2(n5545), .ZN(n5549) );
  INV_X1 U7018 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7450) );
  OR2_X1 U7019 ( .A1(n5574), .A2(n7450), .ZN(n5548) );
  INV_X1 U7020 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6694) );
  AND4_X2 U7021 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n6827)
         );
  NAND2_X1 U7022 ( .A1(n8555), .A2(n8213), .ZN(n5556) );
  INV_X1 U7023 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U7024 ( .A1(n6216), .A2(n8561), .ZN(n5554) );
  XNOR2_X1 U7025 ( .A(n5894), .B(n6958), .ZN(n5557) );
  XNOR2_X1 U7026 ( .A(n5556), .B(n5557), .ZN(n6530) );
  NAND2_X1 U7027 ( .A1(n8205), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U7028 ( .A1(n5552), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5558) );
  XNOR2_X1 U7029 ( .A(n5558), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7030 ( .A1(n6216), .A2(n6699), .ZN(n5559) );
  XNOR2_X1 U7031 ( .A(n6837), .B(n5894), .ZN(n5571) );
  OR2_X1 U7032 ( .A1(n5574), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7033 ( .A1(n5562), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5567) );
  INV_X1 U7034 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6672) );
  OR2_X1 U7035 ( .A1(n5796), .A2(n6672), .ZN(n5566) );
  INV_X1 U7036 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5563) );
  OR2_X1 U7037 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  NAND4_X1 U7038 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(n8554)
         );
  XNOR2_X1 U7039 ( .A(n5571), .B(n5569), .ZN(n6524) );
  INV_X1 U7040 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7041 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  NAND2_X1 U7042 ( .A1(n5562), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5579) );
  INV_X1 U7043 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6673) );
  OR2_X1 U7044 ( .A1(n5796), .A2(n6673), .ZN(n5578) );
  OAI21_X1 U7045 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5573), .ZN(n7016) );
  OR2_X1 U7046 ( .A1(n5574), .A2(n7016), .ZN(n5577) );
  INV_X1 U7047 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5575) );
  OR2_X1 U7048 ( .A1(n5564), .A2(n5575), .ZN(n5576) );
  NOR2_X1 U7049 ( .A1(n6826), .A2(n5970), .ZN(n5591) );
  NAND2_X1 U7050 ( .A1(n8194), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7051 ( .A1(n5580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5581) );
  XNOR2_X1 U7052 ( .A(n5581), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U7053 ( .A1(n6216), .A2(n8575), .ZN(n5582) );
  OAI211_X1 U7054 ( .C1(n6084), .C2(n5523), .A(n5583), .B(n5582), .ZN(n6658)
         );
  XNOR2_X1 U7055 ( .A(n7017), .B(n5894), .ZN(n5592) );
  AND2_X1 U7056 ( .A1(n5591), .A2(n5592), .ZN(n6504) );
  INV_X1 U7057 ( .A(n6504), .ZN(n5584) );
  NAND2_X1 U7058 ( .A1(n5585), .A2(n5584), .ZN(n6048) );
  INV_X1 U7059 ( .A(n5586), .ZN(n5588) );
  INV_X1 U7060 ( .A(n5587), .ZN(n8510) );
  NAND2_X1 U7061 ( .A1(n5588), .A2(n8510), .ZN(n5590) );
  INV_X1 U7062 ( .A(n6052), .ZN(n5595) );
  INV_X1 U7063 ( .A(n5591), .ZN(n5594) );
  INV_X1 U7064 ( .A(n5592), .ZN(n5593) );
  NAND2_X1 U7065 ( .A1(n5594), .A2(n5593), .ZN(n6503) );
  AND2_X1 U7066 ( .A1(n5595), .A2(n6503), .ZN(n6049) );
  AND2_X1 U7067 ( .A1(n6049), .A2(n5596), .ZN(n6057) );
  INV_X1 U7068 ( .A(n6063), .ZN(n5597) );
  AND2_X1 U7069 ( .A1(n6057), .A2(n5597), .ZN(n5598) );
  NAND2_X1 U7070 ( .A1(n6048), .A2(n5598), .ZN(n6062) );
  NAND2_X1 U7071 ( .A1(n5599), .A2(n6062), .ZN(n5616) );
  NAND2_X1 U7072 ( .A1(n5600), .A2(n7434), .ZN(n5601) );
  NAND2_X1 U7073 ( .A1(n5628), .A2(n5601), .ZN(n6574) );
  OR2_X1 U7074 ( .A1(n5574), .A2(n6574), .ZN(n5607) );
  NAND2_X1 U7075 ( .A1(n5562), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5606) );
  INV_X1 U7076 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5602) );
  OR2_X1 U7077 ( .A1(n5796), .A2(n5602), .ZN(n5605) );
  INV_X1 U7078 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5603) );
  OR2_X1 U7079 ( .A1(n5564), .A2(n5603), .ZN(n5604) );
  NAND4_X1 U7080 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n8549)
         );
  NAND2_X1 U7081 ( .A1(n8549), .A2(n8213), .ZN(n5614) );
  NAND2_X1 U7082 ( .A1(n6089), .A2(n8204), .ZN(n5613) );
  NAND2_X1 U7083 ( .A1(n5617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5610) );
  XNOR2_X1 U7084 ( .A(n5610), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6689) );
  INV_X1 U7085 ( .A(n6689), .ZN(n7115) );
  OAI22_X1 U7086 ( .A1(n5807), .A2(n6092), .B1(n6667), .B2(n7115), .ZN(n5611)
         );
  INV_X1 U7087 ( .A(n5611), .ZN(n5612) );
  XNOR2_X1 U7088 ( .A(n7285), .B(n5894), .ZN(n6619) );
  OR2_X1 U7089 ( .A1(n5614), .A2(n6619), .ZN(n5635) );
  NAND2_X1 U7090 ( .A1(n6619), .A2(n5614), .ZN(n5615) );
  AND2_X1 U7091 ( .A1(n5635), .A2(n5615), .ZN(n6568) );
  NAND2_X1 U7092 ( .A1(n5616), .A2(n6568), .ZN(n6618) );
  NAND2_X1 U7093 ( .A1(n6093), .A2(n8204), .ZN(n5625) );
  NOR2_X1 U7094 ( .A1(n5617), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5621) );
  NOR2_X1 U7095 ( .A1(n5621), .A2(n5468), .ZN(n5618) );
  MUX2_X1 U7096 ( .A(n5468), .B(n5618), .S(P2_IR_REG_9__SCAN_IN), .Z(n5619) );
  INV_X1 U7097 ( .A(n5619), .ZN(n5623) );
  INV_X1 U7098 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5620) );
  INV_X1 U7099 ( .A(n5659), .ZN(n5622) );
  AOI22_X1 U7100 ( .A1(n8194), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6216), .B2(
        n6688), .ZN(n5624) );
  XNOR2_X1 U7101 ( .A(n10011), .B(n5894), .ZN(n5637) );
  INV_X1 U7102 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7103 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  NAND2_X1 U7104 ( .A1(n5645), .A2(n5629), .ZN(n7291) );
  OR2_X1 U7105 ( .A1(n5574), .A2(n7291), .ZN(n5634) );
  NAND2_X1 U7106 ( .A1(n5562), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5633) );
  INV_X1 U7107 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7292) );
  OR2_X1 U7108 ( .A1(n5796), .A2(n7292), .ZN(n5632) );
  INV_X1 U7109 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5630) );
  OR2_X1 U7110 ( .A1(n5564), .A2(n5630), .ZN(n5631) );
  NAND4_X1 U7111 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n8548)
         );
  NAND2_X1 U7112 ( .A1(n8548), .A2(n8213), .ZN(n5638) );
  XNOR2_X1 U7113 ( .A(n5637), .B(n5638), .ZN(n6629) );
  AND2_X1 U7114 ( .A1(n6629), .A2(n5635), .ZN(n5636) );
  INV_X1 U7115 ( .A(n5637), .ZN(n5639) );
  NAND2_X1 U7116 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  NAND2_X1 U7117 ( .A1(n6097), .A2(n8204), .ZN(n5643) );
  OR2_X1 U7118 ( .A1(n5659), .A2(n5468), .ZN(n5641) );
  XNOR2_X1 U7119 ( .A(n5641), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6686) );
  AOI22_X1 U7120 ( .A1(n8205), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6216), .B2(
        n6686), .ZN(n5642) );
  NAND2_X1 U7121 ( .A1(n5643), .A2(n5642), .ZN(n9127) );
  XNOR2_X1 U7122 ( .A(n9127), .B(n5644), .ZN(n5652) );
  NAND2_X1 U7123 ( .A1(n5544), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5651) );
  INV_X1 U7124 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6687) );
  OR2_X1 U7125 ( .A1(n5816), .A2(n6687), .ZN(n5650) );
  INV_X1 U7126 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U7127 ( .A1(n5645), .A2(n7463), .ZN(n5646) );
  NAND2_X1 U7128 ( .A1(n5666), .A2(n5646), .ZN(n7568) );
  OR2_X1 U7129 ( .A1(n5574), .A2(n7568), .ZN(n5649) );
  INV_X1 U7130 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5647) );
  OR2_X1 U7131 ( .A1(n5564), .A2(n5647), .ZN(n5648) );
  NOR2_X1 U7132 ( .A1(n7600), .A2(n5970), .ZN(n5653) );
  NAND2_X1 U7133 ( .A1(n5652), .A2(n5653), .ZN(n5657) );
  INV_X1 U7134 ( .A(n5652), .ZN(n6840) );
  INV_X1 U7135 ( .A(n5653), .ZN(n5654) );
  NAND2_X1 U7136 ( .A1(n6840), .A2(n5654), .ZN(n5655) );
  NAND2_X1 U7137 ( .A1(n5657), .A2(n5655), .ZN(n6919) );
  INV_X1 U7138 ( .A(n6919), .ZN(n5656) );
  NAND2_X1 U7139 ( .A1(n6916), .A2(n5657), .ZN(n5676) );
  NAND2_X1 U7140 ( .A1(n6101), .A2(n8204), .ZN(n5663) );
  INV_X1 U7141 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6104) );
  INV_X1 U7142 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5658) );
  OR2_X1 U7143 ( .A1(n5679), .A2(n5468), .ZN(n5660) );
  INV_X1 U7144 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5678) );
  XNOR2_X1 U7145 ( .A(n5660), .B(n5678), .ZN(n6736) );
  OAI22_X1 U7146 ( .A1(n5807), .A2(n6104), .B1(n6667), .B2(n6736), .ZN(n5661)
         );
  INV_X1 U7147 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7148 ( .A1(n5663), .A2(n5662), .ZN(n8652) );
  XNOR2_X1 U7149 ( .A(n8652), .B(n5644), .ZN(n5672) );
  INV_X1 U7150 ( .A(n5564), .ZN(n5831) );
  NAND2_X1 U7151 ( .A1(n5831), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5671) );
  INV_X1 U7152 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6706) );
  OR2_X1 U7153 ( .A1(n5816), .A2(n6706), .ZN(n5670) );
  INV_X1 U7154 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7604) );
  OR2_X1 U7155 ( .A1(n5796), .A2(n7604), .ZN(n5669) );
  INV_X1 U7156 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7157 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  NAND2_X1 U7158 ( .A1(n5685), .A2(n5667), .ZN(n7603) );
  OR2_X1 U7159 ( .A1(n5574), .A2(n7603), .ZN(n5668) );
  NOR2_X1 U7160 ( .A1(n9013), .A2(n5970), .ZN(n5673) );
  NAND2_X1 U7161 ( .A1(n5672), .A2(n5673), .ZN(n5677) );
  INV_X1 U7162 ( .A(n5672), .ZN(n6999) );
  INV_X1 U7163 ( .A(n5673), .ZN(n5674) );
  NAND2_X1 U7164 ( .A1(n6999), .A2(n5674), .ZN(n5675) );
  AND2_X1 U7165 ( .A1(n5677), .A2(n5675), .ZN(n6838) );
  NAND2_X1 U7166 ( .A1(n5676), .A2(n6838), .ZN(n6841) );
  NAND2_X1 U7167 ( .A1(n6841), .A2(n5677), .ZN(n5695) );
  NAND2_X1 U7168 ( .A1(n6111), .A2(n8204), .ZN(n5683) );
  NAND2_X1 U7169 ( .A1(n5679), .A2(n5678), .ZN(n5697) );
  NAND2_X1 U7170 ( .A1(n5697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  XNOR2_X1 U7171 ( .A(n5680), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7246) );
  INV_X1 U7172 ( .A(n7246), .ZN(n6732) );
  OAI22_X1 U7173 ( .A1(n5807), .A2(n6114), .B1(n6667), .B2(n6732), .ZN(n5681)
         );
  INV_X1 U7174 ( .A(n5681), .ZN(n5682) );
  XNOR2_X1 U7175 ( .A(n9121), .B(n5644), .ZN(n5691) );
  NAND2_X1 U7176 ( .A1(n5831), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5690) );
  INV_X1 U7177 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6731) );
  OR2_X1 U7178 ( .A1(n5816), .A2(n6731), .ZN(n5689) );
  INV_X1 U7179 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5684) );
  OR2_X1 U7180 ( .A1(n5796), .A2(n5684), .ZN(n5688) );
  INV_X1 U7181 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U7182 ( .A1(n5685), .A2(n7237), .ZN(n5686) );
  NAND2_X1 U7183 ( .A1(n5703), .A2(n5686), .ZN(n9004) );
  OR2_X1 U7184 ( .A1(n5574), .A2(n9004), .ZN(n5687) );
  NOR2_X1 U7185 ( .A1(n8978), .A2(n5970), .ZN(n5692) );
  NAND2_X1 U7186 ( .A1(n5691), .A2(n5692), .ZN(n5696) );
  INV_X1 U7187 ( .A(n5691), .ZN(n7176) );
  INV_X1 U7188 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7189 ( .A1(n7176), .A2(n5693), .ZN(n5694) );
  AND2_X1 U7190 ( .A1(n5696), .A2(n5694), .ZN(n6997) );
  NAND2_X1 U7191 ( .A1(n5695), .A2(n6997), .ZN(n7000) );
  NAND2_X1 U7192 ( .A1(n7000), .A2(n5696), .ZN(n5713) );
  NAND2_X1 U7193 ( .A1(n6184), .A2(n8204), .ZN(n5701) );
  OR2_X1 U7194 ( .A1(n5697), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7195 ( .A1(n5698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5715) );
  XNOR2_X1 U7196 ( .A(n5715), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6784) );
  INV_X1 U7197 ( .A(n6784), .ZN(n6780) );
  OAI22_X1 U7198 ( .A1(n5807), .A2(n6185), .B1(n6667), .B2(n6780), .ZN(n5699)
         );
  INV_X1 U7199 ( .A(n5699), .ZN(n5700) );
  XNOR2_X1 U7200 ( .A(n9116), .B(n5644), .ZN(n5709) );
  NAND2_X1 U7201 ( .A1(n5831), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5708) );
  INV_X1 U7202 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6779) );
  OR2_X1 U7203 ( .A1(n5816), .A2(n6779), .ZN(n5707) );
  INV_X1 U7204 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5702) );
  OR2_X1 U7205 ( .A1(n5796), .A2(n5702), .ZN(n5706) );
  INV_X1 U7206 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U7207 ( .A1(n5703), .A2(n6743), .ZN(n5704) );
  NAND2_X1 U7208 ( .A1(n5721), .A2(n5704), .ZN(n8988) );
  OR2_X1 U7209 ( .A1(n5574), .A2(n8988), .ZN(n5705) );
  NOR2_X1 U7210 ( .A1(n9015), .A2(n5970), .ZN(n5710) );
  NAND2_X1 U7211 ( .A1(n5709), .A2(n5710), .ZN(n5727) );
  INV_X1 U7212 ( .A(n5709), .ZN(n7610) );
  INV_X1 U7213 ( .A(n5710), .ZN(n5711) );
  NAND2_X1 U7214 ( .A1(n7610), .A2(n5711), .ZN(n5712) );
  AND2_X1 U7215 ( .A1(n5727), .A2(n5712), .ZN(n7174) );
  NAND2_X1 U7216 ( .A1(n5713), .A2(n7174), .ZN(n7177) );
  NAND2_X1 U7217 ( .A1(n6277), .A2(n8204), .ZN(n5718) );
  INV_X1 U7218 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7219 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  NAND2_X1 U7220 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X1 U7221 ( .A(n5734), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7162) );
  AOI22_X1 U7222 ( .A1(n8205), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6216), .B2(
        n7162), .ZN(n5717) );
  XNOR2_X1 U7223 ( .A(n9111), .B(n5644), .ZN(n5729) );
  NAND2_X1 U7224 ( .A1(n5831), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5726) );
  INV_X1 U7225 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7165) );
  OR2_X1 U7226 ( .A1(n5816), .A2(n7165), .ZN(n5725) );
  INV_X1 U7227 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7228 ( .A1(n5796), .A2(n5719), .ZN(n5724) );
  INV_X1 U7229 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U7230 ( .A1(n5721), .A2(n7474), .ZN(n5722) );
  NAND2_X1 U7231 ( .A1(n5742), .A2(n5722), .ZN(n8956) );
  OR2_X1 U7232 ( .A1(n5574), .A2(n8956), .ZN(n5723) );
  NAND2_X1 U7233 ( .A1(n4646), .A2(n8213), .ZN(n5730) );
  XNOR2_X1 U7234 ( .A(n5729), .B(n5730), .ZN(n7620) );
  AND2_X1 U7235 ( .A1(n7620), .A2(n5727), .ZN(n5728) );
  INV_X1 U7236 ( .A(n5729), .ZN(n5731) );
  NAND2_X1 U7237 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  NAND2_X1 U7238 ( .A1(n7613), .A2(n5732), .ZN(n5750) );
  NAND2_X1 U7239 ( .A1(n6323), .A2(n8204), .ZN(n5738) );
  INV_X1 U7240 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7241 ( .A1(n5734), .A2(n5733), .ZN(n5735) );
  NAND2_X1 U7242 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U7243 ( .A(n5736), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7623) );
  AOI22_X1 U7244 ( .A1(n8194), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7623), .B2(
        n6216), .ZN(n5737) );
  XNOR2_X1 U7245 ( .A(n9106), .B(n5644), .ZN(n5748) );
  XNOR2_X1 U7246 ( .A(n5750), .B(n5748), .ZN(n8533) );
  NAND2_X1 U7247 ( .A1(n5831), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5747) );
  INV_X1 U7248 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5739) );
  OR2_X1 U7249 ( .A1(n5816), .A2(n5739), .ZN(n5746) );
  INV_X1 U7250 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8945) );
  OR2_X1 U7251 ( .A1(n5796), .A2(n8945), .ZN(n5745) );
  INV_X1 U7252 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7253 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NAND2_X1 U7254 ( .A1(n5759), .A2(n5743), .ZN(n8944) );
  OR2_X1 U7255 ( .A1(n5574), .A2(n8944), .ZN(n5744) );
  INV_X1 U7256 ( .A(n8908), .ZN(n8967) );
  NAND2_X1 U7257 ( .A1(n8967), .A2(n8213), .ZN(n8531) );
  NAND2_X1 U7258 ( .A1(n8533), .A2(n8531), .ZN(n5752) );
  INV_X1 U7259 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7260 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U7261 ( .A1(n5752), .A2(n5751), .ZN(n8466) );
  NAND2_X1 U7262 ( .A1(n6372), .A2(n8204), .ZN(n5758) );
  NOR2_X1 U7263 ( .A1(n5753), .A2(n5468), .ZN(n5754) );
  MUX2_X1 U7264 ( .A(n5468), .B(n5754), .S(P2_IR_REG_16__SCAN_IN), .Z(n5755)
         );
  INV_X1 U7265 ( .A(n5755), .ZN(n5756) );
  AND2_X1 U7266 ( .A1(n5756), .A2(n5769), .ZN(n7715) );
  AOI22_X1 U7267 ( .A1(n8194), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6216), .B2(
        n7715), .ZN(n5757) );
  XNOR2_X1 U7268 ( .A(n9097), .B(n5644), .ZN(n5765) );
  NAND2_X1 U7269 ( .A1(n5544), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5764) );
  INV_X1 U7270 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9103) );
  OR2_X1 U7271 ( .A1(n5816), .A2(n9103), .ZN(n5763) );
  INV_X1 U7272 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U7273 ( .A1(n5759), .A2(n7440), .ZN(n5760) );
  NAND2_X1 U7274 ( .A1(n5776), .A2(n5760), .ZN(n8915) );
  OR2_X1 U7275 ( .A1(n5574), .A2(n8915), .ZN(n5762) );
  INV_X1 U7276 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9148) );
  OR2_X1 U7277 ( .A1(n5564), .A2(n9148), .ZN(n5761) );
  NAND2_X1 U7278 ( .A1(n8929), .A2(n8213), .ZN(n5766) );
  XNOR2_X1 U7279 ( .A(n5765), .B(n5766), .ZN(n8467) );
  INV_X1 U7280 ( .A(n5765), .ZN(n5767) );
  NAND2_X1 U7281 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  NAND2_X1 U7282 ( .A1(n6453), .A2(n8204), .ZN(n5774) );
  NAND2_X1 U7283 ( .A1(n5769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5770) );
  MUX2_X1 U7284 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5770), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5771) );
  AND2_X1 U7285 ( .A1(n5771), .A2(n4367), .ZN(n8593) );
  INV_X1 U7286 ( .A(n8593), .ZN(n8588) );
  OAI22_X1 U7287 ( .A1(n5807), .A2(n6454), .B1(n6667), .B2(n8588), .ZN(n5772)
         );
  INV_X1 U7288 ( .A(n5772), .ZN(n5773) );
  XNOR2_X1 U7289 ( .A(n9093), .B(n5644), .ZN(n5784) );
  INV_X1 U7290 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U7291 ( .A1(n5776), .A2(n7713), .ZN(n5777) );
  NAND2_X1 U7292 ( .A1(n5793), .A2(n5777), .ZN(n8890) );
  OR2_X1 U7293 ( .A1(n5574), .A2(n8890), .ZN(n5783) );
  NAND2_X1 U7294 ( .A1(n5562), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5782) );
  INV_X1 U7295 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7296 ( .A1(n5796), .A2(n5778), .ZN(n5781) );
  INV_X1 U7297 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7298 ( .A1(n5564), .A2(n5779), .ZN(n5780) );
  NAND4_X1 U7299 ( .A1(n5783), .A2(n5782), .A3(n5781), .A4(n5780), .ZN(n8906)
         );
  AND2_X1 U7300 ( .A1(n8906), .A2(n8213), .ZN(n5785) );
  NAND2_X1 U7301 ( .A1(n5784), .A2(n5785), .ZN(n5788) );
  INV_X1 U7302 ( .A(n5784), .ZN(n8490) );
  INV_X1 U7303 ( .A(n5785), .ZN(n5786) );
  NAND2_X1 U7304 ( .A1(n8490), .A2(n5786), .ZN(n5787) );
  NAND2_X1 U7305 ( .A1(n5788), .A2(n5787), .ZN(n6042) );
  NAND2_X1 U7306 ( .A1(n6491), .A2(n8204), .ZN(n5792) );
  INV_X1 U7307 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7308 ( .A1(n4367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5789) );
  XNOR2_X1 U7309 ( .A(n5789), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8594) );
  INV_X1 U7310 ( .A(n8594), .ZN(n8609) );
  OAI22_X1 U7311 ( .A1(n5807), .A2(n6492), .B1(n6667), .B2(n8609), .ZN(n5790)
         );
  INV_X1 U7312 ( .A(n5790), .ZN(n5791) );
  XNOR2_X1 U7313 ( .A(n9087), .B(n5644), .ZN(n5802) );
  NAND2_X1 U7314 ( .A1(n5562), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5801) );
  INV_X1 U7315 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U7316 ( .A1(n5793), .A2(n8493), .ZN(n5794) );
  AND2_X1 U7317 ( .A1(n5813), .A2(n5794), .ZN(n8861) );
  NAND2_X1 U7318 ( .A1(n5924), .A2(n8861), .ZN(n5800) );
  INV_X1 U7319 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5795) );
  OR2_X1 U7320 ( .A1(n5796), .A2(n5795), .ZN(n5799) );
  INV_X1 U7321 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5797) );
  OR2_X1 U7322 ( .A1(n5564), .A2(n5797), .ZN(n5798) );
  NAND4_X1 U7323 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n8879)
         );
  AND2_X1 U7324 ( .A1(n8879), .A2(n8213), .ZN(n5803) );
  NAND2_X1 U7325 ( .A1(n5802), .A2(n5803), .ZN(n5821) );
  INV_X1 U7326 ( .A(n5802), .ZN(n8435) );
  INV_X1 U7327 ( .A(n5803), .ZN(n5804) );
  NAND2_X1 U7328 ( .A1(n8435), .A2(n5804), .ZN(n5805) );
  NAND2_X1 U7329 ( .A1(n5806), .A2(n8488), .ZN(n8434) );
  NAND2_X1 U7330 ( .A1(n6548), .A2(n8204), .ZN(n5810) );
  OAI22_X1 U7331 ( .A1(n5807), .A2(n8404), .B1(n6667), .B2(n8888), .ZN(n5808)
         );
  INV_X1 U7332 ( .A(n5808), .ZN(n5809) );
  XNOR2_X1 U7333 ( .A(n9083), .B(n5644), .ZN(n5823) );
  INV_X1 U7334 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7335 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7336 ( .A1(n5829), .A2(n5814), .ZN(n8852) );
  NOR2_X1 U7337 ( .A1(n8852), .A2(n5574), .ZN(n5820) );
  INV_X1 U7338 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5815) );
  INV_X1 U7339 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8606) );
  OAI22_X1 U7340 ( .A1(n5816), .A2(n5815), .B1(n5796), .B2(n8606), .ZN(n5819)
         );
  INV_X1 U7341 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5817) );
  NOR2_X1 U7342 ( .A1(n5564), .A2(n5817), .ZN(n5818) );
  NAND2_X1 U7343 ( .A1(n8868), .A2(n8213), .ZN(n5824) );
  XNOR2_X1 U7344 ( .A(n5823), .B(n5824), .ZN(n8443) );
  AND2_X1 U7345 ( .A1(n8443), .A2(n5821), .ZN(n5822) );
  INV_X1 U7346 ( .A(n5823), .ZN(n5825) );
  NAND2_X1 U7347 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  NAND2_X1 U7348 ( .A1(n6631), .A2(n8204), .ZN(n5828) );
  NAND2_X1 U7349 ( .A1(n8205), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5827) );
  XNOR2_X1 U7350 ( .A(n9077), .B(n5644), .ZN(n5835) );
  INV_X1 U7351 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7478) );
  NAND2_X1 U7352 ( .A1(n5829), .A2(n7478), .ZN(n5830) );
  AND2_X1 U7353 ( .A1(n5856), .A2(n5830), .ZN(n8831) );
  NAND2_X1 U7354 ( .A1(n8831), .A2(n5924), .ZN(n5834) );
  AOI22_X1 U7355 ( .A1(n5562), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5544), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7356 ( .A1(n5831), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5832) );
  NOR2_X1 U7357 ( .A1(n8690), .A2(n5970), .ZN(n5836) );
  NAND2_X1 U7358 ( .A1(n5835), .A2(n5836), .ZN(n5840) );
  INV_X1 U7359 ( .A(n5835), .ZN(n8448) );
  INV_X1 U7360 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7361 ( .A1(n8448), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U7362 ( .A1(n5840), .A2(n5838), .ZN(n8475) );
  NAND2_X1 U7363 ( .A1(n8445), .A2(n5840), .ZN(n5847) );
  NAND2_X1 U7364 ( .A1(n6718), .A2(n8204), .ZN(n5842) );
  NAND2_X1 U7365 ( .A1(n8194), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7366 ( .A(n8819), .B(n5644), .ZN(n5848) );
  XNOR2_X1 U7367 ( .A(n5856), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8817) );
  INV_X1 U7368 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7369 ( .A1(n5562), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7370 ( .A1(n5544), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5843) );
  OAI211_X1 U7371 ( .C1(n5845), .C2(n5564), .A(n5844), .B(n5843), .ZN(n5846)
         );
  AOI21_X1 U7372 ( .B1(n8817), .B2(n5924), .A(n5846), .ZN(n8691) );
  NOR2_X1 U7373 ( .A1(n8691), .A2(n5970), .ZN(n5849) );
  XNOR2_X1 U7374 ( .A(n5848), .B(n5849), .ZN(n8446) );
  NAND2_X1 U7375 ( .A1(n5847), .A2(n8446), .ZN(n8449) );
  INV_X1 U7376 ( .A(n5848), .ZN(n5850) );
  NAND2_X1 U7377 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  NAND2_X1 U7378 ( .A1(n6888), .A2(n8204), .ZN(n5853) );
  NAND2_X1 U7379 ( .A1(n8205), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7380 ( .A(n9067), .B(n5894), .ZN(n5862) );
  NAND2_X1 U7381 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5854) );
  INV_X1 U7382 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7498) );
  INV_X1 U7383 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5855) );
  OAI21_X1 U7384 ( .B1(n5856), .B2(n7498), .A(n5855), .ZN(n5857) );
  AND2_X1 U7385 ( .A1(n5875), .A2(n5857), .ZN(n8804) );
  INV_X1 U7386 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7387 ( .A1(n5562), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7388 ( .A1(n5544), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U7389 ( .C1(n5860), .C2(n5564), .A(n5859), .B(n5858), .ZN(n5861)
         );
  AOI21_X1 U7390 ( .B1(n8804), .B2(n5924), .A(n5861), .ZN(n8693) );
  OR2_X1 U7391 ( .A1(n8693), .A2(n5970), .ZN(n8480) );
  INV_X1 U7392 ( .A(n5862), .ZN(n5863) );
  AOI21_X2 U7393 ( .B1(n8481), .B2(n8480), .A(n5865), .ZN(n5887) );
  NAND2_X1 U7394 ( .A1(n7090), .A2(n8204), .ZN(n5867) );
  NAND2_X1 U7395 ( .A1(n8205), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U7396 ( .A(n9062), .B(n5894), .ZN(n5885) );
  XNOR2_X1 U7397 ( .A(n5887), .B(n5885), .ZN(n6000) );
  NAND2_X1 U7398 ( .A1(n7538), .A2(n8204), .ZN(n5869) );
  NAND2_X1 U7399 ( .A1(n8194), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5868) );
  XNOR2_X1 U7400 ( .A(n9057), .B(n5644), .ZN(n5889) );
  XNOR2_X1 U7401 ( .A(n5895), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8772) );
  INV_X1 U7402 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7403 ( .A1(n5562), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7404 ( .A1(n5544), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5871) );
  OAI211_X1 U7405 ( .C1(n5873), .C2(n5564), .A(n5872), .B(n5871), .ZN(n5874)
         );
  AOI21_X1 U7406 ( .B1(n8772), .B2(n5924), .A(n5874), .ZN(n8459) );
  INV_X1 U7407 ( .A(n8459), .ZN(n8796) );
  INV_X1 U7408 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U7409 ( .A1(n5875), .A2(n8427), .ZN(n5876) );
  AND2_X1 U7410 ( .A1(n5895), .A2(n5876), .ZN(n8791) );
  NAND2_X1 U7411 ( .A1(n8791), .A2(n5924), .ZN(n5882) );
  INV_X1 U7412 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7413 ( .A1(n5562), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7414 ( .A1(n5544), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5877) );
  OAI211_X1 U7415 ( .C1(n5879), .C2(n5564), .A(n5878), .B(n5877), .ZN(n5880)
         );
  INV_X1 U7416 ( .A(n5880), .ZN(n5881) );
  NOR2_X1 U7417 ( .A1(n8780), .A2(n5970), .ZN(n6001) );
  NAND2_X1 U7418 ( .A1(n6000), .A2(n5884), .ZN(n5891) );
  OR2_X1 U7419 ( .A1(n8459), .A2(n5970), .ZN(n6005) );
  INV_X1 U7420 ( .A(n6005), .ZN(n5888) );
  INV_X1 U7421 ( .A(n5885), .ZN(n5886) );
  OAI21_X1 U7422 ( .B1(n5888), .B2(n5889), .A(n6002), .ZN(n5890) );
  INV_X1 U7423 ( .A(n5889), .ZN(n6003) );
  NAND2_X1 U7424 ( .A1(n7651), .A2(n8204), .ZN(n5893) );
  NAND2_X1 U7425 ( .A1(n8205), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U7426 ( .A(n9053), .B(n5894), .ZN(n8517) );
  INV_X1 U7427 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6009) );
  INV_X1 U7428 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8461) );
  OAI21_X1 U7429 ( .B1(n5895), .B2(n6009), .A(n8461), .ZN(n5896) );
  AND2_X1 U7430 ( .A1(n5896), .A2(n5908), .ZN(n8764) );
  NAND2_X1 U7431 ( .A1(n8764), .A2(n5924), .ZN(n5902) );
  INV_X1 U7432 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7433 ( .A1(n5562), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7434 ( .A1(n5544), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5897) );
  OAI211_X1 U7435 ( .C1(n5899), .C2(n5564), .A(n5898), .B(n5897), .ZN(n5900)
         );
  INV_X1 U7436 ( .A(n5900), .ZN(n5901) );
  INV_X1 U7437 ( .A(n8781), .ZN(n8695) );
  NAND2_X1 U7438 ( .A1(n8695), .A2(n8213), .ZN(n5903) );
  NOR2_X1 U7439 ( .A1(n8517), .A2(n5903), .ZN(n5904) );
  AOI21_X1 U7440 ( .B1(n8517), .B2(n5903), .A(n5904), .ZN(n8457) );
  NAND2_X1 U7441 ( .A1(n7676), .A2(n8204), .ZN(n5906) );
  NAND2_X1 U7442 ( .A1(n8205), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7443 ( .A(n9048), .B(n5644), .ZN(n5916) );
  INV_X1 U7444 ( .A(n5908), .ZN(n5907) );
  NAND2_X1 U7445 ( .A1(n5907), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5922) );
  INV_X1 U7446 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U7447 ( .A1(n5908), .A2(n8522), .ZN(n5909) );
  NAND2_X1 U7448 ( .A1(n5922), .A2(n5909), .ZN(n8740) );
  OR2_X1 U7449 ( .A1(n8740), .A2(n5574), .ZN(n5915) );
  INV_X1 U7450 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7451 ( .A1(n5562), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7452 ( .A1(n5544), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5910) );
  OAI211_X1 U7453 ( .C1(n5912), .C2(n5564), .A(n5911), .B(n5910), .ZN(n5913)
         );
  INV_X1 U7454 ( .A(n5913), .ZN(n5914) );
  NOR2_X1 U7455 ( .A1(n8546), .A2(n5970), .ZN(n5917) );
  NAND2_X1 U7456 ( .A1(n5916), .A2(n5917), .ZN(n5972) );
  INV_X1 U7457 ( .A(n5916), .ZN(n5971) );
  INV_X1 U7458 ( .A(n5917), .ZN(n5918) );
  NAND2_X1 U7459 ( .A1(n5971), .A2(n5918), .ZN(n5919) );
  NAND2_X1 U7460 ( .A1(n5972), .A2(n5919), .ZN(n8519) );
  NAND2_X1 U7461 ( .A1(n7679), .A2(n8204), .ZN(n5921) );
  NAND2_X1 U7462 ( .A1(n8194), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7463 ( .A(n9042), .B(n5644), .ZN(n5931) );
  INV_X1 U7464 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7371) );
  NAND2_X1 U7465 ( .A1(n5922), .A2(n7371), .ZN(n5923) );
  NAND2_X1 U7466 ( .A1(n8732), .A2(n5924), .ZN(n5930) );
  INV_X1 U7467 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7468 ( .A1(n5562), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7469 ( .A1(n5544), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5925) );
  OAI211_X1 U7470 ( .C1(n5927), .C2(n5564), .A(n5926), .B(n5925), .ZN(n5928)
         );
  INV_X1 U7471 ( .A(n5928), .ZN(n5929) );
  NOR2_X1 U7472 ( .A1(n8545), .A2(n5970), .ZN(n5932) );
  NAND2_X1 U7473 ( .A1(n5931), .A2(n5932), .ZN(n7766) );
  INV_X1 U7474 ( .A(n5931), .ZN(n5934) );
  INV_X1 U7475 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7476 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  INV_X1 U7477 ( .A(n5973), .ZN(n5969) );
  NOR4_X1 U7478 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5939) );
  NOR4_X1 U7479 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5938) );
  NOR4_X1 U7480 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5937) );
  NOR4_X1 U7481 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5936) );
  NAND4_X1 U7482 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n5958)
         );
  NOR2_X1 U7483 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5943) );
  NOR4_X1 U7484 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5942) );
  NOR4_X1 U7485 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5941) );
  NOR4_X1 U7486 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5940) );
  NAND4_X1 U7487 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n5957)
         );
  NAND2_X1 U7488 ( .A1(n5944), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5945) );
  MUX2_X1 U7489 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5945), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5946) );
  NAND2_X1 U7490 ( .A1(n5946), .A2(n4378), .ZN(n7656) );
  NAND2_X1 U7491 ( .A1(n5947), .A2(n5463), .ZN(n5948) );
  NAND2_X1 U7492 ( .A1(n5948), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  INV_X1 U7493 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7494 ( .A1(n5963), .A2(n5962), .ZN(n5949) );
  NAND2_X1 U7495 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7496 ( .A(n7580), .B(P2_B_REG_SCAN_IN), .ZN(n5952) );
  NAND2_X1 U7497 ( .A1(n4378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5953) );
  MUX2_X1 U7498 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5953), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5955) );
  NAND2_X1 U7499 ( .A1(n5955), .A2(n5954), .ZN(n7687) );
  OAI21_X1 U7500 ( .B1(n5958), .B2(n5957), .A(n9969), .ZN(n6499) );
  INV_X1 U7501 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U7502 ( .A1(n9969), .A2(n9976), .ZN(n5959) );
  NAND2_X1 U7503 ( .A1(n7687), .A2(n7656), .ZN(n9974) );
  NAND2_X1 U7504 ( .A1(n5959), .A2(n9974), .ZN(n6467) );
  INV_X1 U7505 ( .A(n6467), .ZN(n5960) );
  AND2_X1 U7506 ( .A1(n7580), .A2(n7687), .ZN(n9973) );
  INV_X1 U7507 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9972) );
  AND2_X1 U7508 ( .A1(n9969), .A2(n9972), .ZN(n5961) );
  XNOR2_X1 U7509 ( .A(n5963), .B(n5962), .ZN(n6215) );
  AND2_X1 U7510 ( .A1(n6816), .A2(n9971), .ZN(n5964) );
  AND2_X1 U7511 ( .A1(n8361), .A2(n8888), .ZN(n5982) );
  INV_X1 U7512 ( .A(n5982), .ZN(n5966) );
  AND2_X2 U7513 ( .A1(n5965), .A2(n5966), .ZN(n9992) );
  NAND2_X1 U7514 ( .A1(n5967), .A2(n5482), .ZN(n6661) );
  INV_X1 U7515 ( .A(n6661), .ZN(n6217) );
  NOR2_X1 U7516 ( .A1(n9992), .A2(n6217), .ZN(n5968) );
  AOI21_X1 U7517 ( .B1(n4334), .B2(n5969), .A(n8518), .ZN(n5975) );
  NOR3_X1 U7518 ( .A1(n5971), .A2(n8546), .A3(n8516), .ZN(n5974) );
  OAI21_X1 U7519 ( .B1(n5975), .B2(n5974), .A(n7767), .ZN(n5999) );
  NOR2_X1 U7520 ( .A1(n5976), .A2(n8361), .ZN(n6819) );
  NAND2_X1 U7521 ( .A1(n5983), .A2(n6819), .ZN(n5978) );
  NAND2_X1 U7522 ( .A1(n8361), .A2(n8623), .ZN(n8389) );
  OR2_X1 U7523 ( .A1(n5976), .A2(n8389), .ZN(n6468) );
  INV_X1 U7524 ( .A(n6468), .ZN(n5977) );
  NAND2_X1 U7525 ( .A1(n6818), .A2(n6816), .ZN(n5979) );
  NAND2_X1 U7526 ( .A1(n5979), .A2(n6468), .ZN(n6463) );
  OR2_X1 U7527 ( .A1(n6661), .A2(n5982), .ZN(n6461) );
  AND3_X1 U7528 ( .A1(n6663), .A2(n6215), .A3(n6461), .ZN(n5980) );
  NAND2_X1 U7529 ( .A1(n6463), .A2(n5980), .ZN(n5981) );
  NAND2_X1 U7530 ( .A1(n5981), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8537) );
  INV_X1 U7531 ( .A(n8537), .ZN(n8526) );
  INV_X1 U7532 ( .A(n5984), .ZN(n6662) );
  NAND2_X1 U7533 ( .A1(n8460), .A2(n8965), .ZN(n8536) );
  NOR2_X1 U7534 ( .A1(n8536), .A2(n8546), .ZN(n5995) );
  NAND2_X1 U7535 ( .A1(n6217), .A2(n5984), .ZN(n9014) );
  NAND2_X1 U7536 ( .A1(n8460), .A2(n8968), .ZN(n8539) );
  INV_X1 U7537 ( .A(n5986), .ZN(n5985) );
  NAND2_X1 U7538 ( .A1(n5985), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8703) );
  INV_X1 U7539 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U7540 ( .A1(n5986), .A2(n7775), .ZN(n5987) );
  NAND2_X1 U7541 ( .A1(n8703), .A2(n5987), .ZN(n8718) );
  OR2_X1 U7542 ( .A1(n8718), .A2(n5574), .ZN(n5993) );
  INV_X1 U7543 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7544 ( .A1(n5562), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7545 ( .A1(n5544), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5988) );
  OAI211_X1 U7546 ( .C1(n5990), .C2(n5564), .A(n5989), .B(n5988), .ZN(n5991)
         );
  INV_X1 U7547 ( .A(n5991), .ZN(n5992) );
  OAI22_X1 U7548 ( .A1(n8539), .A2(n8188), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7371), .ZN(n5994) );
  AOI211_X1 U7549 ( .C1(n8526), .C2(n8732), .A(n5995), .B(n5994), .ZN(n5996)
         );
  INV_X1 U7550 ( .A(n5997), .ZN(n5998) );
  AND2_X1 U7551 ( .A1(n6000), .A2(n6001), .ZN(n8432) );
  NOR2_X1 U7552 ( .A1(n8432), .A2(n6002), .ZN(n6004) );
  XNOR2_X1 U7553 ( .A(n6004), .B(n6003), .ZN(n6006) );
  OAI22_X1 U7554 ( .A1(n6006), .A2(n8518), .B1(n8459), .B2(n8516), .ZN(n6008)
         );
  INV_X1 U7555 ( .A(n9057), .ZN(n8774) );
  NOR2_X1 U7556 ( .A1(n8536), .A2(n8780), .ZN(n6011) );
  OAI22_X1 U7557 ( .A1(n8539), .A2(n8781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6009), .ZN(n6010) );
  AOI211_X1 U7558 ( .C1(n8526), .C2(n8772), .A(n6011), .B(n6010), .ZN(n6012)
         );
  NAND2_X1 U7559 ( .A1(n6015), .A2(n6014), .ZN(P2_U3231) );
  INV_X1 U7560 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7561 ( .A1(n6105), .A2(n6110), .ZN(n6018) );
  INV_X1 U7562 ( .A(n6016), .ZN(n6017) );
  AOI22_X1 U7563 ( .A1(n6018), .A2(n6107), .B1(n6105), .B2(n6017), .ZN(n6019)
         );
  AND2_X1 U7564 ( .A1(n6300), .A2(n6019), .ZN(n6024) );
  AND2_X2 U7565 ( .A1(n6024), .A2(n6020), .ZN(n9952) );
  NAND2_X1 U7566 ( .A1(n6021), .A2(n9952), .ZN(n6023) );
  NAND2_X1 U7567 ( .A1(n6023), .A2(n4745), .ZN(P1_U3520) );
  INV_X1 U7568 ( .A(n6282), .ZN(n9887) );
  NAND2_X1 U7569 ( .A1(n6024), .A2(n9887), .ZN(n6721) );
  NAND2_X1 U7570 ( .A1(n9889), .A2(n9867), .ZN(n6025) );
  OR2_X1 U7571 ( .A1(n6027), .A2(n6284), .ZN(n8083) );
  AND2_X1 U7572 ( .A1(n6381), .A2(n8083), .ZN(n9833) );
  NAND2_X1 U7573 ( .A1(n9884), .A2(n9833), .ZN(n9855) );
  AND2_X1 U7574 ( .A1(n9884), .A2(n9850), .ZN(n9535) );
  INV_X1 U7575 ( .A(n8029), .ZN(n8034) );
  OR2_X1 U7576 ( .A1(n6366), .A2(n6029), .ZN(n9881) );
  INV_X1 U7577 ( .A(n9881), .ZN(n9828) );
  NAND2_X1 U7578 ( .A1(n9884), .A2(n9828), .ZN(n9539) );
  INV_X1 U7579 ( .A(n9880), .ZN(n9826) );
  AOI22_X1 U7580 ( .A1(n9856), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n6030), .B2(
        n9826), .ZN(n6031) );
  OAI21_X1 U7581 ( .B1(n8034), .B2(n9539), .A(n6031), .ZN(n6032) );
  OR2_X1 U7582 ( .A1(n6036), .A2(n6035), .ZN(P1_U3355) );
  INV_X1 U7583 ( .A(n6441), .ZN(n7091) );
  NOR2_X1 U7584 ( .A1(n6442), .A2(n7091), .ZN(n9759) );
  AND2_X2 U7585 ( .A1(n9759), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U7586 ( .A(n6663), .ZN(n6037) );
  NAND2_X1 U7587 ( .A1(n8042), .A2(n6442), .ZN(n6038) );
  NAND2_X1 U7588 ( .A1(n6038), .A2(n6441), .ZN(n6120) );
  NAND2_X1 U7589 ( .A1(n6120), .A2(n6039), .ZN(n9737) );
  NAND2_X1 U7590 ( .A1(n9737), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7591 ( .A(n6040), .ZN(n6041) );
  AOI211_X1 U7592 ( .C1(n6043), .C2(n6042), .A(n8518), .B(n6041), .ZN(n6047)
         );
  INV_X1 U7593 ( .A(n9093), .ZN(n8685) );
  NOR2_X1 U7594 ( .A1(n8685), .A2(n8544), .ZN(n6046) );
  INV_X1 U7595 ( .A(n8879), .ZN(n8687) );
  OAI22_X1 U7596 ( .A1(n8539), .A2(n8687), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7713), .ZN(n6045) );
  OAI22_X1 U7597 ( .A1(n8536), .A2(n8538), .B1(n8537), .B2(n8890), .ZN(n6044)
         );
  OR4_X1 U7598 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(P2_U3230)
         );
  NAND2_X1 U7599 ( .A1(n6058), .A2(n6503), .ZN(n6051) );
  NAND2_X1 U7600 ( .A1(n6058), .A2(n6049), .ZN(n8502) );
  INV_X1 U7601 ( .A(n8502), .ZN(n6050) );
  AOI211_X1 U7602 ( .C1(n6052), .C2(n6051), .A(n8518), .B(n6050), .ZN(n6056)
         );
  NOR2_X1 U7603 ( .A1(n8537), .A2(n6910), .ZN(n6055) );
  OAI22_X1 U7604 ( .A1(n6826), .A2(n8536), .B1(n8539), .B2(n6878), .ZN(n6054)
         );
  OAI22_X1 U7605 ( .A1(n8544), .A2(n10001), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5506), .ZN(n6053) );
  OR4_X1 U7606 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(P2_U3229)
         );
  NAND2_X1 U7607 ( .A1(n6058), .A2(n6057), .ZN(n6060) );
  AND2_X1 U7608 ( .A1(n6060), .A2(n6059), .ZN(n6064) );
  NAND2_X1 U7609 ( .A1(n6062), .A2(n6061), .ZN(n6567) );
  AOI211_X1 U7610 ( .C1(n6064), .C2(n6063), .A(n8518), .B(n6567), .ZN(n6068)
         );
  NOR2_X1 U7611 ( .A1(n8537), .A2(n6882), .ZN(n6067) );
  INV_X1 U7612 ( .A(n8549), .ZN(n7287) );
  OAI22_X1 U7613 ( .A1(n7287), .A2(n8539), .B1(n8536), .B2(n6878), .ZN(n6066)
         );
  OAI22_X1 U7614 ( .A1(n8544), .A2(n10004), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5452), .ZN(n6065) );
  OR4_X1 U7615 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(P2_U3215)
         );
  XNOR2_X1 U7616 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U7617 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7618 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n9731) );
  OAI21_X1 U7619 ( .B1(n6070), .B2(P1_STATE_REG_SCAN_IN), .A(n9731), .ZN(
        P1_U3353) );
  OR2_X1 U7620 ( .A1(n7852), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9667) );
  NAND2_X1 U7621 ( .A1(n7852), .A2(P1_U3084), .ZN(n9665) );
  OAI222_X1 U7622 ( .A1(n9667), .A2(n6071), .B1(n9665), .B2(n6075), .C1(n6312), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  AND2_X1 U7623 ( .A1(n7852), .A2(P2_U3152), .ZN(n9162) );
  INV_X1 U7624 ( .A(n9162), .ZN(n8405) );
  INV_X1 U7625 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6072) );
  INV_X1 U7626 ( .A(n6699), .ZN(n6803) );
  OAI222_X1 U7627 ( .A1(n8405), .A2(n6072), .B1(n9165), .B2(n4332), .C1(
        P2_U3152), .C2(n6803), .ZN(P2_U3355) );
  INV_X1 U7628 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6073) );
  INV_X1 U7629 ( .A(n8561), .ZN(n6671) );
  OAI222_X1 U7630 ( .A1(n8405), .A2(n6073), .B1(n9165), .B2(n6086), .C1(
        P2_U3152), .C2(n6671), .ZN(P2_U3356) );
  INV_X1 U7631 ( .A(n8575), .ZN(n8574) );
  OAI222_X1 U7632 ( .A1(n8405), .A2(n4813), .B1(n9165), .B2(n6084), .C1(
        P2_U3152), .C2(n8574), .ZN(P2_U3354) );
  INV_X1 U7633 ( .A(n6692), .ZN(n7126) );
  OAI222_X1 U7634 ( .A1(n8405), .A2(n6074), .B1(n9165), .B2(n6080), .C1(
        P2_U3152), .C2(n7126), .ZN(P2_U3352) );
  INV_X1 U7635 ( .A(n6702), .ZN(n6815) );
  OAI222_X1 U7636 ( .A1(n8405), .A2(n4826), .B1(n9165), .B2(n6078), .C1(
        P2_U3152), .C2(n6815), .ZN(P2_U3353) );
  INV_X1 U7637 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6076) );
  INV_X1 U7638 ( .A(n7232), .ZN(n6670) );
  OAI222_X1 U7639 ( .A1(n8405), .A2(n6076), .B1(n9165), .B2(n6075), .C1(
        P2_U3152), .C2(n6670), .ZN(P2_U3357) );
  INV_X1 U7640 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6077) );
  INV_X1 U7641 ( .A(n6690), .ZN(n7150) );
  OAI222_X1 U7642 ( .A1(n8405), .A2(n6077), .B1(n9165), .B2(n6082), .C1(
        P2_U3152), .C2(n7150), .ZN(P2_U3351) );
  INV_X1 U7643 ( .A(n9665), .ZN(n7748) );
  INV_X1 U7644 ( .A(n7748), .ZN(n9671) );
  OAI222_X1 U7645 ( .A1(n9667), .A2(n6079), .B1(n9671), .B2(n6078), .C1(n6194), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  OAI222_X1 U7646 ( .A1(n9667), .A2(n6081), .B1(n9671), .B2(n6080), .C1(n6274), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  OAI222_X1 U7647 ( .A1(n9667), .A2(n6083), .B1(n9671), .B2(n6082), .C1(n6207), 
        .C2(P1_U3084), .ZN(P1_U3346) );
  OAI222_X1 U7648 ( .A1(n9667), .A2(n6085), .B1(n9671), .B2(n6084), .C1(n9778), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  INV_X1 U7649 ( .A(n9667), .ZN(n7681) );
  INV_X1 U7650 ( .A(n7681), .ZN(n7753) );
  OAI222_X1 U7651 ( .A1(n7753), .A2(n6087), .B1(n9671), .B2(n6086), .C1(n9754), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  OAI222_X1 U7652 ( .A1(n7753), .A2(n6088), .B1(n9671), .B2(n4332), .C1(n6148), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U7653 ( .A(n6089), .ZN(n6091) );
  OAI222_X1 U7654 ( .A1(n6180), .A2(P1_U3084), .B1(n9665), .B2(n6091), .C1(
        n6090), .C2(n7753), .ZN(P1_U3345) );
  OAI222_X1 U7655 ( .A1(n8405), .A2(n6092), .B1(n9165), .B2(n6091), .C1(
        P2_U3152), .C2(n7115), .ZN(P2_U3350) );
  INV_X1 U7656 ( .A(n6093), .ZN(n6096) );
  INV_X1 U7657 ( .A(n6688), .ZN(n7138) );
  OAI222_X1 U7658 ( .A1(n8405), .A2(n6094), .B1(n9165), .B2(n6096), .C1(n7138), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U7659 ( .A1(P1_U3084), .A2(n6245), .B1(n9665), .B2(n6096), .C1(
        n6095), .C2(n9667), .ZN(P1_U3344) );
  INV_X1 U7660 ( .A(n6224), .ZN(n6257) );
  INV_X1 U7661 ( .A(n6097), .ZN(n6099) );
  OAI222_X1 U7662 ( .A1(P1_U3084), .A2(n6257), .B1(n9665), .B2(n6099), .C1(
        n6098), .C2(n9667), .ZN(P1_U3343) );
  INV_X1 U7663 ( .A(n6686), .ZN(n7103) );
  OAI222_X1 U7664 ( .A1(n8405), .A2(n6100), .B1(n9165), .B2(n6099), .C1(n7103), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7665 ( .A(n6234), .ZN(n6339) );
  INV_X1 U7666 ( .A(n6101), .ZN(n6103) );
  INV_X1 U7667 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6102) );
  OAI222_X1 U7668 ( .A1(P1_U3084), .A2(n6339), .B1(n9665), .B2(n6103), .C1(
        n6102), .C2(n7753), .ZN(P1_U3342) );
  OAI222_X1 U7669 ( .A1(n8405), .A2(n6104), .B1(n9165), .B2(n6103), .C1(n6736), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7670 ( .A(n6105), .ZN(n6106) );
  NAND2_X1 U7671 ( .A1(n6106), .A2(n9889), .ZN(n9886) );
  INV_X1 U7672 ( .A(n9886), .ZN(n6108) );
  OAI21_X1 U7673 ( .B1(n6108), .B2(P1_D_REG_0__SCAN_IN), .A(n6107), .ZN(n6109)
         );
  OAI21_X1 U7674 ( .B1(n9889), .B2(n6110), .A(n6109), .ZN(P1_U3440) );
  INV_X1 U7675 ( .A(n6335), .ZN(n6357) );
  INV_X1 U7676 ( .A(n6111), .ZN(n6113) );
  OAI222_X1 U7677 ( .A1(n6357), .A2(P1_U3084), .B1(n9665), .B2(n6113), .C1(
        n6112), .C2(n9667), .ZN(P1_U3341) );
  OAI222_X1 U7678 ( .A1(n8405), .A2(n6114), .B1(n9165), .B2(n6113), .C1(
        P2_U3152), .C2(n6732), .ZN(P2_U3346) );
  INV_X1 U7679 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6140) );
  OR2_X1 U7680 ( .A1(P1_U3083), .A2(n9759), .ZN(n9782) );
  NOR2_X1 U7681 ( .A1(n9755), .A2(P1_U3084), .ZN(n7680) );
  NAND2_X1 U7682 ( .A1(n6120), .A2(n7680), .ZN(n9299) );
  AND2_X1 U7683 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6449) );
  INV_X1 U7684 ( .A(n6449), .ZN(n6124) );
  INV_X1 U7685 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9957) );
  MUX2_X1 U7686 ( .A(n9957), .B(P1_REG1_REG_3__SCAN_IN), .S(n6148), .Z(n6122)
         );
  INV_X1 U7687 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U7688 ( .A(n9953), .B(P1_REG1_REG_1__SCAN_IN), .S(n6312), .Z(n6305)
         );
  NAND2_X1 U7689 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6306) );
  INV_X1 U7690 ( .A(n6306), .ZN(n6115) );
  NAND2_X1 U7691 ( .A1(n6305), .A2(n6115), .ZN(n6309) );
  INV_X1 U7692 ( .A(n6312), .ZN(n6319) );
  NAND2_X1 U7693 ( .A1(n6319), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7694 ( .A1(n6309), .A2(n6116), .ZN(n9750) );
  XNOR2_X1 U7695 ( .A(n9754), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U7696 ( .A1(n9750), .A2(n9751), .ZN(n9749) );
  INV_X1 U7697 ( .A(n9754), .ZN(n6132) );
  NAND2_X1 U7698 ( .A1(n6132), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7699 ( .A1(n9749), .A2(n6117), .ZN(n6121) );
  OR2_X1 U7700 ( .A1(n4312), .A2(P1_U3084), .ZN(n9730) );
  INV_X1 U7701 ( .A(n9755), .ZN(n6118) );
  NOR2_X1 U7702 ( .A1(n9730), .A2(n6118), .ZN(n6119) );
  NAND2_X1 U7703 ( .A1(n6121), .A2(n6122), .ZN(n6164) );
  OAI211_X1 U7704 ( .C1(n6122), .C2(n6121), .A(n9813), .B(n6164), .ZN(n6123)
         );
  OAI211_X1 U7705 ( .C1(n9808), .C2(n6148), .A(n6124), .B(n6123), .ZN(n6125)
         );
  INV_X1 U7706 ( .A(n6125), .ZN(n6139) );
  INV_X1 U7707 ( .A(n9299), .ZN(n6126) );
  INV_X1 U7708 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6127) );
  MUX2_X1 U7709 ( .A(n6127), .B(P1_REG2_REG_2__SCAN_IN), .S(n9754), .Z(n6131)
         );
  INV_X1 U7710 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6128) );
  MUX2_X1 U7711 ( .A(n6128), .B(P1_REG2_REG_1__SCAN_IN), .S(n6312), .Z(n6129)
         );
  AND2_X1 U7712 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6311) );
  NAND2_X1 U7713 ( .A1(n6129), .A2(n6311), .ZN(n6313) );
  OR2_X1 U7714 ( .A1(n6312), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7715 ( .A1(n6313), .A2(n6130), .ZN(n9744) );
  NAND2_X1 U7716 ( .A1(n6131), .A2(n9744), .ZN(n9745) );
  NAND2_X1 U7717 ( .A1(n6132), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7718 ( .A1(n9745), .A2(n6135), .ZN(n6134) );
  INV_X1 U7719 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6542) );
  MUX2_X1 U7720 ( .A(n6542), .B(P1_REG2_REG_3__SCAN_IN), .S(n6148), .Z(n6133)
         );
  NAND2_X1 U7721 ( .A1(n6134), .A2(n6133), .ZN(n6150) );
  MUX2_X1 U7722 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6542), .S(n6148), .Z(n6136)
         );
  NAND3_X1 U7723 ( .A1(n6136), .A2(n9745), .A3(n6135), .ZN(n6137) );
  NAND3_X1 U7724 ( .A1(n9817), .A2(n6150), .A3(n6137), .ZN(n6138) );
  OAI211_X1 U7725 ( .C1(n6140), .C2(n9782), .A(n6139), .B(n6138), .ZN(P1_U3244) );
  INV_X1 U7726 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6145) );
  INV_X1 U7727 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7728 ( .A1(n5562), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6142) );
  INV_X1 U7729 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8635) );
  OR2_X1 U7730 ( .A1(n5796), .A2(n8635), .ZN(n6141) );
  OAI211_X1 U7731 ( .C1(n5564), .C2(n6143), .A(n6142), .B(n6141), .ZN(n8634)
         );
  NAND2_X1 U7732 ( .A1(n8634), .A2(P2_U3966), .ZN(n6144) );
  OAI21_X1 U7733 ( .B1(n6145), .B2(P2_U3966), .A(n6144), .ZN(P2_U3583) );
  NOR2_X1 U7734 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6160), .ZN(n6155) );
  INV_X1 U7735 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6146) );
  MUX2_X1 U7736 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6146), .S(n6160), .Z(n6147)
         );
  INV_X1 U7737 ( .A(n6147), .ZN(n6210) );
  INV_X1 U7738 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6154) );
  NOR2_X1 U7739 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6167), .ZN(n6153) );
  INV_X1 U7740 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6151) );
  INV_X1 U7741 ( .A(n6148), .ZN(n6162) );
  NAND2_X1 U7742 ( .A1(n6162), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6149) );
  AND2_X1 U7743 ( .A1(n6150), .A2(n6149), .ZN(n9769) );
  MUX2_X1 U7744 ( .A(n6151), .B(P1_REG2_REG_4__SCAN_IN), .S(n9778), .Z(n9768)
         );
  AND2_X1 U7745 ( .A1(n9769), .A2(n9768), .ZN(n9766) );
  AOI21_X1 U7746 ( .B1(n6151), .B2(n9778), .A(n9766), .ZN(n6197) );
  INV_X1 U7747 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6152) );
  MUX2_X1 U7748 ( .A(n6152), .B(P1_REG2_REG_5__SCAN_IN), .S(n6167), .Z(n6196)
         );
  NOR2_X1 U7749 ( .A1(n6197), .A2(n6196), .ZN(n6195) );
  NOR2_X1 U7750 ( .A1(n6153), .A2(n6195), .ZN(n6267) );
  MUX2_X1 U7751 ( .A(n6154), .B(P1_REG2_REG_6__SCAN_IN), .S(n6274), .Z(n6266)
         );
  NAND2_X1 U7752 ( .A1(n6267), .A2(n6266), .ZN(n6265) );
  OAI21_X1 U7753 ( .B1(n6274), .B2(n6154), .A(n6265), .ZN(n6209) );
  NOR2_X1 U7754 ( .A1(n6210), .A2(n6209), .ZN(n6208) );
  NOR2_X1 U7755 ( .A1(n6155), .A2(n6208), .ZN(n6158) );
  INV_X1 U7756 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6156) );
  AOI22_X1 U7757 ( .A1(n6228), .A2(n6156), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6180), .ZN(n6157) );
  NOR2_X1 U7758 ( .A1(n6158), .A2(n6157), .ZN(n6229) );
  AOI21_X1 U7759 ( .B1(n6158), .B2(n6157), .A(n6229), .ZN(n6183) );
  INV_X1 U7760 ( .A(n9817), .ZN(n6314) );
  INV_X1 U7761 ( .A(n9782), .ZN(n9811) );
  NAND2_X1 U7762 ( .A1(n6228), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7763 ( .A1(n6160), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6170) );
  NOR2_X1 U7764 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6160), .ZN(n6159) );
  AOI21_X1 U7765 ( .B1(n6160), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6159), .ZN(
        n6204) );
  INV_X1 U7766 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7767 ( .A1(n6274), .A2(n6168), .ZN(n6169) );
  NAND2_X1 U7768 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6167), .ZN(n6161) );
  OAI21_X1 U7769 ( .B1(n6167), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6161), .ZN(
        n6189) );
  NAND2_X1 U7770 ( .A1(n6162), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6163) );
  AND2_X1 U7771 ( .A1(n6164), .A2(n6163), .ZN(n9773) );
  INV_X1 U7772 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6165) );
  MUX2_X1 U7773 ( .A(n6165), .B(P1_REG1_REG_4__SCAN_IN), .S(n9778), .Z(n9772)
         );
  NAND2_X1 U7774 ( .A1(n9773), .A2(n9772), .ZN(n9771) );
  NAND2_X1 U7775 ( .A1(n9778), .A2(n6165), .ZN(n6166) );
  NAND2_X1 U7776 ( .A1(n9771), .A2(n6166), .ZN(n6190) );
  NOR2_X1 U7777 ( .A1(n6189), .A2(n6190), .ZN(n6188) );
  AOI21_X1 U7778 ( .B1(n6167), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6188), .ZN(
        n6269) );
  MUX2_X1 U7779 ( .A(n6168), .B(P1_REG1_REG_6__SCAN_IN), .S(n6274), .Z(n6270)
         );
  NAND2_X1 U7780 ( .A1(n6269), .A2(n6270), .ZN(n6268) );
  NAND2_X1 U7781 ( .A1(n6169), .A2(n6268), .ZN(n6203) );
  NAND2_X1 U7782 ( .A1(n6204), .A2(n6203), .ZN(n6202) );
  NAND2_X1 U7783 ( .A1(n6170), .A2(n6202), .ZN(n6175) );
  NAND2_X1 U7784 ( .A1(n6174), .A2(n6175), .ZN(n6171) );
  OR2_X1 U7785 ( .A1(n6228), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6172) );
  INV_X1 U7786 ( .A(n6175), .ZN(n6173) );
  NOR2_X1 U7787 ( .A1(n6173), .A2(n6172), .ZN(n6176) );
  OAI22_X1 U7788 ( .A1(n6244), .A2(n6176), .B1(n6175), .B2(n6174), .ZN(n6178)
         );
  INV_X1 U7789 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6177) );
  NOR2_X1 U7790 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6177), .ZN(n6872) );
  AOI21_X1 U7791 ( .B1(n9813), .B2(n6178), .A(n6872), .ZN(n6179) );
  OAI21_X1 U7792 ( .B1(n6180), .B2(n9808), .A(n6179), .ZN(n6181) );
  AOI21_X1 U7793 ( .B1(n9811), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6181), .ZN(
        n6182) );
  OAI21_X1 U7794 ( .B1(n6183), .B2(n6314), .A(n6182), .ZN(P1_U3249) );
  INV_X1 U7795 ( .A(n6184), .ZN(n6187) );
  OAI222_X1 U7796 ( .A1(n8405), .A2(n6185), .B1(n9165), .B2(n6187), .C1(n6780), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7797 ( .A(n6341), .ZN(n6417) );
  OAI222_X1 U7798 ( .A1(P1_U3084), .A2(n6417), .B1(n9665), .B2(n6187), .C1(
        n6186), .C2(n9667), .ZN(P1_U3340) );
  AOI21_X1 U7799 ( .B1(n6190), .B2(n6189), .A(n6188), .ZN(n6192) );
  INV_X1 U7800 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6191) );
  NOR2_X1 U7801 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6191), .ZN(n6772) );
  AOI21_X1 U7802 ( .B1(n9813), .B2(n6192), .A(n6772), .ZN(n6193) );
  OAI21_X1 U7803 ( .B1(n6194), .B2(n9808), .A(n6193), .ZN(n6200) );
  AOI21_X1 U7804 ( .B1(n6197), .B2(n6196), .A(n6195), .ZN(n6198) );
  NOR2_X1 U7805 ( .A1(n6314), .A2(n6198), .ZN(n6199) );
  AOI211_X1 U7806 ( .C1(P1_ADDR_REG_5__SCAN_IN), .C2(n9811), .A(n6200), .B(
        n6199), .ZN(n6201) );
  INV_X1 U7807 ( .A(n6201), .ZN(P1_U3246) );
  OAI21_X1 U7808 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(n6205) );
  AND2_X1 U7809 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6614) );
  AOI21_X1 U7810 ( .B1(n9813), .B2(n6205), .A(n6614), .ZN(n6206) );
  OAI21_X1 U7811 ( .B1(n6207), .B2(n9808), .A(n6206), .ZN(n6213) );
  AOI21_X1 U7812 ( .B1(n6210), .B2(n6209), .A(n6208), .ZN(n6211) );
  NOR2_X1 U7813 ( .A1(n6314), .A2(n6211), .ZN(n6212) );
  AOI211_X1 U7814 ( .C1(P1_ADDR_REG_7__SCAN_IN), .C2(n9811), .A(n6213), .B(
        n6212), .ZN(n6214) );
  INV_X1 U7815 ( .A(n6214), .ZN(P1_U3248) );
  OR2_X1 U7816 ( .A1(n6215), .A2(P2_U3152), .ZN(n8402) );
  INV_X1 U7817 ( .A(n8402), .ZN(n7028) );
  OAI21_X1 U7818 ( .B1(n9971), .B2(n7028), .A(n6216), .ZN(n6219) );
  NAND2_X1 U7819 ( .A1(n9971), .A2(n6217), .ZN(n6218) );
  NOR2_X1 U7820 ( .A1(n8599), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7821 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9678) );
  NOR2_X1 U7822 ( .A1(n6227), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6220) );
  INV_X1 U7823 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7310) );
  AOI22_X1 U7824 ( .A1(n6227), .A2(n7310), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6245), .ZN(n6243) );
  NOR2_X1 U7825 ( .A1(n6244), .A2(n6243), .ZN(n6242) );
  NOR2_X1 U7826 ( .A1(n6220), .A2(n6242), .ZN(n6255) );
  AOI22_X1 U7827 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6257), .B1(n6224), .B2(
        n9678), .ZN(n6254) );
  NOR2_X1 U7828 ( .A1(n6255), .A2(n6254), .ZN(n6253) );
  AOI21_X1 U7829 ( .B1(n9678), .B2(n6257), .A(n6253), .ZN(n6222) );
  INV_X1 U7830 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7650) );
  AOI22_X1 U7831 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6339), .B1(n6234), .B2(
        n7650), .ZN(n6221) );
  NOR2_X1 U7832 ( .A1(n6222), .A2(n6221), .ZN(n6331) );
  AOI21_X1 U7833 ( .B1(n6222), .B2(n6221), .A(n6331), .ZN(n6241) );
  INV_X1 U7834 ( .A(n9813), .ZN(n7059) );
  AND2_X1 U7835 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7279) );
  NOR2_X1 U7836 ( .A1(n9808), .A2(n6339), .ZN(n6223) );
  AOI211_X1 U7837 ( .C1(n9811), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7279), .B(
        n6223), .ZN(n6240) );
  NAND2_X1 U7838 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6224), .ZN(n6233) );
  INV_X1 U7839 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6225) );
  MUX2_X1 U7840 ( .A(n6225), .B(P1_REG2_REG_10__SCAN_IN), .S(n6224), .Z(n6226)
         );
  INV_X1 U7841 ( .A(n6226), .ZN(n6260) );
  NAND2_X1 U7842 ( .A1(n6227), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U7843 ( .A1(n6228), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6230) );
  NOR2_X1 U7844 ( .A1(n6230), .A2(n6229), .ZN(n6249) );
  INV_X1 U7845 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6231) );
  MUX2_X1 U7846 ( .A(n6231), .B(P1_REG2_REG_9__SCAN_IN), .S(n6245), .Z(n6248)
         );
  NAND2_X1 U7847 ( .A1(n6249), .A2(n6248), .ZN(n6247) );
  NAND2_X1 U7848 ( .A1(n6232), .A2(n6247), .ZN(n6261) );
  NAND2_X1 U7849 ( .A1(n6260), .A2(n6261), .ZN(n6259) );
  NAND2_X1 U7850 ( .A1(n6233), .A2(n6259), .ZN(n6236) );
  INV_X1 U7851 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6235) );
  MUX2_X1 U7852 ( .A(n6235), .B(P1_REG2_REG_11__SCAN_IN), .S(n6234), .Z(n6237)
         );
  AND2_X1 U7853 ( .A1(n6236), .A2(n6237), .ZN(n6238) );
  NOR2_X1 U7854 ( .A1(n6237), .A2(n6236), .ZN(n6338) );
  OAI21_X1 U7855 ( .B1(n6238), .B2(n6338), .A(n9817), .ZN(n6239) );
  OAI211_X1 U7856 ( .C1(n6241), .C2(n7059), .A(n6240), .B(n6239), .ZN(P1_U3252) );
  AOI21_X1 U7857 ( .B1(n6244), .B2(n6243), .A(n6242), .ZN(n6252) );
  AND2_X1 U7858 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7157) );
  NOR2_X1 U7859 ( .A1(n9808), .A2(n6245), .ZN(n6246) );
  AOI211_X1 U7860 ( .C1(n9811), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7157), .B(
        n6246), .ZN(n6251) );
  OAI211_X1 U7861 ( .C1(n6249), .C2(n6248), .A(n9817), .B(n6247), .ZN(n6250)
         );
  OAI211_X1 U7862 ( .C1(n6252), .C2(n7059), .A(n6251), .B(n6250), .ZN(P1_U3250) );
  AOI21_X1 U7863 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(n6264) );
  NOR2_X1 U7864 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6256), .ZN(n7086) );
  NOR2_X1 U7865 ( .A1(n9808), .A2(n6257), .ZN(n6258) );
  AOI211_X1 U7866 ( .C1(n9811), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n7086), .B(
        n6258), .ZN(n6263) );
  OAI211_X1 U7867 ( .C1(n6261), .C2(n6260), .A(n9817), .B(n6259), .ZN(n6262)
         );
  OAI211_X1 U7868 ( .C1(n6264), .C2(n7059), .A(n6263), .B(n6262), .ZN(P1_U3251) );
  OAI211_X1 U7869 ( .C1(n6267), .C2(n6266), .A(n9817), .B(n6265), .ZN(n6273)
         );
  OAI21_X1 U7870 ( .B1(n6270), .B2(n6269), .A(n6268), .ZN(n6271) );
  AND2_X1 U7871 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6933) );
  AOI21_X1 U7872 ( .B1(n9813), .B2(n6271), .A(n6933), .ZN(n6272) );
  OAI211_X1 U7873 ( .C1(n9808), .C2(n6274), .A(n6273), .B(n6272), .ZN(n6275)
         );
  AOI21_X1 U7874 ( .B1(n9811), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6275), .ZN(
        n6276) );
  INV_X1 U7875 ( .A(n6276), .ZN(P1_U3247) );
  INV_X1 U7876 ( .A(n6277), .ZN(n6280) );
  INV_X1 U7877 ( .A(n7162), .ZN(n7166) );
  OAI222_X1 U7878 ( .A1(n8405), .A2(n6278), .B1(n9165), .B2(n6280), .C1(n7166), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7879 ( .A(n7048), .ZN(n7033) );
  OAI222_X1 U7880 ( .A1(P1_U3084), .A2(n7033), .B1(n9665), .B2(n6280), .C1(
        n6279), .C2(n7753), .ZN(P1_U3339) );
  NAND2_X1 U7881 ( .A1(n9881), .A2(n8083), .ZN(n6283) );
  OR2_X1 U7882 ( .A1(n6282), .A2(n6281), .ZN(n6438) );
  NAND3_X1 U7883 ( .A1(n6283), .A2(n6438), .A3(n9889), .ZN(n6445) );
  AND2_X1 U7884 ( .A1(n6445), .A2(n6300), .ZN(n9693) );
  NAND2_X1 U7885 ( .A1(n9693), .A2(n9913), .ZN(n9224) );
  AND2_X2 U7886 ( .A1(n6286), .A2(n6442), .ZN(n6395) );
  NAND2_X1 U7887 ( .A1(n9860), .A2(n6395), .ZN(n6288) );
  INV_X1 U7888 ( .A(n6442), .ZN(n6293) );
  NAND2_X1 U7889 ( .A1(n6293), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7890 ( .A1(n6292), .A2(n6395), .ZN(n6295) );
  NAND2_X1 U7891 ( .A1(n6293), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6294) );
  OAI211_X1 U7892 ( .C1(n6367), .C2(n7186), .A(n6295), .B(n6294), .ZN(n6374)
         );
  NAND2_X1 U7893 ( .A1(n6296), .A2(n6374), .ZN(n6376) );
  OAI21_X1 U7894 ( .B1(n6296), .B2(n6374), .A(n6376), .ZN(n9756) );
  INV_X1 U7895 ( .A(n9889), .ZN(n8082) );
  NOR2_X1 U7896 ( .A1(n6438), .A2(n8082), .ZN(n6297) );
  AND2_X1 U7897 ( .A1(n9898), .A2(n8042), .ZN(n6439) );
  INV_X1 U7898 ( .A(n6297), .ZN(n6298) );
  OR2_X1 U7899 ( .A1(n6298), .A2(n8083), .ZN(n6388) );
  AOI22_X1 U7900 ( .A1(n9756), .A2(n9694), .B1(n9222), .B2(n9291), .ZN(n6304)
         );
  INV_X1 U7901 ( .A(n6300), .ZN(n6301) );
  OAI21_X1 U7902 ( .B1(n6438), .B2(n6301), .A(n9224), .ZN(n6413) );
  INV_X1 U7903 ( .A(n6413), .ZN(n6302) );
  NAND2_X1 U7904 ( .A1(n6302), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6303) );
  OAI211_X1 U7905 ( .C1(n9224), .C2(n6367), .A(n6304), .B(n6303), .ZN(P1_U3230) );
  INV_X1 U7906 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6322) );
  INV_X1 U7907 ( .A(n9808), .ZN(n6320) );
  INV_X1 U7908 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9879) );
  INV_X1 U7909 ( .A(n6305), .ZN(n6307) );
  NAND2_X1 U7910 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  NAND3_X1 U7911 ( .A1(n9813), .A2(n6309), .A3(n6308), .ZN(n6310) );
  OAI21_X1 U7912 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9879), .A(n6310), .ZN(n6318) );
  INV_X1 U7913 ( .A(n6311), .ZN(n9757) );
  MUX2_X1 U7914 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6128), .S(n6312), .Z(n6316)
         );
  INV_X1 U7915 ( .A(n6313), .ZN(n6315) );
  AOI211_X1 U7916 ( .C1(n9757), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6317)
         );
  AOI211_X1 U7917 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n6317), .ZN(n6321)
         );
  OAI21_X1 U7918 ( .B1(n9782), .B2(n6322), .A(n6321), .ZN(P1_U3242) );
  INV_X1 U7919 ( .A(n6323), .ZN(n6361) );
  AOI22_X1 U7920 ( .A1(n9784), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7681), .ZN(n6324) );
  OAI21_X1 U7921 ( .B1(n6361), .B2(n9665), .A(n6324), .ZN(P1_U3338) );
  INV_X1 U7922 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7923 ( .A1(n6325), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7924 ( .A1(n5236), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7925 ( .A1(n5328), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6326) );
  NAND3_X1 U7926 ( .A1(n6328), .A2(n6327), .A3(n6326), .ZN(n9309) );
  NAND2_X1 U7927 ( .A1(n9309), .A2(P1_U4006), .ZN(n6329) );
  OAI21_X1 U7928 ( .B1(P1_U4006), .B2(n6330), .A(n6329), .ZN(P1_U3586) );
  INV_X1 U7929 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9724) );
  AOI21_X1 U7930 ( .B1(n7650), .B2(n6339), .A(n6331), .ZN(n6351) );
  AOI22_X1 U7931 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6357), .B1(n6335), .B2(
        n9724), .ZN(n6350) );
  NOR2_X1 U7932 ( .A1(n6351), .A2(n6350), .ZN(n6349) );
  AOI21_X1 U7933 ( .B1(n9724), .B2(n6357), .A(n6349), .ZN(n6333) );
  INV_X1 U7934 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6418) );
  AOI22_X1 U7935 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n6417), .B1(n6341), .B2(
        n6418), .ZN(n6332) );
  NOR2_X1 U7936 ( .A1(n6333), .A2(n6332), .ZN(n6416) );
  AOI21_X1 U7937 ( .B1(n6333), .B2(n6332), .A(n6416), .ZN(n6348) );
  AND2_X1 U7938 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7216) );
  NOR2_X1 U7939 ( .A1(n9808), .A2(n6417), .ZN(n6334) );
  AOI211_X1 U7940 ( .C1(n9811), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7216), .B(
        n6334), .ZN(n6347) );
  NAND2_X1 U7941 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6335), .ZN(n6340) );
  INV_X1 U7942 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6337) );
  INV_X1 U7943 ( .A(n6340), .ZN(n6336) );
  AOI21_X1 U7944 ( .B1(n6337), .B2(n6357), .A(n6336), .ZN(n6353) );
  AOI21_X1 U7945 ( .B1(n6339), .B2(n6235), .A(n6338), .ZN(n6354) );
  NAND2_X1 U7946 ( .A1(n6353), .A2(n6354), .ZN(n6352) );
  NAND2_X1 U7947 ( .A1(n6340), .A2(n6352), .ZN(n6345) );
  INV_X1 U7948 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7949 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6341), .ZN(n6424) );
  INV_X1 U7950 ( .A(n6424), .ZN(n6342) );
  AOI21_X1 U7951 ( .B1(n6343), .B2(n6417), .A(n6342), .ZN(n6344) );
  NAND2_X1 U7952 ( .A1(n6344), .A2(n6345), .ZN(n6423) );
  OAI211_X1 U7953 ( .C1(n6345), .C2(n6344), .A(n9817), .B(n6423), .ZN(n6346)
         );
  OAI211_X1 U7954 ( .C1(n6348), .C2(n7059), .A(n6347), .B(n6346), .ZN(P1_U3254) );
  AOI21_X1 U7955 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n6360) );
  OAI211_X1 U7956 ( .C1(n6354), .C2(n6353), .A(n9817), .B(n6352), .ZN(n6356)
         );
  NAND2_X1 U7957 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6355) );
  OAI211_X1 U7958 ( .C1(n9808), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6358)
         );
  AOI21_X1 U7959 ( .B1(n9811), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n6358), .ZN(
        n6359) );
  OAI21_X1 U7960 ( .B1(n6360), .B2(n7059), .A(n6359), .ZN(P1_U3253) );
  INV_X1 U7961 ( .A(n7623), .ZN(n7629) );
  OAI222_X1 U7962 ( .A1(n8405), .A2(n6362), .B1(n9165), .B2(n6361), .C1(
        P2_U3152), .C2(n7629), .ZN(P2_U3343) );
  INV_X1 U7963 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6369) );
  AND2_X1 U7964 ( .A1(n6367), .A2(n6292), .ZN(n8049) );
  NOR2_X1 U7965 ( .A1(n9869), .A2(n8049), .ZN(n7868) );
  INV_X1 U7966 ( .A(n8083), .ZN(n6364) );
  INV_X1 U7967 ( .A(n6366), .ZN(n6363) );
  NOR3_X1 U7968 ( .A1(n7868), .A2(n6364), .A3(n6363), .ZN(n6365) );
  AOI21_X1 U7969 ( .B1(n9873), .B2(n9291), .A(n6365), .ZN(n6552) );
  OAI21_X1 U7970 ( .B1(n6367), .B2(n6366), .A(n6552), .ZN(n6370) );
  NAND2_X1 U7971 ( .A1(n6370), .A2(n9952), .ZN(n6368) );
  OAI21_X1 U7972 ( .B1(n9952), .B2(n6369), .A(n6368), .ZN(P1_U3454) );
  INV_X1 U7973 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U7974 ( .A1(n6370), .A2(n9968), .ZN(n6371) );
  OAI21_X1 U7975 ( .B1(n9968), .B2(n9740), .A(n6371), .ZN(P1_U3523) );
  INV_X1 U7976 ( .A(n6372), .ZN(n6414) );
  AOI22_X1 U7977 ( .A1(n7715), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9162), .ZN(n6373) );
  OAI21_X1 U7978 ( .B1(n6414), .B2(n9165), .A(n6373), .ZN(P2_U3342) );
  INV_X1 U7979 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U7980 ( .A1(n6375), .A2(n6381), .ZN(n6377) );
  NAND2_X1 U7981 ( .A1(n9291), .A2(n6395), .ZN(n6380) );
  NAND2_X1 U7982 ( .A1(n6378), .A2(n8155), .ZN(n6379) );
  NAND2_X1 U7983 ( .A1(n6380), .A2(n6379), .ZN(n6382) );
  NAND2_X1 U7984 ( .A1(n6384), .A2(n6383), .ZN(n6403) );
  INV_X1 U7985 ( .A(n6383), .ZN(n6386) );
  INV_X1 U7986 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U7987 ( .A1(n6386), .A2(n6385), .ZN(n6404) );
  NAND2_X1 U7988 ( .A1(n6403), .A2(n6404), .ZN(n6387) );
  BUF_X8 U7989 ( .A(n6395), .Z(n8412) );
  AOI22_X1 U7990 ( .A1(n9291), .A2(n8411), .B1(n6378), .B2(n8412), .ZN(n6402)
         );
  XNOR2_X1 U7991 ( .A(n6387), .B(n6402), .ZN(n6393) );
  INV_X1 U7992 ( .A(n6292), .ZN(n6389) );
  OR2_X1 U7993 ( .A1(n6388), .A2(n4312), .ZN(n9271) );
  OAI22_X1 U7994 ( .A1(n6389), .A2(n9271), .B1(n9682), .B2(n4444), .ZN(n6391)
         );
  NOR2_X1 U7995 ( .A1(n6413), .A2(n9879), .ZN(n6390) );
  AOI211_X1 U7996 ( .C1(n9276), .C2(n6378), .A(n6391), .B(n6390), .ZN(n6392)
         );
  OAI21_X1 U7997 ( .B1(n6393), .B2(n9278), .A(n6392), .ZN(P1_U3220) );
  INV_X1 U7998 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7999 ( .A1(n6394), .A2(n8155), .ZN(n6397) );
  NAND2_X1 U8000 ( .A1(n9874), .A2(n6395), .ZN(n6396) );
  NAND2_X1 U8001 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  XNOR2_X1 U8002 ( .A(n6398), .B(n4311), .ZN(n6400) );
  AOI22_X1 U8003 ( .A1(n9874), .A2(n8411), .B1(n6394), .B2(n8412), .ZN(n6399)
         );
  NAND2_X1 U8004 ( .A1(n6400), .A2(n6399), .ZN(n6429) );
  NAND2_X1 U8005 ( .A1(n6403), .A2(n6402), .ZN(n6405) );
  NAND2_X1 U8006 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U8007 ( .A1(n6406), .A2(n4746), .ZN(n6430) );
  OAI21_X1 U8008 ( .B1(n4746), .B2(n6406), .A(n6430), .ZN(n6407) );
  NAND2_X1 U8009 ( .A1(n6407), .A2(n9694), .ZN(n6412) );
  INV_X1 U8010 ( .A(n9291), .ZN(n6409) );
  INV_X1 U8011 ( .A(n9290), .ZN(n6408) );
  OAI22_X1 U8012 ( .A1(n6409), .A2(n9271), .B1(n9682), .B2(n6408), .ZN(n6410)
         );
  AOI21_X1 U8013 ( .B1(n9276), .B2(n6394), .A(n6410), .ZN(n6411) );
  OAI211_X1 U8014 ( .C1(n6413), .C2(n6641), .A(n6412), .B(n6411), .ZN(P1_U3235) );
  INV_X1 U8015 ( .A(n7044), .ZN(n9795) );
  OAI222_X1 U8016 ( .A1(n9667), .A2(n6415), .B1(n9665), .B2(n6414), .C1(
        P1_U3084), .C2(n9795), .ZN(P1_U3337) );
  AOI21_X1 U8017 ( .B1(n6418), .B2(n6417), .A(n6416), .ZN(n6420) );
  INV_X1 U8018 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9718) );
  AOI22_X1 U8019 ( .A1(n7048), .A2(n9718), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n7033), .ZN(n6419) );
  NOR2_X1 U8020 ( .A1(n6420), .A2(n6419), .ZN(n7032) );
  AOI21_X1 U8021 ( .B1(n6420), .B2(n6419), .A(n7032), .ZN(n6428) );
  NOR2_X1 U8022 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6421), .ZN(n7554) );
  NOR2_X1 U8023 ( .A1(n9808), .A2(n7033), .ZN(n6422) );
  AOI211_X1 U8024 ( .C1(n9811), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7554), .B(
        n6422), .ZN(n6427) );
  NAND2_X1 U8025 ( .A1(n6424), .A2(n6423), .ZN(n7047) );
  XNOR2_X1 U8026 ( .A(n7047), .B(n7033), .ZN(n6425) );
  NAND2_X1 U8027 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n6425), .ZN(n7049) );
  OAI211_X1 U8028 ( .C1(n6425), .C2(P1_REG2_REG_14__SCAN_IN), .A(n9817), .B(
        n7049), .ZN(n6426) );
  OAI211_X1 U8029 ( .C1(n6428), .C2(n7059), .A(n6427), .B(n6426), .ZN(P1_U3255) );
  NAND2_X1 U8030 ( .A1(n6430), .A2(n6429), .ZN(n6581) );
  NAND2_X1 U8031 ( .A1(n9290), .A2(n8412), .ZN(n6432) );
  NAND2_X1 U8032 ( .A1(n9905), .A2(n8406), .ZN(n6431) );
  NAND2_X1 U8033 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  XNOR2_X1 U8034 ( .A(n6433), .B(n4311), .ZN(n6435) );
  AOI22_X1 U8035 ( .A1(n9290), .A2(n8411), .B1(n9905), .B2(n8412), .ZN(n6434)
         );
  AND2_X1 U8036 ( .A1(n6435), .A2(n6434), .ZN(n6580) );
  INV_X1 U8037 ( .A(n6580), .ZN(n6436) );
  OR2_X1 U8038 ( .A1(n6435), .A2(n6434), .ZN(n6579) );
  NAND2_X1 U8039 ( .A1(n6436), .A2(n6579), .ZN(n6437) );
  XNOR2_X1 U8040 ( .A(n6581), .B(n6437), .ZN(n6452) );
  NAND2_X1 U8041 ( .A1(n6439), .A2(n6438), .ZN(n6443) );
  NAND4_X1 U8042 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n6444)
         );
  NAND2_X1 U8043 ( .A1(n6444), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6446) );
  INV_X1 U8044 ( .A(n9699), .ZN(n9259) );
  INV_X1 U8045 ( .A(n9271), .ZN(n9685) );
  AOI22_X1 U8046 ( .A1(n9259), .A2(n6447), .B1(n9685), .B2(n9874), .ZN(n6451)
         );
  NOR2_X1 U8047 ( .A1(n9224), .A2(n6544), .ZN(n6448) );
  AOI211_X1 U8048 ( .C1(n9222), .C2(n9845), .A(n6449), .B(n6448), .ZN(n6450)
         );
  OAI211_X1 U8049 ( .C1(n6452), .C2(n9278), .A(n6451), .B(n6450), .ZN(P1_U3216) );
  INV_X1 U8050 ( .A(n6453), .ZN(n6456) );
  OAI222_X1 U8051 ( .A1(n8405), .A2(n6454), .B1(n9165), .B2(n6456), .C1(n8588), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8052 ( .A(n7041), .ZN(n9807) );
  OAI222_X1 U8053 ( .A1(P1_U3084), .A2(n9807), .B1(n9665), .B2(n6456), .C1(
        n6455), .C2(n7753), .ZN(P1_U3336) );
  INV_X1 U8054 ( .A(n6457), .ZN(n6458) );
  AOI21_X1 U8055 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6466) );
  NAND2_X1 U8056 ( .A1(n9971), .A2(n6461), .ZN(n8399) );
  INV_X1 U8057 ( .A(n8399), .ZN(n6462) );
  NAND2_X1 U8058 ( .A1(n6463), .A2(n6462), .ZN(n6532) );
  AOI22_X1 U8059 ( .A1(n8508), .A2(n6990), .B1(n6532), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6465) );
  INV_X1 U8060 ( .A(n8557), .ZN(n6477) );
  OAI22_X1 U8061 ( .A1(n6477), .A2(n9012), .B1(n6827), .B2(n9014), .ZN(n6991)
         );
  NAND2_X1 U8062 ( .A1(n8460), .A2(n6991), .ZN(n6464) );
  OAI211_X1 U8063 ( .C1(n6466), .C2(n8518), .A(n6465), .B(n6464), .ZN(P2_U3224) );
  NAND2_X1 U8064 ( .A1(n6468), .A2(n6467), .ZN(n6495) );
  INV_X1 U8065 ( .A(n6495), .ZN(n6469) );
  NAND2_X1 U8066 ( .A1(n6496), .A2(n6469), .ZN(n6470) );
  NOR2_X1 U8067 ( .A1(n8399), .A2(n6470), .ZN(n6471) );
  AND2_X2 U8068 ( .A1(n6499), .A2(n6471), .ZN(n10017) );
  INV_X1 U8069 ( .A(n6990), .ZN(n9986) );
  NAND2_X1 U8070 ( .A1(n6472), .A2(n6990), .ZN(n8225) );
  NAND2_X1 U8071 ( .A1(n6983), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U8072 ( .A1(n6472), .A2(n9986), .ZN(n6473) );
  NAND2_X1 U8073 ( .A1(n6984), .A2(n6473), .ZN(n6474) );
  NAND2_X1 U8074 ( .A1(n6827), .A2(n6958), .ZN(n8232) );
  NAND2_X1 U8075 ( .A1(n6474), .A2(n8362), .ZN(n6650) );
  OAI21_X1 U8076 ( .B1(n6474), .B2(n8362), .A(n6650), .ZN(n6957) );
  INV_X1 U8077 ( .A(n6957), .ZN(n6489) );
  NAND2_X1 U8078 ( .A1(n8361), .A2(n5482), .ZN(n6475) );
  XNOR2_X1 U8079 ( .A(n5967), .B(n6475), .ZN(n6476) );
  NAND2_X1 U8080 ( .A1(n6476), .A2(n8888), .ZN(n8982) );
  OR2_X1 U8081 ( .A1(n8389), .A2(n5967), .ZN(n10009) );
  NAND2_X1 U8082 ( .A1(n8982), .A2(n10009), .ZN(n10024) );
  NAND2_X1 U8083 ( .A1(n7023), .A2(n8225), .ZN(n6479) );
  NAND2_X1 U8084 ( .A1(n8229), .A2(n8362), .ZN(n6480) );
  NAND2_X1 U8085 ( .A1(n6654), .A2(n6480), .ZN(n6482) );
  NAND2_X1 U8086 ( .A1(n6482), .A2(n8986), .ZN(n6485) );
  AOI22_X1 U8087 ( .A1(n6483), .A2(n8965), .B1(n8968), .B2(n8554), .ZN(n6484)
         );
  NAND2_X1 U8088 ( .A1(n6485), .A2(n6484), .ZN(n6951) );
  INV_X1 U8089 ( .A(n6951), .ZN(n6488) );
  NOR2_X1 U8090 ( .A1(n6990), .A2(n9979), .ZN(n6986) );
  OR2_X1 U8091 ( .A1(n6986), .A2(n6648), .ZN(n6486) );
  NAND2_X1 U8092 ( .A1(n6648), .A2(n6986), .ZN(n6823) );
  AND2_X1 U8093 ( .A1(n6486), .A2(n6823), .ZN(n6956) );
  AOI22_X1 U8094 ( .A1(n6956), .A2(n9993), .B1(n9992), .B2(n6958), .ZN(n6487)
         );
  OAI211_X1 U8095 ( .C1(n6489), .C2(n9125), .A(n6488), .B(n6487), .ZN(n6500)
         );
  NAND2_X1 U8096 ( .A1(n6500), .A2(n10017), .ZN(n6490) );
  OAI21_X1 U8097 ( .B1(n10017), .B2(n5545), .A(n6490), .ZN(P2_U3457) );
  INV_X1 U8098 ( .A(n6491), .ZN(n6494) );
  OAI222_X1 U8099 ( .A1(n8405), .A2(n6492), .B1(n9165), .B2(n6494), .C1(
        P2_U3152), .C2(n8609), .ZN(P2_U3340) );
  INV_X1 U8100 ( .A(n7031), .ZN(n9296) );
  INV_X1 U8101 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6493) );
  OAI222_X1 U8102 ( .A1(n9296), .A2(P1_U3084), .B1(n9671), .B2(n6494), .C1(
        n6493), .C2(n7753), .ZN(P1_U3335) );
  OR2_X1 U8103 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  NOR2_X1 U8104 ( .A1(n8399), .A2(n6497), .ZN(n6498) );
  AND2_X2 U8105 ( .A1(n6499), .A2(n6498), .ZN(n10039) );
  NAND2_X1 U8106 ( .A1(n6500), .A2(n10039), .ZN(n6501) );
  OAI21_X1 U8107 ( .B1(n10039), .B2(n6694), .A(n6501), .ZN(P2_U3522) );
  INV_X1 U8108 ( .A(n6503), .ZN(n6505) );
  NOR2_X1 U8109 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  XNOR2_X1 U8110 ( .A(n6502), .B(n6506), .ZN(n6512) );
  INV_X1 U8111 ( .A(n7016), .ZN(n6510) );
  INV_X1 U8112 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7376) );
  NOR2_X1 U8113 ( .A1(n7376), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8573) );
  INV_X1 U8114 ( .A(n8573), .ZN(n6507) );
  OAI21_X1 U8115 ( .B1(n8544), .B2(n7017), .A(n6507), .ZN(n6509) );
  INV_X1 U8116 ( .A(n8554), .ZN(n8244) );
  INV_X1 U8117 ( .A(n8552), .ZN(n6752) );
  OAI22_X1 U8118 ( .A1(n8244), .A2(n8536), .B1(n8539), .B2(n6752), .ZN(n6508)
         );
  AOI211_X1 U8119 ( .C1(n6510), .C2(n8526), .A(n6509), .B(n6508), .ZN(n6511)
         );
  OAI21_X1 U8120 ( .B1(n6512), .B2(n8518), .A(n6511), .ZN(P2_U3232) );
  INV_X1 U8121 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8171) );
  OR2_X1 U8122 ( .A1(n8703), .A2(n5574), .ZN(n6518) );
  INV_X1 U8123 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8124 ( .A1(n5562), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8125 ( .A1(n5544), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6513) );
  OAI211_X1 U8126 ( .C1(n6515), .C2(n5564), .A(n6514), .B(n6513), .ZN(n6516)
         );
  INV_X1 U8127 ( .A(n6516), .ZN(n6517) );
  INV_X1 U8128 ( .A(n8192), .ZN(n8710) );
  NAND2_X1 U8129 ( .A1(n8710), .A2(P2_U3966), .ZN(n6519) );
  OAI21_X1 U8130 ( .B1(n8171), .B2(P2_U3966), .A(n6519), .ZN(P2_U3581) );
  INV_X1 U8131 ( .A(n9979), .ZN(n6520) );
  NAND2_X1 U8132 ( .A1(n8557), .A2(n6520), .ZN(n8227) );
  INV_X1 U8133 ( .A(n8539), .ZN(n8496) );
  AOI22_X1 U8134 ( .A1(n8496), .A2(n6483), .B1(n9979), .B2(n8508), .ZN(n6523)
         );
  OAI21_X1 U8135 ( .B1(n6520), .B2(n8213), .A(n7023), .ZN(n6521) );
  AOI22_X1 U8136 ( .A1(n8532), .A2(n6521), .B1(n6532), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8137 ( .C1(n8516), .C2(n8227), .A(n6523), .B(n6522), .ZN(P2_U3234) );
  XNOR2_X1 U8138 ( .A(n6525), .B(n6524), .ZN(n6529) );
  INV_X1 U8139 ( .A(n8536), .ZN(n8511) );
  OAI22_X1 U8140 ( .A1(n6837), .A2(n8544), .B1(n8539), .B2(n6826), .ZN(n6526)
         );
  AOI21_X1 U8141 ( .B1(n8511), .B2(n8555), .A(n6526), .ZN(n6528) );
  MUX2_X1 U8142 ( .A(n8537), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6527) );
  OAI211_X1 U8143 ( .C1(n6529), .C2(n8518), .A(n6528), .B(n6527), .ZN(P2_U3220) );
  XNOR2_X1 U8144 ( .A(n6531), .B(n6530), .ZN(n6535) );
  AOI22_X1 U8145 ( .A1(n8511), .A2(n6483), .B1(n8496), .B2(n8554), .ZN(n6534)
         );
  AOI22_X1 U8146 ( .A1(n8508), .A2(n6958), .B1(n6532), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6533) );
  OAI211_X1 U8147 ( .C1(n6535), .C2(n8518), .A(n6534), .B(n6533), .ZN(P2_U3239) );
  XNOR2_X1 U8148 ( .A(n6536), .B(n7865), .ZN(n6541) );
  INV_X1 U8149 ( .A(n6541), .ZN(n9909) );
  NOR2_X1 U8150 ( .A1(n6284), .A2(n9850), .ZN(n6537) );
  NAND2_X1 U8151 ( .A1(n9884), .A2(n6537), .ZN(n6643) );
  INV_X1 U8152 ( .A(n9878), .ZN(n7699) );
  XNOR2_X1 U8153 ( .A(n7803), .B(n7865), .ZN(n6539) );
  INV_X1 U8154 ( .A(n9871), .ZN(n9527) );
  AOI22_X1 U8155 ( .A1(n9875), .A2(n9874), .B1(n9845), .B2(n9873), .ZN(n6538)
         );
  OAI21_X1 U8156 ( .B1(n6539), .B2(n9527), .A(n6538), .ZN(n6540) );
  AOI21_X1 U8157 ( .B1(n7699), .B2(n6541), .A(n6540), .ZN(n9908) );
  MUX2_X1 U8158 ( .A(n6542), .B(n9908), .S(n9884), .Z(n6547) );
  NAND2_X1 U8159 ( .A1(n9535), .A2(n9914), .ZN(n9440) );
  INV_X1 U8160 ( .A(n6639), .ZN(n6543) );
  AOI21_X1 U8161 ( .B1(n9905), .B2(n6543), .A(n5388), .ZN(n9906) );
  OAI22_X1 U8162 ( .A1(n9539), .A2(n6544), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9880), .ZN(n6545) );
  AOI21_X1 U8163 ( .B1(n9504), .B2(n9906), .A(n6545), .ZN(n6546) );
  OAI211_X1 U8164 ( .C1(n9909), .C2(n6643), .A(n6547), .B(n6546), .ZN(P1_U3288) );
  INV_X1 U8165 ( .A(n6548), .ZN(n8403) );
  OAI222_X1 U8166 ( .A1(P1_U3084), .A2(n9850), .B1(n9671), .B2(n8403), .C1(
        n6549), .C2(n7753), .ZN(P1_U3334) );
  AOI22_X1 U8167 ( .A1(n9856), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n9826), .ZN(n6551) );
  INV_X1 U8168 ( .A(n9539), .ZN(n9555) );
  OAI21_X1 U8169 ( .B1(n9504), .B2(n9555), .A(n9860), .ZN(n6550) );
  OAI211_X1 U8170 ( .C1(n6552), .C2(n9856), .A(n6551), .B(n6550), .ZN(P1_U3291) );
  NAND2_X1 U8171 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  XNOR2_X1 U8172 ( .A(n6555), .B(n7864), .ZN(n6560) );
  INV_X1 U8173 ( .A(n6560), .ZN(n9919) );
  XNOR2_X1 U8174 ( .A(n6556), .B(n7864), .ZN(n6558) );
  AOI22_X1 U8175 ( .A1(n9875), .A2(n9290), .B1(n9289), .B2(n9873), .ZN(n6557)
         );
  OAI21_X1 U8176 ( .B1(n6558), .B2(n9527), .A(n6557), .ZN(n6559) );
  AOI21_X1 U8177 ( .B1(n7699), .B2(n6560), .A(n6559), .ZN(n9917) );
  MUX2_X1 U8178 ( .A(n6151), .B(n9917), .S(n9884), .Z(n6566) );
  INV_X1 U8179 ( .A(n9837), .ZN(n6561) );
  AOI21_X1 U8180 ( .B1(n9912), .B2(n6562), .A(n6561), .ZN(n9915) );
  INV_X1 U8181 ( .A(n9223), .ZN(n6563) );
  AOI21_X1 U8182 ( .B1(n9915), .B2(n9504), .A(n6564), .ZN(n6565) );
  OAI211_X1 U8183 ( .C1(n9919), .C2(n6643), .A(n6566), .B(n6565), .ZN(P1_U3287) );
  INV_X1 U8184 ( .A(n6567), .ZN(n6570) );
  INV_X1 U8185 ( .A(n6568), .ZN(n6569) );
  AOI21_X1 U8186 ( .B1(n6570), .B2(n6569), .A(n8518), .ZN(n6573) );
  NOR3_X1 U8187 ( .A1(n8516), .A2(n6571), .A3(n8505), .ZN(n6572) );
  OAI21_X1 U8188 ( .B1(n6573), .B2(n6572), .A(n6618), .ZN(n6578) );
  INV_X1 U8189 ( .A(n6574), .ZN(n6977) );
  INV_X1 U8190 ( .A(n7285), .ZN(n8259) );
  OAI22_X1 U8191 ( .A1(n8544), .A2(n8259), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7434), .ZN(n6576) );
  INV_X1 U8192 ( .A(n8548), .ZN(n7557) );
  OAI22_X1 U8193 ( .A1(n8505), .A2(n8536), .B1(n8539), .B2(n7557), .ZN(n6575)
         );
  AOI211_X1 U8194 ( .C1(n6977), .C2(n8526), .A(n6576), .B(n6575), .ZN(n6577)
         );
  NAND2_X1 U8195 ( .A1(n6578), .A2(n6577), .ZN(P2_U3223) );
  NAND2_X1 U8196 ( .A1(n9845), .A2(n8412), .ZN(n6583) );
  NAND2_X1 U8197 ( .A1(n9912), .A2(n8406), .ZN(n6582) );
  NAND2_X1 U8198 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  XNOR2_X1 U8199 ( .A(n6584), .B(n6381), .ZN(n6585) );
  AOI22_X1 U8200 ( .A1(n9845), .A2(n8411), .B1(n9912), .B2(n8412), .ZN(n6586)
         );
  XNOR2_X1 U8201 ( .A(n6585), .B(n6586), .ZN(n9221) );
  NAND2_X1 U8202 ( .A1(n9289), .A2(n8411), .ZN(n6589) );
  NAND2_X1 U8203 ( .A1(n5015), .A2(n8412), .ZN(n6588) );
  NAND2_X1 U8204 ( .A1(n6589), .A2(n6588), .ZN(n6770) );
  NAND2_X1 U8205 ( .A1(n9289), .A2(n8412), .ZN(n6591) );
  NAND2_X1 U8206 ( .A1(n5015), .A2(n8406), .ZN(n6590) );
  NAND2_X1 U8207 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  XNOR2_X1 U8208 ( .A(n6592), .B(n6381), .ZN(n6600) );
  NAND2_X1 U8209 ( .A1(n9846), .A2(n8412), .ZN(n6594) );
  NAND2_X1 U8210 ( .A1(n6930), .A2(n8406), .ZN(n6593) );
  NAND2_X1 U8211 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  XNOR2_X1 U8212 ( .A(n6595), .B(n6381), .ZN(n6599) );
  NAND2_X1 U8213 ( .A1(n9846), .A2(n8411), .ZN(n6597) );
  NAND2_X1 U8214 ( .A1(n6930), .A2(n8412), .ZN(n6596) );
  NAND2_X1 U8215 ( .A1(n6597), .A2(n6596), .ZN(n6926) );
  AOI22_X1 U8216 ( .A1(n6770), .A2(n6600), .B1(n6599), .B2(n6926), .ZN(n6598)
         );
  OAI21_X1 U8217 ( .B1(n6600), .B2(n6770), .A(n6926), .ZN(n6602) );
  INV_X1 U8218 ( .A(n6599), .ZN(n6927) );
  INV_X1 U8219 ( .A(n6600), .ZN(n6925) );
  NOR2_X1 U8220 ( .A1(n6770), .A2(n6926), .ZN(n6601) );
  AOI22_X1 U8221 ( .A1(n6602), .A2(n6927), .B1(n6925), .B2(n6601), .ZN(n6603)
         );
  NAND2_X1 U8222 ( .A1(n9288), .A2(n8412), .ZN(n6606) );
  NAND2_X1 U8223 ( .A1(n6612), .A2(n8406), .ZN(n6605) );
  NAND2_X1 U8224 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  XNOR2_X1 U8225 ( .A(n6607), .B(n4311), .ZN(n6855) );
  NAND2_X1 U8226 ( .A1(n9288), .A2(n8411), .ZN(n6609) );
  NAND2_X1 U8227 ( .A1(n6612), .A2(n8412), .ZN(n6608) );
  AND2_X1 U8228 ( .A1(n6609), .A2(n6608), .ZN(n6856) );
  XNOR2_X1 U8229 ( .A(n6855), .B(n6856), .ZN(n6610) );
  XNOR2_X1 U8230 ( .A(n6861), .B(n6610), .ZN(n6617) );
  INV_X1 U8231 ( .A(n6722), .ZN(n6611) );
  AOI22_X1 U8232 ( .A1(n9259), .A2(n6611), .B1(n9685), .B2(n9846), .ZN(n6616)
         );
  INV_X1 U8233 ( .A(n9693), .ZN(n6931) );
  NAND2_X1 U8234 ( .A1(n9913), .A2(n6612), .ZN(n9937) );
  NOR2_X1 U8235 ( .A1(n6931), .A2(n9937), .ZN(n6613) );
  AOI211_X1 U8236 ( .C1(n9222), .C2(n9287), .A(n6614), .B(n6613), .ZN(n6615)
         );
  OAI211_X1 U8237 ( .C1(n6617), .C2(n9278), .A(n6616), .B(n6615), .ZN(P1_U3211) );
  INV_X1 U8238 ( .A(n6618), .ZN(n6621) );
  NOR3_X1 U8239 ( .A1(n8516), .A2(n6619), .A3(n7287), .ZN(n6620) );
  AOI21_X1 U8240 ( .B1(n6621), .B2(n8532), .A(n6620), .ZN(n6630) );
  INV_X1 U8241 ( .A(n6622), .ZN(n6627) );
  OAI22_X1 U8242 ( .A1(n7287), .A2(n8536), .B1(n8539), .B2(n7600), .ZN(n6626)
         );
  NOR2_X1 U8243 ( .A1(n5627), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7132) );
  INV_X1 U8244 ( .A(n7132), .ZN(n6624) );
  INV_X1 U8245 ( .A(n10011), .ZN(n7297) );
  NAND2_X1 U8246 ( .A1(n8508), .A2(n7297), .ZN(n6623) );
  OAI211_X1 U8247 ( .C1(n8537), .C2(n7291), .A(n6624), .B(n6623), .ZN(n6625)
         );
  AOI211_X1 U8248 ( .C1(n6627), .C2(n8532), .A(n6626), .B(n6625), .ZN(n6628)
         );
  OAI21_X1 U8249 ( .B1(n6630), .B2(n6629), .A(n6628), .ZN(P2_U3233) );
  INV_X1 U8250 ( .A(n6631), .ZN(n6717) );
  OAI222_X1 U8251 ( .A1(n9165), .A2(n6717), .B1(P2_U3152), .B2(n8361), .C1(
        n6632), .C2(n8405), .ZN(P2_U3338) );
  XOR2_X1 U8252 ( .A(n7866), .B(n8051), .Z(n6638) );
  AOI22_X1 U8253 ( .A1(n9875), .A2(n9291), .B1(n9290), .B2(n9873), .ZN(n6637)
         );
  NAND2_X1 U8254 ( .A1(n6633), .A2(n7866), .ZN(n6634) );
  NAND2_X1 U8255 ( .A1(n6635), .A2(n6634), .ZN(n9902) );
  NAND2_X1 U8256 ( .A1(n9902), .A2(n7699), .ZN(n6636) );
  OAI211_X1 U8257 ( .C1(n6638), .C2(n9527), .A(n6637), .B(n6636), .ZN(n9900)
         );
  AND2_X1 U8258 ( .A1(n9862), .A2(n6394), .ZN(n6640) );
  OR2_X1 U8259 ( .A1(n6640), .A2(n6639), .ZN(n9899) );
  OAI22_X1 U8260 ( .A1(n9884), .A2(n6127), .B1(n6641), .B2(n9880), .ZN(n6642)
         );
  AOI21_X1 U8261 ( .B1(n9555), .B2(n6394), .A(n6642), .ZN(n6645) );
  INV_X1 U8262 ( .A(n6643), .ZN(n7706) );
  NAND2_X1 U8263 ( .A1(n9902), .A2(n7706), .ZN(n6644) );
  OAI211_X1 U8264 ( .C1(n9440), .C2(n9899), .A(n6645), .B(n6644), .ZN(n6646)
         );
  AOI21_X1 U8265 ( .B1(n9900), .B2(n9884), .A(n6646), .ZN(n6647) );
  INV_X1 U8266 ( .A(n6647), .ZN(P1_U3289) );
  INV_X1 U8267 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U8268 ( .A1(n6827), .A2(n6648), .ZN(n6649) );
  NAND2_X1 U8269 ( .A1(n6650), .A2(n6649), .ZN(n6834) );
  NAND2_X1 U8270 ( .A1(n6834), .A2(n8363), .ZN(n6833) );
  NAND2_X1 U8271 ( .A1(n8244), .A2(n6837), .ZN(n6651) );
  NAND2_X1 U8272 ( .A1(n6833), .A2(n6651), .ZN(n6652) );
  NAND2_X1 U8273 ( .A1(n6826), .A2(n6658), .ZN(n8220) );
  INV_X1 U8274 ( .A(n6826), .ZN(n8553) );
  NAND2_X1 U8275 ( .A1(n8553), .A2(n7017), .ZN(n6906) );
  NAND2_X1 U8276 ( .A1(n8220), .A2(n6906), .ZN(n8359) );
  NAND2_X1 U8277 ( .A1(n6652), .A2(n8359), .ZN(n6750) );
  OAI21_X1 U8278 ( .B1(n6652), .B2(n8359), .A(n6750), .ZN(n6653) );
  INV_X1 U8279 ( .A(n6653), .ZN(n7018) );
  INV_X1 U8280 ( .A(n8363), .ZN(n8237) );
  NAND2_X1 U8281 ( .A1(n6824), .A2(n8237), .ZN(n6825) );
  NAND2_X1 U8282 ( .A1(n8244), .A2(n9991), .ZN(n8219) );
  XOR2_X1 U8283 ( .A(n6755), .B(n8359), .Z(n6655) );
  AOI222_X1 U8284 ( .A1(n8986), .A2(n6655), .B1(n8552), .B2(n8968), .C1(n8554), 
        .C2(n8965), .ZN(n7022) );
  AND2_X1 U8285 ( .A1(n6821), .A2(n6658), .ZN(n6657) );
  NOR2_X1 U8286 ( .A1(n6904), .A2(n6657), .ZN(n7014) );
  AOI22_X1 U8287 ( .A1(n7014), .A2(n9993), .B1(n9992), .B2(n6658), .ZN(n6659)
         );
  OAI211_X1 U8288 ( .C1(n9125), .C2(n7018), .A(n7022), .B(n6659), .ZN(n6776)
         );
  NAND2_X1 U8289 ( .A1(n6776), .A2(n10039), .ZN(n6660) );
  OAI21_X1 U8290 ( .B1(n10039), .B2(n8576), .A(n6660), .ZN(P2_U3524) );
  NAND2_X1 U8291 ( .A1(n9971), .A2(n6661), .ZN(n6666) );
  NAND2_X1 U8292 ( .A1(n6662), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7726) );
  OAI21_X1 U8293 ( .B1(n6663), .B2(n7726), .A(n8402), .ZN(n6664) );
  INV_X1 U8294 ( .A(n6664), .ZN(n6665) );
  NAND2_X1 U8295 ( .A1(n6666), .A2(n6665), .ZN(n6668) );
  NAND2_X1 U8296 ( .A1(n6668), .A2(n6667), .ZN(n6707) );
  INV_X2 U8297 ( .A(P2_U3966), .ZN(n8556) );
  NAND2_X1 U8298 ( .A1(n6707), .A2(n8556), .ZN(n6684) );
  INV_X1 U8299 ( .A(n8398), .ZN(n8632) );
  NAND2_X1 U8300 ( .A1(n6684), .A2(n8632), .ZN(n8614) );
  NOR2_X2 U8301 ( .A1(n8614), .A2(n5984), .ZN(n8613) );
  MUX2_X1 U8302 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7604), .S(n6736), .Z(n6669)
         );
  INV_X1 U8303 ( .A(n6669), .ZN(n6683) );
  INV_X1 U8304 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6953) );
  XNOR2_X1 U8305 ( .A(n8561), .B(n6953), .ZN(n8560) );
  MUX2_X1 U8306 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6993), .S(n7232), .Z(n7225)
         );
  NAND3_X1 U8307 ( .A1(n7225), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n7226) );
  OAI21_X1 U8308 ( .B1(n6670), .B2(n6993), .A(n7226), .ZN(n8559) );
  NAND2_X1 U8309 ( .A1(n8560), .A2(n8559), .ZN(n8558) );
  OAI21_X1 U8310 ( .B1(n6953), .B2(n6671), .A(n8558), .ZN(n6799) );
  MUX2_X1 U8311 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6672), .S(n6699), .Z(n6800)
         );
  NAND2_X1 U8312 ( .A1(n6799), .A2(n6800), .ZN(n6798) );
  OAI21_X1 U8313 ( .B1(n6672), .B2(n6803), .A(n6798), .ZN(n8571) );
  MUX2_X1 U8314 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6673), .S(n8575), .Z(n8572)
         );
  NAND2_X1 U8315 ( .A1(n8571), .A2(n8572), .ZN(n8570) );
  OAI21_X1 U8316 ( .B1(n8574), .B2(n6673), .A(n8570), .ZN(n6811) );
  OR2_X1 U8317 ( .A1(n6702), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8318 ( .A1(n6702), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6674) );
  AND2_X1 U8319 ( .A1(n6675), .A2(n6674), .ZN(n6812) );
  INV_X1 U8320 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U8321 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6676), .S(n6692), .Z(n6677)
         );
  INV_X1 U8322 ( .A(n6677), .ZN(n7119) );
  AOI21_X1 U8323 ( .B1(n6692), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7118), .ZN(
        n7143) );
  NAND2_X1 U8324 ( .A1(n6690), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6678) );
  OAI21_X1 U8325 ( .B1(n6690), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6678), .ZN(
        n7142) );
  NOR2_X1 U8326 ( .A1(n7143), .A2(n7142), .ZN(n7141) );
  AOI21_X1 U8327 ( .B1(n6690), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7141), .ZN(
        n7108) );
  NAND2_X1 U8328 ( .A1(n6689), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U8329 ( .B1(n6689), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6679), .ZN(
        n7107) );
  NOR2_X1 U8330 ( .A1(n7108), .A2(n7107), .ZN(n7106) );
  NAND2_X1 U8331 ( .A1(n6688), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6680) );
  OAI21_X1 U8332 ( .B1(n6688), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6680), .ZN(
        n7130) );
  NAND2_X1 U8333 ( .A1(n6686), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6681) );
  OAI21_X1 U8334 ( .B1(n6686), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6681), .ZN(
        n7095) );
  AOI21_X1 U8335 ( .B1(n6686), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7094), .ZN(
        n6682) );
  NAND2_X1 U8336 ( .A1(n6682), .A2(n6683), .ZN(n6737) );
  OAI21_X1 U8337 ( .B1(n6683), .B2(n6682), .A(n6737), .ZN(n6714) );
  NAND2_X1 U8338 ( .A1(n6684), .A2(n5984), .ZN(n8619) );
  NOR2_X1 U8339 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5665), .ZN(n6685) );
  AOI21_X1 U8340 ( .B1(n8599), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6685), .ZN(
        n6712) );
  MUX2_X1 U8341 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6687), .S(n6686), .Z(n7099)
         );
  INV_X1 U8342 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10035) );
  MUX2_X1 U8343 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10035), .S(n6688), .Z(n7134)
         );
  INV_X1 U8344 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7256) );
  MUX2_X1 U8345 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7256), .S(n6689), .Z(n7111)
         );
  NAND2_X1 U8346 ( .A1(n6690), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8347 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6691), .S(n6690), .Z(n7147)
         );
  MUX2_X1 U8348 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6693), .S(n6692), .Z(n7122)
         );
  MUX2_X1 U8349 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6694), .S(n8561), .Z(n8565)
         );
  INV_X1 U8350 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6695) );
  MUX2_X1 U8351 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6695), .S(n7232), .Z(n6697)
         );
  AND2_X1 U8352 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6696) );
  NAND2_X1 U8353 ( .A1(n6697), .A2(n6696), .ZN(n7221) );
  NAND2_X1 U8354 ( .A1(n7232), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8355 ( .A1(n7221), .A2(n6698), .ZN(n8564) );
  NAND2_X1 U8356 ( .A1(n8565), .A2(n8564), .ZN(n8563) );
  NAND2_X1 U8357 ( .A1(n8561), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6794) );
  INV_X1 U8358 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10030) );
  MUX2_X1 U8359 ( .A(n10030), .B(P2_REG1_REG_3__SCAN_IN), .S(n6699), .Z(n6793)
         );
  AOI21_X1 U8360 ( .B1(n8563), .B2(n6794), .A(n6793), .ZN(n8582) );
  AND2_X1 U8361 ( .A1(n6699), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8577) );
  OR2_X1 U8362 ( .A1(n8582), .A2(n8577), .ZN(n6701) );
  MUX2_X1 U8363 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n8576), .S(n8575), .Z(n6700)
         );
  NAND2_X1 U8364 ( .A1(n6701), .A2(n6700), .ZN(n8580) );
  NAND2_X1 U8365 ( .A1(n8575), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6805) );
  INV_X1 U8366 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10032) );
  MUX2_X1 U8367 ( .A(n10032), .B(P2_REG1_REG_5__SCAN_IN), .S(n6702), .Z(n6804)
         );
  AOI21_X1 U8368 ( .B1(n8580), .B2(n6805), .A(n6804), .ZN(n6807) );
  INV_X1 U8369 ( .A(n6807), .ZN(n6704) );
  NAND2_X1 U8370 ( .A1(n6702), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8371 ( .A1(n6704), .A2(n6703), .ZN(n7123) );
  NAND2_X1 U8372 ( .A1(n7122), .A2(n7123), .ZN(n7121) );
  OAI21_X1 U8373 ( .B1(n7126), .B2(n6693), .A(n7121), .ZN(n7146) );
  NAND2_X1 U8374 ( .A1(n7147), .A2(n7146), .ZN(n7145) );
  NAND2_X1 U8375 ( .A1(n6705), .A2(n7145), .ZN(n7112) );
  NAND2_X1 U8376 ( .A1(n7111), .A2(n7112), .ZN(n7110) );
  OAI21_X1 U8377 ( .B1(n7115), .B2(n7256), .A(n7110), .ZN(n7135) );
  NAND2_X1 U8378 ( .A1(n7134), .A2(n7135), .ZN(n7133) );
  OAI21_X1 U8379 ( .B1(n7138), .B2(n10035), .A(n7133), .ZN(n7100) );
  NAND2_X1 U8380 ( .A1(n7099), .A2(n7100), .ZN(n7098) );
  OAI21_X1 U8381 ( .B1(n7103), .B2(n6687), .A(n7098), .ZN(n6710) );
  MUX2_X1 U8382 ( .A(n6706), .B(P2_REG1_REG_11__SCAN_IN), .S(n6736), .Z(n6709)
         );
  INV_X1 U8383 ( .A(n6707), .ZN(n6708) );
  AND2_X1 U8384 ( .A1(n6708), .A2(n8398), .ZN(n8612) );
  NAND2_X1 U8385 ( .A1(n6709), .A2(n6710), .ZN(n6730) );
  OAI211_X1 U8386 ( .C1(n6710), .C2(n6709), .A(n8612), .B(n6730), .ZN(n6711)
         );
  OAI211_X1 U8387 ( .C1(n8619), .C2(n6736), .A(n6712), .B(n6711), .ZN(n6713)
         );
  AOI21_X1 U8388 ( .B1(n8613), .B2(n6714), .A(n6713), .ZN(n6715) );
  INV_X1 U8389 ( .A(n6715), .ZN(P2_U3256) );
  OAI222_X1 U8390 ( .A1(n6029), .A2(P1_U3084), .B1(n9671), .B2(n6717), .C1(
        n6716), .C2(n7753), .ZN(P1_U3333) );
  INV_X1 U8391 ( .A(n6718), .ZN(n7755) );
  INV_X1 U8392 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6719) );
  OAI222_X1 U8393 ( .A1(n9165), .A2(n7755), .B1(P2_U3152), .B2(n8193), .C1(
        n6719), .C2(n8405), .ZN(P2_U3337) );
  XNOR2_X1 U8394 ( .A(n6720), .B(n7869), .ZN(n9941) );
  INV_X1 U8395 ( .A(n9855), .ZN(n9488) );
  OAI211_X1 U8396 ( .C1(n6893), .C2(n6723), .A(n9914), .B(n6943), .ZN(n9938)
         );
  NOR2_X1 U8397 ( .A1(n6721), .A2(n9867), .ZN(n9513) );
  INV_X1 U8398 ( .A(n9513), .ZN(n9559) );
  NOR2_X1 U8399 ( .A1(n9938), .A2(n9559), .ZN(n6725) );
  OAI22_X1 U8400 ( .A1(n9539), .A2(n6723), .B1(n9880), .B2(n6722), .ZN(n6724)
         );
  AOI211_X1 U8401 ( .C1(n9941), .C2(n9488), .A(n6725), .B(n6724), .ZN(n6729)
         );
  XNOR2_X1 U8402 ( .A(n6726), .B(n7869), .ZN(n6727) );
  AOI222_X1 U8403 ( .A1(n9871), .A2(n6727), .B1(n9287), .B2(n9873), .C1(n9846), 
        .C2(n9875), .ZN(n9939) );
  MUX2_X1 U8404 ( .A(n6146), .B(n9939), .S(n9884), .Z(n6728) );
  NAND2_X1 U8405 ( .A1(n6729), .A2(n6728), .ZN(P1_U3284) );
  OAI21_X1 U8406 ( .B1(n6736), .B2(n6706), .A(n6730), .ZN(n7235) );
  MUX2_X1 U8407 ( .A(n6731), .B(P2_REG1_REG_12__SCAN_IN), .S(n7246), .Z(n7236)
         );
  NOR2_X1 U8408 ( .A1(n7235), .A2(n7236), .ZN(n7234) );
  AOI21_X1 U8409 ( .B1(n6732), .B2(n6731), .A(n7234), .ZN(n6734) );
  AOI22_X1 U8410 ( .A1(n6784), .A2(n6779), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n6780), .ZN(n6733) );
  NOR2_X1 U8411 ( .A1(n6734), .A2(n6733), .ZN(n6778) );
  AOI21_X1 U8412 ( .B1(n6734), .B2(n6733), .A(n6778), .ZN(n6748) );
  INV_X1 U8413 ( .A(n8612), .ZN(n8620) );
  NAND2_X1 U8414 ( .A1(n7246), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6735) );
  OAI21_X1 U8415 ( .B1(n7246), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6735), .ZN(
        n7242) );
  INV_X1 U8416 ( .A(n6736), .ZN(n6738) );
  OAI21_X1 U8417 ( .B1(n6738), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6737), .ZN(
        n7243) );
  NOR2_X1 U8418 ( .A1(n7242), .A2(n7243), .ZN(n7241) );
  NOR2_X1 U8419 ( .A1(n6784), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6739) );
  AOI21_X1 U8420 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6784), .A(n6739), .ZN(
        n6740) );
  OAI21_X1 U8421 ( .B1(n6741), .B2(n6740), .A(n6783), .ZN(n6742) );
  NAND2_X1 U8422 ( .A1(n6742), .A2(n8613), .ZN(n6747) );
  INV_X1 U8423 ( .A(n8619), .ZN(n8562) );
  INV_X1 U8424 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6744) );
  OAI22_X1 U8425 ( .A1(n8629), .A2(n6744), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6743), .ZN(n6745) );
  AOI21_X1 U8426 ( .B1(n8562), .B2(n6784), .A(n6745), .ZN(n6746) );
  OAI211_X1 U8427 ( .C1(n6748), .C2(n8620), .A(n6747), .B(n6746), .ZN(P2_U3258) );
  NAND2_X1 U8428 ( .A1(n6826), .A2(n7017), .ZN(n6749) );
  NOR2_X1 U8429 ( .A1(n8552), .A2(n6751), .ZN(n6754) );
  NAND2_X1 U8430 ( .A1(n6752), .A2(n6751), .ZN(n8221) );
  NAND2_X1 U8431 ( .A1(n8552), .A2(n10001), .ZN(n8242) );
  NAND2_X1 U8432 ( .A1(n8221), .A2(n8242), .ZN(n8360) );
  OR2_X1 U8433 ( .A1(n8360), .A2(n6752), .ZN(n6753) );
  NAND2_X1 U8434 ( .A1(n6878), .A2(n4310), .ZN(n8250) );
  NAND2_X1 U8435 ( .A1(n8551), .A2(n6762), .ZN(n8248) );
  NAND2_X1 U8436 ( .A1(n8250), .A2(n8248), .ZN(n8364) );
  XNOR2_X1 U8437 ( .A(n6875), .B(n8364), .ZN(n7013) );
  INV_X1 U8438 ( .A(n8364), .ZN(n6758) );
  NAND2_X1 U8439 ( .A1(n8220), .A2(n8221), .ZN(n8218) );
  INV_X1 U8440 ( .A(n8218), .ZN(n6756) );
  OAI21_X1 U8441 ( .B1(n6758), .B2(n6757), .A(n6968), .ZN(n6761) );
  NAND2_X1 U8442 ( .A1(n8552), .A2(n8965), .ZN(n6759) );
  OAI21_X1 U8443 ( .B1(n8505), .B2(n9014), .A(n6759), .ZN(n6760) );
  AOI21_X1 U8444 ( .B1(n6761), .B2(n8986), .A(n6760), .ZN(n7010) );
  INV_X1 U8445 ( .A(n6880), .ZN(n6763) );
  AOI21_X1 U8446 ( .B1(n4310), .B2(n4376), .A(n6763), .ZN(n7007) );
  AOI22_X1 U8447 ( .A1(n7007), .A2(n9993), .B1(n9992), .B2(n4310), .ZN(n6764)
         );
  OAI211_X1 U8448 ( .C1(n7013), .C2(n9125), .A(n7010), .B(n6764), .ZN(n6766)
         );
  NAND2_X1 U8449 ( .A1(n6766), .A2(n10039), .ZN(n6765) );
  OAI21_X1 U8450 ( .B1(n10039), .B2(n6693), .A(n6765), .ZN(P2_U3526) );
  NAND2_X1 U8451 ( .A1(n6766), .A2(n10017), .ZN(n6767) );
  OAI21_X1 U8452 ( .B1(n10017), .B2(n5488), .A(n6767), .ZN(P2_U3469) );
  XNOR2_X1 U8453 ( .A(n6768), .B(n6925), .ZN(n6769) );
  NOR2_X1 U8454 ( .A1(n6769), .A2(n6770), .ZN(n6924) );
  AOI21_X1 U8455 ( .B1(n6770), .B2(n6769), .A(n6924), .ZN(n6775) );
  AOI22_X1 U8456 ( .A1(n9222), .A2(n9846), .B1(n9685), .B2(n9845), .ZN(n6774)
         );
  AND2_X1 U8457 ( .A1(n9913), .A2(n5015), .ZN(n9925) );
  NOR2_X1 U8458 ( .A1(n9699), .A2(n9838), .ZN(n6771) );
  AOI211_X1 U8459 ( .C1(n9693), .C2(n9925), .A(n6772), .B(n6771), .ZN(n6773)
         );
  OAI211_X1 U8460 ( .C1(n6775), .C2(n9278), .A(n6774), .B(n6773), .ZN(P1_U3225) );
  NAND2_X1 U8461 ( .A1(n6776), .A2(n10017), .ZN(n6777) );
  OAI21_X1 U8462 ( .B1(n10017), .B2(n5575), .A(n6777), .ZN(P2_U3463) );
  AOI21_X1 U8463 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6782) );
  AOI22_X1 U8464 ( .A1(n7162), .A2(n7165), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7166), .ZN(n6781) );
  NOR2_X1 U8465 ( .A1(n6782), .A2(n6781), .ZN(n7164) );
  AOI21_X1 U8466 ( .B1(n6782), .B2(n6781), .A(n7164), .ZN(n6792) );
  AOI22_X1 U8467 ( .A1(n7162), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n5719), .B2(
        n7166), .ZN(n6786) );
  OAI21_X1 U8468 ( .B1(n6786), .B2(n6785), .A(n7161), .ZN(n6787) );
  NAND2_X1 U8469 ( .A1(n6787), .A2(n8613), .ZN(n6791) );
  INV_X1 U8470 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8471 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7614) );
  OAI21_X1 U8472 ( .B1(n8629), .B2(n6788), .A(n7614), .ZN(n6789) );
  AOI21_X1 U8473 ( .B1(n8562), .B2(n7162), .A(n6789), .ZN(n6790) );
  OAI211_X1 U8474 ( .C1(n6792), .C2(n8620), .A(n6791), .B(n6790), .ZN(P2_U3259) );
  INV_X1 U8475 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7378) );
  NOR2_X1 U8476 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7378), .ZN(n6797) );
  AND3_X1 U8477 ( .A1(n8563), .A2(n6794), .A3(n6793), .ZN(n6795) );
  NOR3_X1 U8478 ( .A1(n8620), .A2(n8582), .A3(n6795), .ZN(n6796) );
  AOI211_X1 U8479 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n8599), .A(n6797), .B(
        n6796), .ZN(n6802) );
  OAI211_X1 U8480 ( .C1(n6800), .C2(n6799), .A(n8613), .B(n6798), .ZN(n6801)
         );
  OAI211_X1 U8481 ( .C1(n8619), .C2(n6803), .A(n6802), .B(n6801), .ZN(P2_U3248) );
  NOR2_X1 U8482 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5506), .ZN(n6809) );
  AND3_X1 U8483 ( .A1(n8580), .A2(n6805), .A3(n6804), .ZN(n6806) );
  NOR3_X1 U8484 ( .A1(n8620), .A2(n6807), .A3(n6806), .ZN(n6808) );
  AOI211_X1 U8485 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n8599), .A(n6809), .B(
        n6808), .ZN(n6814) );
  OAI211_X1 U8486 ( .C1(n6812), .C2(n6811), .A(n8613), .B(n6810), .ZN(n6813)
         );
  OAI211_X1 U8487 ( .C1(n8619), .C2(n6815), .A(n6814), .B(n6813), .ZN(P2_U3250) );
  NOR2_X1 U8488 ( .A1(n8399), .A2(n6816), .ZN(n6817) );
  NAND2_X1 U8489 ( .A1(n6818), .A2(n6817), .ZN(n6820) );
  NOR2_X1 U8490 ( .A1(n6820), .A2(n8213), .ZN(n9022) );
  INV_X1 U8491 ( .A(n6821), .ZN(n6822) );
  AOI21_X1 U8492 ( .B1(n9991), .B2(n6823), .A(n6822), .ZN(n9994) );
  OAI22_X1 U8493 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8943), .B1(n6672), .B2(
        n8946), .ZN(n6831) );
  OAI21_X1 U8494 ( .B1(n6824), .B2(n8237), .A(n6825), .ZN(n6829) );
  OAI22_X1 U8495 ( .A1(n6827), .A2(n9012), .B1(n6826), .B2(n9014), .ZN(n6828)
         );
  AOI21_X1 U8496 ( .B1(n6829), .B2(n8986), .A(n6828), .ZN(n9996) );
  NOR2_X1 U8497 ( .A1(n9996), .A2(n9019), .ZN(n6830) );
  AOI211_X1 U8498 ( .C1(n8995), .C2(n9994), .A(n6831), .B(n6830), .ZN(n6836)
         );
  OR2_X1 U8499 ( .A1(n8389), .A2(n8193), .ZN(n6974) );
  NAND2_X1 U8500 ( .A1(n8982), .A2(n6974), .ZN(n6832) );
  OAI21_X1 U8501 ( .B1(n6834), .B2(n8363), .A(n6833), .ZN(n9998) );
  NAND2_X1 U8502 ( .A1(n8940), .A2(n9998), .ZN(n6835) );
  OAI211_X1 U8503 ( .C1(n6837), .C2(n9008), .A(n6836), .B(n6835), .ZN(P2_U3293) );
  INV_X1 U8504 ( .A(n6838), .ZN(n6839) );
  AOI21_X1 U8505 ( .B1(n6916), .B2(n6839), .A(n8518), .ZN(n6843) );
  NOR3_X1 U8506 ( .A1(n8516), .A2(n6840), .A3(n7600), .ZN(n6842) );
  OAI21_X1 U8507 ( .B1(n6843), .B2(n6842), .A(n6841), .ZN(n6847) );
  OAI22_X1 U8508 ( .A1(n8536), .A2(n7600), .B1(n8537), .B2(n7603), .ZN(n6845)
         );
  OAI22_X1 U8509 ( .A1(n8539), .A2(n8978), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5665), .ZN(n6844) );
  AOI211_X1 U8510 ( .C1(n8652), .C2(n8508), .A(n6845), .B(n6844), .ZN(n6846)
         );
  NAND2_X1 U8511 ( .A1(n6847), .A2(n6846), .ZN(P2_U3238) );
  AOI22_X1 U8512 ( .A1(n8613), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n8612), .ZN(n6852) );
  INV_X1 U8513 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8514 ( .A1(n8612), .A2(n6848), .ZN(n6849) );
  OAI211_X1 U8515 ( .C1(n8614), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6849), .B(
        n8619), .ZN(n6850) );
  INV_X1 U8516 ( .A(n6850), .ZN(n6851) );
  MUX2_X1 U8517 ( .A(n6852), .B(n6851), .S(P2_IR_REG_0__SCAN_IN), .Z(n6854) );
  AOI22_X1 U8518 ( .A1(n8599), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n6853) );
  NAND2_X1 U8519 ( .A1(n6854), .A2(n6853), .ZN(P2_U3245) );
  NAND2_X1 U8520 ( .A1(n6947), .A2(n9913), .ZN(n9943) );
  AND2_X1 U8521 ( .A1(n6855), .A2(n6856), .ZN(n6860) );
  INV_X1 U8522 ( .A(n6855), .ZN(n6858) );
  INV_X1 U8523 ( .A(n6856), .ZN(n6857) );
  NAND2_X1 U8524 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  OAI21_X2 U8525 ( .B1(n6861), .B2(n6860), .A(n6859), .ZN(n7065) );
  NAND2_X1 U8526 ( .A1(n9287), .A2(n8412), .ZN(n6863) );
  NAND2_X1 U8527 ( .A1(n6947), .A2(n8406), .ZN(n6862) );
  NAND2_X1 U8528 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  XNOR2_X1 U8529 ( .A(n6864), .B(n6381), .ZN(n7063) );
  NAND2_X1 U8530 ( .A1(n9287), .A2(n8411), .ZN(n6866) );
  NAND2_X1 U8531 ( .A1(n6947), .A2(n8412), .ZN(n6865) );
  NAND2_X1 U8532 ( .A1(n6866), .A2(n6865), .ZN(n7064) );
  XNOR2_X1 U8533 ( .A(n7063), .B(n7064), .ZN(n6867) );
  XNOR2_X1 U8534 ( .A(n7065), .B(n6867), .ZN(n6868) );
  NAND2_X1 U8535 ( .A1(n6868), .A2(n9694), .ZN(n6874) );
  INV_X1 U8536 ( .A(n6869), .ZN(n6945) );
  OAI22_X1 U8537 ( .A1(n9699), .A2(n6945), .B1(n9271), .B2(n6870), .ZN(n6871)
         );
  AOI211_X1 U8538 ( .C1(n9222), .C2(n9286), .A(n6872), .B(n6871), .ZN(n6873)
         );
  OAI211_X1 U8539 ( .C1(n6931), .C2(n9943), .A(n6874), .B(n6873), .ZN(P1_U3219) );
  NAND2_X1 U8540 ( .A1(n8505), .A2(n6879), .ZN(n8255) );
  INV_X1 U8541 ( .A(n8505), .ZN(n8550) );
  NAND2_X1 U8542 ( .A1(n8550), .A2(n10004), .ZN(n8256) );
  NAND2_X1 U8543 ( .A1(n8255), .A2(n8256), .ZN(n8369) );
  XNOR2_X1 U8544 ( .A(n4379), .B(n8369), .ZN(n10008) );
  INV_X1 U8545 ( .A(n10008), .ZN(n6887) );
  NAND2_X1 U8546 ( .A1(n6968), .A2(n8250), .ZN(n6876) );
  XNOR2_X1 U8547 ( .A(n6876), .B(n8369), .ZN(n6877) );
  INV_X1 U8548 ( .A(n8986), .ZN(n9010) );
  OAI222_X1 U8549 ( .A1(n9012), .A2(n6878), .B1(n9014), .B2(n7287), .C1(n6877), 
        .C2(n9010), .ZN(n10006) );
  INV_X1 U8550 ( .A(n9022), .ZN(n8638) );
  NAND2_X1 U8551 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NAND2_X1 U8552 ( .A1(n4760), .A2(n6881), .ZN(n10005) );
  OAI22_X1 U8553 ( .A1(n8638), .A2(n10005), .B1(n6882), .B2(n8943), .ZN(n6883)
         );
  AOI21_X1 U8554 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n9019), .A(n6883), .ZN(
        n6884) );
  OAI21_X1 U8555 ( .B1(n10004), .B2(n9008), .A(n6884), .ZN(n6885) );
  AOI21_X1 U8556 ( .B1(n10006), .B2(n8946), .A(n6885), .ZN(n6886) );
  OAI21_X1 U8557 ( .B1(n9024), .B2(n6887), .A(n6886), .ZN(P2_U3289) );
  INV_X1 U8558 ( .A(n6888), .ZN(n7062) );
  OAI222_X1 U8559 ( .A1(n8405), .A2(n6889), .B1(n9165), .B2(n7062), .C1(n8388), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  XNOR2_X1 U8560 ( .A(n6890), .B(n7911), .ZN(n9929) );
  NOR2_X1 U8561 ( .A1(n9836), .A2(n6891), .ZN(n6892) );
  OR2_X1 U8562 ( .A1(n6893), .A2(n6892), .ZN(n9931) );
  AOI22_X1 U8563 ( .A1(n9555), .A2(n6930), .B1(n6934), .B2(n9826), .ZN(n6894)
         );
  OAI21_X1 U8564 ( .B1(n9931), .B2(n9440), .A(n6894), .ZN(n6901) );
  INV_X1 U8565 ( .A(n8057), .ZN(n7787) );
  OR2_X1 U8566 ( .A1(n6556), .A2(n7787), .ZN(n9841) );
  NAND2_X1 U8567 ( .A1(n7905), .A2(n9840), .ZN(n7903) );
  INV_X1 U8568 ( .A(n7903), .ZN(n7785) );
  NAND2_X1 U8569 ( .A1(n9841), .A2(n7785), .ZN(n6895) );
  NAND2_X1 U8570 ( .A1(n6895), .A2(n7904), .ZN(n6896) );
  XNOR2_X1 U8571 ( .A(n6896), .B(n7911), .ZN(n6897) );
  NAND2_X1 U8572 ( .A1(n6897), .A2(n9871), .ZN(n6899) );
  AOI22_X1 U8573 ( .A1(n9875), .A2(n9289), .B1(n9288), .B2(n9873), .ZN(n6898)
         );
  NAND2_X1 U8574 ( .A1(n6899), .A2(n6898), .ZN(n9933) );
  MUX2_X1 U8575 ( .A(n9933), .B(P1_REG2_REG_6__SCAN_IN), .S(n9856), .Z(n6900)
         );
  AOI211_X1 U8576 ( .C1(n9929), .C2(n9488), .A(n6901), .B(n6900), .ZN(n6902)
         );
  INV_X1 U8577 ( .A(n6902), .ZN(P1_U3285) );
  XNOR2_X1 U8578 ( .A(n6903), .B(n8360), .ZN(n10003) );
  INV_X1 U8579 ( .A(n10003), .ZN(n6915) );
  OAI211_X1 U8580 ( .C1(n10001), .C2(n6904), .A(n4376), .B(n9993), .ZN(n9999)
         );
  INV_X1 U8581 ( .A(n8220), .ZN(n6905) );
  OR2_X1 U8582 ( .A1(n6755), .A2(n6905), .ZN(n6907) );
  NAND2_X1 U8583 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8584 ( .A(n6908), .B(n8360), .ZN(n6909) );
  AOI222_X1 U8585 ( .A1(n8986), .A2(n6909), .B1(n8551), .B2(n8968), .C1(n8553), 
        .C2(n8965), .ZN(n10000) );
  OAI21_X1 U8586 ( .B1(n8623), .B2(n9999), .A(n10000), .ZN(n6913) );
  NOR2_X1 U8587 ( .A1(n9008), .A2(n10001), .ZN(n6912) );
  OAI22_X1 U8588 ( .A1(n8946), .A2(n5509), .B1(n6910), .B2(n8943), .ZN(n6911)
         );
  AOI211_X1 U8589 ( .C1(n6913), .C2(n8946), .A(n6912), .B(n6911), .ZN(n6914)
         );
  OAI21_X1 U8590 ( .B1(n6915), .B2(n9024), .A(n6914), .ZN(P2_U3291) );
  INV_X1 U8591 ( .A(n6916), .ZN(n6917) );
  AOI211_X1 U8592 ( .C1(n6919), .C2(n6918), .A(n8518), .B(n6917), .ZN(n6923)
         );
  INV_X1 U8593 ( .A(n9013), .ZN(n8651) );
  AOI22_X1 U8594 ( .A1(n8511), .A2(n8548), .B1(n8496), .B2(n8651), .ZN(n6921)
         );
  AOI22_X1 U8595 ( .A1(n8508), .A2(n9127), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n6920) );
  OAI211_X1 U8596 ( .C1(n7568), .C2(n8537), .A(n6921), .B(n6920), .ZN(n6922)
         );
  OR2_X1 U8597 ( .A1(n6923), .A2(n6922), .ZN(P2_U3219) );
  AOI21_X1 U8598 ( .B1(n6925), .B2(n6768), .A(n6924), .ZN(n6929) );
  XNOR2_X1 U8599 ( .A(n6927), .B(n6926), .ZN(n6928) );
  XNOR2_X1 U8600 ( .A(n6929), .B(n6928), .ZN(n6937) );
  AOI22_X1 U8601 ( .A1(n9685), .A2(n9289), .B1(n9222), .B2(n9288), .ZN(n6936)
         );
  NAND2_X1 U8602 ( .A1(n9913), .A2(n6930), .ZN(n9930) );
  NOR2_X1 U8603 ( .A1(n6931), .A2(n9930), .ZN(n6932) );
  AOI211_X1 U8604 ( .C1(n6934), .C2(n9259), .A(n6933), .B(n6932), .ZN(n6935)
         );
  OAI211_X1 U8605 ( .C1(n6937), .C2(n9278), .A(n6936), .B(n6935), .ZN(P1_U3237) );
  XNOR2_X1 U8606 ( .A(n6938), .B(n7872), .ZN(n6939) );
  AOI222_X1 U8607 ( .A1(n9871), .A2(n6939), .B1(n9286), .B2(n9873), .C1(n9288), 
        .C2(n9875), .ZN(n9944) );
  INV_X1 U8608 ( .A(n6940), .ZN(n6941) );
  AOI21_X1 U8609 ( .B1(n7872), .B2(n6942), .A(n6941), .ZN(n9949) );
  NAND2_X1 U8610 ( .A1(n6943), .A2(n6947), .ZN(n6944) );
  NAND2_X1 U8611 ( .A1(n7303), .A2(n6944), .ZN(n9945) );
  OAI22_X1 U8612 ( .A1(n9884), .A2(n6156), .B1(n6945), .B2(n9880), .ZN(n6946)
         );
  AOI21_X1 U8613 ( .B1(n9555), .B2(n6947), .A(n6946), .ZN(n6948) );
  OAI21_X1 U8614 ( .B1(n9945), .B2(n9440), .A(n6948), .ZN(n6949) );
  AOI21_X1 U8615 ( .B1(n9949), .B2(n9488), .A(n6949), .ZN(n6950) );
  OAI21_X1 U8616 ( .B1(n9856), .B2(n9944), .A(n6950), .ZN(P1_U3283) );
  NOR2_X1 U8617 ( .A1(n8943), .A2(n7450), .ZN(n6955) );
  NAND2_X1 U8618 ( .A1(n8946), .A2(n6951), .ZN(n6952) );
  OAI21_X1 U8619 ( .B1(n8946), .B2(n6953), .A(n6952), .ZN(n6954) );
  AOI211_X1 U8620 ( .C1(n9022), .C2(n6956), .A(n6955), .B(n6954), .ZN(n6960)
         );
  AOI22_X1 U8621 ( .A1(n8892), .A2(n6958), .B1(n8940), .B2(n6957), .ZN(n6959)
         );
  NAND2_X1 U8622 ( .A1(n6960), .A2(n6959), .ZN(P2_U3294) );
  XNOR2_X1 U8623 ( .A(n8549), .B(n7285), .ZN(n8371) );
  NAND2_X1 U8624 ( .A1(n8505), .A2(n10004), .ZN(n6961) );
  NAND2_X1 U8625 ( .A1(n6962), .A2(n6961), .ZN(n6965) );
  INV_X1 U8626 ( .A(n6965), .ZN(n6963) );
  NAND2_X1 U8627 ( .A1(n6963), .A2(n4408), .ZN(n7283) );
  INV_X1 U8628 ( .A(n7283), .ZN(n6964) );
  AOI21_X1 U8629 ( .B1(n8371), .B2(n6965), .A(n6964), .ZN(n7248) );
  INV_X1 U8630 ( .A(n8982), .ZN(n8883) );
  INV_X1 U8631 ( .A(n8250), .ZN(n6966) );
  NOR2_X1 U8632 ( .A1(n8369), .A2(n6966), .ZN(n6967) );
  NAND2_X1 U8633 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  NAND2_X1 U8634 ( .A1(n6970), .A2(n4408), .ZN(n6971) );
  AOI21_X1 U8635 ( .B1(n7286), .B2(n6971), .A(n9010), .ZN(n6973) );
  OAI22_X1 U8636 ( .A1(n7557), .A2(n9014), .B1(n8505), .B2(n9012), .ZN(n6972)
         );
  AOI211_X1 U8637 ( .C1(n7248), .C2(n8883), .A(n6973), .B(n6972), .ZN(n7251)
         );
  INV_X1 U8638 ( .A(n6974), .ZN(n6975) );
  NAND2_X1 U8639 ( .A1(n8946), .A2(n6975), .ZN(n8992) );
  INV_X1 U8640 ( .A(n8992), .ZN(n6981) );
  AND2_X1 U8641 ( .A1(n4760), .A2(n7285), .ZN(n6976) );
  NOR2_X1 U8642 ( .A1(n7293), .A2(n6976), .ZN(n7249) );
  INV_X1 U8643 ( .A(n8943), .ZN(n9005) );
  AOI22_X1 U8644 ( .A1(n7249), .A2(n8995), .B1(n6977), .B2(n9005), .ZN(n6979)
         );
  NAND2_X1 U8645 ( .A1(n9019), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6978) );
  OAI211_X1 U8646 ( .C1(n8259), .C2(n9008), .A(n6979), .B(n6978), .ZN(n6980)
         );
  AOI21_X1 U8647 ( .B1(n7248), .B2(n6981), .A(n6980), .ZN(n6982) );
  OAI21_X1 U8648 ( .B1(n7251), .B2(n9019), .A(n6982), .ZN(P2_U3288) );
  OAI21_X1 U8649 ( .B1(n6983), .B2(n6985), .A(n6984), .ZN(n9990) );
  INV_X1 U8650 ( .A(n9990), .ZN(n6996) );
  INV_X1 U8651 ( .A(n6986), .ZN(n9984) );
  NAND2_X1 U8652 ( .A1(n9979), .A2(n6990), .ZN(n9983) );
  NAND3_X1 U8653 ( .A1(n8995), .A2(n9984), .A3(n9983), .ZN(n6987) );
  OAI21_X1 U8654 ( .B1(n8943), .B2(n6988), .A(n6987), .ZN(n6989) );
  AOI21_X1 U8655 ( .B1(n8892), .B2(n6990), .A(n6989), .ZN(n6995) );
  XNOR2_X1 U8656 ( .A(n6983), .B(n7023), .ZN(n6992) );
  AOI21_X1 U8657 ( .B1(n6992), .B2(n8986), .A(n6991), .ZN(n9987) );
  MUX2_X1 U8658 ( .A(n6993), .B(n9987), .S(n8946), .Z(n6994) );
  OAI211_X1 U8659 ( .C1(n6996), .C2(n9024), .A(n6995), .B(n6994), .ZN(P2_U3295) );
  INV_X1 U8660 ( .A(n6997), .ZN(n6998) );
  AOI21_X1 U8661 ( .B1(n6841), .B2(n6998), .A(n8518), .ZN(n7002) );
  NOR3_X1 U8662 ( .A1(n8516), .A2(n6999), .A3(n9013), .ZN(n7001) );
  OAI21_X1 U8663 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7006) );
  OAI22_X1 U8664 ( .A1(n8539), .A2(n9015), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7237), .ZN(n7004) );
  OAI22_X1 U8665 ( .A1(n8536), .A2(n9013), .B1(n8537), .B2(n9004), .ZN(n7003)
         );
  AOI211_X1 U8666 ( .C1(n9121), .C2(n8508), .A(n7004), .B(n7003), .ZN(n7005)
         );
  NAND2_X1 U8667 ( .A1(n7006), .A2(n7005), .ZN(P2_U3226) );
  INV_X1 U8668 ( .A(n7007), .ZN(n7008) );
  OAI22_X1 U8669 ( .A1(n7008), .A2(n8638), .B1(n8504), .B2(n8943), .ZN(n7009)
         );
  AOI21_X1 U8670 ( .B1(n8892), .B2(n4310), .A(n7009), .ZN(n7012) );
  MUX2_X1 U8671 ( .A(n6676), .B(n7010), .S(n8946), .Z(n7011) );
  OAI211_X1 U8672 ( .C1(n7013), .C2(n9024), .A(n7012), .B(n7011), .ZN(P2_U3290) );
  NAND2_X1 U8673 ( .A1(n8995), .A2(n7014), .ZN(n7015) );
  OAI21_X1 U8674 ( .B1(n8943), .B2(n7016), .A(n7015), .ZN(n7020) );
  OAI22_X1 U8675 ( .A1(n7018), .A2(n9024), .B1(n7017), .B2(n9008), .ZN(n7019)
         );
  AOI211_X1 U8676 ( .C1(n9019), .C2(P2_REG2_REG_4__SCAN_IN), .A(n7020), .B(
        n7019), .ZN(n7021) );
  OAI21_X1 U8677 ( .B1(n9019), .B2(n7022), .A(n7021), .ZN(P2_U3292) );
  NAND2_X1 U8678 ( .A1(n7023), .A2(n8227), .ZN(n9980) );
  INV_X1 U8679 ( .A(n9980), .ZN(n7027) );
  AOI22_X1 U8680 ( .A1(n9980), .A2(n8986), .B1(n8968), .B2(n6483), .ZN(n9982)
         );
  OAI22_X1 U8681 ( .A1(n9019), .A2(n9982), .B1(n5529), .B2(n8943), .ZN(n7024)
         );
  AOI21_X1 U8682 ( .B1(n9019), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7024), .ZN(
        n7026) );
  OAI21_X1 U8683 ( .B1(n8892), .B2(n9022), .A(n9979), .ZN(n7025) );
  OAI211_X1 U8684 ( .C1(n7027), .C2(n9024), .A(n7026), .B(n7025), .ZN(P2_U3296) );
  INV_X1 U8685 ( .A(n7090), .ZN(n7030) );
  AOI21_X1 U8686 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9162), .A(n7028), .ZN(
        n7029) );
  OAI21_X1 U8687 ( .B1(n7030), .B2(n9165), .A(n7029), .ZN(P2_U3335) );
  INV_X1 U8688 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9293) );
  AOI22_X1 U8689 ( .A1(n7031), .A2(n9293), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9296), .ZN(n7039) );
  INV_X1 U8690 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7037) );
  XNOR2_X1 U8691 ( .A(n9807), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9815) );
  INV_X1 U8692 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7036) );
  XOR2_X1 U8693 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7044), .Z(n9799) );
  AOI21_X1 U8694 ( .B1(n7033), .B2(n9718), .A(n7032), .ZN(n7034) );
  NAND2_X1 U8695 ( .A1(n9784), .A2(n7034), .ZN(n7035) );
  XOR2_X1 U8696 ( .A(n9784), .B(n7034), .Z(n9789) );
  NAND2_X1 U8697 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9789), .ZN(n9788) );
  NAND2_X1 U8698 ( .A1(n7035), .A2(n9788), .ZN(n9800) );
  NAND2_X1 U8699 ( .A1(n9799), .A2(n9800), .ZN(n9798) );
  OAI21_X1 U8700 ( .B1(n9795), .B2(n7036), .A(n9798), .ZN(n9814) );
  NAND2_X1 U8701 ( .A1(n9815), .A2(n9814), .ZN(n9812) );
  OAI21_X1 U8702 ( .B1(n7037), .B2(n9807), .A(n9812), .ZN(n7038) );
  NOR2_X1 U8703 ( .A1(n7039), .A2(n7038), .ZN(n9292) );
  AOI21_X1 U8704 ( .B1(n7039), .B2(n7038), .A(n9292), .ZN(n7060) );
  NAND2_X1 U8705 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9260) );
  OAI21_X1 U8706 ( .B1(n9808), .B2(n9296), .A(n9260), .ZN(n7040) );
  AOI21_X1 U8707 ( .B1(n9811), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n7040), .ZN(
        n7058) );
  NAND2_X1 U8708 ( .A1(n7041), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7054) );
  INV_X1 U8709 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7043) );
  INV_X1 U8710 ( .A(n7054), .ZN(n7042) );
  AOI21_X1 U8711 ( .B1(n7043), .B2(n9807), .A(n7042), .ZN(n9818) );
  NAND2_X1 U8712 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7044), .ZN(n7053) );
  INV_X1 U8713 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7046) );
  INV_X1 U8714 ( .A(n7053), .ZN(n7045) );
  AOI21_X1 U8715 ( .B1(n7046), .B2(n9795), .A(n7045), .ZN(n9802) );
  NAND2_X1 U8716 ( .A1(n7048), .A2(n7047), .ZN(n7050) );
  NAND2_X1 U8717 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8718 ( .A1(n9784), .A2(n7051), .ZN(n7052) );
  XOR2_X1 U8719 ( .A(n9784), .B(n7051), .Z(n9791) );
  NAND2_X1 U8720 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9791), .ZN(n9790) );
  NAND2_X1 U8721 ( .A1(n7052), .A2(n9790), .ZN(n9803) );
  NAND2_X1 U8722 ( .A1(n9802), .A2(n9803), .ZN(n9801) );
  NAND2_X1 U8723 ( .A1(n7053), .A2(n9801), .ZN(n9819) );
  NAND2_X1 U8724 ( .A1(n9818), .A2(n9819), .ZN(n9816) );
  NAND2_X1 U8725 ( .A1(n7054), .A2(n9816), .ZN(n7056) );
  XNOR2_X1 U8726 ( .A(n9296), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8727 ( .A1(n7055), .A2(n7056), .ZN(n9295) );
  OAI211_X1 U8728 ( .C1(n7056), .C2(n7055), .A(n9817), .B(n9295), .ZN(n7057)
         );
  OAI211_X1 U8729 ( .C1(n7060), .C2(n7059), .A(n7058), .B(n7057), .ZN(P1_U3259) );
  OAI222_X1 U8730 ( .A1(P1_U3084), .A2(n5346), .B1(n9671), .B2(n7062), .C1(
        n7061), .C2(n7753), .ZN(P1_U3331) );
  NAND2_X1 U8731 ( .A1(n9827), .A2(n8406), .ZN(n7067) );
  NAND2_X1 U8732 ( .A1(n9286), .A2(n8412), .ZN(n7066) );
  NAND2_X1 U8733 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  XNOR2_X1 U8734 ( .A(n7068), .B(n4311), .ZN(n7070) );
  AOI22_X1 U8735 ( .A1(n9827), .A2(n8412), .B1(n8411), .B2(n9286), .ZN(n7069)
         );
  NAND2_X1 U8736 ( .A1(n7070), .A2(n7069), .ZN(n7203) );
  OR2_X1 U8737 ( .A1(n7070), .A2(n7069), .ZN(n7071) );
  NAND2_X1 U8738 ( .A1(n7203), .A2(n7071), .ZN(n7185) );
  OR2_X1 U8739 ( .A1(n7206), .A2(n7185), .ZN(n7153) );
  NAND2_X1 U8740 ( .A1(n7153), .A2(n7203), .ZN(n7082) );
  NAND2_X1 U8741 ( .A1(n9672), .A2(n8406), .ZN(n7073) );
  NAND2_X1 U8742 ( .A1(n9285), .A2(n8412), .ZN(n7072) );
  NAND2_X1 U8743 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  XNOR2_X1 U8744 ( .A(n7074), .B(n6381), .ZN(n7077) );
  NAND2_X1 U8745 ( .A1(n9672), .A2(n8412), .ZN(n7076) );
  NAND2_X1 U8746 ( .A1(n9285), .A2(n8411), .ZN(n7075) );
  NAND2_X1 U8747 ( .A1(n7076), .A2(n7075), .ZN(n7078) );
  NAND2_X1 U8748 ( .A1(n7077), .A2(n7078), .ZN(n7184) );
  INV_X1 U8749 ( .A(n7077), .ZN(n7080) );
  INV_X1 U8750 ( .A(n7078), .ZN(n7079) );
  NAND2_X1 U8751 ( .A1(n7080), .A2(n7079), .ZN(n7272) );
  NAND2_X1 U8752 ( .A1(n7184), .A2(n7272), .ZN(n7081) );
  XNOR2_X1 U8753 ( .A(n7082), .B(n7081), .ZN(n7089) );
  INV_X1 U8754 ( .A(n7083), .ZN(n7264) );
  OAI22_X1 U8755 ( .A1(n9699), .A2(n7264), .B1(n9271), .B2(n7084), .ZN(n7085)
         );
  AOI211_X1 U8756 ( .C1(n9222), .C2(n9684), .A(n7086), .B(n7085), .ZN(n7088)
         );
  NAND2_X1 U8757 ( .A1(n9276), .A2(n9672), .ZN(n7087) );
  OAI211_X1 U8758 ( .C1(n7089), .C2(n9278), .A(n7088), .B(n7087), .ZN(P1_U3215) );
  NAND2_X1 U8759 ( .A1(n7090), .A2(n7748), .ZN(n7092) );
  NAND2_X1 U8760 ( .A1(n7091), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8086) );
  OAI211_X1 U8761 ( .C1(n7093), .C2(n9667), .A(n7092), .B(n8086), .ZN(P1_U3330) );
  AOI211_X1 U8762 ( .C1(n7096), .C2(n7095), .A(n7094), .B(n7710), .ZN(n7105)
         );
  NOR2_X1 U8763 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7463), .ZN(n7097) );
  AOI21_X1 U8764 ( .B1(n8599), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7097), .ZN(
        n7102) );
  OAI211_X1 U8765 ( .C1(n7100), .C2(n7099), .A(n8612), .B(n7098), .ZN(n7101)
         );
  OAI211_X1 U8766 ( .C1(n8619), .C2(n7103), .A(n7102), .B(n7101), .ZN(n7104)
         );
  OR2_X1 U8767 ( .A1(n7105), .A2(n7104), .ZN(P2_U3255) );
  AOI211_X1 U8768 ( .C1(n7108), .C2(n7107), .A(n7106), .B(n7710), .ZN(n7117)
         );
  NOR2_X1 U8769 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7434), .ZN(n7109) );
  AOI21_X1 U8770 ( .B1(n8599), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7109), .ZN(
        n7114) );
  OAI211_X1 U8771 ( .C1(n7112), .C2(n7111), .A(n8612), .B(n7110), .ZN(n7113)
         );
  OAI211_X1 U8772 ( .C1(n8619), .C2(n7115), .A(n7114), .B(n7113), .ZN(n7116)
         );
  OR2_X1 U8773 ( .A1(n7117), .A2(n7116), .ZN(P2_U3253) );
  AOI211_X1 U8774 ( .C1(n7120), .C2(n7119), .A(n7118), .B(n7710), .ZN(n7128)
         );
  AND2_X1 U8775 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8507) );
  AOI21_X1 U8776 ( .B1(n8599), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8507), .ZN(
        n7125) );
  OAI211_X1 U8777 ( .C1(n7123), .C2(n7122), .A(n8612), .B(n7121), .ZN(n7124)
         );
  OAI211_X1 U8778 ( .C1(n8619), .C2(n7126), .A(n7125), .B(n7124), .ZN(n7127)
         );
  OR2_X1 U8779 ( .A1(n7128), .A2(n7127), .ZN(P2_U3251) );
  AOI211_X1 U8780 ( .C1(n7131), .C2(n7130), .A(n7129), .B(n7710), .ZN(n7140)
         );
  AOI21_X1 U8781 ( .B1(n8599), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7132), .ZN(
        n7137) );
  OAI211_X1 U8782 ( .C1(n7135), .C2(n7134), .A(n8612), .B(n7133), .ZN(n7136)
         );
  OAI211_X1 U8783 ( .C1(n8619), .C2(n7138), .A(n7137), .B(n7136), .ZN(n7139)
         );
  OR2_X1 U8784 ( .A1(n7140), .A2(n7139), .ZN(P2_U3254) );
  AOI211_X1 U8785 ( .C1(n7143), .C2(n7142), .A(n7141), .B(n7710), .ZN(n7152)
         );
  NOR2_X1 U8786 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5452), .ZN(n7144) );
  AOI21_X1 U8787 ( .B1(n8599), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7144), .ZN(
        n7149) );
  OAI211_X1 U8788 ( .C1(n7147), .C2(n7146), .A(n8612), .B(n7145), .ZN(n7148)
         );
  OAI211_X1 U8789 ( .C1(n8619), .C2(n7150), .A(n7149), .B(n7148), .ZN(n7151)
         );
  OR2_X1 U8790 ( .A1(n7152), .A2(n7151), .ZN(P2_U3252) );
  INV_X1 U8791 ( .A(n7153), .ZN(n7154) );
  AOI21_X1 U8792 ( .B1(n7185), .B2(n7206), .A(n7154), .ZN(n7160) );
  INV_X1 U8793 ( .A(n9825), .ZN(n7155) );
  OAI22_X1 U8794 ( .A1(n9699), .A2(n7155), .B1(n9271), .B2(n7306), .ZN(n7156)
         );
  AOI211_X1 U8795 ( .C1(n9222), .C2(n9285), .A(n7157), .B(n7156), .ZN(n7159)
         );
  NAND2_X1 U8796 ( .A1(n9276), .A2(n9827), .ZN(n7158) );
  OAI211_X1 U8797 ( .C1(n7160), .C2(n9278), .A(n7159), .B(n7158), .ZN(P1_U3229) );
  OAI21_X1 U8798 ( .B1(n7162), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7161), .ZN(
        n7628) );
  XNOR2_X1 U8799 ( .A(n7628), .B(n7623), .ZN(n7163) );
  NAND2_X1 U8800 ( .A1(n7163), .A2(n8945), .ZN(n7630) );
  OAI21_X1 U8801 ( .B1(n7163), .B2(n8945), .A(n7630), .ZN(n7172) );
  AOI21_X1 U8802 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7622) );
  XNOR2_X1 U8803 ( .A(n7622), .B(n7629), .ZN(n7167) );
  NAND2_X1 U8804 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7167), .ZN(n7624) );
  OAI211_X1 U8805 ( .C1(n7167), .C2(P2_REG1_REG_15__SCAN_IN), .A(n8612), .B(
        n7624), .ZN(n7170) );
  NOR2_X1 U8806 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5741), .ZN(n7168) );
  AOI21_X1 U8807 ( .B1(n8599), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7168), .ZN(
        n7169) );
  OAI211_X1 U8808 ( .C1(n8619), .C2(n7629), .A(n7170), .B(n7169), .ZN(n7171)
         );
  AOI21_X1 U8809 ( .B1(n8613), .B2(n7172), .A(n7171), .ZN(n7173) );
  INV_X1 U8810 ( .A(n7173), .ZN(P2_U3260) );
  INV_X1 U8811 ( .A(n7174), .ZN(n7175) );
  AOI21_X1 U8812 ( .B1(n7000), .B2(n7175), .A(n8518), .ZN(n7179) );
  NOR3_X1 U8813 ( .A1(n8516), .A2(n7176), .A3(n8978), .ZN(n7178) );
  OAI21_X1 U8814 ( .B1(n7179), .B2(n7178), .A(n7177), .ZN(n7183) );
  OAI22_X1 U8815 ( .A1(n8539), .A2(n8977), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6743), .ZN(n7181) );
  OAI22_X1 U8816 ( .A1(n8536), .A2(n8978), .B1(n8537), .B2(n8988), .ZN(n7180)
         );
  AOI211_X1 U8817 ( .C1(n9116), .C2(n8508), .A(n7181), .B(n7180), .ZN(n7182)
         );
  NAND2_X1 U8818 ( .A1(n7183), .A2(n7182), .ZN(P2_U3236) );
  INV_X1 U8819 ( .A(n7702), .ZN(n9638) );
  INV_X1 U8820 ( .A(n7184), .ZN(n7204) );
  OR2_X1 U8821 ( .A1(n7185), .A2(n7204), .ZN(n7269) );
  INV_X1 U8822 ( .A(n7192), .ZN(n7190) );
  AND2_X1 U8823 ( .A1(n9284), .A2(n8411), .ZN(n7189) );
  AOI21_X1 U8824 ( .B1(n7187), .B2(n6395), .A(n7189), .ZN(n7191) );
  NAND2_X1 U8825 ( .A1(n7190), .A2(n7191), .ZN(n7202) );
  NAND2_X1 U8826 ( .A1(n7641), .A2(n8406), .ZN(n7194) );
  NAND2_X1 U8827 ( .A1(n9684), .A2(n8412), .ZN(n7193) );
  NAND2_X1 U8828 ( .A1(n7194), .A2(n7193), .ZN(n7195) );
  XNOR2_X1 U8829 ( .A(n7195), .B(n4311), .ZN(n7200) );
  INV_X1 U8830 ( .A(n7200), .ZN(n7198) );
  AND2_X1 U8831 ( .A1(n9684), .A2(n8411), .ZN(n7196) );
  AOI21_X1 U8832 ( .B1(n7641), .B2(n8412), .A(n7196), .ZN(n7199) );
  INV_X1 U8833 ( .A(n7199), .ZN(n7197) );
  NAND2_X1 U8834 ( .A1(n7198), .A2(n7197), .ZN(n9686) );
  AND2_X1 U8835 ( .A1(n7275), .A2(n7202), .ZN(n7205) );
  OR2_X1 U8836 ( .A1(n7204), .A2(n7203), .ZN(n7270) );
  AND2_X1 U8837 ( .A1(n9549), .A2(n8411), .ZN(n7207) );
  AOI21_X1 U8838 ( .B1(n7702), .B2(n6395), .A(n7207), .ZN(n7541) );
  NAND2_X1 U8839 ( .A1(n7702), .A2(n8406), .ZN(n7209) );
  NAND2_X1 U8840 ( .A1(n9549), .A2(n8412), .ZN(n7208) );
  NAND2_X1 U8841 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  XNOR2_X1 U8842 ( .A(n7210), .B(n4311), .ZN(n7542) );
  XOR2_X1 U8843 ( .A(n7541), .B(n7542), .Z(n7211) );
  XNOR2_X1 U8844 ( .A(n7545), .B(n7211), .ZN(n7212) );
  NAND2_X1 U8845 ( .A1(n7212), .A2(n9694), .ZN(n7218) );
  INV_X1 U8846 ( .A(n7701), .ZN(n7214) );
  OAI22_X1 U8847 ( .A1(n9699), .A2(n7214), .B1(n9271), .B2(n7213), .ZN(n7215)
         );
  AOI211_X1 U8848 ( .C1(n9222), .C2(n9283), .A(n7216), .B(n7215), .ZN(n7217)
         );
  OAI211_X1 U8849 ( .C1(n9638), .C2(n9224), .A(n7218), .B(n7217), .ZN(P1_U3232) );
  INV_X1 U8850 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7224) );
  MUX2_X1 U8851 ( .A(n6695), .B(P2_REG1_REG_1__SCAN_IN), .S(n7232), .Z(n7219)
         );
  OAI21_X1 U8852 ( .B1(n6848), .B2(n4415), .A(n7219), .ZN(n7220) );
  NAND3_X1 U8853 ( .A1(n8612), .A2(n7221), .A3(n7220), .ZN(n7223) );
  NAND2_X1 U8854 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7222) );
  OAI211_X1 U8855 ( .C1(n8629), .C2(n7224), .A(n7223), .B(n7222), .ZN(n7231)
         );
  NAND2_X1 U8856 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n7229) );
  INV_X1 U8857 ( .A(n7225), .ZN(n7228) );
  INV_X1 U8858 ( .A(n7226), .ZN(n7227) );
  AOI211_X1 U8859 ( .C1(n7229), .C2(n7228), .A(n7227), .B(n7710), .ZN(n7230)
         );
  AOI211_X1 U8860 ( .C1(n8562), .C2(n7232), .A(n7231), .B(n7230), .ZN(n7233)
         );
  INV_X1 U8861 ( .A(n7233), .ZN(P2_U3246) );
  AOI21_X1 U8862 ( .B1(n7236), .B2(n7235), .A(n7234), .ZN(n7240) );
  NOR2_X1 U8863 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7237), .ZN(n7238) );
  AOI21_X1 U8864 ( .B1(n8599), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7238), .ZN(
        n7239) );
  OAI21_X1 U8865 ( .B1(n8620), .B2(n7240), .A(n7239), .ZN(n7245) );
  AOI211_X1 U8866 ( .C1(n7243), .C2(n7242), .A(n7241), .B(n7710), .ZN(n7244)
         );
  AOI211_X1 U8867 ( .C1(n8562), .C2(n7246), .A(n7245), .B(n7244), .ZN(n7247)
         );
  INV_X1 U8868 ( .A(n7247), .ZN(P2_U3257) );
  INV_X1 U8869 ( .A(n7248), .ZN(n7252) );
  AOI22_X1 U8870 ( .A1(n7249), .A2(n9993), .B1(n9992), .B2(n7285), .ZN(n7250)
         );
  OAI211_X1 U8871 ( .C1(n10009), .C2(n7252), .A(n7251), .B(n7250), .ZN(n7254)
         );
  NAND2_X1 U8872 ( .A1(n7254), .A2(n10017), .ZN(n7253) );
  OAI21_X1 U8873 ( .B1(n10017), .B2(n5603), .A(n7253), .ZN(P2_U3475) );
  NAND2_X1 U8874 ( .A1(n7254), .A2(n10039), .ZN(n7255) );
  OAI21_X1 U8875 ( .B1(n10039), .B2(n7256), .A(n7255), .ZN(P2_U3528) );
  INV_X1 U8876 ( .A(n7257), .ZN(n7925) );
  NAND2_X1 U8877 ( .A1(n7258), .A2(n7925), .ZN(n7259) );
  XNOR2_X1 U8878 ( .A(n7259), .B(n7874), .ZN(n7260) );
  AOI222_X1 U8879 ( .A1(n9871), .A2(n7260), .B1(n9684), .B2(n9873), .C1(n9286), 
        .C2(n9875), .ZN(n9674) );
  OAI21_X1 U8880 ( .B1(n7262), .B2(n5085), .A(n7261), .ZN(n9676) );
  AOI21_X1 U8881 ( .B1(n7301), .B2(n9672), .A(n9946), .ZN(n7263) );
  NAND2_X1 U8882 ( .A1(n4377), .A2(n7263), .ZN(n9673) );
  OAI22_X1 U8883 ( .A1(n9884), .A2(n6225), .B1(n7264), .B2(n9880), .ZN(n7265)
         );
  AOI21_X1 U8884 ( .B1(n9555), .B2(n9672), .A(n7265), .ZN(n7266) );
  OAI21_X1 U8885 ( .B1(n9673), .B2(n9559), .A(n7266), .ZN(n7267) );
  AOI21_X1 U8886 ( .B1(n9676), .B2(n9488), .A(n7267), .ZN(n7268) );
  OAI21_X1 U8887 ( .B1(n9674), .B2(n9856), .A(n7268), .ZN(P1_U3281) );
  OR2_X1 U8888 ( .A1(n7206), .A2(n7269), .ZN(n7271) );
  AND2_X1 U8889 ( .A1(n7271), .A2(n7270), .ZN(n7276) );
  NAND2_X1 U8890 ( .A1(n7276), .A2(n7272), .ZN(n7274) );
  AOI21_X1 U8891 ( .B1(n7274), .B2(n7273), .A(n9278), .ZN(n7277) );
  NAND2_X1 U8892 ( .A1(n7276), .A2(n7275), .ZN(n9688) );
  NAND2_X1 U8893 ( .A1(n7277), .A2(n9688), .ZN(n7281) );
  OAI22_X1 U8894 ( .A1(n9699), .A2(n7318), .B1(n9271), .B2(n7307), .ZN(n7278)
         );
  AOI211_X1 U8895 ( .C1(n9222), .C2(n9284), .A(n7279), .B(n7278), .ZN(n7280)
         );
  OAI211_X1 U8896 ( .C1(n7317), .C2(n9224), .A(n7281), .B(n7280), .ZN(P1_U3234) );
  NAND2_X1 U8897 ( .A1(n10011), .A2(n8548), .ZN(n8268) );
  NAND2_X1 U8898 ( .A1(n7297), .A2(n7557), .ZN(n8265) );
  NAND2_X1 U8899 ( .A1(n8549), .A2(n7285), .ZN(n7282) );
  NAND2_X1 U8900 ( .A1(n7283), .A2(n7282), .ZN(n8656) );
  INV_X1 U8901 ( .A(n7558), .ZN(n7284) );
  AOI21_X1 U8902 ( .B1(n8655), .B2(n8656), .A(n7284), .ZN(n10010) );
  NAND2_X1 U8903 ( .A1(n7287), .A2(n7285), .ZN(n8261) );
  XNOR2_X1 U8904 ( .A(n7562), .B(n8655), .ZN(n7289) );
  OAI22_X1 U8905 ( .A1(n7287), .A2(n9012), .B1(n7600), .B2(n9014), .ZN(n7288)
         );
  AOI21_X1 U8906 ( .B1(n7289), .B2(n8986), .A(n7288), .ZN(n7290) );
  OAI21_X1 U8907 ( .B1(n10010), .B2(n8982), .A(n7290), .ZN(n10013) );
  NAND2_X1 U8908 ( .A1(n10013), .A2(n8946), .ZN(n7299) );
  OAI22_X1 U8909 ( .A1(n8946), .A2(n7292), .B1(n7291), .B2(n8943), .ZN(n7296)
         );
  NOR2_X1 U8910 ( .A1(n7293), .A2(n10011), .ZN(n7294) );
  OR2_X1 U8911 ( .A1(n7572), .A2(n7294), .ZN(n10012) );
  NOR2_X1 U8912 ( .A1(n10012), .A2(n8638), .ZN(n7295) );
  AOI211_X1 U8913 ( .C1(n8892), .C2(n7297), .A(n7296), .B(n7295), .ZN(n7298)
         );
  OAI211_X1 U8914 ( .C1(n10010), .C2(n8992), .A(n7299), .B(n7298), .ZN(
        P2_U3287) );
  AND2_X1 U8915 ( .A1(n7925), .A2(n7927), .ZN(n7873) );
  XOR2_X1 U8916 ( .A(n7873), .B(n7300), .Z(n9823) );
  INV_X1 U8917 ( .A(n7301), .ZN(n7302) );
  AOI211_X1 U8918 ( .C1(n9827), .C2(n7303), .A(n9946), .B(n7302), .ZN(n9824)
         );
  XNOR2_X1 U8919 ( .A(n7304), .B(n7873), .ZN(n7305) );
  OAI222_X1 U8920 ( .A1(n9531), .A2(n7307), .B1(n9529), .B2(n7306), .C1(n9527), 
        .C2(n7305), .ZN(n9831) );
  AOI211_X1 U8921 ( .C1(n9913), .C2(n9827), .A(n9824), .B(n9831), .ZN(n7308)
         );
  OAI21_X1 U8922 ( .B1(n9922), .B2(n9823), .A(n7308), .ZN(n7311) );
  NAND2_X1 U8923 ( .A1(n7311), .A2(n9968), .ZN(n7309) );
  OAI21_X1 U8924 ( .B1(n9968), .B2(n7310), .A(n7309), .ZN(P1_U3532) );
  INV_X1 U8925 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U8926 ( .A1(n7311), .A2(n9952), .ZN(n7312) );
  OAI21_X1 U8927 ( .B1(n9952), .B2(n7313), .A(n7312), .ZN(P1_U3481) );
  XNOR2_X1 U8928 ( .A(n7314), .B(n7955), .ZN(n7645) );
  XNOR2_X1 U8929 ( .A(n7589), .B(n7955), .ZN(n7315) );
  AOI222_X1 U8930 ( .A1(n9871), .A2(n7315), .B1(n9284), .B2(n9873), .C1(n9285), 
        .C2(n9875), .ZN(n7644) );
  OR2_X1 U8931 ( .A1(n7644), .A2(n9856), .ZN(n7322) );
  INV_X1 U8932 ( .A(n7583), .ZN(n7316) );
  AOI21_X1 U8933 ( .B1(n7641), .B2(n4377), .A(n7316), .ZN(n7642) );
  NOR2_X1 U8934 ( .A1(n7317), .A2(n9539), .ZN(n7320) );
  OAI22_X1 U8935 ( .A1(n9884), .A2(n6235), .B1(n7318), .B2(n9880), .ZN(n7319)
         );
  AOI211_X1 U8936 ( .C1(n7642), .C2(n9504), .A(n7320), .B(n7319), .ZN(n7321)
         );
  OAI211_X1 U8937 ( .C1(n7645), .C2(n9855), .A(n7322), .B(n7321), .ZN(P1_U3280) );
  INV_X1 U8938 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U8939 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7323) );
  AOI21_X1 U8940 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7323), .ZN(n10046) );
  NOR2_X1 U8941 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7324) );
  AOI21_X1 U8942 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7324), .ZN(n10049) );
  NOR2_X1 U8943 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7325) );
  AOI21_X1 U8944 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7325), .ZN(n10052) );
  NOR2_X1 U8945 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7326) );
  AOI21_X1 U8946 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7326), .ZN(n10055) );
  NOR2_X1 U8947 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7327) );
  AOI21_X1 U8948 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7327), .ZN(n10058) );
  INV_X1 U8949 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U8950 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7333) );
  INV_X1 U8951 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9783) );
  XOR2_X1 U8952 ( .A(n9783), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10086) );
  NAND2_X1 U8953 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7331) );
  XOR2_X1 U8954 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10084) );
  NAND2_X1 U8955 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7329) );
  XNOR2_X1 U8956 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9765), .ZN(n10072) );
  AOI21_X1 U8957 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10040) );
  NAND3_X1 U8958 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10042) );
  OAI21_X1 U8959 ( .B1(n10040), .B2(n7224), .A(n10042), .ZN(n10071) );
  NAND2_X1 U8960 ( .A1(n10072), .A2(n10071), .ZN(n7328) );
  NAND2_X1 U8961 ( .A1(n7329), .A2(n7328), .ZN(n10083) );
  NAND2_X1 U8962 ( .A1(n10084), .A2(n10083), .ZN(n7330) );
  NAND2_X1 U8963 ( .A1(n7331), .A2(n7330), .ZN(n10085) );
  NOR2_X1 U8964 ( .A1(n10086), .A2(n10085), .ZN(n7332) );
  NOR2_X1 U8965 ( .A1(n7333), .A2(n7332), .ZN(n10081) );
  NAND2_X1 U8966 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10081), .ZN(n7334) );
  NOR2_X1 U8967 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10081), .ZN(n10080) );
  AOI21_X1 U8968 ( .B1(n7335), .B2(n7334), .A(n10080), .ZN(n7336) );
  NAND2_X1 U8969 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7336), .ZN(n7338) );
  XOR2_X1 U8970 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7336), .Z(n10079) );
  NAND2_X1 U8971 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10079), .ZN(n7337) );
  NAND2_X1 U8972 ( .A1(n7338), .A2(n7337), .ZN(n7339) );
  NAND2_X1 U8973 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7339), .ZN(n7341) );
  XOR2_X1 U8974 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7339), .Z(n10078) );
  NAND2_X1 U8975 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10078), .ZN(n7340) );
  NAND2_X1 U8976 ( .A1(n7341), .A2(n7340), .ZN(n7342) );
  NAND2_X1 U8977 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7342), .ZN(n7344) );
  XOR2_X1 U8978 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7342), .Z(n10073) );
  NAND2_X1 U8979 ( .A1(n10073), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U8980 ( .A1(n7344), .A2(n7343), .ZN(n7345) );
  AND2_X1 U8981 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7345), .ZN(n7346) );
  XNOR2_X1 U8982 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7345), .ZN(n10070) );
  INV_X1 U8983 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10069) );
  NOR2_X1 U8984 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  NOR2_X1 U8985 ( .A1(n7346), .A2(n10068), .ZN(n10067) );
  NAND2_X1 U8986 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7347) );
  OAI21_X1 U8987 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7347), .ZN(n10066) );
  NOR2_X1 U8988 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  AOI21_X1 U8989 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10065), .ZN(n10064) );
  NAND2_X1 U8990 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7348) );
  OAI21_X1 U8991 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7348), .ZN(n10063) );
  NOR2_X1 U8992 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  AOI21_X1 U8993 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10062), .ZN(n10061) );
  NOR2_X1 U8994 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7349) );
  AOI21_X1 U8995 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7349), .ZN(n10060) );
  NAND2_X1 U8996 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  OAI21_X1 U8997 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10059), .ZN(n10057) );
  NAND2_X1 U8998 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  OAI21_X1 U8999 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10056), .ZN(n10054) );
  NAND2_X1 U9000 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  OAI21_X1 U9001 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10053), .ZN(n10051) );
  NAND2_X1 U9002 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  OAI21_X1 U9003 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10050), .ZN(n10048) );
  NAND2_X1 U9004 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  OAI21_X1 U9005 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10047), .ZN(n10045) );
  NAND2_X1 U9006 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  OAI21_X1 U9007 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10044), .ZN(n10075) );
  NOR2_X1 U9008 ( .A1(n10076), .A2(n10075), .ZN(n7350) );
  NAND2_X1 U9009 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  OAI21_X1 U9010 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7350), .A(n10074), .ZN(
        n7533) );
  AOI22_X1 U9011 ( .A1(n7713), .A2(keyinput_g50), .B1(n7498), .B2(keyinput_g45), .ZN(n7351) );
  OAI221_X1 U9012 ( .B1(n7713), .B2(keyinput_g50), .C1(n7498), .C2(
        keyinput_g45), .A(n7351), .ZN(n7360) );
  INV_X1 U9013 ( .A(SI_30_), .ZN(n7848) );
  AOI22_X1 U9014 ( .A1(n7848), .A2(keyinput_g2), .B1(n7353), .B2(keyinput_g6), 
        .ZN(n7352) );
  OAI221_X1 U9015 ( .B1(n7848), .B2(keyinput_g2), .C1(n7353), .C2(keyinput_g6), 
        .A(n7352), .ZN(n7359) );
  INV_X1 U9016 ( .A(SI_12_), .ZN(n7471) );
  INV_X1 U9017 ( .A(SI_17_), .ZN(n7462) );
  AOI22_X1 U9018 ( .A1(n7471), .A2(keyinput_g20), .B1(n7462), .B2(keyinput_g15), .ZN(n7354) );
  OAI221_X1 U9019 ( .B1(n7471), .B2(keyinput_g20), .C1(n7462), .C2(
        keyinput_g15), .A(n7354), .ZN(n7358) );
  AOI22_X1 U9020 ( .A1(n7356), .A2(keyinput_g7), .B1(keyinput_g49), .B2(n5506), 
        .ZN(n7355) );
  OAI221_X1 U9021 ( .B1(n7356), .B2(keyinput_g7), .C1(n5506), .C2(keyinput_g49), .A(n7355), .ZN(n7357) );
  NOR4_X1 U9022 ( .A1(n7360), .A2(n7359), .A3(n7358), .A4(n7357), .ZN(n7396)
         );
  AOI22_X1 U9023 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n7361) );
  OAI221_X1 U9024 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_15_), .C2(
        keyinput_g17), .A(n7361), .ZN(n7369) );
  INV_X1 U9025 ( .A(SI_14_), .ZN(n7472) );
  AOI22_X1 U9026 ( .A1(n8427), .A2(keyinput_g38), .B1(n7472), .B2(keyinput_g18), .ZN(n7362) );
  OAI221_X1 U9027 ( .B1(n8427), .B2(keyinput_g38), .C1(n7472), .C2(
        keyinput_g18), .A(n7362), .ZN(n7368) );
  XNOR2_X1 U9028 ( .A(SI_2_), .B(keyinput_g30), .ZN(n7366) );
  XNOR2_X1 U9029 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n7365)
         );
  XNOR2_X1 U9030 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n7364) );
  XNOR2_X1 U9031 ( .A(SI_24_), .B(keyinput_g8), .ZN(n7363) );
  NAND4_X1 U9032 ( .A1(n7366), .A2(n7365), .A3(n7364), .A4(n7363), .ZN(n7367)
         );
  NOR3_X1 U9033 ( .A1(n7369), .A2(n7368), .A3(n7367), .ZN(n7395) );
  AOI22_X1 U9034 ( .A1(n7371), .A2(keyinput_g36), .B1(keyinput_g3), .B2(n7836), 
        .ZN(n7370) );
  OAI221_X1 U9035 ( .B1(n7371), .B2(keyinput_g36), .C1(n7836), .C2(keyinput_g3), .A(n7370), .ZN(n7382) );
  AOI22_X1 U9036 ( .A1(n7373), .A2(keyinput_g12), .B1(keyinput_g34), .B2(
        P2_U3152), .ZN(n7372) );
  OAI221_X1 U9037 ( .B1(n7373), .B2(keyinput_g12), .C1(P2_U3152), .C2(
        keyinput_g34), .A(n7372), .ZN(n7381) );
  AOI22_X1 U9038 ( .A1(n7376), .A2(keyinput_g52), .B1(n7375), .B2(keyinput_g21), .ZN(n7374) );
  OAI221_X1 U9039 ( .B1(n7376), .B2(keyinput_g52), .C1(n7375), .C2(
        keyinput_g21), .A(n7374), .ZN(n7380) );
  AOI22_X1 U9040 ( .A1(n5665), .A2(keyinput_g58), .B1(keyinput_g40), .B2(n7378), .ZN(n7377) );
  OAI221_X1 U9041 ( .B1(n5665), .B2(keyinput_g58), .C1(n7378), .C2(
        keyinput_g40), .A(n7377), .ZN(n7379) );
  NOR4_X1 U9042 ( .A1(n7382), .A2(n7381), .A3(n7380), .A4(n7379), .ZN(n7394)
         );
  AOI22_X1 U9043 ( .A1(n8522), .A2(keyinput_g62), .B1(keyinput_g35), .B2(n5452), .ZN(n7383) );
  OAI221_X1 U9044 ( .B1(n8522), .B2(keyinput_g62), .C1(n5452), .C2(
        keyinput_g35), .A(n7383), .ZN(n7392) );
  INV_X1 U9045 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9729) );
  AOI22_X1 U9046 ( .A1(n9729), .A2(keyinput_g0), .B1(n7385), .B2(keyinput_g28), 
        .ZN(n7384) );
  OAI221_X1 U9047 ( .B1(n9729), .B2(keyinput_g0), .C1(n7385), .C2(keyinput_g28), .A(n7384), .ZN(n7391) );
  INV_X1 U9048 ( .A(SI_6_), .ZN(n7433) );
  AOI22_X1 U9049 ( .A1(n7433), .A2(keyinput_g26), .B1(keyinput_g43), .B2(n7434), .ZN(n7386) );
  OAI221_X1 U9050 ( .B1(n7433), .B2(keyinput_g26), .C1(n7434), .C2(
        keyinput_g43), .A(n7386), .ZN(n7390) );
  XOR2_X1 U9051 ( .A(n5627), .B(keyinput_g53), .Z(n7388) );
  XNOR2_X1 U9052 ( .A(SI_1_), .B(keyinput_g31), .ZN(n7387) );
  NAND2_X1 U9053 ( .A1(n7388), .A2(n7387), .ZN(n7389) );
  NOR4_X1 U9054 ( .A1(n7392), .A2(n7391), .A3(n7390), .A4(n7389), .ZN(n7393)
         );
  NAND4_X1 U9055 ( .A1(n7396), .A2(n7395), .A3(n7394), .A4(n7393), .ZN(n7531)
         );
  AOI22_X1 U9056 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(SI_27_), .B2(keyinput_g5), .ZN(n7397) );
  OAI221_X1 U9057 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        SI_27_), .C2(keyinput_g5), .A(n7397), .ZN(n7404) );
  AOI22_X1 U9058 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(SI_22_), .B2(keyinput_g10), .ZN(n7398) );
  OAI221_X1 U9059 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_22_), .C2(keyinput_g10), .A(n7398), .ZN(n7403) );
  AOI22_X1 U9060 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_5_), 
        .B2(keyinput_g27), .ZN(n7399) );
  OAI221_X1 U9061 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(SI_5_), 
        .C2(keyinput_g27), .A(n7399), .ZN(n7402) );
  AOI22_X1 U9062 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_21_), 
        .B2(keyinput_g11), .ZN(n7400) );
  OAI221_X1 U9063 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_21_), .C2(keyinput_g11), .A(n7400), .ZN(n7401) );
  NOR4_X1 U9064 ( .A1(n7404), .A2(n7403), .A3(n7402), .A4(n7401), .ZN(n7431)
         );
  XOR2_X1 U9065 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_g42), .Z(n7411) );
  AOI22_X1 U9066 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(SI_3_), 
        .B2(keyinput_g29), .ZN(n7405) );
  OAI221_X1 U9067 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(SI_3_), .C2(keyinput_g29), .A(n7405), .ZN(n7410) );
  AOI22_X1 U9068 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_23_), .B2(keyinput_g9), .ZN(n7406) );
  OAI221_X1 U9069 ( .B1(SI_28_), .B2(keyinput_g4), .C1(SI_23_), .C2(
        keyinput_g9), .A(n7406), .ZN(n7409) );
  AOI22_X1 U9070 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n7407) );
  OAI221_X1 U9071 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n7407), .ZN(n7408) );
  NOR4_X1 U9072 ( .A1(n7411), .A2(n7410), .A3(n7409), .A4(n7408), .ZN(n7430)
         );
  AOI22_X1 U9073 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_19_), .B2(
        keyinput_g13), .ZN(n7412) );
  OAI221_X1 U9074 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_19_), .C2(
        keyinput_g13), .A(n7412), .ZN(n7419) );
  AOI22_X1 U9075 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n7413) );
  OAI221_X1 U9076 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n7413), .ZN(n7418) );
  AOI22_X1 U9077 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n7414) );
  OAI221_X1 U9078 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(SI_9_), .C2(keyinput_g23), .A(n7414), .ZN(n7417) );
  AOI22_X1 U9079 ( .A1(SI_31_), .A2(keyinput_g1), .B1(SI_16_), .B2(
        keyinput_g16), .ZN(n7415) );
  OAI221_X1 U9080 ( .B1(SI_31_), .B2(keyinput_g1), .C1(SI_16_), .C2(
        keyinput_g16), .A(n7415), .ZN(n7416) );
  NOR4_X1 U9081 ( .A1(n7419), .A2(n7418), .A3(n7417), .A4(n7416), .ZN(n7429)
         );
  AOI22_X1 U9082 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(SI_7_), 
        .B2(keyinput_g25), .ZN(n7420) );
  OAI221_X1 U9083 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(SI_7_), .C2(keyinput_g25), .A(n7420), .ZN(n7427) );
  AOI22_X1 U9084 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n7421) );
  OAI221_X1 U9085 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n7421), .ZN(n7426) );
  AOI22_X1 U9086 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n7422) );
  OAI221_X1 U9087 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n7422), .ZN(n7425) );
  AOI22_X1 U9088 ( .A1(SI_13_), .A2(keyinput_g19), .B1(SI_18_), .B2(
        keyinput_g14), .ZN(n7423) );
  OAI221_X1 U9089 ( .B1(SI_13_), .B2(keyinput_g19), .C1(SI_18_), .C2(
        keyinput_g14), .A(n7423), .ZN(n7424) );
  NOR4_X1 U9090 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n7428)
         );
  NAND4_X1 U9091 ( .A1(n7431), .A2(n7430), .A3(n7429), .A4(n7428), .ZN(n7530)
         );
  XNOR2_X1 U9092 ( .A(SI_8_), .B(keyinput_g24), .ZN(n7529) );
  AOI22_X1 U9093 ( .A1(n7434), .A2(keyinput_f43), .B1(n7433), .B2(keyinput_f26), .ZN(n7432) );
  OAI221_X1 U9094 ( .B1(n7434), .B2(keyinput_f43), .C1(n7433), .C2(
        keyinput_f26), .A(n7432), .ZN(n7444) );
  AOI22_X1 U9095 ( .A1(n8461), .A2(keyinput_f47), .B1(n7436), .B2(keyinput_f22), .ZN(n7435) );
  OAI221_X1 U9096 ( .B1(n8461), .B2(keyinput_f47), .C1(n7436), .C2(
        keyinput_f22), .A(n7435), .ZN(n7443) );
  INV_X1 U9097 ( .A(SI_31_), .ZN(n7853) );
  AOI22_X1 U9098 ( .A1(n7853), .A2(keyinput_f1), .B1(n7438), .B2(keyinput_f16), 
        .ZN(n7437) );
  OAI221_X1 U9099 ( .B1(n7853), .B2(keyinput_f1), .C1(n7438), .C2(keyinput_f16), .A(n7437), .ZN(n7442) );
  AOI22_X1 U9100 ( .A1(n7440), .A2(keyinput_f48), .B1(keyinput_f63), .B2(n5741), .ZN(n7439) );
  OAI221_X1 U9101 ( .B1(n7440), .B2(keyinput_f48), .C1(n5741), .C2(
        keyinput_f63), .A(n7439), .ZN(n7441) );
  NOR4_X1 U9102 ( .A1(n7444), .A2(n7443), .A3(n7442), .A4(n7441), .ZN(n7488)
         );
  AOI22_X1 U9103 ( .A1(n7836), .A2(keyinput_f3), .B1(n5452), .B2(keyinput_f35), 
        .ZN(n7445) );
  OAI221_X1 U9104 ( .B1(n7836), .B2(keyinput_f3), .C1(n5452), .C2(keyinput_f35), .A(n7445), .ZN(n7456) );
  INV_X1 U9105 ( .A(SI_18_), .ZN(n7447) );
  AOI22_X1 U9106 ( .A1(n6743), .A2(keyinput_f56), .B1(n7447), .B2(keyinput_f14), .ZN(n7446) );
  OAI221_X1 U9107 ( .B1(n6743), .B2(keyinput_f56), .C1(n7447), .C2(
        keyinput_f14), .A(n7446), .ZN(n7455) );
  AOI22_X1 U9108 ( .A1(n7450), .A2(keyinput_f59), .B1(n7449), .B2(keyinput_f23), .ZN(n7448) );
  OAI221_X1 U9109 ( .B1(n7450), .B2(keyinput_f59), .C1(n7449), .C2(
        keyinput_f23), .A(n7448), .ZN(n7454) );
  XOR2_X1 U9110 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_f52), .Z(n7452) );
  XNOR2_X1 U9111 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7451) );
  NAND2_X1 U9112 ( .A1(n7452), .A2(n7451), .ZN(n7453) );
  NOR4_X1 U9113 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n7487)
         );
  INV_X1 U9114 ( .A(SI_15_), .ZN(n7458) );
  AOI22_X1 U9115 ( .A1(n5506), .A2(keyinput_f49), .B1(n7458), .B2(keyinput_f17), .ZN(n7457) );
  OAI221_X1 U9116 ( .B1(n5506), .B2(keyinput_f49), .C1(n7458), .C2(
        keyinput_f17), .A(n7457), .ZN(n7469) );
  AOI22_X1 U9117 ( .A1(n5322), .A2(keyinput_f4), .B1(n7460), .B2(keyinput_f25), 
        .ZN(n7459) );
  OAI221_X1 U9118 ( .B1(n5322), .B2(keyinput_f4), .C1(n7460), .C2(keyinput_f25), .A(n7459), .ZN(n7468) );
  AOI22_X1 U9119 ( .A1(n7463), .A2(keyinput_f39), .B1(n7462), .B2(keyinput_f15), .ZN(n7461) );
  OAI221_X1 U9120 ( .B1(n7463), .B2(keyinput_f39), .C1(n7462), .C2(
        keyinput_f15), .A(n7461), .ZN(n7467) );
  XNOR2_X1 U9121 ( .A(SI_0_), .B(keyinput_f32), .ZN(n7465) );
  XNOR2_X1 U9122 ( .A(SI_30_), .B(keyinput_f2), .ZN(n7464) );
  NAND2_X1 U9123 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NOR4_X1 U9124 ( .A1(n7469), .A2(n7468), .A3(n7467), .A4(n7466), .ZN(n7486)
         );
  AOI22_X1 U9125 ( .A1(n7472), .A2(keyinput_f18), .B1(keyinput_f20), .B2(n7471), .ZN(n7470) );
  OAI221_X1 U9126 ( .B1(n7472), .B2(keyinput_f18), .C1(n7471), .C2(
        keyinput_f20), .A(n7470), .ZN(n7484) );
  AOI22_X1 U9127 ( .A1(n7475), .A2(keyinput_f19), .B1(keyinput_f37), .B2(n7474), .ZN(n7473) );
  OAI221_X1 U9128 ( .B1(n7475), .B2(keyinput_f19), .C1(n7474), .C2(
        keyinput_f37), .A(n7473), .ZN(n7483) );
  AOI22_X1 U9129 ( .A1(n7478), .A2(keyinput_f55), .B1(n7477), .B2(keyinput_f5), 
        .ZN(n7476) );
  OAI221_X1 U9130 ( .B1(n7478), .B2(keyinput_f55), .C1(n7477), .C2(keyinput_f5), .A(n7476), .ZN(n7482) );
  XNOR2_X1 U9131 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n7480) );
  XNOR2_X1 U9132 ( .A(SI_21_), .B(keyinput_f11), .ZN(n7479) );
  NAND2_X1 U9133 ( .A1(n7480), .A2(n7479), .ZN(n7481) );
  NOR4_X1 U9134 ( .A1(n7484), .A2(n7483), .A3(n7482), .A4(n7481), .ZN(n7485)
         );
  NAND4_X1 U9135 ( .A1(n7488), .A2(n7487), .A3(n7486), .A4(n7485), .ZN(n7527)
         );
  AOI22_X1 U9136 ( .A1(SI_3_), .A2(keyinput_f29), .B1(SI_5_), .B2(keyinput_f27), .ZN(n7489) );
  OAI221_X1 U9137 ( .B1(SI_3_), .B2(keyinput_f29), .C1(SI_5_), .C2(
        keyinput_f27), .A(n7489), .ZN(n7496) );
  AOI22_X1 U9138 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n7490) );
  OAI221_X1 U9139 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n7490), .ZN(n7495) );
  AOI22_X1 U9140 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n7491) );
  OAI221_X1 U9141 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n7491), .ZN(n7494) );
  AOI22_X1 U9142 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n7492) );
  OAI221_X1 U9143 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n7492), .ZN(n7493) );
  NOR4_X1 U9144 ( .A1(n7496), .A2(n7495), .A3(n7494), .A4(n7493), .ZN(n7524)
         );
  XOR2_X1 U9145 ( .A(P2_U3152), .B(keyinput_f34), .Z(n7504) );
  AOI22_X1 U9146 ( .A1(SI_25_), .A2(keyinput_f7), .B1(n7498), .B2(keyinput_f45), .ZN(n7497) );
  OAI221_X1 U9147 ( .B1(SI_25_), .B2(keyinput_f7), .C1(n7498), .C2(
        keyinput_f45), .A(n7497), .ZN(n7503) );
  AOI22_X1 U9148 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n7499) );
  OAI221_X1 U9149 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n7499), .ZN(n7502) );
  AOI22_X1 U9150 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n7500) );
  OAI221_X1 U9151 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_26_), .C2(
        keyinput_f6), .A(n7500), .ZN(n7501) );
  NOR4_X1 U9152 ( .A1(n7504), .A2(n7503), .A3(n7502), .A4(n7501), .ZN(n7523)
         );
  AOI22_X1 U9153 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(SI_23_), 
        .B2(keyinput_f9), .ZN(n7505) );
  OAI221_X1 U9154 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(SI_23_), .C2(keyinput_f9), .A(n7505), .ZN(n7512) );
  AOI22_X1 U9155 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(SI_20_), 
        .B2(keyinput_f12), .ZN(n7506) );
  OAI221_X1 U9156 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(SI_20_), .C2(keyinput_f12), .A(n7506), .ZN(n7511) );
  AOI22_X1 U9157 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n7507) );
  OAI221_X1 U9158 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n7507), .ZN(n7510) );
  AOI22_X1 U9159 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n7508) );
  OAI221_X1 U9160 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n7508), .ZN(n7509) );
  NOR4_X1 U9161 ( .A1(n7512), .A2(n7511), .A3(n7510), .A4(n7509), .ZN(n7522)
         );
  AOI22_X1 U9162 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(SI_19_), .B2(keyinput_f13), .ZN(n7513) );
  OAI221_X1 U9163 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        SI_19_), .C2(keyinput_f13), .A(n7513), .ZN(n7520) );
  AOI22_X1 U9164 ( .A1(SI_4_), .A2(keyinput_f28), .B1(SI_24_), .B2(keyinput_f8), .ZN(n7514) );
  OAI221_X1 U9165 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_24_), .C2(
        keyinput_f8), .A(n7514), .ZN(n7519) );
  AOI22_X1 U9166 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(SI_2_), 
        .B2(keyinput_f30), .ZN(n7515) );
  OAI221_X1 U9167 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(SI_2_), 
        .C2(keyinput_f30), .A(n7515), .ZN(n7518) );
  AOI22_X1 U9168 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(SI_22_), .B2(keyinput_f10), .ZN(n7516) );
  OAI221_X1 U9169 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        SI_22_), .C2(keyinput_f10), .A(n7516), .ZN(n7517) );
  NOR4_X1 U9170 ( .A1(n7520), .A2(n7519), .A3(n7518), .A4(n7517), .ZN(n7521)
         );
  NAND4_X1 U9171 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n7526)
         );
  NAND2_X1 U9172 ( .A1(SI_8_), .A2(keyinput_f24), .ZN(n7525) );
  OAI221_X1 U9173 ( .B1(n7527), .B2(n7526), .C1(SI_8_), .C2(keyinput_f24), .A(
        n7525), .ZN(n7528) );
  OAI211_X1 U9174 ( .C1(n7531), .C2(n7530), .A(n7529), .B(n7528), .ZN(n7532)
         );
  XNOR2_X1 U9175 ( .A(n7533), .B(n7532), .ZN(n7537) );
  NOR2_X1 U9176 ( .A1(n7534), .A2(n7535), .ZN(n7536) );
  XNOR2_X1 U9177 ( .A(n7537), .B(n7536), .ZN(ADD_1071_U4) );
  INV_X1 U9178 ( .A(n7538), .ZN(n7578) );
  OAI222_X1 U9179 ( .A1(n7540), .A2(P1_U3084), .B1(n9671), .B2(n7578), .C1(
        n7539), .C2(n9667), .ZN(P1_U3329) );
  AND2_X1 U9180 ( .A1(n7542), .A2(n7541), .ZN(n7544) );
  OR2_X1 U9181 ( .A1(n7542), .A2(n7541), .ZN(n7543) );
  NAND2_X1 U9182 ( .A1(n9556), .A2(n8406), .ZN(n7547) );
  NAND2_X1 U9183 ( .A1(n9283), .A2(n8412), .ZN(n7546) );
  NAND2_X1 U9184 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  XNOR2_X1 U9185 ( .A(n7548), .B(n4311), .ZN(n7659) );
  AND2_X1 U9186 ( .A1(n9283), .A2(n8411), .ZN(n7549) );
  AOI21_X1 U9187 ( .B1(n9556), .B2(n8412), .A(n7549), .ZN(n7660) );
  XNOR2_X1 U9188 ( .A(n7659), .B(n7660), .ZN(n7550) );
  XNOR2_X1 U9189 ( .A(n7658), .B(n7550), .ZN(n7551) );
  NAND2_X1 U9190 ( .A1(n7551), .A2(n9694), .ZN(n7556) );
  INV_X1 U9191 ( .A(n9554), .ZN(n7552) );
  OAI22_X1 U9192 ( .A1(n9699), .A2(n7552), .B1(n9682), .B2(n9517), .ZN(n7553)
         );
  AOI211_X1 U9193 ( .C1(n9685), .C2(n9549), .A(n7554), .B(n7553), .ZN(n7555)
         );
  OAI211_X1 U9194 ( .C1(n9714), .C2(n9224), .A(n7556), .B(n7555), .ZN(P1_U3213) );
  NAND2_X1 U9195 ( .A1(n10011), .A2(n7557), .ZN(n8659) );
  NAND2_X1 U9196 ( .A1(n7558), .A2(n8659), .ZN(n7559) );
  NAND2_X1 U9197 ( .A1(n9127), .A2(n7600), .ZN(n8266) );
  OR2_X1 U9198 ( .A1(n7559), .A2(n8658), .ZN(n8998) );
  NAND2_X1 U9199 ( .A1(n7559), .A2(n8658), .ZN(n7560) );
  NAND2_X1 U9200 ( .A1(n8998), .A2(n7560), .ZN(n9130) );
  OR2_X1 U9201 ( .A1(n9130), .A2(n8982), .ZN(n7567) );
  INV_X1 U9202 ( .A(n8265), .ZN(n7561) );
  AOI21_X1 U9203 ( .B1(n7562), .B2(n8268), .A(n7561), .ZN(n7563) );
  NAND2_X1 U9204 ( .A1(n7563), .A2(n8658), .ZN(n7598) );
  OAI211_X1 U9205 ( .C1(n7563), .C2(n8658), .A(n7598), .B(n8986), .ZN(n7565)
         );
  AOI22_X1 U9206 ( .A1(n8651), .A2(n8968), .B1(n8965), .B2(n8548), .ZN(n7564)
         );
  AND2_X1 U9207 ( .A1(n7565), .A2(n7564), .ZN(n7566) );
  NAND2_X1 U9208 ( .A1(n7567), .A2(n7566), .ZN(n9132) );
  INV_X1 U9209 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7569) );
  OAI22_X1 U9210 ( .A1(n8946), .A2(n7569), .B1(n7568), .B2(n8943), .ZN(n7570)
         );
  AOI21_X1 U9211 ( .B1(n8892), .B2(n9127), .A(n7570), .ZN(n7575) );
  INV_X1 U9212 ( .A(n9127), .ZN(n7571) );
  OR2_X1 U9213 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  AND2_X1 U9214 ( .A1(n7601), .A2(n7573), .ZN(n9128) );
  NAND2_X1 U9215 ( .A1(n9128), .A2(n9022), .ZN(n7574) );
  OAI211_X1 U9216 ( .C1(n9130), .C2(n8992), .A(n7575), .B(n7574), .ZN(n7576)
         );
  AOI21_X1 U9217 ( .B1(n8946), .B2(n9132), .A(n7576), .ZN(n7577) );
  INV_X1 U9218 ( .A(n7577), .ZN(P2_U3286) );
  INV_X1 U9219 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7579) );
  OAI222_X1 U9220 ( .A1(P2_U3152), .A2(n7580), .B1(n8405), .B2(n7579), .C1(
        n9165), .C2(n7578), .ZN(P2_U3334) );
  XNOR2_X1 U9221 ( .A(n7581), .B(n7878), .ZN(n9719) );
  INV_X1 U9222 ( .A(n4756), .ZN(n7582) );
  AOI211_X1 U9223 ( .C1(n7187), .C2(n7583), .A(n9946), .B(n7582), .ZN(n9721)
         );
  INV_X1 U9224 ( .A(n7187), .ZN(n9692) );
  NOR2_X1 U9225 ( .A1(n9692), .A2(n9539), .ZN(n7585) );
  OAI22_X1 U9226 ( .A1(n9884), .A2(n6337), .B1(n9698), .B2(n9880), .ZN(n7584)
         );
  AOI211_X1 U9227 ( .C1(n9721), .C2(n9513), .A(n7585), .B(n7584), .ZN(n7596)
         );
  INV_X1 U9228 ( .A(n7586), .ZN(n7588) );
  OAI21_X1 U9229 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7591) );
  INV_X1 U9230 ( .A(n7878), .ZN(n7590) );
  XNOR2_X1 U9231 ( .A(n7591), .B(n7590), .ZN(n7592) );
  NAND2_X1 U9232 ( .A1(n7592), .A2(n9871), .ZN(n7594) );
  AOI22_X1 U9233 ( .A1(n9875), .A2(n9684), .B1(n9549), .B2(n9873), .ZN(n7593)
         );
  NAND2_X1 U9234 ( .A1(n7594), .A2(n7593), .ZN(n9720) );
  NAND2_X1 U9235 ( .A1(n9720), .A2(n9884), .ZN(n7595) );
  OAI211_X1 U9236 ( .C1(n9719), .C2(n9855), .A(n7596), .B(n7595), .ZN(P1_U3279) );
  OR2_X1 U9237 ( .A1(n8652), .A2(n9013), .ZN(n8276) );
  NAND2_X1 U9238 ( .A1(n8652), .A2(n9013), .ZN(n8274) );
  NAND2_X1 U9239 ( .A1(n8276), .A2(n8274), .ZN(n8664) );
  INV_X1 U9240 ( .A(n7600), .ZN(n8547) );
  NAND2_X1 U9241 ( .A1(n9127), .A2(n8547), .ZN(n8653) );
  NAND2_X1 U9242 ( .A1(n8998), .A2(n8653), .ZN(n7597) );
  XOR2_X1 U9243 ( .A(n8664), .B(n7597), .Z(n10025) );
  INV_X1 U9244 ( .A(n10025), .ZN(n7609) );
  XOR2_X1 U9245 ( .A(n8173), .B(n8664), .Z(n7599) );
  OAI222_X1 U9246 ( .A1(n9014), .A2(n8978), .B1(n9012), .B2(n7600), .C1(n9010), 
        .C2(n7599), .ZN(n10022) );
  INV_X1 U9247 ( .A(n7601), .ZN(n7602) );
  INV_X1 U9248 ( .A(n8652), .ZN(n10019) );
  OAI21_X1 U9249 ( .B1(n7602), .B2(n10019), .A(n9003), .ZN(n10021) );
  OAI22_X1 U9250 ( .A1(n8946), .A2(n7604), .B1(n7603), .B2(n8943), .ZN(n7605)
         );
  AOI21_X1 U9251 ( .B1(n8892), .B2(n8652), .A(n7605), .ZN(n7606) );
  OAI21_X1 U9252 ( .B1(n10021), .B2(n8638), .A(n7606), .ZN(n7607) );
  AOI21_X1 U9253 ( .B1(n10022), .B2(n8946), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9254 ( .B1(n7609), .B2(n9024), .A(n7608), .ZN(P2_U3285) );
  INV_X1 U9255 ( .A(n7177), .ZN(n7612) );
  NOR3_X1 U9256 ( .A1(n7610), .A2(n9015), .A3(n8516), .ZN(n7611) );
  AOI21_X1 U9257 ( .B1(n7612), .B2(n8532), .A(n7611), .ZN(n7621) );
  NOR2_X1 U9258 ( .A1(n7613), .A2(n8518), .ZN(n7618) );
  AND2_X1 U9259 ( .A1(n8508), .A2(n9111), .ZN(n7617) );
  OAI21_X1 U9260 ( .B1(n8539), .B2(n8908), .A(n7614), .ZN(n7616) );
  OAI22_X1 U9261 ( .A1(n8536), .A2(n9015), .B1(n8537), .B2(n8956), .ZN(n7615)
         );
  NOR4_X1 U9262 ( .A1(n7618), .A2(n7617), .A3(n7616), .A4(n7615), .ZN(n7619)
         );
  OAI21_X1 U9263 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(P2_U3217) );
  NAND2_X1 U9264 ( .A1(n7623), .A2(n7622), .ZN(n7625) );
  NAND2_X1 U9265 ( .A1(n7625), .A2(n7624), .ZN(n7627) );
  XNOR2_X1 U9266 ( .A(n7715), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7626) );
  NOR2_X1 U9267 ( .A1(n7626), .A2(n7627), .ZN(n7716) );
  AOI21_X1 U9268 ( .B1(n7627), .B2(n7626), .A(n7716), .ZN(n7640) );
  NAND2_X1 U9269 ( .A1(n7629), .A2(n7628), .ZN(n7631) );
  NAND2_X1 U9270 ( .A1(n7631), .A2(n7630), .ZN(n7634) );
  NAND2_X1 U9271 ( .A1(n7715), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7632) );
  OAI21_X1 U9272 ( .B1(n7715), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7632), .ZN(
        n7633) );
  NOR2_X1 U9273 ( .A1(n7633), .A2(n7634), .ZN(n7708) );
  AOI211_X1 U9274 ( .C1(n7634), .C2(n7633), .A(n7708), .B(n7710), .ZN(n7635)
         );
  INV_X1 U9275 ( .A(n7635), .ZN(n7639) );
  INV_X1 U9276 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9277 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8468) );
  OAI21_X1 U9278 ( .B1(n8629), .B2(n7636), .A(n8468), .ZN(n7637) );
  AOI21_X1 U9279 ( .B1(n8562), .B2(n7715), .A(n7637), .ZN(n7638) );
  OAI211_X1 U9280 ( .C1(n7640), .C2(n8620), .A(n7639), .B(n7638), .ZN(P2_U3261) );
  INV_X1 U9281 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7647) );
  AOI22_X1 U9282 ( .A1(n7642), .A2(n9914), .B1(n9913), .B2(n7641), .ZN(n7643)
         );
  OAI211_X1 U9283 ( .C1(n7645), .C2(n9922), .A(n7644), .B(n7643), .ZN(n7648)
         );
  NAND2_X1 U9284 ( .A1(n7648), .A2(n9952), .ZN(n7646) );
  OAI21_X1 U9285 ( .B1(n9952), .B2(n7647), .A(n7646), .ZN(P1_U3487) );
  NAND2_X1 U9286 ( .A1(n7648), .A2(n9968), .ZN(n7649) );
  OAI21_X1 U9287 ( .B1(n9968), .B2(n7650), .A(n7649), .ZN(P1_U3534) );
  INV_X1 U9288 ( .A(n7651), .ZN(n7655) );
  OAI222_X1 U9289 ( .A1(P1_U3084), .A2(n7653), .B1(n9671), .B2(n7655), .C1(
        n7652), .C2(n7753), .ZN(P1_U3328) );
  OAI222_X1 U9290 ( .A1(n7656), .A2(P2_U3152), .B1(n9165), .B2(n7655), .C1(
        n7654), .C2(n8405), .ZN(P2_U3333) );
  NAND2_X1 U9291 ( .A1(n7659), .A2(n7660), .ZN(n7657) );
  NAND2_X1 U9292 ( .A1(n7658), .A2(n7657), .ZN(n7664) );
  INV_X1 U9293 ( .A(n7659), .ZN(n7662) );
  INV_X1 U9294 ( .A(n7660), .ZN(n7661) );
  NAND2_X1 U9295 ( .A1(n7662), .A2(n7661), .ZN(n7663) );
  NAND2_X1 U9296 ( .A1(n9635), .A2(n8406), .ZN(n7666) );
  NAND2_X1 U9297 ( .A1(n9548), .A2(n8412), .ZN(n7665) );
  NAND2_X1 U9298 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  XNOR2_X1 U9299 ( .A(n7667), .B(n6381), .ZN(n7728) );
  NAND2_X1 U9300 ( .A1(n9635), .A2(n8412), .ZN(n7669) );
  NAND2_X1 U9301 ( .A1(n9548), .A2(n8411), .ZN(n7668) );
  NAND2_X1 U9302 ( .A1(n7669), .A2(n7668), .ZN(n7729) );
  XNOR2_X1 U9303 ( .A(n7728), .B(n7729), .ZN(n7670) );
  XNOR2_X1 U9304 ( .A(n7730), .B(n7670), .ZN(n7671) );
  NAND2_X1 U9305 ( .A1(n7671), .A2(n9694), .ZN(n7675) );
  AND2_X1 U9306 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9787) );
  INV_X1 U9307 ( .A(n9536), .ZN(n7672) );
  OAI22_X1 U9308 ( .A1(n9699), .A2(n7672), .B1(n9682), .B2(n9530), .ZN(n7673)
         );
  AOI211_X1 U9309 ( .C1(n9685), .C2(n9283), .A(n9787), .B(n7673), .ZN(n7674)
         );
  OAI211_X1 U9310 ( .C1(n9540), .C2(n9224), .A(n7675), .B(n7674), .ZN(P1_U3239) );
  INV_X1 U9311 ( .A(n7676), .ZN(n7685) );
  OAI222_X1 U9312 ( .A1(n7678), .A2(P1_U3084), .B1(n9671), .B2(n7685), .C1(
        n7677), .C2(n7753), .ZN(P1_U3327) );
  INV_X1 U9313 ( .A(n7679), .ZN(n7684) );
  AOI21_X1 U9314 ( .B1(n7681), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7680), .ZN(
        n7682) );
  OAI21_X1 U9315 ( .B1(n7684), .B2(n9665), .A(n7682), .ZN(P1_U3326) );
  AOI22_X1 U9316 ( .A1(n8632), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9162), .ZN(n7683) );
  OAI21_X1 U9317 ( .B1(n7684), .B2(n9165), .A(n7683), .ZN(P2_U3331) );
  OAI222_X1 U9318 ( .A1(P2_U3152), .A2(n7687), .B1(n8405), .B2(n7686), .C1(
        n9165), .C2(n7685), .ZN(P2_U3332) );
  XNOR2_X1 U9319 ( .A(n7689), .B(n7880), .ZN(n9641) );
  NAND2_X1 U9320 ( .A1(n7690), .A2(n7943), .ZN(n7692) );
  INV_X1 U9321 ( .A(n7880), .ZN(n7691) );
  NAND2_X1 U9322 ( .A1(n7692), .A2(n7691), .ZN(n7694) );
  NAND2_X1 U9323 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9324 ( .A1(n7695), .A2(n9871), .ZN(n7697) );
  AOI22_X1 U9325 ( .A1(n9875), .A2(n9284), .B1(n9283), .B2(n9873), .ZN(n7696)
         );
  NAND2_X1 U9326 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  AOI21_X1 U9327 ( .B1(n9641), .B2(n7699), .A(n7698), .ZN(n9643) );
  AND2_X1 U9328 ( .A1(n4756), .A2(n7702), .ZN(n7700) );
  OR2_X1 U9329 ( .A1(n7700), .A2(n9553), .ZN(n9639) );
  AOI22_X1 U9330 ( .A1(n9856), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7701), .B2(
        n9826), .ZN(n7704) );
  NAND2_X1 U9331 ( .A1(n7702), .A2(n9555), .ZN(n7703) );
  OAI211_X1 U9332 ( .C1(n9639), .C2(n9440), .A(n7704), .B(n7703), .ZN(n7705)
         );
  AOI21_X1 U9333 ( .B1(n9641), .B2(n7706), .A(n7705), .ZN(n7707) );
  OAI21_X1 U9334 ( .B1(n9643), .B2(n9856), .A(n7707), .ZN(P1_U3278) );
  NAND2_X1 U9335 ( .A1(n8593), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7709) );
  OAI21_X1 U9336 ( .B1(n8593), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7709), .ZN(
        n7711) );
  AOI211_X1 U9337 ( .C1(n7712), .C2(n7711), .A(n8592), .B(n7710), .ZN(n7724)
         );
  NOR2_X1 U9338 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7713), .ZN(n7714) );
  AOI21_X1 U9339 ( .B1(n8599), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7714), .ZN(
        n7722) );
  XNOR2_X1 U9340 ( .A(n8588), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7720) );
  OR2_X1 U9341 ( .A1(n7715), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7718) );
  INV_X1 U9342 ( .A(n7716), .ZN(n7717) );
  AND2_X1 U9343 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  NAND2_X1 U9344 ( .A1(n7720), .A2(n7719), .ZN(n8587) );
  OAI211_X1 U9345 ( .C1(n7720), .C2(n7719), .A(n8612), .B(n8587), .ZN(n7721)
         );
  OAI211_X1 U9346 ( .C1(n8619), .C2(n8588), .A(n7722), .B(n7721), .ZN(n7723)
         );
  OR2_X1 U9347 ( .A1(n7724), .A2(n7723), .ZN(P2_U3262) );
  INV_X1 U9348 ( .A(n7768), .ZN(n7727) );
  NAND2_X1 U9349 ( .A1(n9162), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7725) );
  OAI211_X1 U9350 ( .C1(n7727), .C2(n9165), .A(n7726), .B(n7725), .ZN(P2_U3330) );
  NAND2_X1 U9351 ( .A1(n9630), .A2(n8406), .ZN(n7732) );
  NAND2_X1 U9352 ( .A1(n9499), .A2(n8412), .ZN(n7731) );
  NAND2_X1 U9353 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  XNOR2_X1 U9354 ( .A(n7733), .B(n4311), .ZN(n7735) );
  AND2_X1 U9355 ( .A1(n9499), .A2(n8411), .ZN(n7734) );
  AOI21_X1 U9356 ( .B1(n9630), .B2(n8412), .A(n7734), .ZN(n7736) );
  NAND2_X1 U9357 ( .A1(n7735), .A2(n7736), .ZN(n8089) );
  INV_X1 U9358 ( .A(n7735), .ZN(n7738) );
  INV_X1 U9359 ( .A(n7736), .ZN(n7737) );
  NAND2_X1 U9360 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U9361 ( .A1(n8089), .A2(n7739), .ZN(n7742) );
  INV_X1 U9362 ( .A(n8090), .ZN(n7741) );
  AOI21_X1 U9363 ( .B1(n7740), .B2(n7742), .A(n7741), .ZN(n7747) );
  INV_X1 U9364 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9365 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7743), .ZN(n9797) );
  OAI22_X1 U9366 ( .A1(n9682), .A2(n9518), .B1(n9699), .B2(n9510), .ZN(n7744)
         );
  AOI211_X1 U9367 ( .C1(n9685), .C2(n9548), .A(n9797), .B(n7744), .ZN(n7746)
         );
  NAND2_X1 U9368 ( .A1(n9630), .A2(n9276), .ZN(n7745) );
  OAI211_X1 U9369 ( .C1(n7747), .C2(n9278), .A(n7746), .B(n7745), .ZN(P1_U3224) );
  NAND2_X1 U9370 ( .A1(n7768), .A2(n7748), .ZN(n7749) );
  OAI211_X1 U9371 ( .C1(n7753), .C2(n7750), .A(n7749), .B(n9730), .ZN(P1_U3325) );
  INV_X1 U9372 ( .A(n8189), .ZN(n8172) );
  AOI22_X1 U9373 ( .A1(n7751), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9162), .ZN(n7752) );
  OAI21_X1 U9374 ( .B1(n8172), .B2(n9165), .A(n7752), .ZN(P2_U3329) );
  OAI222_X1 U9375 ( .A1(n5343), .A2(P1_U3084), .B1(n9671), .B2(n7755), .C1(
        n7754), .C2(n7753), .ZN(P1_U3332) );
  XOR2_X1 U9376 ( .A(n7756), .B(n7887), .Z(n9585) );
  AOI21_X1 U9377 ( .B1(n5293), .B2(n9382), .A(n9356), .ZN(n9582) );
  AOI22_X1 U9378 ( .A1(n9856), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9197), .B2(
        n9826), .ZN(n7757) );
  OAI21_X1 U9379 ( .B1(n4614), .B2(n9539), .A(n7757), .ZN(n7764) );
  NAND2_X1 U9380 ( .A1(n9376), .A2(n7993), .ZN(n7758) );
  XOR2_X1 U9381 ( .A(n7887), .B(n7758), .Z(n7762) );
  NAND2_X1 U9382 ( .A1(n9282), .A2(n9873), .ZN(n7760) );
  NAND2_X1 U9383 ( .A1(n9403), .A2(n9875), .ZN(n7759) );
  AOI211_X1 U9384 ( .C1(n9504), .C2(n9582), .A(n7764), .B(n7763), .ZN(n7765)
         );
  OAI21_X1 U9385 ( .B1(n9585), .B2(n9855), .A(n7765), .ZN(P1_U3266) );
  NAND2_X1 U9386 ( .A1(n7767), .A2(n7766), .ZN(n7774) );
  NAND2_X1 U9387 ( .A1(n7768), .A2(n8204), .ZN(n7770) );
  NAND2_X1 U9388 ( .A1(n8194), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U9389 ( .A1(n8725), .A2(n8213), .ZN(n7771) );
  XNOR2_X1 U9390 ( .A(n7771), .B(n5644), .ZN(n7772) );
  XNOR2_X1 U9391 ( .A(n9036), .B(n7772), .ZN(n7773) );
  XNOR2_X1 U9392 ( .A(n7774), .B(n7773), .ZN(n7779) );
  OAI22_X1 U9393 ( .A1(n8539), .A2(n8192), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7775), .ZN(n7777) );
  OAI22_X1 U9394 ( .A1(n8536), .A2(n8545), .B1(n8537), .B2(n8718), .ZN(n7776)
         );
  AOI211_X1 U9395 ( .C1(n9036), .C2(n8508), .A(n7777), .B(n7776), .ZN(n7778)
         );
  OAI21_X1 U9396 ( .B1(n7779), .B2(n8518), .A(n7778), .ZN(P2_U3222) );
  INV_X1 U9397 ( .A(n8023), .ZN(n7780) );
  AOI21_X1 U9398 ( .B1(n8034), .B2(n9325), .A(n7780), .ZN(n8068) );
  INV_X1 U9399 ( .A(n8068), .ZN(n7844) );
  AND2_X1 U9400 ( .A1(n7917), .A2(n7781), .ZN(n7914) );
  NAND2_X1 U9401 ( .A1(n7914), .A2(n7782), .ZN(n8056) );
  NAND2_X1 U9402 ( .A1(n9840), .A2(n7783), .ZN(n7784) );
  NOR2_X1 U9403 ( .A1(n8056), .A2(n7784), .ZN(n8062) );
  INV_X1 U9404 ( .A(n8054), .ZN(n7786) );
  OAI21_X1 U9405 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n7789) );
  INV_X1 U9406 ( .A(n7914), .ZN(n7788) );
  AOI21_X1 U9407 ( .B1(n7789), .B2(n8058), .A(n7788), .ZN(n7802) );
  INV_X1 U9408 ( .A(n9431), .ZN(n7790) );
  NAND2_X1 U9409 ( .A1(n7819), .A2(n7790), .ZN(n7791) );
  AND2_X1 U9410 ( .A1(n7791), .A2(n7979), .ZN(n7792) );
  NAND2_X1 U9411 ( .A1(n7792), .A2(n9400), .ZN(n7823) );
  INV_X1 U9412 ( .A(n7823), .ZN(n7793) );
  NAND3_X1 U9413 ( .A1(n7793), .A2(n7995), .A3(n7970), .ZN(n7817) );
  AND2_X1 U9414 ( .A1(n7818), .A2(n7863), .ZN(n7900) );
  INV_X1 U9415 ( .A(n7900), .ZN(n7815) );
  NAND2_X1 U9416 ( .A1(n9556), .A2(n9528), .ZN(n7809) );
  NAND2_X1 U9417 ( .A1(n7809), .A2(n7794), .ZN(n7940) );
  INV_X1 U9418 ( .A(n7940), .ZN(n7798) );
  INV_X1 U9419 ( .A(n7952), .ZN(n7795) );
  NOR2_X1 U9420 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  AND3_X1 U9421 ( .A1(n7942), .A2(n7798), .A3(n7797), .ZN(n7804) );
  NAND2_X1 U9422 ( .A1(n7924), .A2(n7916), .ZN(n7913) );
  INV_X1 U9423 ( .A(n7913), .ZN(n7799) );
  NAND3_X1 U9424 ( .A1(n7804), .A2(n7964), .A3(n7799), .ZN(n7800) );
  OR2_X1 U9425 ( .A1(n7815), .A2(n7800), .ZN(n7801) );
  OR2_X1 U9426 ( .A1(n7817), .A2(n7801), .ZN(n8059) );
  AOI211_X1 U9427 ( .C1(n8062), .C2(n7803), .A(n7802), .B(n8059), .ZN(n7828)
         );
  INV_X1 U9428 ( .A(n7804), .ZN(n7807) );
  AND2_X1 U9429 ( .A1(n7927), .A2(n7923), .ZN(n7805) );
  NAND2_X1 U9430 ( .A1(n7928), .A2(n7805), .ZN(n7953) );
  INV_X1 U9431 ( .A(n7953), .ZN(n7806) );
  OR2_X1 U9432 ( .A1(n7807), .A2(n7806), .ZN(n7812) );
  NAND2_X1 U9433 ( .A1(n7930), .A2(n7808), .ZN(n7945) );
  NAND2_X1 U9434 ( .A1(n7945), .A2(n7809), .ZN(n7937) );
  OAI21_X1 U9435 ( .B1(n7940), .B2(n7943), .A(n7937), .ZN(n7810) );
  NAND2_X1 U9436 ( .A1(n7810), .A2(n7942), .ZN(n7811) );
  NAND4_X1 U9437 ( .A1(n7812), .A2(n7941), .A3(n7965), .A4(n7811), .ZN(n7813)
         );
  NAND2_X1 U9438 ( .A1(n7813), .A2(n7964), .ZN(n7814) );
  OR2_X1 U9439 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  OR2_X1 U9440 ( .A1(n7817), .A2(n7816), .ZN(n7827) );
  NOR2_X1 U9441 ( .A1(n9588), .A2(n9198), .ZN(n7996) );
  INV_X1 U9442 ( .A(n7996), .ZN(n7826) );
  AND2_X1 U9443 ( .A1(n7970), .A2(n7818), .ZN(n7975) );
  INV_X1 U9444 ( .A(n7975), .ZN(n7821) );
  AND2_X1 U9445 ( .A1(n7822), .A2(n7819), .ZN(n7984) );
  NAND2_X1 U9446 ( .A1(n7978), .A2(n7898), .ZN(n7973) );
  INV_X1 U9447 ( .A(n7973), .ZN(n7820) );
  OAI211_X1 U9448 ( .C1(n7899), .C2(n7821), .A(n7984), .B(n7820), .ZN(n7824)
         );
  NAND2_X1 U9449 ( .A1(n7823), .A2(n7822), .ZN(n7985) );
  NAND3_X1 U9450 ( .A1(n7824), .A2(n7995), .A3(n7985), .ZN(n7825) );
  NAND4_X1 U9451 ( .A1(n7827), .A2(n7826), .A3(n7825), .A4(n7991), .ZN(n8063)
         );
  OAI21_X1 U9452 ( .B1(n7828), .B2(n8063), .A(n9361), .ZN(n7829) );
  NAND3_X1 U9453 ( .A1(n7829), .A2(n8066), .A3(n8020), .ZN(n7843) );
  NAND2_X1 U9454 ( .A1(n8020), .A2(n7830), .ZN(n7831) );
  NAND3_X1 U9455 ( .A1(n8024), .A2(n8019), .A3(n7831), .ZN(n7832) );
  INV_X1 U9456 ( .A(n9325), .ZN(n8033) );
  AOI22_X1 U9457 ( .A1(n8068), .A2(n7832), .B1(n8033), .B2(n8029), .ZN(n8070)
         );
  INV_X1 U9458 ( .A(n7835), .ZN(n7837) );
  NAND2_X1 U9459 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  MUX2_X1 U9460 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7852), .Z(n7847) );
  XNOR2_X1 U9461 ( .A(n7847), .B(n7848), .ZN(n7845) );
  NAND2_X1 U9462 ( .A1(n9161), .A2(n7859), .ZN(n7841) );
  INV_X1 U9463 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9668) );
  OR2_X1 U9464 ( .A1(n7857), .A2(n9668), .ZN(n7840) );
  AOI21_X1 U9465 ( .B1(n9309), .B2(n9280), .A(n9566), .ZN(n8030) );
  INV_X1 U9466 ( .A(n8030), .ZN(n7842) );
  OAI211_X1 U9467 ( .C1(n7844), .C2(n7843), .A(n8070), .B(n7842), .ZN(n7860)
         );
  NAND2_X1 U9468 ( .A1(n9566), .A2(n9280), .ZN(n8072) );
  INV_X1 U9469 ( .A(n7847), .ZN(n7849) );
  NAND2_X1 U9470 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  MUX2_X1 U9471 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7852), .Z(n7854) );
  XNOR2_X1 U9472 ( .A(n7854), .B(n7853), .ZN(n7855) );
  NOR2_X1 U9473 ( .A1(n7857), .A2(n6145), .ZN(n7858) );
  AOI21_X1 U9474 ( .B1(n9309), .B2(n8072), .A(n9701), .ZN(n8028) );
  INV_X1 U9475 ( .A(n8028), .ZN(n8037) );
  INV_X1 U9476 ( .A(n9701), .ZN(n7862) );
  INV_X1 U9477 ( .A(n9309), .ZN(n7861) );
  AOI211_X1 U9478 ( .C1(n7860), .C2(n8037), .A(n5343), .B(n8071), .ZN(n7896)
         );
  NAND2_X1 U9479 ( .A1(n7862), .A2(n7861), .ZN(n8074) );
  INV_X1 U9480 ( .A(n7990), .ZN(n9401) );
  NAND2_X1 U9481 ( .A1(n7978), .A2(n9431), .ZN(n9454) );
  AND2_X1 U9482 ( .A1(n9475), .A2(n7863), .ZN(n9498) );
  NOR2_X1 U9483 ( .A1(n7865), .A2(n7864), .ZN(n7867) );
  NAND4_X1 U9484 ( .A1(n7868), .A2(n7867), .A3(n9842), .A4(n7866), .ZN(n7871)
         );
  NAND2_X1 U9485 ( .A1(n9870), .A2(n7911), .ZN(n7870) );
  NOR3_X1 U9486 ( .A1(n7871), .A2(n7870), .A3(n7869), .ZN(n7875) );
  NAND4_X1 U9487 ( .A1(n7875), .A2(n7874), .A3(n7873), .A4(n7872), .ZN(n7877)
         );
  INV_X1 U9488 ( .A(n7955), .ZN(n7876) );
  NOR2_X1 U9489 ( .A1(n7877), .A2(n7876), .ZN(n7879) );
  NAND3_X1 U9490 ( .A1(n7880), .A2(n7879), .A3(n7878), .ZN(n7881) );
  OR3_X1 U9491 ( .A1(n9525), .A2(n9544), .A3(n7881), .ZN(n7882) );
  NOR2_X1 U9492 ( .A1(n9514), .A2(n7882), .ZN(n7883) );
  NAND4_X1 U9493 ( .A1(n9469), .A2(n9498), .A3(n9486), .A4(n7883), .ZN(n7884)
         );
  NOR2_X1 U9494 ( .A1(n9454), .A2(n7884), .ZN(n7885) );
  NAND4_X1 U9495 ( .A1(n9401), .A2(n9420), .A3(n5264), .A4(n7885), .ZN(n7886)
         );
  NOR3_X1 U9496 ( .A1(n7887), .A2(n9378), .A3(n7886), .ZN(n7889) );
  NAND2_X1 U9497 ( .A1(n8015), .A2(n7888), .ZN(n9365) );
  AND2_X1 U9498 ( .A1(n7889), .A2(n9365), .ZN(n7890) );
  AND4_X1 U9499 ( .A1(n7891), .A2(n9323), .A3(n8067), .A4(n7890), .ZN(n7893)
         );
  INV_X1 U9500 ( .A(n9566), .ZN(n9314) );
  XNOR2_X1 U9501 ( .A(n9314), .B(n9280), .ZN(n7892) );
  NAND4_X1 U9502 ( .A1(n8040), .A2(n8074), .A3(n7893), .A4(n7892), .ZN(n7894)
         );
  NAND2_X1 U9503 ( .A1(n7894), .A2(n5343), .ZN(n8041) );
  INV_X1 U9504 ( .A(n8041), .ZN(n7895) );
  NOR2_X1 U9505 ( .A1(n7896), .A2(n7895), .ZN(n8044) );
  AND2_X1 U9506 ( .A1(n7898), .A2(n7897), .ZN(n7972) );
  MUX2_X1 U9507 ( .A(n7900), .B(n7899), .S(n8032), .Z(n7969) );
  NAND3_X1 U9508 ( .A1(n6556), .A2(n9840), .A3(n8032), .ZN(n7901) );
  OAI21_X1 U9509 ( .B1(n9841), .B2(n8032), .A(n7901), .ZN(n7902) );
  NAND2_X1 U9510 ( .A1(n7902), .A2(n9842), .ZN(n7910) );
  NAND2_X1 U9511 ( .A1(n7903), .A2(n7904), .ZN(n7908) );
  NAND2_X1 U9512 ( .A1(n7904), .A2(n8057), .ZN(n7906) );
  NAND2_X1 U9513 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  MUX2_X1 U9514 ( .A(n7908), .B(n7907), .S(n8032), .Z(n7909) );
  NAND2_X1 U9515 ( .A1(n7910), .A2(n7909), .ZN(n7912) );
  NAND2_X1 U9516 ( .A1(n7912), .A2(n7911), .ZN(n7920) );
  AOI21_X1 U9517 ( .B1(n7920), .B2(n7914), .A(n7913), .ZN(n7922) );
  AND2_X1 U9518 ( .A1(n7916), .A2(n7915), .ZN(n7919) );
  INV_X1 U9519 ( .A(n7917), .ZN(n7918) );
  AOI21_X1 U9520 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7921) );
  MUX2_X1 U9521 ( .A(n7922), .B(n7921), .S(n8032), .Z(n7954) );
  NAND2_X1 U9522 ( .A1(n7954), .A2(n7923), .ZN(n7926) );
  NAND3_X1 U9523 ( .A1(n7926), .A2(n7925), .A3(n7924), .ZN(n7929) );
  NAND3_X1 U9524 ( .A1(n7929), .A2(n7928), .A3(n7927), .ZN(n7936) );
  NAND2_X1 U9525 ( .A1(n7940), .A2(n7930), .ZN(n7931) );
  NAND2_X1 U9526 ( .A1(n7942), .A2(n7931), .ZN(n7947) );
  NAND4_X1 U9527 ( .A1(n7933), .A2(n7955), .A3(n7932), .A4(n8032), .ZN(n7934)
         );
  NOR2_X1 U9528 ( .A1(n7947), .A2(n7934), .ZN(n7935) );
  NAND2_X1 U9529 ( .A1(n7936), .A2(n7935), .ZN(n7963) );
  NAND2_X1 U9530 ( .A1(n7937), .A2(n7941), .ZN(n7958) );
  INV_X1 U9531 ( .A(n7938), .ZN(n7939) );
  INV_X1 U9532 ( .A(n8032), .ZN(n7997) );
  OAI21_X1 U9533 ( .B1(n7940), .B2(n7939), .A(n7997), .ZN(n7950) );
  MUX2_X1 U9534 ( .A(n7942), .B(n7941), .S(n8032), .Z(n7949) );
  INV_X1 U9535 ( .A(n7943), .ZN(n7944) );
  NOR2_X1 U9536 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  OR3_X1 U9537 ( .A1(n7947), .A2(n7997), .A3(n7946), .ZN(n7948) );
  OAI211_X1 U9538 ( .C1(n7958), .C2(n7950), .A(n7949), .B(n7948), .ZN(n7951)
         );
  NOR2_X1 U9539 ( .A1(n7951), .A2(n9514), .ZN(n7962) );
  OAI21_X1 U9540 ( .B1(n7954), .B2(n7953), .A(n7952), .ZN(n7960) );
  NAND3_X1 U9541 ( .A1(n7956), .A2(n7955), .A3(n7997), .ZN(n7957) );
  NOR2_X1 U9542 ( .A1(n7958), .A2(n7957), .ZN(n7959) );
  NAND2_X1 U9543 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  NAND3_X1 U9544 ( .A1(n7963), .A2(n7962), .A3(n7961), .ZN(n7967) );
  MUX2_X1 U9545 ( .A(n7965), .B(n7964), .S(n8032), .Z(n7966) );
  NAND3_X1 U9546 ( .A1(n7967), .A2(n9498), .A3(n7966), .ZN(n7968) );
  NAND2_X1 U9547 ( .A1(n7969), .A2(n7968), .ZN(n7974) );
  NAND2_X1 U9548 ( .A1(n9431), .A2(n7970), .ZN(n7971) );
  AOI21_X1 U9549 ( .B1(n7972), .B2(n7974), .A(n7971), .ZN(n7977) );
  AOI21_X1 U9550 ( .B1(n7975), .B2(n7974), .A(n7973), .ZN(n7976) );
  MUX2_X1 U9551 ( .A(n7977), .B(n7976), .S(n8032), .Z(n7983) );
  INV_X1 U9552 ( .A(n7978), .ZN(n7980) );
  OAI21_X1 U9553 ( .B1(n7983), .B2(n7980), .A(n7979), .ZN(n7982) );
  AOI21_X1 U9554 ( .B1(n7982), .B2(n7984), .A(n7981), .ZN(n7989) );
  INV_X1 U9555 ( .A(n7983), .ZN(n7987) );
  INV_X1 U9556 ( .A(n7984), .ZN(n7986) );
  OAI21_X1 U9557 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n7988) );
  MUX2_X1 U9558 ( .A(n7989), .B(n7988), .S(n8032), .Z(n8002) );
  OR2_X1 U9559 ( .A1(n9378), .A2(n7990), .ZN(n8001) );
  INV_X1 U9560 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U9561 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  NAND2_X1 U9562 ( .A1(n9403), .A2(n8032), .ZN(n7998) );
  OR2_X1 U9563 ( .A1(n9588), .A2(n7998), .ZN(n7999) );
  OAI211_X1 U9564 ( .C1(n8002), .C2(n8001), .A(n8000), .B(n7999), .ZN(n8016)
         );
  NAND2_X1 U9565 ( .A1(n9577), .A2(n9362), .ZN(n8003) );
  NAND2_X1 U9566 ( .A1(n8019), .A2(n8003), .ZN(n8006) );
  NAND2_X1 U9567 ( .A1(n8010), .A2(n9282), .ZN(n8004) );
  NAND2_X1 U9568 ( .A1(n8020), .A2(n8004), .ZN(n8005) );
  MUX2_X1 U9569 ( .A(n8006), .B(n8005), .S(n8032), .Z(n8007) );
  OAI21_X1 U9570 ( .B1(n9345), .B2(n8016), .A(n8007), .ZN(n8018) );
  NAND2_X1 U9571 ( .A1(n9362), .A2(n9348), .ZN(n8008) );
  NAND2_X1 U9572 ( .A1(n8009), .A2(n8008), .ZN(n8013) );
  NOR2_X1 U9573 ( .A1(n8010), .A2(n9282), .ZN(n8011) );
  NOR2_X1 U9574 ( .A1(n8011), .A2(n9577), .ZN(n8012) );
  MUX2_X1 U9575 ( .A(n8013), .B(n8012), .S(n8032), .Z(n8014) );
  OAI21_X1 U9576 ( .B1(n8016), .B2(n8015), .A(n8014), .ZN(n8017) );
  NAND2_X1 U9577 ( .A1(n8018), .A2(n8017), .ZN(n8022) );
  MUX2_X1 U9578 ( .A(n8020), .B(n8019), .S(n8032), .Z(n8021) );
  NAND2_X1 U9579 ( .A1(n8022), .A2(n4752), .ZN(n8026) );
  MUX2_X1 U9580 ( .A(n8024), .B(n8023), .S(n8032), .Z(n8025) );
  NAND2_X1 U9581 ( .A1(n8026), .A2(n8025), .ZN(n8035) );
  INV_X1 U9582 ( .A(n8035), .ZN(n8027) );
  NOR2_X1 U9583 ( .A1(n8034), .A2(n8032), .ZN(n8031) );
  AOI211_X1 U9584 ( .C1(n9325), .C2(n8032), .A(n8031), .B(n8030), .ZN(n8038)
         );
  NAND3_X1 U9585 ( .A1(n8035), .A2(n8034), .A3(n8033), .ZN(n8036) );
  NAND3_X1 U9586 ( .A1(n8038), .A2(n8037), .A3(n8036), .ZN(n8039) );
  OAI21_X1 U9587 ( .B1(n8046), .B2(n8042), .A(n8041), .ZN(n8043) );
  NOR3_X1 U9588 ( .A1(n8071), .A2(n5377), .A3(n5343), .ZN(n8045) );
  NAND2_X1 U9589 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  AOI21_X1 U9590 ( .B1(n9893), .B2(n9291), .A(n5343), .ZN(n8053) );
  INV_X1 U9591 ( .A(n8049), .ZN(n8052) );
  AOI211_X1 U9592 ( .C1(n8053), .C2(n8052), .A(n4965), .B(n8051), .ZN(n8055)
         );
  OAI21_X1 U9593 ( .B1(n8055), .B2(n4753), .A(n8054), .ZN(n8061) );
  AOI21_X1 U9594 ( .B1(n8058), .B2(n8057), .A(n8056), .ZN(n8060) );
  AOI211_X1 U9595 ( .C1(n8062), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8064)
         );
  OAI21_X1 U9596 ( .B1(n8064), .B2(n8063), .A(n9361), .ZN(n8065) );
  NAND4_X1 U9597 ( .A1(n8068), .A2(n8067), .A3(n8066), .A4(n8065), .ZN(n8069)
         );
  OAI211_X1 U9598 ( .C1(n9566), .C2(n9280), .A(n8070), .B(n8069), .ZN(n8073)
         );
  AOI21_X1 U9599 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8076) );
  INV_X1 U9600 ( .A(n8074), .ZN(n8075) );
  NOR2_X1 U9601 ( .A1(n8076), .A2(n8075), .ZN(n8077) );
  XNOR2_X1 U9602 ( .A(n8077), .B(n9867), .ZN(n8078) );
  NAND2_X1 U9603 ( .A1(n8078), .A2(n6029), .ZN(n8079) );
  NOR4_X1 U9604 ( .A1(n8083), .A2(n4312), .A3(n8082), .A4(n9755), .ZN(n8085)
         );
  OAI21_X1 U9605 ( .B1(n5377), .B2(n8086), .A(P1_B_REG_SCAN_IN), .ZN(n8084) );
  OAI22_X1 U9606 ( .A1(n8087), .A2(n8086), .B1(n8085), .B2(n8084), .ZN(
        P1_U3240) );
  AOI22_X1 U9607 ( .A1(n9588), .A2(n6395), .B1(n8411), .B2(n9403), .ZN(n8141)
         );
  AOI22_X1 U9608 ( .A1(n9588), .A2(n8406), .B1(n8412), .B2(n9403), .ZN(n8088)
         );
  XNOR2_X1 U9609 ( .A(n8088), .B(n6381), .ZN(n8140) );
  NAND2_X1 U9610 ( .A1(n9623), .A2(n8406), .ZN(n8092) );
  NAND2_X1 U9611 ( .A1(n9478), .A2(n8412), .ZN(n8091) );
  NAND2_X1 U9612 ( .A1(n8092), .A2(n8091), .ZN(n8093) );
  XNOR2_X1 U9613 ( .A(n8093), .B(n6381), .ZN(n8095) );
  AND2_X1 U9614 ( .A1(n9478), .A2(n8411), .ZN(n8094) );
  AOI21_X1 U9615 ( .B1(n9623), .B2(n8412), .A(n8094), .ZN(n8096) );
  XNOR2_X1 U9616 ( .A(n8095), .B(n8096), .ZN(n9206) );
  INV_X1 U9617 ( .A(n8095), .ZN(n8097) );
  NAND2_X1 U9618 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U9619 ( .A1(n9618), .A2(n8155), .ZN(n8100) );
  NAND2_X1 U9620 ( .A1(n9500), .A2(n8412), .ZN(n8099) );
  NAND2_X1 U9621 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  XNOR2_X1 U9622 ( .A(n8101), .B(n4311), .ZN(n8104) );
  INV_X1 U9623 ( .A(n8104), .ZN(n8102) );
  AND2_X1 U9624 ( .A1(n9500), .A2(n8411), .ZN(n8103) );
  NAND2_X1 U9625 ( .A1(n9254), .A2(n9255), .ZN(n9253) );
  NAND2_X1 U9626 ( .A1(n9611), .A2(n8155), .ZN(n8107) );
  NAND2_X1 U9627 ( .A1(n9479), .A2(n8412), .ZN(n8106) );
  NAND2_X1 U9628 ( .A1(n8107), .A2(n8106), .ZN(n8108) );
  XNOR2_X1 U9629 ( .A(n8108), .B(n6381), .ZN(n8110) );
  AND2_X1 U9630 ( .A1(n9479), .A2(n8411), .ZN(n8109) );
  AOI21_X1 U9631 ( .B1(n9611), .B2(n8412), .A(n8109), .ZN(n8111) );
  XNOR2_X1 U9632 ( .A(n8110), .B(n8111), .ZN(n9177) );
  INV_X1 U9633 ( .A(n8110), .ZN(n8112) );
  NAND2_X1 U9634 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  NAND2_X1 U9635 ( .A1(n9606), .A2(n8155), .ZN(n8115) );
  NAND2_X1 U9636 ( .A1(n9470), .A2(n8412), .ZN(n8114) );
  NAND2_X1 U9637 ( .A1(n8115), .A2(n8114), .ZN(n8116) );
  XNOR2_X1 U9638 ( .A(n8116), .B(n6381), .ZN(n8119) );
  NAND2_X1 U9639 ( .A1(n9606), .A2(n8412), .ZN(n8118) );
  NAND2_X1 U9640 ( .A1(n9470), .A2(n8411), .ZN(n8117) );
  NAND2_X1 U9641 ( .A1(n8118), .A2(n8117), .ZN(n8120) );
  NAND2_X1 U9642 ( .A1(n8119), .A2(n8120), .ZN(n9231) );
  INV_X1 U9643 ( .A(n8119), .ZN(n8122) );
  INV_X1 U9644 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U9645 ( .A1(n8122), .A2(n8121), .ZN(n9233) );
  NAND2_X1 U9646 ( .A1(n9601), .A2(n8155), .ZN(n8124) );
  NAND2_X1 U9647 ( .A1(n9455), .A2(n8412), .ZN(n8123) );
  NAND2_X1 U9648 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  XNOR2_X1 U9649 ( .A(n8125), .B(n6381), .ZN(n8127) );
  AND2_X1 U9650 ( .A1(n9455), .A2(n8411), .ZN(n8126) );
  AOI21_X1 U9651 ( .B1(n9601), .B2(n8412), .A(n8126), .ZN(n8128) );
  XNOR2_X1 U9652 ( .A(n8127), .B(n8128), .ZN(n9185) );
  INV_X1 U9653 ( .A(n8127), .ZN(n8129) );
  NAND2_X1 U9654 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  AND2_X1 U9655 ( .A1(n9435), .A2(n8411), .ZN(n8132) );
  AOI21_X1 U9656 ( .B1(n9597), .B2(n8412), .A(n8132), .ZN(n8136) );
  NAND2_X1 U9657 ( .A1(n9597), .A2(n8155), .ZN(n8134) );
  NAND2_X1 U9658 ( .A1(n9435), .A2(n8412), .ZN(n8133) );
  NAND2_X1 U9659 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  XNOR2_X1 U9660 ( .A(n8135), .B(n6381), .ZN(n9244) );
  AOI22_X1 U9661 ( .A1(n9591), .A2(n8406), .B1(n8412), .B2(n9421), .ZN(n8137)
         );
  XOR2_X1 U9662 ( .A(n6381), .B(n8137), .Z(n8138) );
  AOI22_X1 U9663 ( .A1(n9591), .A2(n6395), .B1(n8411), .B2(n9421), .ZN(n9168)
         );
  XNOR2_X1 U9664 ( .A(n8140), .B(n8141), .ZN(n9213) );
  AOI22_X1 U9665 ( .A1(n5293), .A2(n6395), .B1(n8411), .B2(n9367), .ZN(n8145)
         );
  NAND2_X1 U9666 ( .A1(n5293), .A2(n8155), .ZN(n8143) );
  NAND2_X1 U9667 ( .A1(n9367), .A2(n8412), .ZN(n8142) );
  NAND2_X1 U9668 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  XNOR2_X1 U9669 ( .A(n8144), .B(n6381), .ZN(n8147) );
  XOR2_X1 U9670 ( .A(n8145), .B(n8147), .Z(n9195) );
  INV_X1 U9671 ( .A(n8145), .ZN(n8146) );
  NAND2_X1 U9672 ( .A1(n9577), .A2(n8155), .ZN(n8149) );
  NAND2_X1 U9673 ( .A1(n9282), .A2(n8412), .ZN(n8148) );
  NAND2_X1 U9674 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  XNOR2_X1 U9675 ( .A(n8150), .B(n6381), .ZN(n8154) );
  NAND2_X1 U9676 ( .A1(n9577), .A2(n8412), .ZN(n8152) );
  NAND2_X1 U9677 ( .A1(n9282), .A2(n8411), .ZN(n8151) );
  NAND2_X1 U9678 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  NAND2_X1 U9679 ( .A1(n8154), .A2(n8153), .ZN(n9268) );
  NOR2_X1 U9680 ( .A1(n8154), .A2(n8153), .ZN(n9267) );
  NAND2_X1 U9681 ( .A1(n9572), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U9682 ( .A1(n9366), .A2(n8412), .ZN(n8156) );
  NAND2_X1 U9683 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  XNOR2_X1 U9684 ( .A(n8158), .B(n4311), .ZN(n8161) );
  AND2_X1 U9685 ( .A1(n9366), .A2(n8411), .ZN(n8159) );
  AOI21_X1 U9686 ( .B1(n9572), .B2(n8412), .A(n8159), .ZN(n8160) );
  NAND2_X1 U9687 ( .A1(n8161), .A2(n8160), .ZN(n8420) );
  OAI21_X1 U9688 ( .B1(n8161), .B2(n8160), .A(n8420), .ZN(n8162) );
  OAI21_X1 U9689 ( .B1(n8426), .B2(n8164), .A(n9694), .ZN(n8169) );
  NOR2_X1 U9690 ( .A1(n9682), .A2(n9347), .ZN(n8167) );
  INV_X1 U9691 ( .A(n9342), .ZN(n8165) );
  OAI22_X1 U9692 ( .A1(n9699), .A2(n8165), .B1(n9271), .B2(n9348), .ZN(n8166)
         );
  AOI211_X1 U9693 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3084), .A(n8167), 
        .B(n8166), .ZN(n8168) );
  OAI211_X1 U9694 ( .C1(n9344), .C2(n9224), .A(n8169), .B(n8168), .ZN(P1_U3212) );
  OAI222_X1 U9695 ( .A1(n8172), .A2(n9671), .B1(n9667), .B2(n8171), .C1(
        P1_U3084), .C2(n8170), .ZN(P1_U3324) );
  INV_X1 U9696 ( .A(n9011), .ZN(n8176) );
  NAND2_X1 U9697 ( .A1(n9121), .A2(n8978), .ZN(n8279) );
  INV_X1 U9698 ( .A(n8289), .ZN(n8175) );
  NAND2_X1 U9699 ( .A1(n9106), .A2(n8908), .ZN(n8288) );
  NAND2_X1 U9700 ( .A1(n8289), .A2(n8288), .ZN(n8938) );
  INV_X1 U9701 ( .A(n8938), .ZN(n8927) );
  INV_X1 U9702 ( .A(n8283), .ZN(n8174) );
  NAND2_X1 U9703 ( .A1(n9116), .A2(n9015), .ZN(n8960) );
  OR2_X1 U9704 ( .A1(n8174), .A2(n8961), .ZN(n8923) );
  AND2_X1 U9705 ( .A1(n8927), .A2(n8923), .ZN(n8924) );
  NOR2_X1 U9706 ( .A1(n8175), .A2(n8924), .ZN(n8179) );
  OR2_X1 U9707 ( .A1(n9097), .A2(n8538), .ZN(n8292) );
  XNOR2_X1 U9708 ( .A(n9116), .B(n9015), .ZN(n8980) );
  INV_X1 U9709 ( .A(n8980), .ZN(n8975) );
  AND2_X1 U9710 ( .A1(n8975), .A2(n8283), .ZN(n8922) );
  AND2_X1 U9711 ( .A1(n8922), .A2(n8289), .ZN(n8177) );
  AND2_X1 U9712 ( .A1(n8177), .A2(n8921), .ZN(n8178) );
  NAND2_X1 U9713 ( .A1(n9097), .A2(n8538), .ZN(n8291) );
  XNOR2_X1 U9714 ( .A(n9093), .B(n8906), .ZN(n8873) );
  INV_X1 U9715 ( .A(n8873), .ZN(n8877) );
  INV_X1 U9716 ( .A(n8906), .ZN(n8686) );
  OR2_X1 U9717 ( .A1(n9093), .A2(n8686), .ZN(n8295) );
  OAI21_X1 U9718 ( .B1(n8878), .B2(n8877), .A(n8295), .ZN(n8864) );
  OR2_X1 U9719 ( .A1(n9087), .A2(n8687), .ZN(n8306) );
  NAND2_X1 U9720 ( .A1(n9087), .A2(n8687), .ZN(n8301) );
  NAND2_X1 U9721 ( .A1(n8306), .A2(n8301), .ZN(n8856) );
  NAND2_X1 U9722 ( .A1(n8865), .A2(n8301), .ZN(n8846) );
  INV_X1 U9723 ( .A(n8868), .ZN(n8688) );
  OR2_X1 U9724 ( .A1(n9083), .A2(n8688), .ZN(n8307) );
  NAND2_X1 U9725 ( .A1(n9083), .A2(n8688), .ZN(n8835) );
  NAND2_X1 U9726 ( .A1(n8307), .A2(n8835), .ZN(n8844) );
  INV_X1 U9727 ( .A(n8844), .ZN(n8847) );
  NAND2_X1 U9728 ( .A1(n9077), .A2(n8690), .ZN(n8312) );
  NAND2_X1 U9729 ( .A1(n8310), .A2(n8312), .ZN(n8828) );
  INV_X1 U9730 ( .A(n8835), .ZN(n8180) );
  NOR2_X1 U9731 ( .A1(n8828), .A2(n8180), .ZN(n8181) );
  OR2_X1 U9732 ( .A1(n9072), .A2(n8691), .ZN(n8314) );
  NAND2_X1 U9733 ( .A1(n9072), .A2(n8691), .ZN(n8807) );
  NAND2_X1 U9734 ( .A1(n8314), .A2(n8807), .ZN(n8813) );
  OR2_X1 U9735 ( .A1(n9067), .A2(n8693), .ZN(n8315) );
  NAND2_X1 U9736 ( .A1(n9067), .A2(n8693), .ZN(n8305) );
  NAND2_X1 U9737 ( .A1(n8315), .A2(n8305), .ZN(n8694) );
  INV_X1 U9738 ( .A(n8807), .ZN(n8182) );
  NOR2_X1 U9739 ( .A1(n8694), .A2(n8182), .ZN(n8183) );
  INV_X1 U9740 ( .A(n8315), .ZN(n8304) );
  XNOR2_X1 U9741 ( .A(n9062), .B(n8780), .ZN(n8788) );
  OR2_X1 U9742 ( .A1(n9057), .A2(n8459), .ZN(n8217) );
  NAND2_X1 U9743 ( .A1(n9057), .A2(n8459), .ZN(n8319) );
  AND2_X1 U9744 ( .A1(n9062), .A2(n8780), .ZN(n8322) );
  NOR2_X1 U9745 ( .A1(n8769), .A2(n8322), .ZN(n8184) );
  XNOR2_X1 U9746 ( .A(n9053), .B(n8781), .ZN(n8758) );
  INV_X1 U9747 ( .A(n8758), .ZN(n8381) );
  OR2_X1 U9748 ( .A1(n9053), .A2(n8781), .ZN(n8328) );
  NAND2_X1 U9749 ( .A1(n9048), .A2(n8546), .ZN(n8331) );
  NAND2_X1 U9750 ( .A1(n9036), .A2(n8188), .ZN(n8341) );
  INV_X1 U9751 ( .A(n8714), .ZN(n8383) );
  NAND2_X1 U9752 ( .A1(n8189), .A2(n8204), .ZN(n8191) );
  NAND2_X1 U9753 ( .A1(n8194), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U9754 ( .A1(n9029), .A2(n8192), .ZN(n8348) );
  INV_X1 U9755 ( .A(n8700), .ZN(n8645) );
  NAND2_X1 U9756 ( .A1(n8643), .A2(n8645), .ZN(n8644) );
  NOR2_X1 U9757 ( .A1(n8634), .A2(n8193), .ZN(n8201) );
  NAND2_X1 U9758 ( .A1(n9161), .A2(n8204), .ZN(n8196) );
  NAND2_X1 U9759 ( .A1(n8194), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8195) );
  INV_X1 U9760 ( .A(n8348), .ZN(n8197) );
  AOI21_X1 U9761 ( .B1(n8201), .B2(n8639), .A(n8197), .ZN(n8203) );
  INV_X1 U9762 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U9763 ( .A1(n5544), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U9764 ( .A1(n5562), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8198) );
  OAI211_X1 U9765 ( .C1(n5564), .C2(n8200), .A(n8199), .B(n8198), .ZN(n8646)
         );
  INV_X1 U9766 ( .A(n8646), .ZN(n8208) );
  NOR2_X1 U9767 ( .A1(n8639), .A2(n8208), .ZN(n8214) );
  INV_X1 U9768 ( .A(n8201), .ZN(n8202) );
  AOI22_X1 U9769 ( .A1(n8644), .A2(n8203), .B1(n8214), .B2(n8202), .ZN(n8210)
         );
  NAND2_X1 U9770 ( .A1(n9157), .A2(n8204), .ZN(n8207) );
  NAND2_X1 U9771 ( .A1(n8205), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8206) );
  INV_X1 U9772 ( .A(n8634), .ZN(n8209) );
  NAND2_X1 U9773 ( .A1(n8639), .A2(n8208), .ZN(n8350) );
  NAND2_X1 U9774 ( .A1(n8353), .A2(n8350), .ZN(n8386) );
  NAND2_X1 U9775 ( .A1(n9025), .A2(n8209), .ZN(n8352) );
  OAI21_X1 U9776 ( .B1(n8210), .B2(n8386), .A(n8352), .ZN(n8211) );
  INV_X1 U9777 ( .A(n8386), .ZN(n8216) );
  INV_X1 U9778 ( .A(n8214), .ZN(n8351) );
  NAND2_X1 U9779 ( .A1(n8352), .A2(n8351), .ZN(n8385) );
  INV_X1 U9780 ( .A(n8385), .ZN(n8215) );
  OR2_X1 U9781 ( .A1(n8392), .A2(n8888), .ZN(n8354) );
  MUX2_X1 U9782 ( .A(n8216), .B(n8215), .S(n8354), .Z(n8358) );
  MUX2_X1 U9783 ( .A(n8319), .B(n8217), .S(n8354), .Z(n8327) );
  INV_X1 U9784 ( .A(n8354), .ZN(n8346) );
  MUX2_X1 U9785 ( .A(n4404), .B(n8218), .S(n8346), .Z(n8236) );
  AND2_X1 U9786 ( .A1(n8220), .A2(n8219), .ZN(n8222) );
  OAI211_X1 U9787 ( .C1(n8236), .C2(n8222), .A(n8250), .B(n8221), .ZN(n8223)
         );
  NAND2_X1 U9788 ( .A1(n8223), .A2(n8354), .ZN(n8241) );
  NAND2_X1 U9789 ( .A1(n6478), .A2(n8227), .ZN(n8224) );
  NAND3_X1 U9790 ( .A1(n8232), .A2(n8225), .A3(n8224), .ZN(n8226) );
  NAND2_X1 U9791 ( .A1(n8226), .A2(n8230), .ZN(n8235) );
  NAND3_X1 U9792 ( .A1(n6478), .A2(n8227), .A3(n5482), .ZN(n8228) );
  NAND2_X1 U9793 ( .A1(n8229), .A2(n8228), .ZN(n8231) );
  NAND2_X1 U9794 ( .A1(n8231), .A2(n8230), .ZN(n8233) );
  NAND2_X1 U9795 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  MUX2_X1 U9796 ( .A(n8235), .B(n8234), .S(n8354), .Z(n8238) );
  INV_X1 U9797 ( .A(n8236), .ZN(n8247) );
  NAND3_X1 U9798 ( .A1(n8238), .A2(n8247), .A3(n8237), .ZN(n8240) );
  INV_X1 U9799 ( .A(n8248), .ZN(n8239) );
  AOI21_X1 U9800 ( .B1(n8241), .B2(n8240), .A(n8239), .ZN(n8254) );
  INV_X1 U9801 ( .A(n8242), .ZN(n8246) );
  OAI21_X1 U9802 ( .B1(n8244), .B2(n9991), .A(n8243), .ZN(n8245) );
  OAI21_X1 U9803 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8249) );
  AOI21_X1 U9804 ( .B1(n8249), .B2(n8248), .A(n8354), .ZN(n8253) );
  NOR2_X1 U9805 ( .A1(n8250), .A2(n8354), .ZN(n8251) );
  NOR2_X1 U9806 ( .A1(n8251), .A2(n8369), .ZN(n8252) );
  OAI21_X1 U9807 ( .B1(n8254), .B2(n8253), .A(n8252), .ZN(n8258) );
  MUX2_X1 U9808 ( .A(n8256), .B(n8255), .S(n8354), .Z(n8257) );
  NAND2_X1 U9809 ( .A1(n8259), .A2(n8549), .ZN(n8260) );
  MUX2_X1 U9810 ( .A(n8261), .B(n8260), .S(n8346), .Z(n8262) );
  NAND2_X1 U9811 ( .A1(n8266), .A2(n8265), .ZN(n8263) );
  NAND2_X1 U9812 ( .A1(n8263), .A2(n8354), .ZN(n8264) );
  NAND2_X1 U9813 ( .A1(n8274), .A2(n8266), .ZN(n8271) );
  INV_X1 U9814 ( .A(n8266), .ZN(n8269) );
  OAI211_X1 U9815 ( .C1(n8269), .C2(n8268), .A(n8276), .B(n8267), .ZN(n8270)
         );
  MUX2_X1 U9816 ( .A(n8271), .B(n8270), .S(n8354), .Z(n8272) );
  NAND3_X1 U9817 ( .A1(n8277), .A2(n8279), .A3(n8274), .ZN(n8275) );
  NAND2_X1 U9818 ( .A1(n8277), .A2(n8276), .ZN(n8280) );
  INV_X1 U9819 ( .A(n8921), .ZN(n8278) );
  INV_X1 U9820 ( .A(n9015), .ZN(n8966) );
  MUX2_X1 U9821 ( .A(n8966), .B(n9116), .S(n8354), .Z(n8281) );
  NAND2_X1 U9822 ( .A1(n9116), .A2(n8966), .ZN(n8951) );
  NAND2_X1 U9823 ( .A1(n8281), .A2(n8951), .ZN(n8282) );
  NAND2_X1 U9824 ( .A1(n8963), .A2(n8282), .ZN(n8286) );
  MUX2_X1 U9825 ( .A(n8284), .B(n8283), .S(n8354), .Z(n8285) );
  AOI21_X1 U9826 ( .B1(n8286), .B2(n8285), .A(n8938), .ZN(n8287) );
  NAND2_X1 U9827 ( .A1(n8292), .A2(n8291), .ZN(n8904) );
  INV_X1 U9828 ( .A(n8904), .ZN(n8377) );
  MUX2_X1 U9829 ( .A(n8289), .B(n8288), .S(n8346), .Z(n8290) );
  MUX2_X1 U9830 ( .A(n8292), .B(n8291), .S(n8354), .Z(n8293) );
  NAND3_X1 U9831 ( .A1(n8294), .A2(n8873), .A3(n8293), .ZN(n8300) );
  OAI21_X1 U9832 ( .B1(n8685), .B2(n8906), .A(n8301), .ZN(n8297) );
  INV_X1 U9833 ( .A(n8295), .ZN(n8296) );
  MUX2_X1 U9834 ( .A(n8297), .B(n8296), .S(n8354), .Z(n8298) );
  INV_X1 U9835 ( .A(n8298), .ZN(n8299) );
  NAND3_X1 U9836 ( .A1(n8300), .A2(n8306), .A3(n8299), .ZN(n8308) );
  NAND2_X1 U9837 ( .A1(n8308), .A2(n8301), .ZN(n8302) );
  NAND2_X1 U9838 ( .A1(n8302), .A2(n8307), .ZN(n8303) );
  NAND3_X1 U9839 ( .A1(n8308), .A2(n8307), .A3(n8306), .ZN(n8309) );
  NAND2_X1 U9840 ( .A1(n8309), .A2(n8835), .ZN(n8311) );
  NAND2_X1 U9841 ( .A1(n8311), .A2(n8310), .ZN(n8313) );
  NAND3_X1 U9842 ( .A1(n8313), .A2(n8312), .A3(n8807), .ZN(n8316) );
  NAND4_X1 U9843 ( .A1(n8316), .A2(n8346), .A3(n8315), .A4(n8314), .ZN(n8317)
         );
  NAND3_X1 U9844 ( .A1(n8318), .A2(n8317), .A3(n4541), .ZN(n8325) );
  OAI21_X1 U9845 ( .B1(n8780), .B2(n9062), .A(n8776), .ZN(n8321) );
  NAND2_X1 U9846 ( .A1(n8319), .A2(n8354), .ZN(n8320) );
  NAND2_X1 U9847 ( .A1(n8321), .A2(n8320), .ZN(n8323) );
  INV_X1 U9848 ( .A(n8322), .ZN(n8777) );
  NAND2_X1 U9849 ( .A1(n8334), .A2(n8328), .ZN(n8329) );
  NAND2_X1 U9850 ( .A1(n8329), .A2(n8346), .ZN(n8330) );
  AND2_X1 U9851 ( .A1(n9053), .A2(n8781), .ZN(n8332) );
  OAI21_X1 U9852 ( .B1(n8742), .B2(n8332), .A(n8354), .ZN(n8333) );
  INV_X1 U9853 ( .A(n8728), .ZN(n8724) );
  INV_X1 U9854 ( .A(n8334), .ZN(n8335) );
  OR3_X1 U9855 ( .A1(n9042), .A2(n8545), .A3(n8354), .ZN(n8337) );
  NAND3_X1 U9856 ( .A1(n8338), .A2(n8343), .A3(n8337), .ZN(n8342) );
  NAND2_X1 U9857 ( .A1(n9042), .A2(n8545), .ZN(n8339) );
  AOI21_X1 U9858 ( .B1(n8341), .B2(n8339), .A(n8346), .ZN(n8340) );
  AOI21_X1 U9859 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8345) );
  NOR2_X1 U9860 ( .A1(n8343), .A2(n8346), .ZN(n8344) );
  MUX2_X1 U9861 ( .A(n8348), .B(n8347), .S(n8346), .Z(n8349) );
  INV_X1 U9862 ( .A(n8352), .ZN(n8356) );
  INV_X1 U9863 ( .A(n8353), .ZN(n8355) );
  MUX2_X1 U9864 ( .A(n8356), .B(n8355), .S(n8354), .Z(n8357) );
  INV_X1 U9865 ( .A(n8828), .ZN(n8836) );
  INV_X1 U9866 ( .A(n8856), .ZN(n8866) );
  NOR2_X1 U9867 ( .A1(n8359), .A2(n9980), .ZN(n8368) );
  NOR2_X1 U9868 ( .A1(n8360), .A2(n6983), .ZN(n8367) );
  NOR2_X1 U9869 ( .A1(n8362), .A2(n8361), .ZN(n8366) );
  NOR2_X1 U9870 ( .A1(n8364), .A2(n8363), .ZN(n8365) );
  NAND4_X1 U9871 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8370)
         );
  NOR2_X1 U9872 ( .A1(n8370), .A2(n8369), .ZN(n8372) );
  NAND4_X1 U9873 ( .A1(n8372), .A2(n8655), .A3(n8658), .A4(n8371), .ZN(n8373)
         );
  NOR2_X1 U9874 ( .A1(n8373), .A2(n8664), .ZN(n8374) );
  NAND4_X1 U9875 ( .A1(n8963), .A2(n8666), .A3(n8374), .A4(n8975), .ZN(n8375)
         );
  NOR2_X1 U9876 ( .A1(n8938), .A2(n8375), .ZN(n8376) );
  NAND4_X1 U9877 ( .A1(n8866), .A2(n8377), .A3(n8376), .A4(n8873), .ZN(n8378)
         );
  NOR2_X1 U9878 ( .A1(n8378), .A2(n8844), .ZN(n8379) );
  NAND4_X1 U9879 ( .A1(n4546), .A2(n8836), .A3(n4635), .A4(n8379), .ZN(n8380)
         );
  NOR4_X1 U9880 ( .A1(n8742), .A2(n8788), .A3(n8769), .A4(n8380), .ZN(n8382)
         );
  NAND4_X1 U9881 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8724), .ZN(n8384)
         );
  XNOR2_X1 U9882 ( .A(n8387), .B(n8623), .ZN(n8390) );
  OAI22_X1 U9883 ( .A1(n8390), .A2(n5482), .B1(n8389), .B2(n8388), .ZN(n8391)
         );
  INV_X1 U9884 ( .A(n8391), .ZN(n8395) );
  INV_X1 U9885 ( .A(n8392), .ZN(n8393) );
  NAND2_X1 U9886 ( .A1(n8396), .A2(n8393), .ZN(n8394) );
  OAI21_X1 U9887 ( .B1(n8396), .B2(n8395), .A(n8394), .ZN(n8397) );
  NOR3_X1 U9888 ( .A1(n8399), .A2(n8398), .A3(n9012), .ZN(n8401) );
  OAI21_X1 U9889 ( .B1(n8402), .B2(n5967), .A(P2_B_REG_SCAN_IN), .ZN(n8400) );
  OAI222_X1 U9890 ( .A1(n8405), .A2(n8404), .B1(n9165), .B2(n8403), .C1(n8888), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9891 ( .A1(n9330), .A2(n8406), .ZN(n8408) );
  NAND2_X1 U9892 ( .A1(n9281), .A2(n8412), .ZN(n8407) );
  NAND2_X1 U9893 ( .A1(n8408), .A2(n8407), .ZN(n8410) );
  XNOR2_X1 U9894 ( .A(n8410), .B(n4311), .ZN(n8416) );
  INV_X1 U9895 ( .A(n8411), .ZN(n8414) );
  NAND2_X1 U9896 ( .A1(n9330), .A2(n8412), .ZN(n8413) );
  OAI21_X1 U9897 ( .B1(n9347), .B2(n8414), .A(n8413), .ZN(n8415) );
  XNOR2_X1 U9898 ( .A(n8416), .B(n8415), .ZN(n8417) );
  INV_X1 U9899 ( .A(n8417), .ZN(n8421) );
  NAND3_X1 U9900 ( .A1(n8421), .A2(n9694), .A3(n8420), .ZN(n8425) );
  AOI22_X1 U9901 ( .A1(n9685), .A2(n9366), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8419) );
  NAND2_X1 U9902 ( .A1(n9222), .A2(n9325), .ZN(n8418) );
  OAI211_X1 U9903 ( .C1(n9699), .C2(n9331), .A(n8419), .B(n8418), .ZN(n8423)
         );
  NOR3_X1 U9904 ( .A1(n8421), .A2(n8420), .A3(n9278), .ZN(n8422) );
  AOI211_X1 U9905 ( .C1(n9276), .C2(n9330), .A(n8423), .B(n8422), .ZN(n8424)
         );
  INV_X1 U9906 ( .A(n8516), .ZN(n8530) );
  AOI22_X1 U9907 ( .A1(n6000), .A2(n8532), .B1(n8530), .B2(n4549), .ZN(n8433)
         );
  OAI22_X1 U9908 ( .A1(n8539), .A2(n8459), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8427), .ZN(n8430) );
  INV_X1 U9909 ( .A(n8791), .ZN(n8428) );
  OAI22_X1 U9910 ( .A1(n8536), .A2(n8693), .B1(n8537), .B2(n8428), .ZN(n8429)
         );
  AOI211_X1 U9911 ( .C1(n9062), .C2(n8508), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9912 ( .B1(n8433), .B2(n8432), .A(n8431), .ZN(P2_U3218) );
  INV_X1 U9913 ( .A(n8434), .ZN(n8437) );
  NOR3_X1 U9914 ( .A1(n8435), .A2(n8687), .A3(n8516), .ZN(n8436) );
  AOI21_X1 U9915 ( .B1(n8437), .B2(n8532), .A(n8436), .ZN(n8444) );
  NAND2_X1 U9916 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8626) );
  OAI22_X1 U9917 ( .A1(n8690), .A2(n9014), .B1(n8687), .B2(n9012), .ZN(n8848)
         );
  NAND2_X1 U9918 ( .A1(n8460), .A2(n8848), .ZN(n8438) );
  OAI211_X1 U9919 ( .C1(n8537), .C2(n8852), .A(n8626), .B(n8438), .ZN(n8441)
         );
  NOR2_X1 U9920 ( .A1(n8439), .A2(n8518), .ZN(n8440) );
  AOI211_X1 U9921 ( .C1(n9083), .C2(n8508), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI21_X1 U9922 ( .B1(n8444), .B2(n8443), .A(n8442), .ZN(P2_U3221) );
  INV_X1 U9923 ( .A(n8446), .ZN(n8447) );
  AOI21_X1 U9924 ( .B1(n8445), .B2(n8447), .A(n8518), .ZN(n8451) );
  NOR3_X1 U9925 ( .A1(n8448), .A2(n8690), .A3(n8516), .ZN(n8450) );
  OAI21_X1 U9926 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8455) );
  INV_X1 U9927 ( .A(n8693), .ZN(n8822) );
  AOI22_X1 U9928 ( .A1(n8496), .A2(n8822), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8454) );
  INV_X1 U9929 ( .A(n8690), .ZN(n8821) );
  AOI22_X1 U9930 ( .A1(n8511), .A2(n8821), .B1(n8526), .B2(n8817), .ZN(n8453)
         );
  NAND2_X1 U9931 ( .A1(n9072), .A2(n8508), .ZN(n8452) );
  NAND4_X1 U9932 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(
        P2_U3225) );
  INV_X1 U9933 ( .A(n9053), .ZN(n8757) );
  OAI211_X1 U9934 ( .C1(n8458), .C2(n8457), .A(n8456), .B(n8532), .ZN(n8465)
         );
  OAI22_X1 U9935 ( .A1(n8546), .A2(n9014), .B1(n8459), .B2(n9012), .ZN(n8760)
         );
  INV_X1 U9936 ( .A(n8760), .ZN(n8462) );
  INV_X1 U9937 ( .A(n8460), .ZN(n8523) );
  OAI22_X1 U9938 ( .A1(n8462), .A2(n8523), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8461), .ZN(n8463) );
  AOI21_X1 U9939 ( .B1(n8764), .B2(n8526), .A(n8463), .ZN(n8464) );
  OAI211_X1 U9940 ( .C1(n8757), .C2(n8544), .A(n8465), .B(n8464), .ZN(P2_U3227) );
  XOR2_X1 U9941 ( .A(n8466), .B(n8467), .Z(n8472) );
  OAI21_X1 U9942 ( .B1(n8536), .B2(n8908), .A(n8468), .ZN(n8470) );
  OAI22_X1 U9943 ( .A1(n8539), .A2(n8686), .B1(n8537), .B2(n8915), .ZN(n8469)
         );
  AOI211_X1 U9944 ( .C1(n9097), .C2(n8508), .A(n8470), .B(n8469), .ZN(n8471)
         );
  OAI21_X1 U9945 ( .B1(n8472), .B2(n8518), .A(n8471), .ZN(P2_U3228) );
  INV_X1 U9946 ( .A(n8445), .ZN(n8473) );
  AOI211_X1 U9947 ( .C1(n8475), .C2(n8474), .A(n8518), .B(n8473), .ZN(n8479)
         );
  INV_X1 U9948 ( .A(n9077), .ZN(n8833) );
  INV_X1 U9949 ( .A(n8691), .ZN(n8838) );
  AOI22_X1 U9950 ( .A1(n8496), .A2(n8838), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8477) );
  AOI22_X1 U9951 ( .A1(n8511), .A2(n8868), .B1(n8526), .B2(n8831), .ZN(n8476)
         );
  OAI211_X1 U9952 ( .C1(n8833), .C2(n8544), .A(n8477), .B(n8476), .ZN(n8478)
         );
  OR2_X1 U9953 ( .A1(n8479), .A2(n8478), .ZN(P2_U3235) );
  NAND2_X1 U9954 ( .A1(n8530), .A2(n8822), .ZN(n8483) );
  NAND2_X1 U9955 ( .A1(n8532), .A2(n8480), .ZN(n8482) );
  MUX2_X1 U9956 ( .A(n8483), .B(n8482), .S(n8481), .Z(n8487) );
  AOI22_X1 U9957 ( .A1(n8511), .A2(n8838), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8486) );
  AOI22_X1 U9958 ( .A1(n8496), .A2(n4549), .B1(n8526), .B2(n8804), .ZN(n8485)
         );
  NAND2_X1 U9959 ( .A1(n9067), .A2(n8508), .ZN(n8484) );
  NAND4_X1 U9960 ( .A1(n8487), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(
        P2_U3237) );
  INV_X1 U9961 ( .A(n8488), .ZN(n8489) );
  AOI21_X1 U9962 ( .B1(n6040), .B2(n8489), .A(n8518), .ZN(n8492) );
  NOR3_X1 U9963 ( .A1(n8490), .A2(n8686), .A3(n8516), .ZN(n8491) );
  OAI21_X1 U9964 ( .B1(n8492), .B2(n8491), .A(n8434), .ZN(n8498) );
  NOR2_X1 U9965 ( .A1(n8493), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8598) );
  INV_X1 U9966 ( .A(n8861), .ZN(n8494) );
  OAI22_X1 U9967 ( .A1(n8536), .A2(n8686), .B1(n8537), .B2(n8494), .ZN(n8495)
         );
  AOI211_X1 U9968 ( .C1(n8496), .C2(n8868), .A(n8598), .B(n8495), .ZN(n8497)
         );
  OAI211_X1 U9969 ( .C1(n8863), .C2(n8544), .A(n8498), .B(n8497), .ZN(P2_U3240) );
  NAND2_X1 U9970 ( .A1(n8502), .A2(n8500), .ZN(n8501) );
  OAI21_X1 U9971 ( .B1(n8499), .B2(n8502), .A(n8501), .ZN(n8503) );
  NAND2_X1 U9972 ( .A1(n8503), .A2(n8532), .ZN(n8515) );
  OAI22_X1 U9973 ( .A1(n8539), .A2(n8505), .B1(n8537), .B2(n8504), .ZN(n8506)
         );
  NOR3_X1 U9974 ( .A1(n8516), .A2(n8510), .A3(n8499), .ZN(n8512) );
  OAI21_X1 U9975 ( .B1(n8512), .B2(n8511), .A(n8552), .ZN(n8513) );
  NAND3_X1 U9976 ( .A1(n8515), .A2(n8514), .A3(n8513), .ZN(P2_U3241) );
  INV_X1 U9977 ( .A(n9048), .ZN(n8630) );
  NOR3_X1 U9978 ( .A1(n8517), .A2(n8781), .A3(n8516), .ZN(n8521) );
  AOI21_X1 U9979 ( .B1(n8456), .B2(n8519), .A(n8518), .ZN(n8520) );
  OAI21_X1 U9980 ( .B1(n8521), .B2(n8520), .A(n4334), .ZN(n8529) );
  INV_X1 U9981 ( .A(n8740), .ZN(n8527) );
  OAI22_X1 U9982 ( .A1(n8545), .A2(n9014), .B1(n8781), .B2(n9012), .ZN(n8745)
         );
  INV_X1 U9983 ( .A(n8745), .ZN(n8524) );
  OAI22_X1 U9984 ( .A1(n8524), .A2(n8523), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8522), .ZN(n8525) );
  AOI21_X1 U9985 ( .B1(n8527), .B2(n8526), .A(n8525), .ZN(n8528) );
  OAI211_X1 U9986 ( .C1(n8630), .C2(n8544), .A(n8529), .B(n8528), .ZN(P2_U3242) );
  INV_X1 U9987 ( .A(n9106), .ZN(n8942) );
  NAND2_X1 U9988 ( .A1(n8530), .A2(n8967), .ZN(n8535) );
  NAND2_X1 U9989 ( .A1(n8532), .A2(n8531), .ZN(n8534) );
  MUX2_X1 U9990 ( .A(n8535), .B(n8534), .S(n8533), .Z(n8543) );
  NOR2_X1 U9991 ( .A1(n8536), .A2(n8977), .ZN(n8541) );
  OAI22_X1 U9992 ( .A1(n8539), .A2(n8538), .B1(n8537), .B2(n8944), .ZN(n8540)
         );
  AOI211_X1 U9993 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(P2_U3152), .A(n8541), 
        .B(n8540), .ZN(n8542) );
  OAI211_X1 U9994 ( .C1(n8942), .C2(n8544), .A(n8543), .B(n8542), .ZN(P2_U3243) );
  MUX2_X1 U9995 ( .A(n8646), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8556), .Z(
        P2_U3582) );
  MUX2_X1 U9996 ( .A(n8725), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8556), .Z(
        P2_U3580) );
  INV_X1 U9997 ( .A(n8545), .ZN(n8711) );
  MUX2_X1 U9998 ( .A(n8711), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8556), .Z(
        P2_U3579) );
  INV_X1 U9999 ( .A(n8546), .ZN(n8726) );
  MUX2_X1 U10000 ( .A(n8726), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8556), .Z(
        P2_U3578) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8695), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8796), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n4549), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8822), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8838), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10006 ( .A(n8821), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8556), .Z(
        P2_U3572) );
  MUX2_X1 U10007 ( .A(n8868), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8556), .Z(
        P2_U3571) );
  MUX2_X1 U10008 ( .A(n8879), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8556), .Z(
        P2_U3570) );
  MUX2_X1 U10009 ( .A(n8906), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8556), .Z(
        P2_U3569) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8929), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8967), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n4646), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10013 ( .A(n8966), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8556), .Z(
        P2_U3565) );
  INV_X1 U10014 ( .A(n8978), .ZN(n8670) );
  MUX2_X1 U10015 ( .A(n8670), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8556), .Z(
        P2_U3564) );
  MUX2_X1 U10016 ( .A(n8651), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8556), .Z(
        P2_U3563) );
  MUX2_X1 U10017 ( .A(n8547), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8556), .Z(
        P2_U3562) );
  MUX2_X1 U10018 ( .A(n8548), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8556), .Z(
        P2_U3561) );
  MUX2_X1 U10019 ( .A(n8549), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8556), .Z(
        P2_U3560) );
  MUX2_X1 U10020 ( .A(n8550), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8556), .Z(
        P2_U3559) );
  MUX2_X1 U10021 ( .A(n8551), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8556), .Z(
        P2_U3558) );
  MUX2_X1 U10022 ( .A(n8552), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8556), .Z(
        P2_U3557) );
  MUX2_X1 U10023 ( .A(n8553), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8556), .Z(
        P2_U3556) );
  MUX2_X1 U10024 ( .A(n8554), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8556), .Z(
        P2_U3555) );
  MUX2_X1 U10025 ( .A(n8555), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8556), .Z(
        P2_U3554) );
  MUX2_X1 U10026 ( .A(n6483), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8556), .Z(
        P2_U3553) );
  MUX2_X1 U10027 ( .A(n8557), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8556), .Z(
        P2_U3552) );
  OAI211_X1 U10028 ( .C1(n8560), .C2(n8559), .A(n8613), .B(n8558), .ZN(n8569)
         );
  AOI22_X1 U10029 ( .A1(n8599), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8568) );
  NAND2_X1 U10030 ( .A1(n8562), .A2(n8561), .ZN(n8567) );
  OAI211_X1 U10031 ( .C1(n8565), .C2(n8564), .A(n8612), .B(n8563), .ZN(n8566)
         );
  NAND4_X1 U10032 ( .A1(n8569), .A2(n8568), .A3(n8567), .A4(n8566), .ZN(
        P2_U3247) );
  OAI211_X1 U10033 ( .C1(n8572), .C2(n8571), .A(n8613), .B(n8570), .ZN(n8586)
         );
  AOI21_X1 U10034 ( .B1(n8599), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8573), .ZN(
        n8585) );
  OR2_X1 U10035 ( .A1(n8619), .A2(n8574), .ZN(n8584) );
  MUX2_X1 U10036 ( .A(n8576), .B(P2_REG1_REG_4__SCAN_IN), .S(n8575), .Z(n8579)
         );
  INV_X1 U10037 ( .A(n8577), .ZN(n8578) );
  NAND2_X1 U10038 ( .A1(n8579), .A2(n8578), .ZN(n8581) );
  OAI211_X1 U10039 ( .C1(n8582), .C2(n8581), .A(n8612), .B(n8580), .ZN(n8583)
         );
  NAND4_X1 U10040 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(
        P2_U3249) );
  INV_X1 U10041 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8589) );
  OAI21_X1 U10042 ( .B1(n8589), .B2(n8588), .A(n8587), .ZN(n8591) );
  INV_X1 U10043 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8610) );
  AOI22_X1 U10044 ( .A1(n8594), .A2(n8610), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8609), .ZN(n8590) );
  NOR2_X1 U10045 ( .A1(n8591), .A2(n8590), .ZN(n8608) );
  AOI21_X1 U10046 ( .B1(n8591), .B2(n8590), .A(n8608), .ZN(n8602) );
  NAND2_X1 U10047 ( .A1(n8595), .A2(n5795), .ZN(n8605) );
  OAI21_X1 U10048 ( .B1(n8595), .B2(n5795), .A(n8605), .ZN(n8596) );
  NAND2_X1 U10049 ( .A1(n8596), .A2(n8613), .ZN(n8601) );
  NOR2_X1 U10050 ( .A1(n8619), .A2(n8609), .ZN(n8597) );
  AOI211_X1 U10051 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n8599), .A(n8598), .B(
        n8597), .ZN(n8600) );
  OAI211_X1 U10052 ( .C1(n8602), .C2(n8620), .A(n8601), .B(n8600), .ZN(
        P2_U3263) );
  INV_X1 U10053 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10054 ( .A1(n8603), .A2(n8609), .ZN(n8604) );
  NAND2_X1 U10055 ( .A1(n8605), .A2(n8604), .ZN(n8607) );
  XOR2_X1 U10056 ( .A(n8607), .B(n8606), .Z(n8615) );
  AOI21_X1 U10057 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8611) );
  XOR2_X1 U10058 ( .A(n8611), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8621) );
  AOI22_X1 U10059 ( .A1(n8615), .A2(n8613), .B1(n8612), .B2(n8621), .ZN(n8625)
         );
  INV_X1 U10060 ( .A(n8614), .ZN(n8617) );
  INV_X1 U10061 ( .A(n8615), .ZN(n8616) );
  NAND2_X1 U10062 ( .A1(n8617), .A2(n8616), .ZN(n8618) );
  OAI211_X1 U10063 ( .C1(n8621), .C2(n8620), .A(n8619), .B(n8618), .ZN(n8622)
         );
  INV_X1 U10064 ( .A(n8622), .ZN(n8624) );
  MUX2_X1 U10065 ( .A(n8625), .B(n8624), .S(n8623), .Z(n8627) );
  OAI211_X1 U10066 ( .C1(n8629), .C2(n8628), .A(n8627), .B(n8626), .ZN(
        P2_U3264) );
  INV_X1 U10067 ( .A(n9116), .ZN(n8991) );
  INV_X1 U10068 ( .A(n9111), .ZN(n8959) );
  INV_X1 U10069 ( .A(n9067), .ZN(n8806) );
  NAND2_X1 U10070 ( .A1(n8702), .A2(n9708), .ZN(n8631) );
  AND2_X1 U10071 ( .A1(n8632), .A2(P2_B_REG_SCAN_IN), .ZN(n8633) );
  NOR2_X1 U10072 ( .A1(n9014), .A2(n8633), .ZN(n8647) );
  NAND2_X1 U10073 ( .A1(n8634), .A2(n8647), .ZN(n9707) );
  NOR2_X1 U10074 ( .A1(n9019), .A2(n9707), .ZN(n8640) );
  NOR2_X1 U10075 ( .A1(n8946), .A2(n8635), .ZN(n8636) );
  AOI211_X1 U10076 ( .C1(n9025), .C2(n8892), .A(n8640), .B(n8636), .ZN(n8637)
         );
  OAI21_X1 U10077 ( .B1(n9027), .B2(n8638), .A(n8637), .ZN(P2_U3265) );
  XNOR2_X1 U10078 ( .A(n8702), .B(n8639), .ZN(n9710) );
  NAND2_X1 U10079 ( .A1(n9710), .A2(n8995), .ZN(n8642) );
  AOI21_X1 U10080 ( .B1(n9019), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8640), .ZN(
        n8641) );
  OAI211_X1 U10081 ( .C1(n9708), .C2(n9008), .A(n8642), .B(n8641), .ZN(
        P2_U3266) );
  OAI21_X1 U10082 ( .B1(n8645), .B2(n8643), .A(n8644), .ZN(n8650) );
  AOI22_X1 U10083 ( .A1(n8725), .A2(n8965), .B1(n8647), .B2(n8646), .ZN(n8648)
         );
  INV_X1 U10084 ( .A(n8648), .ZN(n8649) );
  AOI21_X1 U10085 ( .B1(n8650), .B2(n8986), .A(n8649), .ZN(n9031) );
  INV_X1 U10086 ( .A(n9062), .ZN(n8793) );
  NAND2_X1 U10087 ( .A1(n8652), .A2(n8651), .ZN(n8663) );
  AND2_X1 U10088 ( .A1(n8653), .A2(n8663), .ZN(n8997) );
  INV_X1 U10089 ( .A(n8666), .ZN(n8654) );
  NAND2_X1 U10090 ( .A1(n8997), .A2(n8654), .ZN(n8662) );
  OR2_X1 U10091 ( .A1(n8655), .A2(n8662), .ZN(n8657) );
  NOR2_X1 U10092 ( .A1(n8657), .A2(n8656), .ZN(n8669) );
  INV_X1 U10093 ( .A(n8658), .ZN(n8660) );
  AND2_X1 U10094 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  OR2_X1 U10095 ( .A1(n8662), .A2(n8661), .ZN(n8668) );
  INV_X1 U10096 ( .A(n8663), .ZN(n8665) );
  OR2_X1 U10097 ( .A1(n8665), .A2(n8664), .ZN(n8999) );
  OR2_X1 U10098 ( .A1(n8666), .A2(n8999), .ZN(n8667) );
  OR2_X1 U10099 ( .A1(n9111), .A2(n4646), .ZN(n8675) );
  AND2_X1 U10100 ( .A1(n8980), .A2(n8675), .ZN(n8932) );
  OR2_X1 U10101 ( .A1(n9106), .A2(n8967), .ZN(n8679) );
  AND2_X1 U10102 ( .A1(n8932), .A2(n8679), .ZN(n8897) );
  OR2_X1 U10103 ( .A1(n9121), .A2(n8670), .ZN(n8895) );
  AND2_X1 U10104 ( .A1(n8897), .A2(n8895), .ZN(n8672) );
  NAND2_X1 U10105 ( .A1(n9097), .A2(n8929), .ZN(n8680) );
  INV_X1 U10106 ( .A(n8680), .ZN(n8671) );
  AND2_X1 U10107 ( .A1(n8672), .A2(n8674), .ZN(n8673) );
  NAND2_X1 U10108 ( .A1(n8896), .A2(n8673), .ZN(n8684) );
  INV_X1 U10109 ( .A(n8674), .ZN(n8682) );
  INV_X1 U10110 ( .A(n8675), .ZN(n8678) );
  INV_X1 U10111 ( .A(n8951), .ZN(n8676) );
  NOR2_X1 U10112 ( .A1(n8963), .A2(n8676), .ZN(n8677) );
  OR2_X1 U10113 ( .A1(n8678), .A2(n8677), .ZN(n8933) );
  AND2_X1 U10114 ( .A1(n8898), .A2(n8680), .ZN(n8681) );
  NAND2_X1 U10115 ( .A1(n8684), .A2(n8683), .ZN(n8874) );
  NAND2_X1 U10116 ( .A1(n8845), .A2(n8844), .ZN(n8843) );
  INV_X1 U10117 ( .A(n9083), .ZN(n8689) );
  NAND2_X1 U10118 ( .A1(n8843), .A2(n4749), .ZN(n8829) );
  NAND2_X1 U10119 ( .A1(n8829), .A2(n8828), .ZN(n8827) );
  NAND2_X1 U10120 ( .A1(n8827), .A2(n4748), .ZN(n8814) );
  NAND2_X1 U10121 ( .A1(n8819), .A2(n8691), .ZN(n8692) );
  OAI22_X1 U10122 ( .A1(n8770), .A2(n8776), .B1(n8796), .B2(n9057), .ZN(n8755)
         );
  NAND2_X1 U10123 ( .A1(n8755), .A2(n8758), .ZN(n8754) );
  NAND2_X1 U10124 ( .A1(n8754), .A2(n8696), .ZN(n8738) );
  NAND2_X1 U10125 ( .A1(n8715), .A2(n8714), .ZN(n8713) );
  NAND2_X1 U10126 ( .A1(n8713), .A2(n8699), .ZN(n8701) );
  XNOR2_X1 U10127 ( .A(n8701), .B(n8700), .ZN(n9028) );
  NAND2_X1 U10128 ( .A1(n9028), .A2(n8940), .ZN(n8708) );
  AOI21_X1 U10129 ( .B1(n9029), .B2(n8716), .A(n8702), .ZN(n9030) );
  INV_X1 U10130 ( .A(n8703), .ZN(n8704) );
  AOI22_X1 U10131 ( .A1(n9019), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8704), .B2(
        n9005), .ZN(n8705) );
  OAI21_X1 U10132 ( .B1(n4735), .B2(n9008), .A(n8705), .ZN(n8706) );
  AOI21_X1 U10133 ( .B1(n9030), .B2(n9022), .A(n8706), .ZN(n8707) );
  OAI211_X1 U10134 ( .C1(n9031), .C2(n9019), .A(n8708), .B(n8707), .ZN(
        P2_U3267) );
  XNOR2_X1 U10135 ( .A(n8709), .B(n8714), .ZN(n8712) );
  AOI222_X2 U10136 ( .A1(n8986), .A2(n8712), .B1(n8711), .B2(n8965), .C1(n8710), .C2(n8968), .ZN(n9039) );
  OAI21_X1 U10137 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n9035) );
  NAND2_X1 U10138 ( .A1(n9035), .A2(n8940), .ZN(n8723) );
  INV_X1 U10139 ( .A(n8716), .ZN(n8717) );
  AOI21_X1 U10140 ( .B1(n9036), .B2(n8730), .A(n8717), .ZN(n9037) );
  INV_X1 U10141 ( .A(n8718), .ZN(n8719) );
  AOI22_X1 U10142 ( .A1(n9019), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8719), .B2(
        n9005), .ZN(n8720) );
  OAI21_X1 U10143 ( .B1(n4737), .B2(n9008), .A(n8720), .ZN(n8721) );
  AOI21_X1 U10144 ( .B1(n9037), .B2(n8995), .A(n8721), .ZN(n8722) );
  OAI211_X1 U10145 ( .C1(n9019), .C2(n9039), .A(n8723), .B(n8722), .ZN(
        P2_U3268) );
  OAI21_X1 U10146 ( .B1(n8729), .B2(n8728), .A(n8727), .ZN(n9041) );
  NAND2_X1 U10147 ( .A1(n9041), .A2(n8940), .ZN(n8736) );
  INV_X1 U10148 ( .A(n8730), .ZN(n8731) );
  AOI21_X1 U10149 ( .B1(n9042), .B2(n8747), .A(n8731), .ZN(n9043) );
  AOI22_X1 U10150 ( .A1(n9019), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8732), .B2(
        n9005), .ZN(n8733) );
  OAI21_X1 U10151 ( .B1(n8698), .B2(n9008), .A(n8733), .ZN(n8734) );
  AOI21_X1 U10152 ( .B1(n9043), .B2(n8995), .A(n8734), .ZN(n8735) );
  OAI211_X1 U10153 ( .C1(n9019), .C2(n9045), .A(n8736), .B(n8735), .ZN(
        P2_U3269) );
  OAI21_X1 U10154 ( .B1(n8738), .B2(n8742), .A(n8737), .ZN(n8739) );
  INV_X1 U10155 ( .A(n8739), .ZN(n9051) );
  INV_X1 U10156 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8741) );
  OAI22_X1 U10157 ( .A1(n8946), .A2(n8741), .B1(n8740), .B2(n8943), .ZN(n8752)
         );
  OAI21_X1 U10158 ( .B1(n8744), .B2(n8186), .A(n8743), .ZN(n8746) );
  AOI21_X1 U10159 ( .B1(n8746), .B2(n8986), .A(n8745), .ZN(n9050) );
  INV_X1 U10160 ( .A(n8762), .ZN(n8749) );
  INV_X1 U10161 ( .A(n9993), .ZN(n10020) );
  INV_X1 U10162 ( .A(n8747), .ZN(n8748) );
  AOI211_X1 U10163 ( .C1(n9048), .C2(n8749), .A(n10020), .B(n8748), .ZN(n9047)
         );
  NAND2_X1 U10164 ( .A1(n9047), .A2(n8888), .ZN(n8750) );
  AOI21_X1 U10165 ( .B1(n9050), .B2(n8750), .A(n9019), .ZN(n8751) );
  AOI211_X1 U10166 ( .C1(n8892), .C2(n9048), .A(n8752), .B(n8751), .ZN(n8753)
         );
  OAI21_X1 U10167 ( .B1(n9051), .B2(n9024), .A(n8753), .ZN(P2_U3270) );
  OAI21_X1 U10168 ( .B1(n8755), .B2(n8758), .A(n8754), .ZN(n8756) );
  INV_X1 U10169 ( .A(n8756), .ZN(n9056) );
  NOR2_X1 U10170 ( .A1(n8757), .A2(n9008), .ZN(n8767) );
  XNOR2_X1 U10171 ( .A(n8759), .B(n8758), .ZN(n8761) );
  AOI21_X1 U10172 ( .B1(n8761), .B2(n8986), .A(n8760), .ZN(n9055) );
  INV_X1 U10173 ( .A(n8771), .ZN(n8763) );
  AOI211_X1 U10174 ( .C1(n9053), .C2(n8763), .A(n10020), .B(n8762), .ZN(n9052)
         );
  AOI22_X1 U10175 ( .A1(n9052), .A2(n8888), .B1(n9005), .B2(n8764), .ZN(n8765)
         );
  AOI21_X1 U10176 ( .B1(n9055), .B2(n8765), .A(n9019), .ZN(n8766) );
  AOI211_X1 U10177 ( .C1(n9019), .C2(P2_REG2_REG_25__SCAN_IN), .A(n8767), .B(
        n8766), .ZN(n8768) );
  OAI21_X1 U10178 ( .B1(n9056), .B2(n9024), .A(n8768), .ZN(P2_U3271) );
  XNOR2_X1 U10179 ( .A(n8770), .B(n8769), .ZN(n9061) );
  AOI21_X1 U10180 ( .B1(n9057), .B2(n8790), .A(n8771), .ZN(n9058) );
  AOI22_X1 U10181 ( .A1(n9019), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8772), .B2(
        n9005), .ZN(n8773) );
  OAI21_X1 U10182 ( .B1(n8774), .B2(n9008), .A(n8773), .ZN(n8785) );
  INV_X1 U10183 ( .A(n8775), .ZN(n8779) );
  AOI21_X1 U10184 ( .B1(n8794), .B2(n8777), .A(n8776), .ZN(n8778) );
  NOR3_X1 U10185 ( .A1(n8779), .A2(n8778), .A3(n9010), .ZN(n8783) );
  OAI22_X1 U10186 ( .A1(n8781), .A2(n9014), .B1(n8780), .B2(n9012), .ZN(n8782)
         );
  NOR2_X1 U10187 ( .A1(n8783), .A2(n8782), .ZN(n9060) );
  NOR2_X1 U10188 ( .A1(n9060), .A2(n9019), .ZN(n8784) );
  AOI211_X1 U10189 ( .C1(n9058), .C2(n8995), .A(n8785), .B(n8784), .ZN(n8786)
         );
  OAI21_X1 U10190 ( .B1(n9061), .B2(n9024), .A(n8786), .ZN(P2_U3272) );
  OAI21_X1 U10191 ( .B1(n8789), .B2(n8788), .A(n8787), .ZN(n9066) );
  AOI21_X1 U10192 ( .B1(n9062), .B2(n8802), .A(n4739), .ZN(n9063) );
  AOI22_X1 U10193 ( .A1(n9019), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8791), .B2(
        n9005), .ZN(n8792) );
  OAI21_X1 U10194 ( .B1(n8793), .B2(n9008), .A(n8792), .ZN(n8799) );
  OAI21_X1 U10195 ( .B1(n8795), .B2(n4541), .A(n8794), .ZN(n8797) );
  AOI222_X1 U10196 ( .A1(n8986), .A2(n8797), .B1(n8822), .B2(n8965), .C1(n8796), .C2(n8968), .ZN(n9065) );
  NOR2_X1 U10197 ( .A1(n9065), .A2(n9019), .ZN(n8798) );
  AOI211_X1 U10198 ( .C1(n9063), .C2(n9022), .A(n8799), .B(n8798), .ZN(n8800)
         );
  OAI21_X1 U10199 ( .B1(n9066), .B2(n9024), .A(n8800), .ZN(P2_U3273) );
  XNOR2_X1 U10200 ( .A(n8801), .B(n4546), .ZN(n9071) );
  INV_X1 U10201 ( .A(n8815), .ZN(n8803) );
  AOI21_X1 U10202 ( .B1(n9067), .B2(n8803), .A(n4740), .ZN(n9068) );
  AOI22_X1 U10203 ( .A1(n9019), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8804), .B2(
        n9005), .ZN(n8805) );
  OAI21_X1 U10204 ( .B1(n8806), .B2(n9008), .A(n8805), .ZN(n8811) );
  NAND2_X1 U10205 ( .A1(n8820), .A2(n8807), .ZN(n8808) );
  XNOR2_X1 U10206 ( .A(n8808), .B(n4546), .ZN(n8809) );
  AOI222_X1 U10207 ( .A1(n8986), .A2(n8809), .B1(n8838), .B2(n8965), .C1(n4549), .C2(n8968), .ZN(n9070) );
  NOR2_X1 U10208 ( .A1(n9070), .A2(n9019), .ZN(n8810) );
  AOI211_X1 U10209 ( .C1(n9068), .C2(n8995), .A(n8811), .B(n8810), .ZN(n8812)
         );
  OAI21_X1 U10210 ( .B1(n9071), .B2(n9024), .A(n8812), .ZN(P2_U3274) );
  XNOR2_X1 U10211 ( .A(n8814), .B(n8813), .ZN(n9076) );
  INV_X1 U10212 ( .A(n8830), .ZN(n8816) );
  AOI21_X1 U10213 ( .B1(n9072), .B2(n8816), .A(n8815), .ZN(n9073) );
  AOI22_X1 U10214 ( .A1(n9019), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8817), .B2(
        n9005), .ZN(n8818) );
  OAI21_X1 U10215 ( .B1(n8819), .B2(n9008), .A(n8818), .ZN(n8825) );
  OAI21_X1 U10216 ( .B1(n4347), .B2(n4635), .A(n8820), .ZN(n8823) );
  AOI222_X1 U10217 ( .A1(n8986), .A2(n8823), .B1(n8822), .B2(n8968), .C1(n8821), .C2(n8965), .ZN(n9075) );
  NOR2_X1 U10218 ( .A1(n9075), .A2(n9019), .ZN(n8824) );
  AOI211_X1 U10219 ( .C1(n9073), .C2(n9022), .A(n8825), .B(n8824), .ZN(n8826)
         );
  OAI21_X1 U10220 ( .B1(n9076), .B2(n9024), .A(n8826), .ZN(P2_U3275) );
  OAI21_X1 U10221 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n9081) );
  AOI21_X1 U10222 ( .B1(n9077), .B2(n4754), .A(n8830), .ZN(n9078) );
  AOI22_X1 U10223 ( .A1(n9019), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8831), .B2(
        n9005), .ZN(n8832) );
  OAI21_X1 U10224 ( .B1(n8833), .B2(n9008), .A(n8832), .ZN(n8841) );
  NAND2_X1 U10225 ( .A1(n8834), .A2(n8835), .ZN(n8837) );
  XNOR2_X1 U10226 ( .A(n8837), .B(n8836), .ZN(n8839) );
  AOI222_X1 U10227 ( .A1(n8986), .A2(n8839), .B1(n8838), .B2(n8968), .C1(n8868), .C2(n8965), .ZN(n9080) );
  NOR2_X1 U10228 ( .A1(n9080), .A2(n9019), .ZN(n8840) );
  AOI211_X1 U10229 ( .C1(n9078), .C2(n8995), .A(n8841), .B(n8840), .ZN(n8842)
         );
  OAI21_X1 U10230 ( .B1(n9081), .B2(n9024), .A(n8842), .ZN(P2_U3276) );
  OAI21_X1 U10231 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n9086) );
  AOI22_X1 U10232 ( .A1(n9083), .A2(n8892), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9019), .ZN(n8855) );
  OAI21_X1 U10233 ( .B1(n8847), .B2(n8846), .A(n8834), .ZN(n8849) );
  AOI21_X1 U10234 ( .B1(n8849), .B2(n8986), .A(n8848), .ZN(n9085) );
  INV_X1 U10235 ( .A(n4754), .ZN(n8850) );
  AOI211_X1 U10236 ( .C1(n9083), .C2(n8858), .A(n10020), .B(n8850), .ZN(n9082)
         );
  NAND2_X1 U10237 ( .A1(n9082), .A2(n8888), .ZN(n8851) );
  OAI211_X1 U10238 ( .C1(n8943), .C2(n8852), .A(n9085), .B(n8851), .ZN(n8853)
         );
  NAND2_X1 U10239 ( .A1(n8853), .A2(n8946), .ZN(n8854) );
  OAI211_X1 U10240 ( .C1(n9086), .C2(n9024), .A(n8855), .B(n8854), .ZN(
        P2_U3277) );
  XNOR2_X1 U10241 ( .A(n8857), .B(n8856), .ZN(n9091) );
  INV_X1 U10242 ( .A(n8887), .ZN(n8860) );
  INV_X1 U10243 ( .A(n8858), .ZN(n8859) );
  AOI21_X1 U10244 ( .B1(n9087), .B2(n8860), .A(n8859), .ZN(n9088) );
  AOI22_X1 U10245 ( .A1(n9019), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8861), .B2(
        n9005), .ZN(n8862) );
  OAI21_X1 U10246 ( .B1(n8863), .B2(n9008), .A(n8862), .ZN(n8871) );
  INV_X1 U10247 ( .A(n8864), .ZN(n8867) );
  OAI21_X1 U10248 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8869) );
  AOI222_X1 U10249 ( .A1(n8986), .A2(n8869), .B1(n8868), .B2(n8968), .C1(n8906), .C2(n8965), .ZN(n9090) );
  NOR2_X1 U10250 ( .A1(n9090), .A2(n9019), .ZN(n8870) );
  AOI211_X1 U10251 ( .C1(n9088), .C2(n8995), .A(n8871), .B(n8870), .ZN(n8872)
         );
  OAI21_X1 U10252 ( .B1(n9091), .B2(n9024), .A(n8872), .ZN(P2_U3278) );
  AND2_X1 U10253 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  OR2_X1 U10254 ( .A1(n8876), .A2(n8875), .ZN(n8884) );
  INV_X1 U10255 ( .A(n8884), .ZN(n9096) );
  XNOR2_X1 U10256 ( .A(n8878), .B(n8877), .ZN(n8881) );
  AOI22_X1 U10257 ( .A1(n8929), .A2(n8965), .B1(n8968), .B2(n8879), .ZN(n8880)
         );
  OAI21_X1 U10258 ( .B1(n8881), .B2(n9010), .A(n8880), .ZN(n8882) );
  AOI21_X1 U10259 ( .B1(n8884), .B2(n8883), .A(n8882), .ZN(n9095) );
  NAND2_X1 U10260 ( .A1(n8914), .A2(n9093), .ZN(n8885) );
  NAND2_X1 U10261 ( .A1(n8885), .A2(n9993), .ZN(n8886) );
  NOR2_X1 U10262 ( .A1(n8887), .A2(n8886), .ZN(n9092) );
  NAND2_X1 U10263 ( .A1(n9092), .A2(n8888), .ZN(n8889) );
  OAI211_X1 U10264 ( .C1(n8943), .C2(n8890), .A(n9095), .B(n8889), .ZN(n8891)
         );
  NAND2_X1 U10265 ( .A1(n8891), .A2(n8946), .ZN(n8894) );
  AOI22_X1 U10266 ( .A1(n9093), .A2(n8892), .B1(n9019), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8893) );
  OAI211_X1 U10267 ( .C1(n9096), .C2(n8992), .A(n8894), .B(n8893), .ZN(
        P2_U3279) );
  NAND2_X1 U10268 ( .A1(n8981), .A2(n8897), .ZN(n8899) );
  NAND2_X1 U10269 ( .A1(n8899), .A2(n8898), .ZN(n8901) );
  NAND2_X1 U10270 ( .A1(n8901), .A2(n8904), .ZN(n8900) );
  OAI21_X1 U10271 ( .B1(n8901), .B2(n8904), .A(n8900), .ZN(n9100) );
  OR2_X1 U10272 ( .A1(n9100), .A2(n8982), .ZN(n8912) );
  NAND2_X1 U10273 ( .A1(n8903), .A2(n8902), .ZN(n8905) );
  XNOR2_X1 U10274 ( .A(n8905), .B(n8904), .ZN(n8910) );
  NAND2_X1 U10275 ( .A1(n8906), .A2(n8968), .ZN(n8907) );
  OAI21_X1 U10276 ( .B1(n8908), .B2(n9012), .A(n8907), .ZN(n8909) );
  AOI21_X1 U10277 ( .B1(n8910), .B2(n8986), .A(n8909), .ZN(n8911) );
  NAND2_X1 U10278 ( .A1(n8912), .A2(n8911), .ZN(n9102) );
  NAND2_X1 U10279 ( .A1(n9102), .A2(n8946), .ZN(n8920) );
  NAND2_X1 U10280 ( .A1(n8941), .A2(n9097), .ZN(n8913) );
  AND2_X1 U10281 ( .A1(n8914), .A2(n8913), .ZN(n9098) );
  NOR2_X1 U10282 ( .A1(n4726), .A2(n9008), .ZN(n8918) );
  INV_X1 U10283 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8916) );
  OAI22_X1 U10284 ( .A1(n8946), .A2(n8916), .B1(n8915), .B2(n8943), .ZN(n8917)
         );
  AOI211_X1 U10285 ( .C1(n9098), .C2(n8995), .A(n8918), .B(n8917), .ZN(n8919)
         );
  OAI211_X1 U10286 ( .C1(n8992), .C2(n9100), .A(n8920), .B(n8919), .ZN(
        P2_U3280) );
  AND2_X1 U10287 ( .A1(n9017), .A2(n8921), .ZN(n8976) );
  NAND2_X1 U10288 ( .A1(n8976), .A2(n8922), .ZN(n8925) );
  AND2_X1 U10289 ( .A1(n8925), .A2(n8923), .ZN(n8928) );
  NAND2_X1 U10290 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  OAI211_X1 U10291 ( .C1(n8928), .C2(n8927), .A(n8926), .B(n8986), .ZN(n8931)
         );
  AOI22_X1 U10292 ( .A1(n8965), .A2(n4646), .B1(n8929), .B2(n8968), .ZN(n8930)
         );
  NAND2_X1 U10293 ( .A1(n8981), .A2(n8932), .ZN(n8936) );
  AND2_X1 U10294 ( .A1(n8936), .A2(n8933), .ZN(n8939) );
  INV_X1 U10295 ( .A(n8934), .ZN(n8935) );
  NAND2_X1 U10296 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  OAI21_X1 U10297 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n9105) );
  NAND2_X1 U10298 ( .A1(n9105), .A2(n8940), .ZN(n8950) );
  AOI21_X1 U10299 ( .B1(n9106), .B2(n8953), .A(n4727), .ZN(n9107) );
  NOR2_X1 U10300 ( .A1(n8942), .A2(n9008), .ZN(n8948) );
  OAI22_X1 U10301 ( .A1(n8946), .A2(n8945), .B1(n8944), .B2(n8943), .ZN(n8947)
         );
  AOI211_X1 U10302 ( .C1(n9107), .C2(n8995), .A(n8948), .B(n8947), .ZN(n8949)
         );
  OAI211_X1 U10303 ( .C1(n9019), .C2(n9109), .A(n8950), .B(n8949), .ZN(
        P2_U3281) );
  NAND2_X1 U10304 ( .A1(n8981), .A2(n8980), .ZN(n8979) );
  NAND2_X1 U10305 ( .A1(n8979), .A2(n8951), .ZN(n8952) );
  XOR2_X1 U10306 ( .A(n8963), .B(n8952), .Z(n9115) );
  INV_X1 U10307 ( .A(n8987), .ZN(n8955) );
  INV_X1 U10308 ( .A(n8953), .ZN(n8954) );
  AOI21_X1 U10309 ( .B1(n9111), .B2(n8955), .A(n8954), .ZN(n9112) );
  INV_X1 U10310 ( .A(n8956), .ZN(n8957) );
  AOI22_X1 U10311 ( .A1(n9019), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8957), .B2(
        n9005), .ZN(n8958) );
  OAI21_X1 U10312 ( .B1(n8959), .B2(n9008), .A(n8958), .ZN(n8972) );
  NAND2_X1 U10313 ( .A1(n8976), .A2(n8975), .ZN(n8974) );
  AND2_X1 U10314 ( .A1(n8974), .A2(n8960), .ZN(n8964) );
  NAND2_X1 U10315 ( .A1(n8974), .A2(n8961), .ZN(n8962) );
  OAI211_X1 U10316 ( .C1(n8964), .C2(n8963), .A(n8962), .B(n8986), .ZN(n8970)
         );
  AOI22_X1 U10317 ( .A1(n8968), .A2(n8967), .B1(n8966), .B2(n8965), .ZN(n8969)
         );
  NOR2_X1 U10318 ( .A1(n9114), .A2(n9019), .ZN(n8971) );
  AOI211_X1 U10319 ( .C1(n9112), .C2(n9022), .A(n8972), .B(n8971), .ZN(n8973)
         );
  OAI21_X1 U10320 ( .B1(n9024), .B2(n9115), .A(n8973), .ZN(P2_U3282) );
  OAI21_X1 U10321 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8985) );
  OAI22_X1 U10322 ( .A1(n8978), .A2(n9012), .B1(n8977), .B2(n9014), .ZN(n8984)
         );
  OAI21_X1 U10323 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n9120) );
  NOR2_X1 U10324 ( .A1(n9120), .A2(n8982), .ZN(n8983) );
  AOI211_X1 U10325 ( .C1(n8986), .C2(n8985), .A(n8984), .B(n8983), .ZN(n9119)
         );
  AOI21_X1 U10326 ( .B1(n9116), .B2(n4733), .A(n8987), .ZN(n9117) );
  INV_X1 U10327 ( .A(n8988), .ZN(n8989) );
  AOI22_X1 U10328 ( .A1(n9019), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8989), .B2(
        n9005), .ZN(n8990) );
  OAI21_X1 U10329 ( .B1(n8991), .B2(n9008), .A(n8990), .ZN(n8994) );
  NOR2_X1 U10330 ( .A1(n9120), .A2(n8992), .ZN(n8993) );
  AOI211_X1 U10331 ( .C1(n9117), .C2(n8995), .A(n8994), .B(n8993), .ZN(n8996)
         );
  OAI21_X1 U10332 ( .B1(n9119), .B2(n9019), .A(n8996), .ZN(P2_U3283) );
  NAND2_X1 U10333 ( .A1(n8998), .A2(n8997), .ZN(n9000) );
  AND2_X1 U10334 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  XNOR2_X1 U10335 ( .A(n9001), .B(n8654), .ZN(n9126) );
  AOI21_X1 U10336 ( .B1(n9121), .B2(n9003), .A(n9002), .ZN(n9122) );
  INV_X1 U10337 ( .A(n9121), .ZN(n9009) );
  INV_X1 U10338 ( .A(n9004), .ZN(n9006) );
  AOI22_X1 U10339 ( .A1(n9019), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9006), .B2(
        n9005), .ZN(n9007) );
  OAI21_X1 U10340 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9021) );
  AOI21_X1 U10341 ( .B1(n9011), .B2(n8654), .A(n9010), .ZN(n9018) );
  OAI22_X1 U10342 ( .A1(n9015), .A2(n9014), .B1(n9013), .B2(n9012), .ZN(n9016)
         );
  AOI21_X1 U10343 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9124) );
  NOR2_X1 U10344 ( .A1(n9124), .A2(n9019), .ZN(n9020) );
  AOI211_X1 U10345 ( .C1(n9122), .C2(n9022), .A(n9021), .B(n9020), .ZN(n9023)
         );
  OAI21_X1 U10346 ( .B1(n9024), .B2(n9126), .A(n9023), .ZN(P2_U3284) );
  NAND2_X1 U10347 ( .A1(n9025), .A2(n9992), .ZN(n9026) );
  OAI211_X1 U10348 ( .C1(n9027), .C2(n10020), .A(n9707), .B(n9026), .ZN(n9134)
         );
  MUX2_X1 U10349 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9134), .S(n10039), .Z(
        P2_U3551) );
  NAND2_X1 U10350 ( .A1(n9028), .A2(n10024), .ZN(n9034) );
  AOI22_X1 U10351 ( .A1(n9030), .A2(n9993), .B1(n9992), .B2(n9029), .ZN(n9032)
         );
  NAND2_X1 U10352 ( .A1(n9034), .A2(n9033), .ZN(n9135) );
  MUX2_X1 U10353 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9135), .S(n10039), .Z(
        P2_U3549) );
  INV_X1 U10354 ( .A(n9035), .ZN(n9040) );
  AOI22_X1 U10355 ( .A1(n9037), .A2(n9993), .B1(n9992), .B2(n9036), .ZN(n9038)
         );
  OAI211_X1 U10356 ( .C1(n9040), .C2(n9125), .A(n9039), .B(n9038), .ZN(n9136)
         );
  MUX2_X1 U10357 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9136), .S(n10039), .Z(
        P2_U3548) );
  INV_X1 U10358 ( .A(n9041), .ZN(n9046) );
  AOI22_X1 U10359 ( .A1(n9043), .A2(n9993), .B1(n9992), .B2(n9042), .ZN(n9044)
         );
  OAI211_X1 U10360 ( .C1(n9046), .C2(n9125), .A(n9045), .B(n9044), .ZN(n9137)
         );
  MUX2_X1 U10361 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9137), .S(n10039), .Z(
        P2_U3547) );
  AOI21_X1 U10362 ( .B1(n9992), .B2(n9048), .A(n9047), .ZN(n9049) );
  OAI211_X1 U10363 ( .C1(n9051), .C2(n9125), .A(n9050), .B(n9049), .ZN(n9138)
         );
  MUX2_X1 U10364 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9138), .S(n10039), .Z(
        P2_U3546) );
  AOI21_X1 U10365 ( .B1(n9992), .B2(n9053), .A(n9052), .ZN(n9054) );
  OAI211_X1 U10366 ( .C1(n9056), .C2(n9125), .A(n9055), .B(n9054), .ZN(n9139)
         );
  MUX2_X1 U10367 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9139), .S(n10039), .Z(
        P2_U3545) );
  AOI22_X1 U10368 ( .A1(n9058), .A2(n9993), .B1(n9992), .B2(n9057), .ZN(n9059)
         );
  OAI211_X1 U10369 ( .C1(n9061), .C2(n9125), .A(n9060), .B(n9059), .ZN(n9140)
         );
  MUX2_X1 U10370 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9140), .S(n10039), .Z(
        P2_U3544) );
  AOI22_X1 U10371 ( .A1(n9063), .A2(n9993), .B1(n9992), .B2(n9062), .ZN(n9064)
         );
  OAI211_X1 U10372 ( .C1(n9066), .C2(n9125), .A(n9065), .B(n9064), .ZN(n9141)
         );
  MUX2_X1 U10373 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9141), .S(n10039), .Z(
        P2_U3543) );
  AOI22_X1 U10374 ( .A1(n9068), .A2(n9993), .B1(n9992), .B2(n9067), .ZN(n9069)
         );
  OAI211_X1 U10375 ( .C1(n9071), .C2(n9125), .A(n9070), .B(n9069), .ZN(n9142)
         );
  MUX2_X1 U10376 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9142), .S(n10039), .Z(
        P2_U3542) );
  AOI22_X1 U10377 ( .A1(n9073), .A2(n9993), .B1(n9992), .B2(n9072), .ZN(n9074)
         );
  OAI211_X1 U10378 ( .C1(n9076), .C2(n9125), .A(n9075), .B(n9074), .ZN(n9143)
         );
  MUX2_X1 U10379 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9143), .S(n10039), .Z(
        P2_U3541) );
  AOI22_X1 U10380 ( .A1(n9078), .A2(n9993), .B1(n9992), .B2(n9077), .ZN(n9079)
         );
  OAI211_X1 U10381 ( .C1(n9081), .C2(n9125), .A(n9080), .B(n9079), .ZN(n9144)
         );
  MUX2_X1 U10382 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9144), .S(n10039), .Z(
        P2_U3540) );
  AOI21_X1 U10383 ( .B1(n9992), .B2(n9083), .A(n9082), .ZN(n9084) );
  OAI211_X1 U10384 ( .C1(n9086), .C2(n9125), .A(n9085), .B(n9084), .ZN(n9145)
         );
  MUX2_X1 U10385 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9145), .S(n10039), .Z(
        P2_U3539) );
  AOI22_X1 U10386 ( .A1(n9088), .A2(n9993), .B1(n9992), .B2(n9087), .ZN(n9089)
         );
  OAI211_X1 U10387 ( .C1(n9091), .C2(n9125), .A(n9090), .B(n9089), .ZN(n9146)
         );
  MUX2_X1 U10388 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9146), .S(n10039), .Z(
        P2_U3538) );
  AOI21_X1 U10389 ( .B1(n9992), .B2(n9093), .A(n9092), .ZN(n9094) );
  OAI211_X1 U10390 ( .C1(n9096), .C2(n10009), .A(n9095), .B(n9094), .ZN(n9147)
         );
  MUX2_X1 U10391 ( .A(n9147), .B(P2_REG1_REG_17__SCAN_IN), .S(n10037), .Z(
        P2_U3537) );
  AOI22_X1 U10392 ( .A1(n9098), .A2(n9993), .B1(n9992), .B2(n9097), .ZN(n9099)
         );
  OAI21_X1 U10393 ( .B1(n9100), .B2(n10009), .A(n9099), .ZN(n9101) );
  NOR2_X1 U10394 ( .A1(n9102), .A2(n9101), .ZN(n9149) );
  MUX2_X1 U10395 ( .A(n9149), .B(n9103), .S(n10037), .Z(n9104) );
  INV_X1 U10396 ( .A(n9104), .ZN(P2_U3536) );
  INV_X1 U10397 ( .A(n9105), .ZN(n9110) );
  AOI22_X1 U10398 ( .A1(n9107), .A2(n9993), .B1(n9992), .B2(n9106), .ZN(n9108)
         );
  OAI211_X1 U10399 ( .C1(n9110), .C2(n9125), .A(n9109), .B(n9108), .ZN(n9151)
         );
  MUX2_X1 U10400 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9151), .S(n10039), .Z(
        P2_U3535) );
  AOI22_X1 U10401 ( .A1(n9112), .A2(n9993), .B1(n9992), .B2(n9111), .ZN(n9113)
         );
  OAI211_X1 U10402 ( .C1(n9115), .C2(n9125), .A(n9114), .B(n9113), .ZN(n9152)
         );
  MUX2_X1 U10403 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9152), .S(n10039), .Z(
        P2_U3534) );
  AOI22_X1 U10404 ( .A1(n9117), .A2(n9993), .B1(n9992), .B2(n9116), .ZN(n9118)
         );
  OAI211_X1 U10405 ( .C1(n10009), .C2(n9120), .A(n9119), .B(n9118), .ZN(n9153)
         );
  MUX2_X1 U10406 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9153), .S(n10039), .Z(
        P2_U3533) );
  AOI22_X1 U10407 ( .A1(n9122), .A2(n9993), .B1(n9992), .B2(n9121), .ZN(n9123)
         );
  OAI211_X1 U10408 ( .C1(n9126), .C2(n9125), .A(n9124), .B(n9123), .ZN(n9154)
         );
  MUX2_X1 U10409 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9154), .S(n10039), .Z(
        P2_U3532) );
  AOI22_X1 U10410 ( .A1(n9128), .A2(n9993), .B1(n9992), .B2(n9127), .ZN(n9129)
         );
  OAI21_X1 U10411 ( .B1(n9130), .B2(n10009), .A(n9129), .ZN(n9131) );
  NOR2_X1 U10412 ( .A1(n9132), .A2(n9131), .ZN(n9155) );
  MUX2_X1 U10413 ( .A(n6687), .B(n9155), .S(n10039), .Z(n9133) );
  INV_X1 U10414 ( .A(n9133), .ZN(P2_U3530) );
  MUX2_X1 U10415 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9134), .S(n10017), .Z(
        P2_U3519) );
  MUX2_X1 U10416 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9135), .S(n10017), .Z(
        P2_U3517) );
  MUX2_X1 U10417 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9136), .S(n10017), .Z(
        P2_U3516) );
  MUX2_X1 U10418 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9137), .S(n10017), .Z(
        P2_U3515) );
  MUX2_X1 U10419 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9138), .S(n10017), .Z(
        P2_U3514) );
  MUX2_X1 U10420 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9139), .S(n10017), .Z(
        P2_U3513) );
  MUX2_X1 U10421 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9140), .S(n10017), .Z(
        P2_U3512) );
  MUX2_X1 U10422 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9141), .S(n10017), .Z(
        P2_U3511) );
  MUX2_X1 U10423 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9142), .S(n10017), .Z(
        P2_U3510) );
  MUX2_X1 U10424 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9143), .S(n10017), .Z(
        P2_U3509) );
  MUX2_X1 U10425 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9144), .S(n10017), .Z(
        P2_U3508) );
  MUX2_X1 U10426 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9145), .S(n10017), .Z(
        P2_U3507) );
  MUX2_X1 U10427 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9146), .S(n10017), .Z(
        P2_U3505) );
  MUX2_X1 U10428 ( .A(n9147), .B(P2_REG0_REG_17__SCAN_IN), .S(n10026), .Z(
        P2_U3502) );
  MUX2_X1 U10429 ( .A(n9149), .B(n9148), .S(n10026), .Z(n9150) );
  INV_X1 U10430 ( .A(n9150), .ZN(P2_U3499) );
  MUX2_X1 U10431 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9151), .S(n10017), .Z(
        P2_U3496) );
  MUX2_X1 U10432 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9152), .S(n10017), .Z(
        P2_U3493) );
  MUX2_X1 U10433 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9153), .S(n10017), .Z(
        P2_U3490) );
  MUX2_X1 U10434 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9154), .S(n10017), .Z(
        P2_U3487) );
  MUX2_X1 U10435 ( .A(n5647), .B(n9155), .S(n10017), .Z(n9156) );
  INV_X1 U10436 ( .A(n9156), .ZN(P2_U3481) );
  INV_X1 U10437 ( .A(n9157), .ZN(n9666) );
  NOR4_X1 U10438 ( .A1(n9158), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5468), .A4(
        P2_U3152), .ZN(n9159) );
  AOI21_X1 U10439 ( .B1(n9162), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9159), .ZN(
        n9160) );
  OAI21_X1 U10440 ( .B1(n9666), .B2(n9165), .A(n9160), .ZN(P2_U3327) );
  INV_X1 U10441 ( .A(n9161), .ZN(n9670) );
  AOI22_X1 U10442 ( .A1(n9163), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9162), .ZN(n9164) );
  OAI21_X1 U10443 ( .B1(n9670), .B2(n9165), .A(n9164), .ZN(P2_U3328) );
  MUX2_X1 U10444 ( .A(n9166), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10445 ( .A1(n4341), .A2(n9167), .ZN(n9169) );
  XNOR2_X1 U10446 ( .A(n9169), .B(n9168), .ZN(n9174) );
  INV_X1 U10447 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9170) );
  OAI22_X1 U10448 ( .A1(n9682), .A2(n9198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9170), .ZN(n9172) );
  OAI22_X1 U10449 ( .A1(n9699), .A2(n9395), .B1(n9188), .B2(n9271), .ZN(n9171)
         );
  AOI211_X1 U10450 ( .C1(n9591), .C2(n9276), .A(n9172), .B(n9171), .ZN(n9173)
         );
  OAI21_X1 U10451 ( .B1(n9174), .B2(n9278), .A(n9173), .ZN(P1_U3214) );
  OAI21_X1 U10452 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9178) );
  NAND2_X1 U10453 ( .A1(n9178), .A2(n9694), .ZN(n9184) );
  NOR2_X1 U10454 ( .A1(n9179), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9306) );
  INV_X1 U10455 ( .A(n9465), .ZN(n9181) );
  OAI22_X1 U10456 ( .A1(n9699), .A2(n9181), .B1(n9271), .B2(n9180), .ZN(n9182)
         );
  AOI211_X1 U10457 ( .C1(n9222), .C2(n9470), .A(n9306), .B(n9182), .ZN(n9183)
         );
  OAI211_X1 U10458 ( .C1(n9467), .C2(n9224), .A(n9184), .B(n9183), .ZN(
        P1_U3217) );
  XOR2_X1 U10459 ( .A(n9186), .B(n9185), .Z(n9193) );
  OAI22_X1 U10460 ( .A1(n9188), .A2(n9682), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9187), .ZN(n9191) );
  OAI22_X1 U10461 ( .A1(n9699), .A2(n9437), .B1(n9271), .B2(n9189), .ZN(n9190)
         );
  AOI211_X1 U10462 ( .C1(n9601), .C2(n9276), .A(n9191), .B(n9190), .ZN(n9192)
         );
  OAI21_X1 U10463 ( .B1(n9193), .B2(n9278), .A(n9192), .ZN(P1_U3221) );
  XOR2_X1 U10464 ( .A(n9195), .B(n9194), .Z(n9203) );
  OAI22_X1 U10465 ( .A1(n9682), .A2(n9348), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9196), .ZN(n9201) );
  INV_X1 U10466 ( .A(n9197), .ZN(n9199) );
  OAI22_X1 U10467 ( .A1(n9699), .A2(n9199), .B1(n9271), .B2(n9198), .ZN(n9200)
         );
  AOI211_X1 U10468 ( .C1(n5293), .C2(n9276), .A(n9201), .B(n9200), .ZN(n9202)
         );
  OAI21_X1 U10469 ( .B1(n9203), .B2(n9278), .A(n9202), .ZN(P1_U3223) );
  INV_X1 U10470 ( .A(n9623), .ZN(n9496) );
  OAI21_X1 U10471 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9207) );
  NAND2_X1 U10472 ( .A1(n9207), .A2(n9694), .ZN(n9210) );
  AND2_X1 U10473 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9810) );
  OAI22_X1 U10474 ( .A1(n9699), .A2(n9493), .B1(n9271), .B2(n9530), .ZN(n9208)
         );
  AOI211_X1 U10475 ( .C1(n9222), .C2(n9500), .A(n9810), .B(n9208), .ZN(n9209)
         );
  OAI211_X1 U10476 ( .C1(n9496), .C2(n9224), .A(n9210), .B(n9209), .ZN(
        P1_U3226) );
  AOI21_X1 U10477 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9218) );
  INV_X1 U10478 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9214) );
  OAI22_X1 U10479 ( .A1(n9682), .A2(n9381), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9214), .ZN(n9216) );
  OAI22_X1 U10480 ( .A1(n9380), .A2(n9271), .B1(n9699), .B2(n9384), .ZN(n9215)
         );
  AOI211_X1 U10481 ( .C1(n9588), .C2(n9276), .A(n9216), .B(n9215), .ZN(n9217)
         );
  OAI21_X1 U10482 ( .B1(n9218), .B2(n9278), .A(n9217), .ZN(P1_U3227) );
  OAI211_X1 U10483 ( .C1(n9219), .C2(n9221), .A(n9220), .B(n9694), .ZN(n9228)
         );
  AOI22_X1 U10484 ( .A1(n9259), .A2(n9223), .B1(n9222), .B2(n9289), .ZN(n9227)
         );
  AND2_X1 U10485 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9774) );
  AOI211_X1 U10486 ( .C1(n9685), .C2(n9290), .A(n9774), .B(n9225), .ZN(n9226)
         );
  NAND3_X1 U10487 ( .A1(n9228), .A2(n9227), .A3(n9226), .ZN(P1_U3228) );
  INV_X1 U10488 ( .A(n9229), .ZN(n9234) );
  AOI21_X1 U10489 ( .B1(n9231), .B2(n9233), .A(n9230), .ZN(n9232) );
  AOI21_X1 U10490 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9240) );
  OAI22_X1 U10491 ( .A1(n9682), .A2(n9248), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9235), .ZN(n9238) );
  INV_X1 U10492 ( .A(n9450), .ZN(n9236) );
  OAI22_X1 U10493 ( .A1(n9699), .A2(n9236), .B1(n9271), .B2(n9262), .ZN(n9237)
         );
  AOI211_X1 U10494 ( .C1(n9606), .C2(n9276), .A(n9238), .B(n9237), .ZN(n9239)
         );
  OAI21_X1 U10495 ( .B1(n9240), .B2(n9278), .A(n9239), .ZN(P1_U3231) );
  INV_X1 U10496 ( .A(n9241), .ZN(n9245) );
  OR2_X1 U10497 ( .A1(n9242), .A2(n9241), .ZN(n9243) );
  AOI22_X1 U10498 ( .A1(n9246), .A2(n9245), .B1(n9244), .B2(n9243), .ZN(n9252)
         );
  INV_X1 U10499 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9247) );
  OAI22_X1 U10500 ( .A1(n9380), .A2(n9682), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9247), .ZN(n9250) );
  OAI22_X1 U10501 ( .A1(n9699), .A2(n9415), .B1(n9271), .B2(n9248), .ZN(n9249)
         );
  AOI211_X1 U10502 ( .C1(n9597), .C2(n9276), .A(n9250), .B(n9249), .ZN(n9251)
         );
  OAI21_X1 U10503 ( .B1(n9252), .B2(n9278), .A(n9251), .ZN(P1_U3233) );
  INV_X1 U10504 ( .A(n9253), .ZN(n9258) );
  AOI21_X1 U10505 ( .B1(n9254), .B2(n9257), .A(n9255), .ZN(n9256) );
  AOI21_X1 U10506 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9265) );
  AOI22_X1 U10507 ( .A1(n9259), .A2(n9482), .B1(n9685), .B2(n9478), .ZN(n9261)
         );
  OAI211_X1 U10508 ( .C1(n9262), .C2(n9682), .A(n9261), .B(n9260), .ZN(n9263)
         );
  AOI21_X1 U10509 ( .B1(n9618), .B2(n9276), .A(n9263), .ZN(n9264) );
  OAI21_X1 U10510 ( .B1(n9265), .B2(n9278), .A(n9264), .ZN(P1_U3236) );
  NAND2_X1 U10511 ( .A1(n4662), .A2(n9268), .ZN(n9269) );
  XNOR2_X1 U10512 ( .A(n9266), .B(n9269), .ZN(n9279) );
  OAI22_X1 U10513 ( .A1(n9271), .A2(n9381), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9270), .ZN(n9275) );
  INV_X1 U10514 ( .A(n9358), .ZN(n9273) );
  OAI22_X1 U10515 ( .A1(n9699), .A2(n9273), .B1(n9682), .B2(n9272), .ZN(n9274)
         );
  AOI211_X1 U10516 ( .C1(n9577), .C2(n9276), .A(n9275), .B(n9274), .ZN(n9277)
         );
  OAI21_X1 U10517 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(P1_U3238) );
  MUX2_X1 U10518 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9280), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10519 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9325), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9281), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10521 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9366), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10522 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9282), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10523 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9367), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9403), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9421), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9435), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9455), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9470), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10529 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9479), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9500), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9478), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9499), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10533 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9548), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9283), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9549), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9284), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9684), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9285), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9286), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9288), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9846), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9289), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9845), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9290), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9874), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9291), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6292), .S(P1_U4006), .Z(
        P1_U3555) );
  AOI21_X1 U10549 ( .B1(n9293), .B2(n9296), .A(n9292), .ZN(n9294) );
  XOR2_X1 U10550 ( .A(n9294), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9303) );
  INV_X1 U10551 ( .A(n9303), .ZN(n9301) );
  INV_X1 U10552 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9297) );
  OAI21_X1 U10553 ( .B1(n9297), .B2(n9296), .A(n9295), .ZN(n9298) );
  XOR2_X1 U10554 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9298), .Z(n9302) );
  OAI21_X1 U10555 ( .B1(n9302), .B2(n9299), .A(n9808), .ZN(n9300) );
  AOI21_X1 U10556 ( .B1(n9301), .B2(n9813), .A(n9300), .ZN(n9305) );
  AOI22_X1 U10557 ( .A1(n9303), .A2(n9813), .B1(n9817), .B2(n9302), .ZN(n9304)
         );
  MUX2_X1 U10558 ( .A(n9305), .B(n9304), .S(n9850), .Z(n9308) );
  AOI21_X1 U10559 ( .B1(n9811), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9306), .ZN(
        n9307) );
  NAND2_X1 U10560 ( .A1(n9308), .A2(n9307), .ZN(P1_U3260) );
  NAND2_X1 U10561 ( .A1(n9703), .A2(n9504), .ZN(n9312) );
  NAND2_X1 U10562 ( .A1(n9310), .A2(n9309), .ZN(n9700) );
  NOR2_X1 U10563 ( .A1(n9856), .A2(n9700), .ZN(n9316) );
  AOI21_X1 U10564 ( .B1(n9856), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9316), .ZN(
        n9311) );
  OAI211_X1 U10565 ( .C1(n9701), .C2(n9539), .A(n9312), .B(n9311), .ZN(
        P1_U3261) );
  INV_X1 U10566 ( .A(n9313), .ZN(n9315) );
  NAND2_X1 U10567 ( .A1(n9315), .A2(n9314), .ZN(n9564) );
  NAND3_X1 U10568 ( .A1(n9564), .A2(n9504), .A3(n9563), .ZN(n9318) );
  AOI21_X1 U10569 ( .B1(n9856), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9316), .ZN(
        n9317) );
  OAI211_X1 U10570 ( .C1(n9566), .C2(n9539), .A(n9318), .B(n9317), .ZN(
        P1_U3262) );
  AND2_X1 U10571 ( .A1(n9319), .A2(n9323), .ZN(n9321) );
  OAI211_X1 U10572 ( .C1(n9324), .C2(n9323), .A(n9322), .B(n9871), .ZN(n9327)
         );
  AOI22_X1 U10573 ( .A1(n9875), .A2(n9366), .B1(n9325), .B2(n9873), .ZN(n9326)
         );
  NAND2_X1 U10574 ( .A1(n9327), .A2(n9326), .ZN(n9569) );
  NAND2_X1 U10575 ( .A1(n9339), .A2(n9330), .ZN(n9328) );
  NAND2_X1 U10576 ( .A1(n9329), .A2(n9328), .ZN(n9567) );
  NOR2_X1 U10577 ( .A1(n9567), .A2(n9440), .ZN(n9335) );
  INV_X1 U10578 ( .A(n9331), .ZN(n9332) );
  AOI22_X1 U10579 ( .A1(n9856), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9332), .B2(
        n9826), .ZN(n9333) );
  OAI21_X1 U10580 ( .B1(n4516), .B2(n9539), .A(n9333), .ZN(n9334) );
  AOI211_X1 U10581 ( .C1(n9569), .C2(n9884), .A(n9335), .B(n9334), .ZN(n9336)
         );
  OAI21_X1 U10582 ( .B1(n9571), .B2(n9855), .A(n9336), .ZN(P1_U3263) );
  XNOR2_X1 U10583 ( .A(n9337), .B(n9345), .ZN(n9576) );
  INV_X1 U10584 ( .A(n9338), .ZN(n9341) );
  INV_X1 U10585 ( .A(n9339), .ZN(n9340) );
  AOI21_X1 U10586 ( .B1(n9572), .B2(n9341), .A(n9340), .ZN(n9573) );
  AOI22_X1 U10587 ( .A1(n9856), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9342), .B2(
        n9826), .ZN(n9343) );
  OAI21_X1 U10588 ( .B1(n9344), .B2(n9539), .A(n9343), .ZN(n9353) );
  AOI21_X1 U10589 ( .B1(n9346), .B2(n9345), .A(n9527), .ZN(n9351) );
  OAI22_X1 U10590 ( .A1(n9348), .A2(n9529), .B1(n9347), .B2(n9531), .ZN(n9349)
         );
  AOI21_X1 U10591 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9575) );
  NOR2_X1 U10592 ( .A1(n9575), .A2(n9856), .ZN(n9352) );
  AOI211_X1 U10593 ( .C1(n9573), .C2(n9504), .A(n9353), .B(n9352), .ZN(n9354)
         );
  OAI21_X1 U10594 ( .B1(n9576), .B2(n9855), .A(n9354), .ZN(P1_U3264) );
  XOR2_X1 U10595 ( .A(n9365), .B(n9355), .Z(n9581) );
  INV_X1 U10596 ( .A(n9356), .ZN(n9357) );
  AOI21_X1 U10597 ( .B1(n9577), .B2(n9357), .A(n9338), .ZN(n9578) );
  AOI22_X1 U10598 ( .A1(n9856), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9358), .B2(
        n9826), .ZN(n9359) );
  OAI21_X1 U10599 ( .B1(n9360), .B2(n9539), .A(n9359), .ZN(n9373) );
  NAND2_X1 U10600 ( .A1(n9376), .A2(n9361), .ZN(n9363) );
  NAND2_X1 U10601 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  XOR2_X1 U10602 ( .A(n9365), .B(n9364), .Z(n9371) );
  NAND2_X1 U10603 ( .A1(n9367), .A2(n9875), .ZN(n9368) );
  AOI211_X1 U10604 ( .C1(n9504), .C2(n9578), .A(n9373), .B(n9372), .ZN(n9374)
         );
  OAI21_X1 U10605 ( .B1(n9581), .B2(n9855), .A(n9374), .ZN(P1_U3265) );
  XNOR2_X1 U10606 ( .A(n9375), .B(n9378), .ZN(n9590) );
  AOI22_X1 U10607 ( .A1(n9588), .A2(n9555), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9856), .ZN(n9388) );
  AOI21_X1 U10608 ( .B1(n9378), .B2(n9377), .A(n5371), .ZN(n9379) );
  OAI222_X1 U10609 ( .A1(n9531), .A2(n9381), .B1(n9529), .B2(n9380), .C1(n9527), .C2(n9379), .ZN(n9586) );
  INV_X1 U10610 ( .A(n9382), .ZN(n9383) );
  AOI211_X1 U10611 ( .C1(n9588), .C2(n9393), .A(n9946), .B(n9383), .ZN(n9587)
         );
  INV_X1 U10612 ( .A(n9587), .ZN(n9385) );
  OAI22_X1 U10613 ( .A1(n9385), .A2(n9867), .B1(n9880), .B2(n9384), .ZN(n9386)
         );
  OAI21_X1 U10614 ( .B1(n9586), .B2(n9386), .A(n9884), .ZN(n9387) );
  OAI211_X1 U10615 ( .C1(n9590), .C2(n9855), .A(n9388), .B(n9387), .ZN(
        P1_U3267) );
  OR2_X1 U10616 ( .A1(n9487), .A2(n9389), .ZN(n9391) );
  AND2_X1 U10617 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  XNOR2_X1 U10618 ( .A(n9392), .B(n9401), .ZN(n9595) );
  INV_X1 U10619 ( .A(n9393), .ZN(n9394) );
  AOI21_X1 U10620 ( .B1(n9591), .B2(n9412), .A(n9394), .ZN(n9592) );
  INV_X1 U10621 ( .A(n9591), .ZN(n9398) );
  INV_X1 U10622 ( .A(n9395), .ZN(n9396) );
  AOI22_X1 U10623 ( .A1(n9856), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9396), .B2(
        n9826), .ZN(n9397) );
  OAI21_X1 U10624 ( .B1(n9398), .B2(n9539), .A(n9397), .ZN(n9406) );
  NAND2_X1 U10625 ( .A1(n9399), .A2(n9400), .ZN(n9402) );
  XNOR2_X1 U10626 ( .A(n9402), .B(n9401), .ZN(n9404) );
  AOI222_X1 U10627 ( .A1(n9871), .A2(n9404), .B1(n9403), .B2(n9873), .C1(n9435), .C2(n9875), .ZN(n9594) );
  NOR2_X1 U10628 ( .A1(n9594), .A2(n9856), .ZN(n9405) );
  AOI211_X1 U10629 ( .C1(n9592), .C2(n9504), .A(n9406), .B(n9405), .ZN(n9407)
         );
  OAI21_X1 U10630 ( .B1(n9595), .B2(n9855), .A(n9407), .ZN(P1_U3268) );
  OR2_X1 U10631 ( .A1(n9487), .A2(n9408), .ZN(n9410) );
  NAND2_X1 U10632 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  XOR2_X1 U10633 ( .A(n9420), .B(n9411), .Z(n9600) );
  INV_X1 U10634 ( .A(n9438), .ZN(n9414) );
  INV_X1 U10635 ( .A(n9412), .ZN(n9413) );
  AOI211_X1 U10636 ( .C1(n9597), .C2(n9414), .A(n9946), .B(n9413), .ZN(n9596)
         );
  INV_X1 U10637 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10638 ( .A1(n9856), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9416), .B2(
        n9826), .ZN(n9417) );
  OAI21_X1 U10639 ( .B1(n9418), .B2(n9539), .A(n9417), .ZN(n9424) );
  OAI21_X1 U10640 ( .B1(n9420), .B2(n9419), .A(n9399), .ZN(n9422) );
  AOI222_X1 U10641 ( .A1(n9871), .A2(n9422), .B1(n9455), .B2(n9875), .C1(n9421), .C2(n9873), .ZN(n9599) );
  NOR2_X1 U10642 ( .A1(n9599), .A2(n9856), .ZN(n9423) );
  AOI211_X1 U10643 ( .C1(n9596), .C2(n9535), .A(n9424), .B(n9423), .ZN(n9425)
         );
  OAI21_X1 U10644 ( .B1(n9855), .B2(n9600), .A(n9425), .ZN(P1_U3269) );
  OR2_X1 U10645 ( .A1(n9487), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U10646 ( .A1(n9428), .A2(n9427), .ZN(n9429) );
  XNOR2_X1 U10647 ( .A(n9429), .B(n9430), .ZN(n9605) );
  NAND3_X1 U10648 ( .A1(n9432), .A2(n9431), .A3(n9430), .ZN(n9433) );
  NAND2_X1 U10649 ( .A1(n9434), .A2(n9433), .ZN(n9436) );
  AOI222_X1 U10650 ( .A1(n9871), .A2(n9436), .B1(n9435), .B2(n9873), .C1(n9470), .C2(n9875), .ZN(n9604) );
  OAI21_X1 U10651 ( .B1(n9437), .B2(n9880), .A(n9604), .ZN(n9443) );
  AOI21_X1 U10652 ( .B1(n9601), .B2(n9449), .A(n9438), .ZN(n9602) );
  INV_X1 U10653 ( .A(n9602), .ZN(n9441) );
  AOI22_X1 U10654 ( .A1(n9601), .A2(n9555), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9856), .ZN(n9439) );
  OAI21_X1 U10655 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9442) );
  AOI21_X1 U10656 ( .B1(n9443), .B2(n9884), .A(n9442), .ZN(n9444) );
  OAI21_X1 U10657 ( .B1(n9605), .B2(n9855), .A(n9444), .ZN(P1_U3270) );
  OR2_X1 U10658 ( .A1(n9487), .A2(n9445), .ZN(n9447) );
  NAND2_X1 U10659 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  XNOR2_X1 U10660 ( .A(n9448), .B(n9454), .ZN(n9610) );
  AOI21_X1 U10661 ( .B1(n9606), .B2(n9463), .A(n4521), .ZN(n9607) );
  INV_X1 U10662 ( .A(n9606), .ZN(n9452) );
  AOI22_X1 U10663 ( .A1(n9856), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9450), .B2(
        n9826), .ZN(n9451) );
  OAI21_X1 U10664 ( .B1(n9452), .B2(n9539), .A(n9451), .ZN(n9458) );
  XOR2_X1 U10665 ( .A(n9454), .B(n9453), .Z(n9456) );
  AOI222_X1 U10666 ( .A1(n9871), .A2(n9456), .B1(n9455), .B2(n9873), .C1(n9479), .C2(n9875), .ZN(n9609) );
  NOR2_X1 U10667 ( .A1(n9609), .A2(n9856), .ZN(n9457) );
  AOI211_X1 U10668 ( .C1(n9607), .C2(n9504), .A(n9458), .B(n9457), .ZN(n9459)
         );
  OAI21_X1 U10669 ( .B1(n9855), .B2(n9610), .A(n9459), .ZN(P1_U3271) );
  OR2_X1 U10670 ( .A1(n9487), .A2(n9486), .ZN(n9617) );
  NAND2_X1 U10671 ( .A1(n9617), .A2(n9460), .ZN(n9461) );
  XOR2_X1 U10672 ( .A(n9469), .B(n9461), .Z(n9615) );
  INV_X1 U10673 ( .A(n9462), .ZN(n9464) );
  AOI21_X1 U10674 ( .B1(n9611), .B2(n9464), .A(n4517), .ZN(n9612) );
  AOI22_X1 U10675 ( .A1(n9856), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9465), .B2(
        n9826), .ZN(n9466) );
  OAI21_X1 U10676 ( .B1(n9467), .B2(n9539), .A(n9466), .ZN(n9473) );
  XNOR2_X1 U10677 ( .A(n9468), .B(n9469), .ZN(n9471) );
  AOI222_X1 U10678 ( .A1(n9871), .A2(n9471), .B1(n9470), .B2(n9873), .C1(n9500), .C2(n9875), .ZN(n9614) );
  NOR2_X1 U10679 ( .A1(n9614), .A2(n9856), .ZN(n9472) );
  AOI211_X1 U10680 ( .C1(n9612), .C2(n9504), .A(n9473), .B(n9472), .ZN(n9474)
         );
  OAI21_X1 U10681 ( .B1(n9855), .B2(n9615), .A(n9474), .ZN(P1_U3272) );
  NAND2_X1 U10682 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  XOR2_X1 U10683 ( .A(n9486), .B(n9477), .Z(n9480) );
  AOI222_X1 U10684 ( .A1(n9871), .A2(n9480), .B1(n9479), .B2(n9873), .C1(n9478), .C2(n9875), .ZN(n9621) );
  INV_X1 U10685 ( .A(n9492), .ZN(n9481) );
  AOI21_X1 U10686 ( .B1(n9618), .B2(n9481), .A(n9462), .ZN(n9619) );
  AOI22_X1 U10687 ( .A1(n9856), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9482), .B2(
        n9826), .ZN(n9483) );
  OAI21_X1 U10688 ( .B1(n9484), .B2(n9539), .A(n9483), .ZN(n9485) );
  AOI21_X1 U10689 ( .B1(n9619), .B2(n9504), .A(n9485), .ZN(n9490) );
  NAND2_X1 U10690 ( .A1(n9487), .A2(n9486), .ZN(n9616) );
  NAND3_X1 U10691 ( .A1(n9617), .A2(n9616), .A3(n9488), .ZN(n9489) );
  OAI211_X1 U10692 ( .C1(n9621), .C2(n9856), .A(n9490), .B(n9489), .ZN(
        P1_U3273) );
  XOR2_X1 U10693 ( .A(n9498), .B(n9491), .Z(n9627) );
  AOI21_X1 U10694 ( .B1(n9623), .B2(n9507), .A(n9492), .ZN(n9624) );
  INV_X1 U10695 ( .A(n9493), .ZN(n9494) );
  AOI22_X1 U10696 ( .A1(n9856), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9494), .B2(
        n9826), .ZN(n9495) );
  OAI21_X1 U10697 ( .B1(n9496), .B2(n9539), .A(n9495), .ZN(n9503) );
  XOR2_X1 U10698 ( .A(n9497), .B(n9498), .Z(n9501) );
  AOI222_X1 U10699 ( .A1(n9871), .A2(n9501), .B1(n9500), .B2(n9873), .C1(n9499), .C2(n9875), .ZN(n9626) );
  NOR2_X1 U10700 ( .A1(n9626), .A2(n9856), .ZN(n9502) );
  AOI211_X1 U10701 ( .C1(n9624), .C2(n9504), .A(n9503), .B(n9502), .ZN(n9505)
         );
  OAI21_X1 U10702 ( .B1(n9855), .B2(n9627), .A(n9505), .ZN(P1_U3274) );
  XNOR2_X1 U10703 ( .A(n9506), .B(n9514), .ZN(n9632) );
  INV_X1 U10704 ( .A(n9507), .ZN(n9508) );
  AOI211_X1 U10705 ( .C1(n9630), .C2(n9533), .A(n9946), .B(n9508), .ZN(n9629)
         );
  INV_X1 U10706 ( .A(n9630), .ZN(n9509) );
  NOR2_X1 U10707 ( .A1(n9509), .A2(n9539), .ZN(n9512) );
  OAI22_X1 U10708 ( .A1(n9884), .A2(n7046), .B1(n9510), .B2(n9880), .ZN(n9511)
         );
  AOI211_X1 U10709 ( .C1(n9629), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9520)
         );
  XNOR2_X1 U10710 ( .A(n9515), .B(n9514), .ZN(n9516) );
  OAI222_X1 U10711 ( .A1(n9531), .A2(n9518), .B1(n9529), .B2(n9517), .C1(n9516), .C2(n9527), .ZN(n9628) );
  NAND2_X1 U10712 ( .A1(n9628), .A2(n9884), .ZN(n9519) );
  OAI211_X1 U10713 ( .C1(n9632), .C2(n9855), .A(n9520), .B(n9519), .ZN(
        P1_U3275) );
  XOR2_X1 U10714 ( .A(n9521), .B(n9525), .Z(n9637) );
  INV_X1 U10715 ( .A(n9522), .ZN(n9523) );
  AOI21_X1 U10716 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9526) );
  OAI222_X1 U10717 ( .A1(n9531), .A2(n9530), .B1(n9529), .B2(n9528), .C1(n9527), .C2(n9526), .ZN(n9633) );
  INV_X1 U10718 ( .A(n9532), .ZN(n9552) );
  INV_X1 U10719 ( .A(n9533), .ZN(n9534) );
  AOI211_X1 U10720 ( .C1(n9635), .C2(n9552), .A(n9946), .B(n9534), .ZN(n9634)
         );
  NAND2_X1 U10721 ( .A1(n9634), .A2(n9535), .ZN(n9538) );
  AOI22_X1 U10722 ( .A1(n9856), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9536), .B2(
        n9826), .ZN(n9537) );
  OAI211_X1 U10723 ( .C1(n9540), .C2(n9539), .A(n9538), .B(n9537), .ZN(n9541)
         );
  AOI21_X1 U10724 ( .B1(n9633), .B2(n9884), .A(n9541), .ZN(n9542) );
  OAI21_X1 U10725 ( .B1(n9637), .B2(n9855), .A(n9542), .ZN(P1_U3276) );
  XOR2_X1 U10726 ( .A(n9543), .B(n9544), .Z(n9717) );
  INV_X1 U10727 ( .A(n9717), .ZN(n9562) );
  INV_X1 U10728 ( .A(n9544), .ZN(n9545) );
  XNOR2_X1 U10729 ( .A(n9546), .B(n9545), .ZN(n9547) );
  NAND2_X1 U10730 ( .A1(n9547), .A2(n9871), .ZN(n9551) );
  AOI22_X1 U10731 ( .A1(n9875), .A2(n9549), .B1(n9548), .B2(n9873), .ZN(n9550)
         );
  NAND2_X1 U10732 ( .A1(n9551), .A2(n9550), .ZN(n9716) );
  OAI211_X1 U10733 ( .C1(n9714), .C2(n9553), .A(n9552), .B(n9914), .ZN(n9713)
         );
  AOI22_X1 U10734 ( .A1(n9856), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9554), .B2(
        n9826), .ZN(n9558) );
  NAND2_X1 U10735 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  OAI211_X1 U10736 ( .C1(n9713), .C2(n9559), .A(n9558), .B(n9557), .ZN(n9560)
         );
  AOI21_X1 U10737 ( .B1(n9716), .B2(n9884), .A(n9560), .ZN(n9561) );
  OAI21_X1 U10738 ( .B1(n9562), .B2(n9855), .A(n9561), .ZN(P1_U3277) );
  NAND3_X1 U10739 ( .A1(n9564), .A2(n9914), .A3(n9563), .ZN(n9565) );
  OAI211_X1 U10740 ( .C1(n9566), .C2(n9898), .A(n9565), .B(n9700), .ZN(n9644)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9644), .S(n9968), .Z(
        P1_U3553) );
  OAI22_X1 U10742 ( .A1(n9567), .A2(n9946), .B1(n4516), .B2(n9898), .ZN(n9568)
         );
  NOR2_X1 U10743 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  OAI21_X1 U10744 ( .B1(n9571), .B2(n9922), .A(n9570), .ZN(n9645) );
  MUX2_X1 U10745 ( .A(n9645), .B(P1_REG1_REG_28__SCAN_IN), .S(n9965), .Z(
        P1_U3551) );
  AOI22_X1 U10746 ( .A1(n9573), .A2(n9914), .B1(n9913), .B2(n9572), .ZN(n9574)
         );
  OAI211_X1 U10747 ( .C1(n9576), .C2(n9922), .A(n9575), .B(n9574), .ZN(n9646)
         );
  MUX2_X1 U10748 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9646), .S(n9968), .Z(
        P1_U3550) );
  AOI22_X1 U10749 ( .A1(n9578), .A2(n9914), .B1(n9913), .B2(n9577), .ZN(n9579)
         );
  OAI211_X1 U10750 ( .C1(n9581), .C2(n9922), .A(n9580), .B(n9579), .ZN(n9647)
         );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9647), .S(n9968), .Z(
        P1_U3549) );
  AOI22_X1 U10752 ( .A1(n9582), .A2(n9914), .B1(n9913), .B2(n5293), .ZN(n9583)
         );
  OAI211_X1 U10753 ( .C1(n9585), .C2(n9922), .A(n9584), .B(n9583), .ZN(n9648)
         );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9648), .S(n9968), .Z(
        P1_U3548) );
  AOI211_X1 U10755 ( .C1(n9913), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9589)
         );
  OAI21_X1 U10756 ( .B1(n9922), .B2(n9590), .A(n9589), .ZN(n9649) );
  MUX2_X1 U10757 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9649), .S(n9968), .Z(
        P1_U3547) );
  AOI22_X1 U10758 ( .A1(n9592), .A2(n9914), .B1(n9913), .B2(n9591), .ZN(n9593)
         );
  OAI211_X1 U10759 ( .C1(n9595), .C2(n9922), .A(n9594), .B(n9593), .ZN(n9650)
         );
  MUX2_X1 U10760 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9650), .S(n9968), .Z(
        P1_U3546) );
  AOI21_X1 U10761 ( .B1(n9913), .B2(n9597), .A(n9596), .ZN(n9598) );
  OAI211_X1 U10762 ( .C1(n9600), .C2(n9922), .A(n9599), .B(n9598), .ZN(n9651)
         );
  MUX2_X1 U10763 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9651), .S(n9968), .Z(
        P1_U3545) );
  AOI22_X1 U10764 ( .A1(n9602), .A2(n9914), .B1(n9913), .B2(n9601), .ZN(n9603)
         );
  OAI211_X1 U10765 ( .C1(n9605), .C2(n9922), .A(n9604), .B(n9603), .ZN(n9652)
         );
  MUX2_X1 U10766 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9652), .S(n9968), .Z(
        P1_U3544) );
  AOI22_X1 U10767 ( .A1(n9607), .A2(n9914), .B1(n9913), .B2(n9606), .ZN(n9608)
         );
  OAI211_X1 U10768 ( .C1(n9610), .C2(n9922), .A(n9609), .B(n9608), .ZN(n9653)
         );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9653), .S(n9968), .Z(
        P1_U3543) );
  AOI22_X1 U10770 ( .A1(n9612), .A2(n9914), .B1(n9913), .B2(n9611), .ZN(n9613)
         );
  OAI211_X1 U10771 ( .C1(n9615), .C2(n9922), .A(n9614), .B(n9613), .ZN(n9654)
         );
  MUX2_X1 U10772 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9654), .S(n9968), .Z(
        P1_U3542) );
  INV_X1 U10773 ( .A(n9922), .ZN(n9948) );
  NAND3_X1 U10774 ( .A1(n9617), .A2(n9616), .A3(n9948), .ZN(n9622) );
  AOI22_X1 U10775 ( .A1(n9619), .A2(n9914), .B1(n9913), .B2(n9618), .ZN(n9620)
         );
  NAND3_X1 U10776 ( .A1(n9622), .A2(n9621), .A3(n9620), .ZN(n9655) );
  MUX2_X1 U10777 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9655), .S(n9968), .Z(
        P1_U3541) );
  AOI22_X1 U10778 ( .A1(n9624), .A2(n9914), .B1(n9913), .B2(n9623), .ZN(n9625)
         );
  OAI211_X1 U10779 ( .C1(n9627), .C2(n9922), .A(n9626), .B(n9625), .ZN(n9656)
         );
  MUX2_X1 U10780 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9656), .S(n9968), .Z(
        P1_U3540) );
  AOI211_X1 U10781 ( .C1(n9913), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9631)
         );
  OAI21_X1 U10782 ( .B1(n9922), .B2(n9632), .A(n9631), .ZN(n9657) );
  MUX2_X1 U10783 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9657), .S(n9968), .Z(
        P1_U3539) );
  AOI211_X1 U10784 ( .C1(n9913), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9636)
         );
  OAI21_X1 U10785 ( .B1(n9922), .B2(n9637), .A(n9636), .ZN(n9658) );
  MUX2_X1 U10786 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9658), .S(n9968), .Z(
        P1_U3538) );
  INV_X1 U10787 ( .A(n9918), .ZN(n9903) );
  OAI22_X1 U10788 ( .A1(n9639), .A2(n9946), .B1(n9638), .B2(n9898), .ZN(n9640)
         );
  AOI21_X1 U10789 ( .B1(n9641), .B2(n9903), .A(n9640), .ZN(n9642) );
  NAND2_X1 U10790 ( .A1(n9643), .A2(n9642), .ZN(n9659) );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9659), .S(n9968), .Z(
        P1_U3536) );
  MUX2_X1 U10792 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9644), .S(n9952), .Z(
        P1_U3521) );
  MUX2_X1 U10793 ( .A(n9645), .B(P1_REG0_REG_28__SCAN_IN), .S(n9950), .Z(
        P1_U3519) );
  MUX2_X1 U10794 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9646), .S(n9952), .Z(
        P1_U3518) );
  MUX2_X1 U10795 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9647), .S(n9952), .Z(
        P1_U3517) );
  MUX2_X1 U10796 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9648), .S(n9952), .Z(
        P1_U3516) );
  MUX2_X1 U10797 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9649), .S(n9952), .Z(
        P1_U3515) );
  MUX2_X1 U10798 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9650), .S(n9952), .Z(
        P1_U3514) );
  MUX2_X1 U10799 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9651), .S(n9952), .Z(
        P1_U3513) );
  MUX2_X1 U10800 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9652), .S(n9952), .Z(
        P1_U3512) );
  MUX2_X1 U10801 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9653), .S(n9952), .Z(
        P1_U3511) );
  MUX2_X1 U10802 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9654), .S(n9952), .Z(
        P1_U3510) );
  MUX2_X1 U10803 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9655), .S(n9952), .Z(
        P1_U3508) );
  MUX2_X1 U10804 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9656), .S(n9952), .Z(
        P1_U3505) );
  MUX2_X1 U10805 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9657), .S(n9952), .Z(
        P1_U3502) );
  MUX2_X1 U10806 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9658), .S(n9952), .Z(
        P1_U3499) );
  MUX2_X1 U10807 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9659), .S(n9952), .Z(
        P1_U3493) );
  INV_X1 U10808 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9660) );
  NAND3_X1 U10809 ( .A1(n9660), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9661) );
  OAI22_X1 U10810 ( .A1(n9662), .A2(n9661), .B1(n6145), .B2(n9667), .ZN(n9663)
         );
  INV_X1 U10811 ( .A(n9663), .ZN(n9664) );
  OAI21_X1 U10812 ( .B1(n9666), .B2(n9665), .A(n9664), .ZN(P1_U3322) );
  OAI222_X1 U10813 ( .A1(n9671), .A2(n9670), .B1(n9669), .B2(P1_U3084), .C1(
        n9668), .C2(n9667), .ZN(P1_U3323) );
  OAI211_X1 U10814 ( .C1(n4514), .C2(n9898), .A(n9674), .B(n9673), .ZN(n9675)
         );
  AOI21_X1 U10815 ( .B1(n9948), .B2(n9676), .A(n9675), .ZN(n9679) );
  INV_X1 U10816 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10817 ( .A1(n9952), .A2(n9679), .B1(n9677), .B2(n9950), .ZN(
        P1_U3484) );
  AOI22_X1 U10818 ( .A1(n9968), .A2(n9679), .B1(n9678), .B2(n9965), .ZN(
        P1_U3533) );
  INV_X1 U10819 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9680) );
  OAI22_X1 U10820 ( .A1(n9682), .A2(n9681), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9680), .ZN(n9683) );
  AOI21_X1 U10821 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9697) );
  AND2_X1 U10822 ( .A1(n9688), .A2(n9686), .ZN(n9690) );
  NAND2_X1 U10823 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  OAI21_X1 U10824 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9695) );
  NOR2_X1 U10825 ( .A1(n9692), .A2(n9898), .ZN(n9722) );
  AOI22_X1 U10826 ( .A1(n9695), .A2(n9694), .B1(n9693), .B2(n9722), .ZN(n9696)
         );
  OAI211_X1 U10827 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(
        P1_U3222) );
  OAI21_X1 U10828 ( .B1(n9701), .B2(n9898), .A(n9700), .ZN(n9702) );
  INV_X1 U10829 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U10830 ( .A1(n9968), .A2(n9706), .B1(n9704), .B2(n9965), .ZN(
        P1_U3554) );
  INV_X1 U10831 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9705) );
  AOI22_X1 U10832 ( .A1(n9952), .A2(n9706), .B1(n9705), .B2(n9950), .ZN(
        P1_U3522) );
  INV_X1 U10833 ( .A(n9992), .ZN(n10018) );
  OAI21_X1 U10834 ( .B1(n9708), .B2(n10018), .A(n9707), .ZN(n9709) );
  AOI21_X1 U10835 ( .B1(n9710), .B2(n9993), .A(n9709), .ZN(n9712) );
  INV_X1 U10836 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9711) );
  AOI22_X1 U10837 ( .A1(n10039), .A2(n9712), .B1(n9711), .B2(n10037), .ZN(
        P2_U3550) );
  AOI22_X1 U10838 ( .A1(n10017), .A2(n9712), .B1(n8200), .B2(n10026), .ZN(
        P2_U3518) );
  OAI21_X1 U10839 ( .B1(n9714), .B2(n9898), .A(n9713), .ZN(n9715) );
  AOI211_X1 U10840 ( .C1(n9717), .C2(n9948), .A(n9716), .B(n9715), .ZN(n9726)
         );
  AOI22_X1 U10841 ( .A1(n9968), .A2(n9726), .B1(n9718), .B2(n9965), .ZN(
        P1_U3537) );
  NOR2_X1 U10842 ( .A1(n9719), .A2(n9922), .ZN(n9723) );
  NOR4_X1 U10843 ( .A1(n9723), .A2(n9722), .A3(n9721), .A4(n9720), .ZN(n9728)
         );
  AOI22_X1 U10844 ( .A1(n9968), .A2(n9728), .B1(n9724), .B2(n9965), .ZN(
        P1_U3535) );
  INV_X1 U10845 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10846 ( .A1(n9952), .A2(n9726), .B1(n9725), .B2(n9950), .ZN(
        P1_U3496) );
  INV_X1 U10847 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9727) );
  AOI22_X1 U10848 ( .A1(n9952), .A2(n9728), .B1(n9727), .B2(n9950), .ZN(
        P1_U3490) );
  XOR2_X1 U10849 ( .A(n9729), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10850 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9743) );
  INV_X1 U10851 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9738) );
  NOR2_X1 U10852 ( .A1(n9755), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9734) );
  OR2_X1 U10853 ( .A1(n9730), .A2(n9734), .ZN(n9732) );
  NAND2_X1 U10854 ( .A1(n9732), .A2(n9731), .ZN(n9758) );
  AOI21_X1 U10855 ( .B1(n9755), .B2(n9740), .A(P1_IR_REG_0__SCAN_IN), .ZN(
        n9733) );
  OR3_X1 U10856 ( .A1(n9734), .A2(n4312), .A3(n9733), .ZN(n9735) );
  NAND2_X1 U10857 ( .A1(n9758), .A2(n9735), .ZN(n9736) );
  OAI22_X1 U10858 ( .A1(n9782), .A2(n9738), .B1(n9737), .B2(n9736), .ZN(n9739)
         );
  INV_X1 U10859 ( .A(n9739), .ZN(n9742) );
  NAND3_X1 U10860 ( .A1(n9813), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9740), .ZN(
        n9741) );
  OAI211_X1 U10861 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9743), .A(n9742), .B(
        n9741), .ZN(P1_U3241) );
  INV_X1 U10862 ( .A(n9744), .ZN(n9748) );
  MUX2_X1 U10863 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6127), .S(n9754), .Z(n9747)
         );
  INV_X1 U10864 ( .A(n9745), .ZN(n9746) );
  AOI21_X1 U10865 ( .B1(n9748), .B2(n9747), .A(n9746), .ZN(n9763) );
  NAND2_X1 U10866 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9753) );
  OAI211_X1 U10867 ( .C1(n9751), .C2(n9750), .A(n9813), .B(n9749), .ZN(n9752)
         );
  OAI211_X1 U10868 ( .C1(n9808), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9762)
         );
  MUX2_X1 U10869 ( .A(n9757), .B(n9756), .S(n9755), .Z(n9760) );
  OAI211_X1 U10870 ( .C1(n9760), .C2(n4312), .A(n9759), .B(n9758), .ZN(n9780)
         );
  INV_X1 U10871 ( .A(n9780), .ZN(n9761) );
  AOI211_X1 U10872 ( .C1(n9817), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9764)
         );
  OAI21_X1 U10873 ( .B1(n9782), .B2(n9765), .A(n9764), .ZN(P1_U3243) );
  INV_X1 U10874 ( .A(n9766), .ZN(n9767) );
  OAI21_X1 U10875 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9770) );
  NAND2_X1 U10876 ( .A1(n9817), .A2(n9770), .ZN(n9777) );
  OAI21_X1 U10877 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9775) );
  AOI21_X1 U10878 ( .B1(n9813), .B2(n9775), .A(n9774), .ZN(n9776) );
  OAI211_X1 U10879 ( .C1(n9808), .C2(n9778), .A(n9777), .B(n9776), .ZN(n9779)
         );
  INV_X1 U10880 ( .A(n9779), .ZN(n9781) );
  OAI211_X1 U10881 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(
        P1_U3245) );
  INV_X1 U10882 ( .A(n9784), .ZN(n9785) );
  NOR2_X1 U10883 ( .A1(n9808), .A2(n9785), .ZN(n9786) );
  AOI211_X1 U10884 ( .C1(n9811), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9787), .B(
        n9786), .ZN(n9794) );
  OAI211_X1 U10885 ( .C1(n9789), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9813), .B(
        n9788), .ZN(n9793) );
  OAI211_X1 U10886 ( .C1(n9791), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9817), .B(
        n9790), .ZN(n9792) );
  NAND3_X1 U10887 ( .A1(n9794), .A2(n9793), .A3(n9792), .ZN(P1_U3256) );
  NOR2_X1 U10888 ( .A1(n9808), .A2(n9795), .ZN(n9796) );
  AOI211_X1 U10889 ( .C1(n9811), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9797), .B(
        n9796), .ZN(n9806) );
  OAI211_X1 U10890 ( .C1(n9800), .C2(n9799), .A(n9813), .B(n9798), .ZN(n9805)
         );
  OAI211_X1 U10891 ( .C1(n9803), .C2(n9802), .A(n9817), .B(n9801), .ZN(n9804)
         );
  NAND3_X1 U10892 ( .A1(n9806), .A2(n9805), .A3(n9804), .ZN(P1_U3257) );
  NOR2_X1 U10893 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  AOI211_X1 U10894 ( .C1(n9811), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9810), .B(
        n9809), .ZN(n9822) );
  OAI211_X1 U10895 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9821)
         );
  OAI211_X1 U10896 ( .C1(n9819), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9820)
         );
  NAND3_X1 U10897 ( .A1(n9822), .A2(n9821), .A3(n9820), .ZN(P1_U3258) );
  INV_X1 U10898 ( .A(n9823), .ZN(n9834) );
  INV_X1 U10899 ( .A(n9824), .ZN(n9830) );
  AOI22_X1 U10900 ( .A1(n9828), .A2(n9827), .B1(n9826), .B2(n9825), .ZN(n9829)
         );
  OAI21_X1 U10901 ( .B1(n9830), .B2(n9867), .A(n9829), .ZN(n9832) );
  AOI211_X1 U10902 ( .C1(n9834), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9835)
         );
  AOI22_X1 U10903 ( .A1(n9856), .A2(n6231), .B1(n9835), .B2(n9884), .ZN(
        P1_U3282) );
  AOI211_X1 U10904 ( .C1(n5015), .C2(n9837), .A(n9946), .B(n9836), .ZN(n9924)
         );
  OAI22_X1 U10905 ( .A1(n9839), .A2(n9881), .B1(n9880), .B2(n9838), .ZN(n9849)
         );
  NAND2_X1 U10906 ( .A1(n9841), .A2(n9840), .ZN(n9843) );
  INV_X1 U10907 ( .A(n9842), .ZN(n9853) );
  XNOR2_X1 U10908 ( .A(n9843), .B(n9853), .ZN(n9844) );
  NAND2_X1 U10909 ( .A1(n9844), .A2(n9871), .ZN(n9848) );
  AOI22_X1 U10910 ( .A1(n9873), .A2(n9846), .B1(n9845), .B2(n9875), .ZN(n9847)
         );
  NAND2_X1 U10911 ( .A1(n9848), .A2(n9847), .ZN(n9926) );
  AOI211_X1 U10912 ( .C1(n9924), .C2(n9850), .A(n9849), .B(n9926), .ZN(n9857)
         );
  INV_X1 U10913 ( .A(n9851), .ZN(n9854) );
  OAI21_X1 U10914 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9923) );
  OAI22_X1 U10915 ( .A1(n9857), .A2(n9856), .B1(n9923), .B2(n9855), .ZN(n9858)
         );
  INV_X1 U10916 ( .A(n9858), .ZN(n9859) );
  OAI21_X1 U10917 ( .B1(n6152), .B2(n9884), .A(n9859), .ZN(P1_U3286) );
  NAND2_X1 U10918 ( .A1(n6378), .A2(n9860), .ZN(n9861) );
  AND3_X1 U10919 ( .A1(n9862), .A2(n9914), .A3(n9861), .ZN(n9891) );
  OR2_X1 U10920 ( .A1(n9865), .A2(n9864), .ZN(n9866) );
  NAND2_X1 U10921 ( .A1(n9863), .A2(n9866), .ZN(n9890) );
  NOR2_X1 U10922 ( .A1(n9890), .A2(n6284), .ZN(n9868) );
  MUX2_X1 U10923 ( .A(n9891), .B(n9868), .S(n9867), .Z(n9883) );
  XNOR2_X1 U10924 ( .A(n9870), .B(n9869), .ZN(n9872) );
  NAND2_X1 U10925 ( .A1(n9872), .A2(n9871), .ZN(n9877) );
  AOI22_X1 U10926 ( .A1(n9875), .A2(n6292), .B1(n9874), .B2(n9873), .ZN(n9876)
         );
  OAI211_X1 U10927 ( .C1(n9878), .C2(n9890), .A(n9877), .B(n9876), .ZN(n9894)
         );
  OAI22_X1 U10928 ( .A1(n9893), .A2(n9881), .B1(n9880), .B2(n9879), .ZN(n9882)
         );
  NOR3_X1 U10929 ( .A1(n9883), .A2(n9894), .A3(n9882), .ZN(n9885) );
  AOI22_X1 U10930 ( .A1(n9856), .A2(n6128), .B1(n9885), .B2(n9884), .ZN(
        P1_U3290) );
  AND2_X1 U10931 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9886), .ZN(P1_U3292) );
  AND2_X1 U10932 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9886), .ZN(P1_U3293) );
  AND2_X1 U10933 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9886), .ZN(P1_U3294) );
  AND2_X1 U10934 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9886), .ZN(P1_U3295) );
  AND2_X1 U10935 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9886), .ZN(P1_U3296) );
  AND2_X1 U10936 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9886), .ZN(P1_U3297) );
  AND2_X1 U10937 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9886), .ZN(P1_U3298) );
  AND2_X1 U10938 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9886), .ZN(P1_U3299) );
  AND2_X1 U10939 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9886), .ZN(P1_U3300) );
  AND2_X1 U10940 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9886), .ZN(P1_U3301) );
  AND2_X1 U10941 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9886), .ZN(P1_U3302) );
  AND2_X1 U10942 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9886), .ZN(P1_U3303) );
  AND2_X1 U10943 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9886), .ZN(P1_U3304) );
  AND2_X1 U10944 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9886), .ZN(P1_U3305) );
  AND2_X1 U10945 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9886), .ZN(P1_U3306) );
  AND2_X1 U10946 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9886), .ZN(P1_U3307) );
  AND2_X1 U10947 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9886), .ZN(P1_U3308) );
  AND2_X1 U10948 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9886), .ZN(P1_U3309) );
  AND2_X1 U10949 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9886), .ZN(P1_U3310) );
  AND2_X1 U10950 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9886), .ZN(P1_U3311) );
  AND2_X1 U10951 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9886), .ZN(P1_U3312) );
  AND2_X1 U10952 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9886), .ZN(P1_U3313) );
  AND2_X1 U10953 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9886), .ZN(P1_U3314) );
  AND2_X1 U10954 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9886), .ZN(P1_U3315) );
  AND2_X1 U10955 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9886), .ZN(P1_U3316) );
  AND2_X1 U10956 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9886), .ZN(P1_U3317) );
  AND2_X1 U10957 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9886), .ZN(P1_U3318) );
  AND2_X1 U10958 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9886), .ZN(P1_U3319) );
  AND2_X1 U10959 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9886), .ZN(P1_U3320) );
  AND2_X1 U10960 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9886), .ZN(P1_U3321) );
  NAND2_X1 U10961 ( .A1(n9887), .A2(n9889), .ZN(n9888) );
  OAI21_X1 U10962 ( .B1(n5420), .B2(n9889), .A(n9888), .ZN(P1_U3441) );
  INV_X1 U10963 ( .A(n9890), .ZN(n9896) );
  INV_X1 U10964 ( .A(n9891), .ZN(n9892) );
  OAI21_X1 U10965 ( .B1(n9893), .B2(n9898), .A(n9892), .ZN(n9895) );
  AOI211_X1 U10966 ( .C1(n9903), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9954)
         );
  INV_X1 U10967 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10968 ( .A1(n9952), .A2(n9954), .B1(n9897), .B2(n9950), .ZN(
        P1_U3457) );
  AOI211_X1 U10969 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9956)
         );
  INV_X1 U10970 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10971 ( .A1(n9952), .A2(n9956), .B1(n9904), .B2(n9950), .ZN(
        P1_U3460) );
  AOI22_X1 U10972 ( .A1(n9906), .A2(n9914), .B1(n9913), .B2(n9905), .ZN(n9907)
         );
  OAI211_X1 U10973 ( .C1(n9909), .C2(n9918), .A(n9908), .B(n9907), .ZN(n9910)
         );
  INV_X1 U10974 ( .A(n9910), .ZN(n9958) );
  INV_X1 U10975 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10976 ( .A1(n9952), .A2(n9958), .B1(n9911), .B2(n9950), .ZN(
        P1_U3463) );
  AOI22_X1 U10977 ( .A1(n9915), .A2(n9914), .B1(n9913), .B2(n9912), .ZN(n9916)
         );
  OAI211_X1 U10978 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  INV_X1 U10979 ( .A(n9920), .ZN(n9959) );
  INV_X1 U10980 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9921) );
  AOI22_X1 U10981 ( .A1(n9952), .A2(n9959), .B1(n9921), .B2(n9950), .ZN(
        P1_U3466) );
  NOR2_X1 U10982 ( .A1(n9923), .A2(n9922), .ZN(n9927) );
  NOR4_X1 U10983 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9961)
         );
  INV_X1 U10984 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10985 ( .A1(n9952), .A2(n9961), .B1(n9928), .B2(n9950), .ZN(
        P1_U3469) );
  NAND2_X1 U10986 ( .A1(n9929), .A2(n9948), .ZN(n9935) );
  OAI21_X1 U10987 ( .B1(n9931), .B2(n9946), .A(n9930), .ZN(n9932) );
  NOR2_X1 U10988 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  AND2_X1 U10989 ( .A1(n9935), .A2(n9934), .ZN(n9962) );
  INV_X1 U10990 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U10991 ( .A1(n9952), .A2(n9962), .B1(n9936), .B2(n9950), .ZN(
        P1_U3472) );
  NAND3_X1 U10992 ( .A1(n9939), .A2(n9938), .A3(n9937), .ZN(n9940) );
  AOI21_X1 U10993 ( .B1(n9948), .B2(n9941), .A(n9940), .ZN(n9964) );
  INV_X1 U10994 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U10995 ( .A1(n9952), .A2(n9964), .B1(n9942), .B2(n9950), .ZN(
        P1_U3475) );
  OAI211_X1 U10996 ( .C1(n9946), .C2(n9945), .A(n9944), .B(n9943), .ZN(n9947)
         );
  AOI21_X1 U10997 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9967) );
  INV_X1 U10998 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U10999 ( .A1(n9952), .A2(n9967), .B1(n9951), .B2(n9950), .ZN(
        P1_U3478) );
  AOI22_X1 U11000 ( .A1(n9968), .A2(n9954), .B1(n9953), .B2(n9965), .ZN(
        P1_U3524) );
  INV_X1 U11001 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9955) );
  AOI22_X1 U11002 ( .A1(n9968), .A2(n9956), .B1(n9955), .B2(n9965), .ZN(
        P1_U3525) );
  AOI22_X1 U11003 ( .A1(n9968), .A2(n9958), .B1(n9957), .B2(n9965), .ZN(
        P1_U3526) );
  AOI22_X1 U11004 ( .A1(n9968), .A2(n9959), .B1(n6165), .B2(n9965), .ZN(
        P1_U3527) );
  INV_X1 U11005 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11006 ( .A1(n9968), .A2(n9961), .B1(n9960), .B2(n9965), .ZN(
        P1_U3528) );
  AOI22_X1 U11007 ( .A1(n9968), .A2(n9962), .B1(n6168), .B2(n9965), .ZN(
        P1_U3529) );
  INV_X1 U11008 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11009 ( .A1(n9968), .A2(n9964), .B1(n9963), .B2(n9965), .ZN(
        P1_U3530) );
  INV_X1 U11010 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9966) );
  AOI22_X1 U11011 ( .A1(n9968), .A2(n9967), .B1(n9966), .B2(n9965), .ZN(
        P1_U3531) );
  INV_X1 U11012 ( .A(n9969), .ZN(n9970) );
  AND2_X1 U11013 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9975), .ZN(P2_U3297) );
  AND2_X1 U11014 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9975), .ZN(P2_U3298) );
  AND2_X1 U11015 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9975), .ZN(P2_U3299) );
  AND2_X1 U11016 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9975), .ZN(P2_U3300) );
  AND2_X1 U11017 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9975), .ZN(P2_U3301) );
  AND2_X1 U11018 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9975), .ZN(P2_U3302) );
  AND2_X1 U11019 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9975), .ZN(P2_U3303) );
  AND2_X1 U11020 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9975), .ZN(P2_U3304) );
  AND2_X1 U11021 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9975), .ZN(P2_U3305) );
  AND2_X1 U11022 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9975), .ZN(P2_U3306) );
  AND2_X1 U11023 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9975), .ZN(P2_U3307) );
  AND2_X1 U11024 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9975), .ZN(P2_U3308) );
  AND2_X1 U11025 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9975), .ZN(P2_U3309) );
  AND2_X1 U11026 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9975), .ZN(P2_U3310) );
  AND2_X1 U11027 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9975), .ZN(P2_U3311) );
  AND2_X1 U11028 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9975), .ZN(P2_U3312) );
  AND2_X1 U11029 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9975), .ZN(P2_U3313) );
  AND2_X1 U11030 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9975), .ZN(P2_U3314) );
  AND2_X1 U11031 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9975), .ZN(P2_U3315) );
  AND2_X1 U11032 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9975), .ZN(P2_U3316) );
  AND2_X1 U11033 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9975), .ZN(P2_U3317) );
  AND2_X1 U11034 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9975), .ZN(P2_U3318) );
  AND2_X1 U11035 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9975), .ZN(P2_U3319) );
  AND2_X1 U11036 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9975), .ZN(P2_U3320) );
  AND2_X1 U11037 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9975), .ZN(P2_U3321) );
  AND2_X1 U11038 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9975), .ZN(P2_U3322) );
  AND2_X1 U11039 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9975), .ZN(P2_U3323) );
  AND2_X1 U11040 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9975), .ZN(P2_U3324) );
  AND2_X1 U11041 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9975), .ZN(P2_U3325) );
  AND2_X1 U11042 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9975), .ZN(P2_U3326) );
  AOI22_X1 U11043 ( .A1(n9978), .A2(n9973), .B1(n9972), .B2(n9975), .ZN(
        P2_U3437) );
  INV_X1 U11044 ( .A(n9974), .ZN(n9977) );
  AOI22_X1 U11045 ( .A1(n9978), .A2(n9977), .B1(n9976), .B2(n9975), .ZN(
        P2_U3438) );
  AOI22_X1 U11046 ( .A1(n9980), .A2(n10024), .B1(n5965), .B2(n9979), .ZN(n9981) );
  AND2_X1 U11047 ( .A1(n9982), .A2(n9981), .ZN(n10028) );
  AOI22_X1 U11048 ( .A1(n10017), .A2(n10028), .B1(n5531), .B2(n10026), .ZN(
        P2_U3451) );
  NAND3_X1 U11049 ( .A1(n9984), .A2(n9993), .A3(n9983), .ZN(n9985) );
  OAI21_X1 U11050 ( .B1(n9986), .B2(n10018), .A(n9985), .ZN(n9989) );
  INV_X1 U11051 ( .A(n9987), .ZN(n9988) );
  AOI211_X1 U11052 ( .C1(n10024), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10029) );
  AOI22_X1 U11053 ( .A1(n10017), .A2(n10029), .B1(n5517), .B2(n10026), .ZN(
        P2_U3454) );
  AOI22_X1 U11054 ( .A1(n9994), .A2(n9993), .B1(n9992), .B2(n9991), .ZN(n9995)
         );
  NAND2_X1 U11055 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  AOI21_X1 U11056 ( .B1(n10024), .B2(n9998), .A(n9997), .ZN(n10031) );
  AOI22_X1 U11057 ( .A1(n10017), .A2(n10031), .B1(n5563), .B2(n10026), .ZN(
        P2_U3460) );
  OAI211_X1 U11058 ( .C1(n10001), .C2(n10018), .A(n10000), .B(n9999), .ZN(
        n10002) );
  AOI21_X1 U11059 ( .B1(n10024), .B2(n10003), .A(n10002), .ZN(n10033) );
  AOI22_X1 U11060 ( .A1(n10017), .A2(n10033), .B1(n5510), .B2(n10026), .ZN(
        P2_U3466) );
  OAI22_X1 U11061 ( .A1(n10005), .A2(n10020), .B1(n10004), .B2(n10018), .ZN(
        n10007) );
  AOI211_X1 U11062 ( .C1(n10008), .C2(n10024), .A(n10007), .B(n10006), .ZN(
        n10034) );
  AOI22_X1 U11063 ( .A1(n10017), .A2(n10034), .B1(n5455), .B2(n10026), .ZN(
        P2_U3472) );
  INV_X1 U11064 ( .A(n10009), .ZN(n10016) );
  INV_X1 U11065 ( .A(n10010), .ZN(n10015) );
  OAI22_X1 U11066 ( .A1(n10012), .A2(n10020), .B1(n10011), .B2(n10018), .ZN(
        n10014) );
  AOI211_X1 U11067 ( .C1(n10016), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10036) );
  AOI22_X1 U11068 ( .A1(n10017), .A2(n10036), .B1(n5630), .B2(n10026), .ZN(
        P2_U3478) );
  OAI22_X1 U11069 ( .A1(n10021), .A2(n10020), .B1(n10019), .B2(n10018), .ZN(
        n10023) );
  AOI211_X1 U11070 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10038) );
  INV_X1 U11071 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11072 ( .A1(n10017), .A2(n10038), .B1(n10027), .B2(n10026), .ZN(
        P2_U3484) );
  AOI22_X1 U11073 ( .A1(n10039), .A2(n10028), .B1(n6848), .B2(n10037), .ZN(
        P2_U3520) );
  AOI22_X1 U11074 ( .A1(n10039), .A2(n10029), .B1(n6695), .B2(n10037), .ZN(
        P2_U3521) );
  AOI22_X1 U11075 ( .A1(n10039), .A2(n10031), .B1(n10030), .B2(n10037), .ZN(
        P2_U3523) );
  AOI22_X1 U11076 ( .A1(n10039), .A2(n10033), .B1(n10032), .B2(n10037), .ZN(
        P2_U3525) );
  AOI22_X1 U11077 ( .A1(n10039), .A2(n10034), .B1(n6691), .B2(n10037), .ZN(
        P2_U3527) );
  AOI22_X1 U11078 ( .A1(n10039), .A2(n10036), .B1(n10035), .B2(n10037), .ZN(
        P2_U3529) );
  AOI22_X1 U11079 ( .A1(n10039), .A2(n10038), .B1(n6706), .B2(n10037), .ZN(
        P2_U3531) );
  INV_X1 U11080 ( .A(n10040), .ZN(n10041) );
  NAND2_X1 U11081 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  XOR2_X1 U11082 ( .A(n7224), .B(n10043), .Z(ADD_1071_U5) );
  XOR2_X1 U11083 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11084 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(ADD_1071_U56) );
  OAI21_X1 U11085 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(ADD_1071_U57) );
  OAI21_X1 U11086 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(ADD_1071_U58) );
  OAI21_X1 U11087 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U59) );
  OAI21_X1 U11088 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(ADD_1071_U60) );
  OAI21_X1 U11089 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(ADD_1071_U61) );
  AOI21_X1 U11090 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(ADD_1071_U62) );
  AOI21_X1 U11091 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(ADD_1071_U63) );
  AOI21_X1 U11092 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(ADD_1071_U47) );
  XOR2_X1 U11093 ( .A(n10072), .B(n10071), .Z(ADD_1071_U54) );
  XOR2_X1 U11094 ( .A(n10073), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11095 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n10077) );
  XNOR2_X1 U11096 ( .A(n10077), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11097 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10078), .Z(ADD_1071_U49) );
  XOR2_X1 U11098 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10079), .Z(ADD_1071_U50) );
  AOI21_X1 U11099 ( .B1(n10081), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10080), .ZN(
        n10082) );
  XOR2_X1 U11100 ( .A(n10082), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11101 ( .A(n10084), .B(n10083), .Z(ADD_1071_U53) );
  XNOR2_X1 U11102 ( .A(n10086), .B(n10085), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4833 ( .A(n5540), .Z(n6667) );
  CLKBUF_X1 U4838 ( .A(n4959), .Z(n6325) );
  CLKBUF_X1 U4891 ( .A(n4955), .Z(n5039) );
  CLKBUF_X1 U4945 ( .A(n8509), .Z(n4310) );
  CLKBUF_X1 U5117 ( .A(n5378), .Z(n4312) );
endmodule

