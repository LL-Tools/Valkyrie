

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4374, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486;

  NAND2_X1 U4879 ( .A1(n7405), .A2(n9637), .ZN(n7131) );
  AND2_X1 U4880 ( .A1(n7563), .A2(n10074), .ZN(n7300) );
  BUF_X2 U4881 ( .A(n6465), .Z(n6622) );
  CLKBUF_X2 U4882 ( .A(n6379), .Z(n6201) );
  CLKBUF_X2 U4883 ( .A(n8190), .Z(n4379) );
  OR2_X1 U4884 ( .A1(n5996), .A2(n5825), .ZN(n5959) );
  NAND4_X1 U4885 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n8448)
         );
  NAND2_X2 U4886 ( .A1(n6641), .A2(n6728), .ZN(n6132) );
  XNOR2_X1 U4888 ( .A(n6040), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6611) );
  INV_X1 U4889 ( .A(n7649), .ZN(n5978) );
  NAND2_X1 U4890 ( .A1(n5648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U4891 ( .A1(n5114), .A2(n8138), .ZN(n6686) );
  NAND2_X1 U4892 ( .A1(n5105), .A2(n5104), .ZN(n8138) );
  BUF_X1 U4893 ( .A(n5131), .Z(n4524) );
  INV_X1 U4894 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U4895 ( .A1(n4668), .A2(n4667), .ZN(n8034) );
  NAND2_X1 U4896 ( .A1(n8693), .A2(n8692), .ZN(n8682) );
  NAND2_X1 U4897 ( .A1(n7168), .A2(n7167), .ZN(n8190) );
  INV_X1 U4898 ( .A(n5959), .ZN(n5939) );
  NAND2_X1 U4901 ( .A1(n8242), .A2(n7188), .ZN(n8358) );
  INV_X2 U4902 ( .A(n6686), .ZN(n6718) );
  AND2_X1 U4903 ( .A1(n6686), .A2(n4380), .ZN(n5186) );
  AND2_X1 U4904 ( .A1(n5207), .A2(n5206), .ZN(n10074) );
  NAND2_X1 U4905 ( .A1(n5302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5303) );
  INV_X1 U4906 ( .A(n7129), .ZN(n6634) );
  INV_X1 U4907 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U4908 ( .A1(n5305), .A2(n5304), .ZN(n7796) );
  OAI22_X1 U4909 ( .A1(n8673), .A2(n8684), .B1(n8680), .B2(n8695), .ZN(n8659)
         );
  NOR3_X1 U4910 ( .A1(n8959), .A2(n8958), .A3(n8957), .ZN(n8962) );
  BUF_X1 U4911 ( .A(n6096), .Z(n7076) );
  OR2_X1 U4913 ( .A1(n9470), .A2(n9692), .ZN(n9471) );
  INV_X2 U4915 ( .A(n7131), .ZN(n9679) );
  OR2_X1 U4916 ( .A1(n5994), .A2(n5971), .ZN(n4374) );
  MUX2_X2 U4917 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n6026) );
  AND2_X1 U4918 ( .A1(n5617), .A2(n4407), .ZN(n5620) );
  OR2_X1 U4919 ( .A1(n5617), .A2(n8890), .ZN(n5624) );
  XNOR2_X2 U4920 ( .A(n5303), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7287) );
  XNOR2_X1 U4921 ( .A(n5627), .B(n5626), .ZN(n7649) );
  OAI21_X2 U4922 ( .B1(n4728), .B2(n4727), .A(n4724), .ZN(n9344) );
  OR2_X4 U4923 ( .A1(n6890), .A2(n6641), .ZN(n7129) );
  BUF_X4 U4924 ( .A(n6159), .Z(n4377) );
  INV_X1 U4925 ( .A(n6139), .ZN(n6159) );
  AOI211_X2 U4926 ( .C1(n9934), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9723)
         );
  XNOR2_X1 U4928 ( .A(n6038), .B(n6037), .ZN(n9332) );
  XNOR2_X2 U4929 ( .A(n5273), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8482) );
  XNOR2_X2 U4930 ( .A(n6212), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6910) );
  AND2_X4 U4931 ( .A1(n4581), .A2(n4580), .ZN(n4380) );
  INV_X1 U4932 ( .A(n5598), .ZN(n5131) );
  NAND2_X1 U4933 ( .A1(n8174), .A2(n5061), .ZN(n8225) );
  NAND2_X1 U4934 ( .A1(n8617), .A2(n5046), .ZN(n8598) );
  NAND2_X1 U4935 ( .A1(n9593), .A2(n9223), .ZN(n9575) );
  CLKBUF_X1 U4936 ( .A(n8128), .Z(n4384) );
  NAND2_X1 U4937 ( .A1(n4639), .A2(n6211), .ZN(n7353) );
  NAND2_X1 U4938 ( .A1(n6353), .A2(n6352), .ZN(n9764) );
  NAND2_X1 U4939 ( .A1(n5383), .A2(n5382), .ZN(n5704) );
  AND2_X1 U4940 ( .A1(n8270), .A2(n7175), .ZN(n8125) );
  AND2_X1 U4941 ( .A1(n7069), .A2(n6108), .ZN(n6127) );
  INV_X2 U4942 ( .A(n7144), .ZN(n9966) );
  INV_X2 U4943 ( .A(n6946), .ZN(n7497) );
  INV_X1 U4944 ( .A(n10016), .ZN(n8239) );
  NAND2_X1 U4945 ( .A1(n9364), .A2(n7473), .ZN(n9295) );
  INV_X2 U4946 ( .A(n6379), .ZN(n6163) );
  INV_X1 U4947 ( .A(n9157), .ZN(n9164) );
  AND4_X1 U4948 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n7668)
         );
  INV_X2 U4949 ( .A(n7122), .ZN(n7456) );
  NAND2_X1 U4950 ( .A1(n5103), .A2(n5083), .ZN(n5104) );
  OR2_X1 U4951 ( .A1(n6024), .A2(n4984), .ZN(n4405) );
  INV_X2 U4952 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X2 U4953 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U4954 ( .A1(n5769), .A2(n5768), .ZN(n6004) );
  AND2_X1 U4955 ( .A1(n8563), .A2(n5767), .ZN(n5768) );
  NOR2_X1 U4956 ( .A1(n8407), .A2(n8201), .ZN(n8199) );
  AOI21_X1 U4957 ( .B1(n8571), .B2(n10020), .A(n8570), .ZN(n8795) );
  OAI21_X1 U4958 ( .B1(n4491), .B2(n5970), .A(n5969), .ZN(n5994) );
  OAI21_X1 U4959 ( .B1(n5819), .B2(n5990), .A(n5967), .ZN(n5820) );
  AND2_X1 U4960 ( .A1(n4881), .A2(n4879), .ZN(n8407) );
  AOI21_X1 U4961 ( .B1(n5966), .B2(n5965), .A(n5964), .ZN(n4491) );
  AND2_X1 U4962 ( .A1(n4774), .A2(n4392), .ZN(n8913) );
  AND2_X1 U4963 ( .A1(n9161), .A2(n9160), .ZN(n4728) );
  AND2_X1 U4964 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  NAND2_X1 U4965 ( .A1(n8960), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U4966 ( .A1(n8225), .A2(n8182), .ZN(n8339) );
  AOI21_X1 U4967 ( .B1(n9492), .B2(n9656), .A(n9491), .ZN(n9713) );
  OR2_X1 U4968 ( .A1(n8094), .A2(n8095), .ZN(n8922) );
  AOI21_X1 U4969 ( .B1(n9535), .B2(n9656), .A(n4536), .ZN(n9728) );
  NAND2_X1 U4970 ( .A1(n4616), .A2(n6522), .ZN(n9007) );
  AND2_X1 U4971 ( .A1(n9165), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U4972 ( .A1(n9214), .A2(n9219), .ZN(n9691) );
  NAND2_X1 U4973 ( .A1(n8051), .A2(n8050), .ZN(n8217) );
  NAND2_X1 U4974 ( .A1(n4548), .A2(n8016), .ZN(n9625) );
  INV_X1 U4975 ( .A(n4857), .ZN(n7901) );
  INV_X1 U4976 ( .A(n4837), .ZN(n4836) );
  OAI211_X1 U4977 ( .C1(n4719), .C2(n5707), .A(n4401), .B(n4714), .ZN(n8673)
         );
  NAND2_X1 U4978 ( .A1(n5479), .A2(n5478), .ZN(n8822) );
  NAND2_X1 U4979 ( .A1(n6506), .A2(n6505), .ZN(n9731) );
  NAND2_X1 U4980 ( .A1(n7353), .A2(n7350), .ZN(n4888) );
  INV_X1 U4981 ( .A(n8700), .ZN(n8834) );
  NAND2_X1 U4982 ( .A1(n6491), .A2(n6490), .ZN(n9736) );
  NOR2_X1 U4983 ( .A1(n9374), .A2(n4785), .ZN(n9377) );
  AND2_X1 U4984 ( .A1(n5441), .A2(n5440), .ZN(n8700) );
  NAND2_X1 U4985 ( .A1(n4490), .A2(n5426), .ZN(n8838) );
  OAI211_X1 U4986 ( .C1(n7612), .C2(n5699), .A(n5067), .B(n5698), .ZN(n7750)
         );
  NAND2_X1 U4987 ( .A1(n6165), .A2(n6164), .ZN(n7087) );
  NAND2_X1 U4988 ( .A1(n5409), .A2(n5408), .ZN(n8842) );
  NAND2_X1 U4989 ( .A1(n6369), .A2(n6368), .ZN(n9672) );
  NAND2_X1 U4990 ( .A1(n6387), .A2(n6386), .ZN(n9774) );
  NAND2_X1 U4991 ( .A1(n5350), .A2(n5349), .ZN(n8854) );
  XNOR2_X1 U4992 ( .A(n5402), .B(n5401), .ZN(n7039) );
  XNOR2_X1 U4993 ( .A(n5422), .B(n5416), .ZN(n7023) );
  OAI21_X1 U4994 ( .B1(n5422), .B2(n5416), .A(n5417), .ZN(n5402) );
  NAND2_X1 U4995 ( .A1(n6296), .A2(n6295), .ZN(n7792) );
  INV_X1 U4996 ( .A(n5693), .ZN(n7619) );
  NAND2_X1 U4997 ( .A1(n6126), .A2(n6127), .ZN(n7071) );
  NAND2_X1 U4998 ( .A1(n6313), .A2(n6312), .ZN(n9779) );
  NAND2_X1 U4999 ( .A1(n5346), .A2(n5345), .ZN(n5373) );
  AND2_X1 U5000 ( .A1(n7138), .A2(n5009), .ZN(n7401) );
  NAND2_X1 U5001 ( .A1(n7551), .A2(n5863), .ZN(n7557) );
  NAND2_X1 U5002 ( .A1(n5253), .A2(n5252), .ZN(n10088) );
  NAND2_X1 U5003 ( .A1(n5275), .A2(n5274), .ZN(n10095) );
  NAND2_X1 U5004 ( .A1(n6238), .A2(n6237), .ZN(n9795) );
  OR2_X1 U5005 ( .A1(n8448), .A2(n7556), .ZN(n7551) );
  XNOR2_X1 U5006 ( .A(n5222), .B(n5238), .ZN(n6752) );
  NAND2_X1 U5007 ( .A1(n6199), .A2(n6198), .ZN(n7144) );
  AND2_X1 U5008 ( .A1(n5192), .A2(n5191), .ZN(n7556) );
  NAND2_X1 U5009 ( .A1(n5124), .A2(n5123), .ZN(n5854) );
  CLKBUF_X3 U5010 ( .A(n6121), .Z(n6465) );
  XNOR2_X1 U5011 ( .A(n5202), .B(n5185), .ZN(n6737) );
  AND4_X1 U5012 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(n7741)
         );
  BUF_X2 U5013 ( .A(n7668), .Z(n4388) );
  CLKBUF_X1 U5014 ( .A(n6924), .Z(n7052) );
  NAND4_X1 U5015 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n10018)
         );
  NAND4_X1 U5016 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n9364)
         );
  AND4_X1 U5017 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n7667)
         );
  AND4_X1 U5018 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n7080)
         );
  INV_X1 U5019 ( .A(n10057), .ZN(n7534) );
  AND2_X2 U5020 ( .A1(n6778), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U5021 ( .A(n9933), .ZN(n6935) );
  NAND3_X1 U5022 ( .A1(n10045), .A2(n7729), .A3(n7166), .ZN(n7168) );
  AOI21_X1 U5023 ( .B1(n4454), .B2(n5058), .A(n4400), .ZN(n4598) );
  BUF_X2 U5024 ( .A(n4377), .Z(n6578) );
  AND2_X1 U5025 ( .A1(n4768), .A2(n4767), .ZN(n4766) );
  CLKBUF_X1 U5026 ( .A(n5678), .Z(n5996) );
  INV_X2 U5027 ( .A(n9055), .ZN(n9064) );
  NOR2_X1 U5028 ( .A1(n6820), .A2(n4811), .ZN(n4810) );
  OAI21_X1 U5029 ( .B1(n5289), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  XNOR2_X1 U5030 ( .A(n5622), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5677) );
  INV_X2 U5031 ( .A(n6783), .ZN(n6453) );
  OR2_X1 U5032 ( .A1(n5250), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U5033 ( .A(n6080), .B(n6079), .ZN(n9281) );
  OAI21_X1 U5034 ( .B1(n6078), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U5035 ( .A1(n5621), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5622) );
  OAI21_X1 U5036 ( .B1(n6063), .B2(P1_IR_REG_28__SCAN_IN), .A(n6062), .ZN(
        n6067) );
  NAND2_X1 U5037 ( .A1(n5104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U5038 ( .A1(n6033), .A2(n6032), .ZN(n6078) );
  OR2_X1 U5039 ( .A1(n6058), .A2(n6061), .ZN(n6023) );
  OAI21_X1 U5040 ( .B1(n6614), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U5041 ( .A1(n4405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6060) );
  NAND2_X2 U5042 ( .A1(n4380), .A2(P1_U3084), .ZN(n9840) );
  NOR2_X1 U5043 ( .A1(n5458), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5617) );
  AND3_X1 U5044 ( .A1(n4958), .A2(n6016), .A3(n4957), .ZN(n6039) );
  AND3_X1 U5045 ( .A1(n6029), .A2(n6196), .A3(n6030), .ZN(n6350) );
  AND2_X1 U5046 ( .A1(n4955), .A2(n4954), .ZN(n4953) );
  NAND2_X1 U5047 ( .A1(n5097), .A2(n9447), .ZN(n4581) );
  NAND2_X1 U5048 ( .A1(n5099), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4580) );
  AND2_X1 U5049 ( .A1(n4751), .A2(n4407), .ZN(n4750) );
  AND4_X1 U5050 ( .A1(n6021), .A2(n6045), .A3(n6041), .A4(n6020), .ZN(n6022)
         );
  AND4_X1 U5051 ( .A1(n5080), .A2(n5656), .A3(n5668), .A4(n5618), .ZN(n5082)
         );
  AND2_X1 U5052 ( .A1(n5078), .A2(n5077), .ZN(n5405) );
  INV_X1 U5053 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6041) );
  INV_X1 U5054 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6037) );
  INV_X1 U5055 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5656) );
  INV_X4 U5056 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5057 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5098) );
  NOR2_X1 U5058 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5077) );
  INV_X1 U5059 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6365) );
  INV_X1 U5060 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10416) );
  INV_X1 U5061 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U5062 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6011) );
  INV_X1 U5063 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10441) );
  INV_X1 U5064 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6179) );
  OR2_X2 U5065 ( .A1(n5678), .A2(n5677), .ZN(n10045) );
  INV_X1 U5066 ( .A(n5678), .ZN(n5716) );
  INV_X1 U5067 ( .A(n5677), .ZN(n7729) );
  NAND2_X2 U5068 ( .A1(n5179), .A2(n5842), .ZN(n7550) );
  NAND2_X2 U5069 ( .A1(n8358), .A2(n4884), .ZN(n8397) );
  NAND2_X2 U5070 ( .A1(n8397), .A2(n7199), .ZN(n8396) );
  AND2_X1 U5071 ( .A1(n5082), .A2(n5079), .ZN(n4749) );
  BUF_X4 U5072 ( .A(n5186), .Z(n5582) );
  NOR2_X4 U5073 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5117) );
  NAND2_X2 U5074 ( .A1(n6618), .A2(n9332), .ZN(n6889) );
  AND2_X2 U5075 ( .A1(n6076), .A2(n6036), .ZN(n6618) );
  NOR2_X2 U5076 ( .A1(n5086), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8888) );
  NAND2_X2 U5077 ( .A1(n8396), .A2(n4885), .ZN(n7314) );
  NAND2_X2 U5078 ( .A1(n7903), .A2(n7902), .ZN(n7964) );
  XNOR2_X1 U5079 ( .A(n7189), .B(n7190), .ZN(n8360) );
  INV_X4 U5080 ( .A(n5254), .ZN(n5786) );
  NAND2_X1 U5081 ( .A1(n8125), .A2(n8124), .ZN(n8123) );
  NAND2_X2 U5082 ( .A1(n7966), .A2(n7965), .ZN(n8051) );
  NAND2_X1 U5083 ( .A1(n7823), .A2(n7706), .ZN(n7824) );
  INV_X2 U5084 ( .A(n5254), .ZN(n5444) );
  INV_X2 U5085 ( .A(n6132), .ZN(n6121) );
  CLKBUF_X1 U5086 ( .A(n7158), .Z(n4381) );
  AOI21_X1 U5087 ( .B1(n4384), .B2(n9222), .A(n5059), .ZN(n4382) );
  OAI21_X1 U5088 ( .B1(n7158), .B2(n9261), .A(n9300), .ZN(n4385) );
  XNOR2_X1 U5089 ( .A(n6060), .B(n6059), .ZN(n4386) );
  AOI21_X1 U5090 ( .B1(n8128), .B2(n9222), .A(n5059), .ZN(n9594) );
  OAI21_X1 U5091 ( .B1(n8034), .B2(n4967), .A(n4965), .ZN(n8128) );
  NAND2_X1 U5092 ( .A1(n7133), .A2(n9265), .ZN(n7158) );
  OAI21_X1 U5093 ( .B1(n7158), .B2(n9261), .A(n9300), .ZN(n7422) );
  XNOR2_X1 U5094 ( .A(n6060), .B(n6059), .ZN(n6070) );
  NAND2_X1 U5095 ( .A1(n7668), .A2(n7076), .ZN(n9289) );
  NAND2_X1 U5097 ( .A1(n7074), .A2(n9933), .ZN(n9293) );
  NOR2_X1 U5098 ( .A1(n6309), .A2(n6015), .ZN(n6029) );
  NOR2_X1 U5099 ( .A1(n9365), .A2(n7457), .ZN(n6938) );
  NAND4_X2 U5100 ( .A1(n6106), .A2(n6103), .A3(n6104), .A4(n6105), .ZN(n9365)
         );
  CLKBUF_X1 U5101 ( .A(n6174), .Z(n4389) );
  BUF_X4 U5102 ( .A(n6174), .Z(n4390) );
  BUF_X4 U5103 ( .A(n6174), .Z(n4391) );
  AND2_X2 U5104 ( .A1(n4386), .A2(n9832), .ZN(n6174) );
  MUX2_X1 U5105 ( .A(n9128), .B(n9127), .S(n9157), .Z(n9136) );
  NAND2_X1 U5106 ( .A1(n5398), .A2(n5397), .ZN(n5419) );
  INV_X1 U5107 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5299) );
  OR2_X1 U5108 ( .A1(n7893), .A2(n7969), .ZN(n5891) );
  NAND2_X1 U5109 ( .A1(n9700), .A2(n8148), .ZN(n9461) );
  OR2_X1 U5110 ( .A1(n9700), .A2(n8148), .ZN(n9460) );
  OR2_X1 U5111 ( .A1(n9706), .A2(n8026), .ZN(n9274) );
  NAND2_X1 U5112 ( .A1(n9505), .A2(n9143), .ZN(n9485) );
  OR2_X1 U5113 ( .A1(n9715), .A2(n9518), .ZN(n9484) );
  NOR2_X1 U5114 ( .A1(n4979), .A2(n8018), .ZN(n4976) );
  NOR2_X1 U5115 ( .A1(n8017), .A2(n4423), .ZN(n4979) );
  OR2_X1 U5116 ( .A1(n4672), .A2(n4670), .ZN(n4667) );
  NAND2_X1 U5117 ( .A1(n7938), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U5118 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  OR2_X1 U5119 ( .A1(n9795), .A2(n7659), .ZN(n9078) );
  NAND2_X1 U5120 ( .A1(n4584), .A2(n4586), .ZN(n5592) );
  INV_X1 U5121 ( .A(n4587), .ZN(n4586) );
  OAI21_X1 U5122 ( .B1(n4909), .B2(n4588), .A(n5735), .ZN(n4587) );
  AOI21_X1 U5123 ( .B1(n6078), .B2(P1_IR_REG_31__SCAN_IN), .A(n4893), .ZN(
        n4892) );
  NAND2_X1 U5124 ( .A1(n4894), .A2(n6034), .ZN(n4893) );
  NAND2_X1 U5125 ( .A1(n4895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U5126 ( .A1(n5265), .A2(n5247), .ZN(n5266) );
  NOR2_X1 U5127 ( .A1(n6963), .A2(n10038), .ZN(n6976) );
  INV_X1 U5128 ( .A(n5791), .ZN(n5790) );
  BUF_X1 U5129 ( .A(n5272), .Z(n4689) );
  INV_X1 U5130 ( .A(n10038), .ZN(n6717) );
  INV_X1 U5131 ( .A(n9059), .ZN(n6650) );
  NAND2_X1 U5132 ( .A1(n9139), .A2(n9247), .ZN(n4735) );
  INV_X1 U5133 ( .A(n5045), .ZN(n5000) );
  INV_X1 U5134 ( .A(n7502), .ZN(n5006) );
  NAND2_X1 U5135 ( .A1(n5473), .A2(n5472), .ZN(n5490) );
  INV_X1 U5136 ( .A(n5370), .ZN(n4597) );
  NAND2_X1 U5137 ( .A1(n5269), .A2(n5268), .ZN(n5285) );
  INV_X1 U5138 ( .A(SI_9_), .ZN(n5268) );
  NOR2_X1 U5139 ( .A1(n4648), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U5140 ( .A1(n4433), .A2(n4417), .ZN(n4928) );
  OAI21_X1 U5141 ( .B1(n4706), .B2(n4705), .A(n4450), .ZN(n4703) );
  NOR2_X1 U5142 ( .A1(n5709), .A2(n4413), .ZN(n4709) );
  OR2_X1 U5143 ( .A1(n8812), .A2(n8282), .ZN(n5929) );
  INV_X1 U5144 ( .A(n5922), .ZN(n4838) );
  INV_X1 U5145 ( .A(n5706), .ZN(n5036) );
  OR2_X1 U5146 ( .A1(n8858), .A2(n8208), .ZN(n5839) );
  NAND2_X1 U5147 ( .A1(n7635), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U5148 ( .A1(n4830), .A2(n5889), .ZN(n4651) );
  NAND2_X1 U5149 ( .A1(n7864), .A2(n5881), .ZN(n4830) );
  OR2_X1 U5150 ( .A1(n7796), .A2(n9999), .ZN(n5887) );
  NOR2_X2 U5151 ( .A1(n7301), .A2(n10088), .ZN(n7624) );
  OR2_X1 U5152 ( .A1(n8777), .A2(n8265), .ZN(n5960) );
  AND3_X2 U5153 ( .A1(n4687), .A2(n4416), .A3(n4749), .ZN(n5103) );
  AND2_X1 U5154 ( .A1(n4750), .A2(n5406), .ZN(n4687) );
  AND2_X1 U5155 ( .A1(n7877), .A2(n7874), .ZN(n6327) );
  INV_X1 U5156 ( .A(n6070), .ZN(n6068) );
  INV_X1 U5157 ( .A(n4810), .ZN(n4804) );
  INV_X1 U5158 ( .A(n9691), .ZN(n9464) );
  INV_X1 U5159 ( .A(n9274), .ZN(n4678) );
  NAND2_X1 U5160 ( .A1(n4995), .A2(n4406), .ZN(n4994) );
  NAND2_X1 U5161 ( .A1(n9172), .A2(n9316), .ZN(n4995) );
  NAND2_X1 U5162 ( .A1(n4503), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6582) );
  OR2_X1 U5163 ( .A1(n9722), .A2(n8963), .ZN(n9249) );
  INV_X1 U5164 ( .A(n4999), .ZN(n4998) );
  OAI21_X1 U5165 ( .B1(n9555), .B2(n5000), .A(n8022), .ZN(n4999) );
  OR2_X1 U5166 ( .A1(n9731), .A2(n9564), .ZN(n8022) );
  NOR2_X1 U5167 ( .A1(n4447), .A2(n4983), .ZN(n4982) );
  INV_X1 U5168 ( .A(n7839), .ZN(n4983) );
  INV_X1 U5169 ( .A(n9186), .ZN(n7153) );
  NAND2_X1 U5170 ( .A1(n7506), .A2(n4424), .ZN(n7519) );
  AND2_X1 U5171 ( .A1(n4378), .A2(n9281), .ZN(n6891) );
  AOI21_X1 U5172 ( .B1(n4994), .B2(n4996), .A(n4992), .ZN(n4991) );
  INV_X1 U5173 ( .A(n4405), .ZN(n6065) );
  NAND2_X1 U5174 ( .A1(n5743), .A2(n5742), .ZN(n5776) );
  AND2_X1 U5175 ( .A1(n5741), .A2(n5740), .ZN(n5743) );
  OR2_X1 U5176 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  NAND2_X1 U5177 ( .A1(n5523), .A2(n5510), .ZN(n5524) );
  NAND2_X1 U5178 ( .A1(n5454), .A2(n5453), .ZN(n5492) );
  NAND2_X1 U5179 ( .A1(n4591), .A2(n4398), .ZN(n5454) );
  OR2_X1 U5180 ( .A1(n5416), .A2(n5418), .ZN(n5421) );
  OR2_X1 U5181 ( .A1(n5418), .A2(n5417), .ZN(n5420) );
  OAI21_X2 U5182 ( .B1(n5373), .B2(n4597), .A(n5372), .ZN(n5422) );
  AOI21_X1 U5183 ( .B1(n4768), .B2(n4764), .A(n4763), .ZN(n4762) );
  INV_X1 U5184 ( .A(n5337), .ZN(n4763) );
  INV_X1 U5185 ( .A(n5298), .ZN(n4772) );
  INV_X1 U5186 ( .A(n5316), .ZN(n5319) );
  XNOR2_X1 U5187 ( .A(n5317), .B(SI_11_), .ZN(n5316) );
  NAND2_X1 U5188 ( .A1(n5291), .A2(n5290), .ZN(n7696) );
  NAND2_X1 U5189 ( .A1(n6768), .A2(n5272), .ZN(n5291) );
  OR2_X1 U5190 ( .A1(n5480), .A2(n8368), .ZN(n5515) );
  OR2_X1 U5191 ( .A1(n5276), .A2(n7828), .ZN(n5307) );
  NAND2_X1 U5192 ( .A1(n5968), .A2(n5962), .ZN(n5990) );
  AOI21_X1 U5193 ( .B1(n8557), .B2(n5763), .A(n5634), .ZN(n8543) );
  AOI21_X1 U5194 ( .B1(n8574), .B2(n5763), .A(n5589), .ZN(n8196) );
  AND2_X1 U5195 ( .A1(n5486), .A2(n5485), .ZN(n8283) );
  AND2_X1 U5196 ( .A1(n5615), .A2(n5614), .ZN(n8410) );
  OR2_X1 U5197 ( .A1(n8203), .A2(n5609), .ZN(n5615) );
  NAND2_X1 U5198 ( .A1(n5713), .A2(n5712), .ZN(n8564) );
  INV_X1 U5199 ( .A(n8799), .ZN(n5711) );
  NAND2_X1 U5200 ( .A1(n4846), .A2(n4844), .ZN(n8582) );
  INV_X1 U5201 ( .A(n4845), .ZN(n4844) );
  NAND2_X1 U5202 ( .A1(n8609), .A2(n4847), .ZN(n4846) );
  OAI21_X1 U5203 ( .B1(n4848), .B2(n5975), .A(n5933), .ZN(n4845) );
  AND2_X1 U5204 ( .A1(n8842), .A2(n8750), .ZN(n5706) );
  NAND2_X1 U5205 ( .A1(n4694), .A2(n5702), .ZN(n4690) );
  NAND2_X1 U5206 ( .A1(n5329), .A2(n5328), .ZN(n7893) );
  NAND2_X1 U5207 ( .A1(n6794), .A2(n4689), .ZN(n5329) );
  OR2_X1 U5208 ( .A1(n7696), .A2(n7830), .ZN(n5885) );
  AND2_X1 U5209 ( .A1(n6974), .A2(n5635), .ZN(n10015) );
  AND2_X1 U5210 ( .A1(n8799), .A2(n10096), .ZN(n4854) );
  OR2_X1 U5211 ( .A1(n6968), .A2(n5670), .ZN(n10038) );
  NAND2_X1 U5212 ( .A1(n4626), .A2(n4622), .ZN(n4619) );
  OR2_X1 U5213 ( .A1(n7048), .A2(n6617), .ZN(n6645) );
  AOI21_X1 U5214 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6813), .A(n7027), .ZN(
        n6863) );
  XNOR2_X1 U5215 ( .A(n4779), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9441) );
  OR2_X1 U5216 ( .A1(n9435), .A2(n4780), .ZN(n4779) );
  AND2_X1 U5217 ( .A1(n9437), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U5218 ( .A1(n9052), .A2(n9051), .ZN(n9449) );
  NAND2_X1 U5219 ( .A1(n9066), .A2(n9065), .ZN(n9692) );
  NAND3_X1 U5220 ( .A1(n9519), .A2(n5015), .A3(n4395), .ZN(n9470) );
  NAND2_X1 U5221 ( .A1(n9171), .A2(n4406), .ZN(n4996) );
  INV_X1 U5222 ( .A(n4994), .ZN(n4993) );
  AND2_X1 U5223 ( .A1(n6631), .A2(n6630), .ZN(n8148) );
  OR2_X1 U5224 ( .A1(n6654), .A2(n6647), .ZN(n6631) );
  NOR2_X1 U5225 ( .A1(n9316), .A2(n4963), .ZN(n4962) );
  AOI21_X1 U5226 ( .B1(n9511), .B2(n4419), .A(n4564), .ZN(n9479) );
  NAND2_X1 U5227 ( .A1(n4452), .A2(n4565), .ZN(n4564) );
  OR2_X1 U5228 ( .A1(n9725), .A2(n9517), .ZN(n9247) );
  NAND2_X1 U5229 ( .A1(n4546), .A2(n4971), .ZN(n9583) );
  NOR2_X1 U5230 ( .A1(n4972), .A2(n4430), .ZN(n4971) );
  NAND2_X1 U5231 ( .A1(n9625), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5232 ( .A1(n9625), .A2(n4973), .ZN(n4977) );
  INV_X1 U5233 ( .A(n4968), .ZN(n4967) );
  AOI21_X1 U5234 ( .B1(n4968), .B2(n9652), .A(n4966), .ZN(n4965) );
  AND2_X1 U5235 ( .A1(n8035), .A2(n9221), .ZN(n4968) );
  NAND2_X1 U5236 ( .A1(n7938), .A2(n9196), .ZN(n4673) );
  NAND2_X1 U5237 ( .A1(n6896), .A2(n6895), .ZN(n9656) );
  INV_X1 U5238 ( .A(n9633), .ZN(n9660) );
  NAND2_X1 U5239 ( .A1(n6280), .A2(n6279), .ZN(n9790) );
  NAND2_X1 U5240 ( .A1(n6364), .A2(n6039), .ZN(n6612) );
  OAI21_X1 U5241 ( .B1(n5492), .B2(n4414), .A(n5053), .ZN(n5506) );
  NAND2_X1 U5242 ( .A1(n5242), .A2(n5241), .ZN(n4545) );
  NAND2_X1 U5243 ( .A1(n8263), .A2(n4577), .ZN(n8262) );
  OR2_X1 U5244 ( .A1(n8260), .A2(n8259), .ZN(n4577) );
  NAND2_X1 U5245 ( .A1(n7062), .A2(n7063), .ZN(n7061) );
  INV_X1 U5246 ( .A(n9532), .ZN(n9725) );
  OR2_X1 U5247 ( .A1(n9939), .A2(n7114), .ZN(n9637) );
  NAND2_X1 U5248 ( .A1(n5892), .A2(n4736), .ZN(n4739) );
  AND2_X1 U5249 ( .A1(n5889), .A2(n5891), .ZN(n4736) );
  AND4_X1 U5250 ( .A1(n5882), .A2(n5939), .A3(n5881), .A4(n5880), .ZN(n5883)
         );
  AND2_X1 U5251 ( .A1(n7976), .A2(n5905), .ZN(n4526) );
  AOI21_X1 U5252 ( .B1(n9114), .B2(n9157), .A(n9652), .ZN(n4732) );
  NAND2_X1 U5253 ( .A1(n9115), .A2(n9164), .ZN(n4733) );
  INV_X1 U5254 ( .A(n7328), .ZN(n4700) );
  INV_X1 U5255 ( .A(n7557), .ZN(n4699) );
  AOI21_X1 U5256 ( .B1(n9173), .B2(n9072), .A(n9071), .ZN(n9073) );
  INV_X1 U5257 ( .A(n4598), .ZN(n4596) );
  INV_X1 U5258 ( .A(n8566), .ZN(n5940) );
  INV_X1 U5259 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5072) );
  INV_X1 U5260 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5071) );
  OAI21_X1 U5261 ( .B1(n4380), .B2(n4583), .A(n4582), .ZN(n5183) );
  NAND2_X1 U5262 ( .A1(n4380), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U5263 ( .A1(n5169), .A2(n5170), .ZN(n5173) );
  INV_X1 U5264 ( .A(n5428), .ZN(n5427) );
  NOR2_X1 U5265 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  AND2_X1 U5266 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5308) );
  OR2_X1 U5267 ( .A1(n4840), .A2(n5801), .ZN(n4839) );
  NOR2_X1 U5268 ( .A1(n4841), .A2(n4843), .ZN(n4840) );
  NAND2_X1 U5269 ( .A1(n5824), .A2(n5802), .ZN(n4653) );
  NOR2_X1 U5270 ( .A1(n5989), .A2(n5988), .ZN(n4926) );
  NAND2_X1 U5271 ( .A1(n5566), .A2(n4608), .ZN(n5607) );
  INV_X1 U5272 ( .A(n5567), .ZN(n5566) );
  OR2_X1 U5273 ( .A1(n8801), .A2(n8232), .ZN(n5933) );
  OR2_X1 U5274 ( .A1(n8822), .A2(n8283), .ZN(n5926) );
  OR2_X1 U5275 ( .A1(n8838), .A2(n8732), .ZN(n5836) );
  NOR2_X1 U5276 ( .A1(n5704), .A2(n8854), .ZN(n4937) );
  NAND2_X1 U5277 ( .A1(n5047), .A2(n4649), .ZN(n5395) );
  NAND2_X1 U5278 ( .A1(n4459), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U5279 ( .A1(n5386), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5410) );
  INV_X1 U5280 ( .A(n5388), .ZN(n5386) );
  OR2_X1 U5281 ( .A1(n5704), .A2(n8731), .ZN(n5909) );
  INV_X1 U5282 ( .A(n5307), .ZN(n5309) );
  NOR2_X1 U5283 ( .A1(n5315), .A2(n4832), .ZN(n4831) );
  INV_X1 U5284 ( .A(n5885), .ZN(n4832) );
  OR2_X1 U5285 ( .A1(n10095), .A2(n9997), .ZN(n5888) );
  OR2_X2 U5286 ( .A1(n8618), .A2(n8801), .ZN(n8601) );
  AND2_X1 U5287 ( .A1(n5406), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5288 ( .A1(n8890), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U5289 ( .A1(n5083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4824) );
  NOR2_X1 U5290 ( .A1(n6542), .A2(n10432), .ZN(n4503) );
  INV_X1 U5291 ( .A(n6856), .ZN(n4808) );
  INV_X1 U5292 ( .A(n4487), .ZN(n4807) );
  INV_X1 U5293 ( .A(n6912), .ZN(n4803) );
  INV_X1 U5294 ( .A(n4410), .ZN(n4811) );
  OAI211_X1 U5295 ( .C1(n9461), .C2(n9464), .A(n4681), .B(n9656), .ZN(n4680)
         );
  NAND2_X1 U5296 ( .A1(n9464), .A2(n4682), .ZN(n4681) );
  AND2_X1 U5297 ( .A1(n9462), .A2(n9461), .ZN(n4682) );
  AND2_X1 U5298 ( .A1(n9074), .A2(n9484), .ZN(n9312) );
  OR2_X1 U5299 ( .A1(n6582), .A2(n6581), .ZN(n6624) );
  AND2_X1 U5300 ( .A1(n9116), .A2(n4981), .ZN(n4973) );
  OR2_X1 U5301 ( .A1(n9764), .A2(n8991), .ZN(n9235) );
  AOI21_X1 U5302 ( .B1(n4672), .B2(n4671), .A(n4670), .ZN(n4665) );
  NAND2_X1 U5303 ( .A1(n4499), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6391) );
  INV_X1 U5304 ( .A(n6389), .ZN(n4499) );
  OR2_X1 U5305 ( .A1(n9774), .A2(n9043), .ZN(n9231) );
  NAND2_X1 U5306 ( .A1(n6050), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6339) );
  INV_X1 U5307 ( .A(n6315), .ZN(n6050) );
  NAND2_X1 U5308 ( .A1(n4442), .A2(n7597), .ZN(n4555) );
  INV_X1 U5309 ( .A(n4555), .ZN(n4551) );
  NAND2_X1 U5310 ( .A1(n4498), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6298) );
  INV_X1 U5311 ( .A(n6281), .ZN(n4498) );
  INV_X1 U5312 ( .A(n5002), .ZN(n5001) );
  OAI21_X1 U5313 ( .B1(n7153), .B2(n5004), .A(n5007), .ZN(n5002) );
  OR2_X1 U5314 ( .A1(n9795), .A2(n9356), .ZN(n5007) );
  NAND2_X1 U5315 ( .A1(n6049), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6256) );
  INV_X1 U5316 ( .A(n6254), .ZN(n6049) );
  AND3_X1 U5317 ( .A1(n6935), .A2(n7497), .A3(n7675), .ZN(n7138) );
  NAND2_X1 U5318 ( .A1(n4991), .A2(n4993), .ZN(n4988) );
  OR2_X1 U5319 ( .A1(n9692), .A2(n9067), .ZN(n9214) );
  INV_X1 U5320 ( .A(SI_10_), .ZN(n10365) );
  AOI21_X1 U5321 ( .B1(n4933), .B2(n4932), .A(n4480), .ZN(n4931) );
  INV_X1 U5322 ( .A(n5775), .ZN(n4932) );
  OR2_X1 U5323 ( .A1(n5596), .A2(n5595), .ZN(n5738) );
  NAND2_X1 U5324 ( .A1(n5505), .A2(n5504), .ZN(n4920) );
  NAND2_X1 U5325 ( .A1(n5490), .A2(n5475), .ZN(n5489) );
  NAND2_X1 U5326 ( .A1(n6350), .A2(n6031), .ZN(n6414) );
  INV_X1 U5327 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5328 ( .A1(n5419), .A2(n5400), .ZN(n5418) );
  NAND2_X1 U5329 ( .A1(n5337), .A2(n5323), .ZN(n5338) );
  AOI21_X1 U5330 ( .B1(n4769), .B2(n4771), .A(n4458), .ZN(n4768) );
  INV_X1 U5331 ( .A(n5054), .ZN(n4769) );
  NAND2_X1 U5332 ( .A1(n4723), .A2(n4902), .ZN(n5297) );
  AOI21_X1 U5333 ( .B1(n4904), .B2(n4906), .A(n4903), .ZN(n4902) );
  INV_X1 U5334 ( .A(n5285), .ZN(n4903) );
  INV_X1 U5335 ( .A(n5239), .ZN(n4655) );
  NOR2_X1 U5336 ( .A1(n5266), .A2(n4908), .ZN(n4907) );
  INV_X1 U5337 ( .A(n5241), .ZN(n4908) );
  NAND2_X1 U5338 ( .A1(n5235), .A2(n5062), .ZN(n4657) );
  NAND2_X1 U5339 ( .A1(n5173), .A2(n5172), .ZN(n5182) );
  OR2_X1 U5340 ( .A1(n5226), .A2(n10227), .ZN(n5257) );
  NAND2_X1 U5341 ( .A1(n5427), .A2(n4612), .ZN(n5462) );
  NAND2_X1 U5342 ( .A1(n4870), .A2(n4872), .ZN(n4866) );
  NOR2_X1 U5343 ( .A1(n8366), .A2(n4869), .ZN(n4868) );
  INV_X1 U5344 ( .A(n4870), .ZN(n4869) );
  OR2_X1 U5345 ( .A1(n5410), .A2(n10333), .ZN(n5428) );
  AOI21_X1 U5346 ( .B1(n4873), .B2(n4871), .A(n4472), .ZN(n4870) );
  AOI21_X1 U5347 ( .B1(n4862), .B2(n7710), .A(n4861), .ZN(n4860) );
  INV_X1 U5348 ( .A(n7803), .ZN(n4861) );
  INV_X1 U5349 ( .A(n7710), .ZN(n4863) );
  NAND2_X1 U5350 ( .A1(n5309), .A2(n5308), .ZN(n5330) );
  NAND2_X1 U5351 ( .A1(n8080), .A2(n8065), .ZN(n8066) );
  AND2_X1 U5352 ( .A1(n5522), .A2(n5521), .ZN(n8282) );
  AND2_X1 U5353 ( .A1(n5406), .A2(n5159), .ZN(n5174) );
  INV_X1 U5354 ( .A(n5174), .ZN(n5187) );
  OR2_X1 U5355 ( .A1(n7340), .A2(n7341), .ZN(n7338) );
  OR2_X1 U5356 ( .A1(n8512), .A2(n8513), .ZN(n4568) );
  AND2_X1 U5357 ( .A1(n5722), .A2(n4939), .ZN(n8162) );
  AND2_X1 U5358 ( .A1(n8773), .A2(n4941), .ZN(n4939) );
  AOI21_X1 U5359 ( .B1(n8777), .B2(n4408), .A(n10113), .ZN(n8550) );
  INV_X1 U5360 ( .A(n4942), .ZN(n4940) );
  NAND2_X1 U5361 ( .A1(n5953), .A2(n5954), .ZN(n8541) );
  NAND2_X1 U5362 ( .A1(n5026), .A2(n5025), .ZN(n8542) );
  AOI21_X1 U5363 ( .B1(n5028), .B2(n5030), .A(n4449), .ZN(n5025) );
  NAND2_X1 U5364 ( .A1(n5830), .A2(n8599), .ZN(n4848) );
  OR2_X1 U5365 ( .A1(n8586), .A2(n5609), .ZN(n5574) );
  INV_X1 U5366 ( .A(n4701), .ZN(n8616) );
  OAI21_X1 U5367 ( .B1(n8659), .B2(n4704), .A(n4702), .ZN(n4701) );
  OR2_X1 U5368 ( .A1(n4708), .A2(n4705), .ZN(n4704) );
  INV_X1 U5369 ( .A(n4703), .ZN(n4702) );
  NAND2_X1 U5370 ( .A1(n8641), .A2(n5929), .ZN(n8609) );
  NOR2_X1 U5371 ( .A1(n8609), .A2(n8615), .ZN(n8610) );
  AND2_X1 U5372 ( .A1(n5500), .A2(n5499), .ZN(n8638) );
  NAND2_X1 U5373 ( .A1(n4511), .A2(n4705), .ZN(n8641) );
  INV_X1 U5374 ( .A(n8635), .ZN(n4511) );
  AND2_X1 U5375 ( .A1(n5539), .A2(n5538), .ZN(n8639) );
  NAND2_X1 U5376 ( .A1(n8647), .A2(n8634), .ZN(n8628) );
  AOI21_X1 U5377 ( .B1(n4836), .B2(n4838), .A(n4835), .ZN(n4834) );
  INV_X1 U5378 ( .A(n5923), .ZN(n4835) );
  AND2_X1 U5379 ( .A1(n5721), .A2(n8650), .ZN(n8647) );
  INV_X1 U5380 ( .A(n5986), .ZN(n8653) );
  NOR2_X2 U5381 ( .A1(n8660), .A2(n8822), .ZN(n5721) );
  NAND2_X1 U5382 ( .A1(n8682), .A2(n5470), .ZN(n8683) );
  INV_X1 U5383 ( .A(n5708), .ZN(n8684) );
  AND2_X1 U5384 ( .A1(n5468), .A2(n5467), .ZN(n8695) );
  AND2_X1 U5385 ( .A1(n8681), .A2(n5918), .ZN(n8692) );
  NOR2_X1 U5386 ( .A1(n5035), .A2(n4718), .ZN(n4717) );
  AND2_X1 U5387 ( .A1(n5034), .A2(n4720), .ZN(n4719) );
  INV_X1 U5388 ( .A(n5035), .ZN(n4721) );
  INV_X1 U5389 ( .A(n8725), .ZN(n5038) );
  NAND2_X1 U5390 ( .A1(n5836), .A2(n5834), .ZN(n8711) );
  NAND2_X1 U5391 ( .A1(n5837), .A2(n8705), .ZN(n8729) );
  AND2_X1 U5392 ( .A1(n8726), .A2(n8729), .ZN(n8725) );
  OR2_X1 U5393 ( .A1(n8854), .A2(n8048), .ZN(n8745) );
  OR2_X1 U5394 ( .A1(n5365), .A2(n5351), .ZN(n5388) );
  NAND2_X1 U5395 ( .A1(n4696), .A2(n5701), .ZN(n4694) );
  NAND2_X1 U5396 ( .A1(n5031), .A2(n4697), .ZN(n4696) );
  INV_X1 U5397 ( .A(n7749), .ZN(n4697) );
  NAND2_X1 U5398 ( .A1(n4695), .A2(n5031), .ZN(n4692) );
  NOR2_X1 U5399 ( .A1(n7893), .A2(n4945), .ZN(n4944) );
  INV_X1 U5400 ( .A(n4946), .ZN(n4945) );
  AOI22_X1 U5401 ( .A1(n7287), .A2(n6718), .B1(n5582), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U5402 ( .A1(n6773), .A2(n4689), .ZN(n5305) );
  NAND2_X1 U5403 ( .A1(n7635), .A2(n5884), .ZN(n5296) );
  AND4_X1 U5404 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n7830)
         );
  OR2_X1 U5405 ( .A1(n5715), .A2(n5635), .ZN(n10000) );
  NAND2_X1 U5406 ( .A1(n10022), .A2(n10021), .ZN(n7321) );
  INV_X1 U5407 ( .A(n10020), .ZN(n9995) );
  INV_X1 U5408 ( .A(n10000), .ZN(n10017) );
  NAND2_X1 U5409 ( .A1(n8542), .A2(n8541), .ZN(n8783) );
  NAND2_X1 U5410 ( .A1(n5606), .A2(n5605), .ZN(n8788) );
  NAND2_X1 U5411 ( .A1(n8899), .A2(n4689), .ZN(n5606) );
  NAND2_X1 U5412 ( .A1(n5584), .A2(n5583), .ZN(n8793) );
  NOR2_X1 U5413 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5017) );
  OR2_X1 U5414 ( .A1(n5358), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5348) );
  NOR2_X1 U5415 ( .A1(n5187), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5416 ( .A1(n4528), .A2(n10348), .ZN(n5324) );
  INV_X1 U5417 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n10348) );
  INV_X1 U5418 ( .A(n7351), .ZN(n4887) );
  OR2_X1 U5419 ( .A1(n6432), .A2(n4624), .ZN(n4623) );
  INV_X1 U5420 ( .A(n4503), .ZN(n6567) );
  XNOR2_X1 U5421 ( .A(n6361), .B(n7129), .ZN(n6403) );
  NAND2_X1 U5422 ( .A1(n6333), .A2(n7873), .ZN(n5041) );
  INV_X1 U5423 ( .A(n6432), .ZN(n4627) );
  NAND2_X1 U5424 ( .A1(n8985), .A2(n6432), .ZN(n4620) );
  NAND2_X1 U5425 ( .A1(n6171), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6216) );
  OR2_X1 U5426 ( .A1(n6562), .A2(n6563), .ZN(n4777) );
  AND2_X1 U5427 ( .A1(n9682), .A2(n9452), .ZN(n9208) );
  AND2_X1 U5428 ( .A1(n6548), .A2(n6547), .ZN(n8963) );
  AOI21_X1 U5429 ( .B1(n9558), .B2(n6510), .A(n6495), .ZN(n9349) );
  XNOR2_X1 U5430 ( .A(n6823), .B(n6810), .ZN(n9878) );
  INV_X1 U5431 ( .A(n6862), .ZN(n4781) );
  INV_X1 U5432 ( .A(n6863), .ZN(n4782) );
  NAND2_X1 U5433 ( .A1(n6989), .A2(n4783), .ZN(n6876) );
  OR2_X1 U5434 ( .A1(n6992), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4783) );
  NOR2_X1 U5435 ( .A1(n6913), .A2(n6914), .ZN(n7006) );
  OR2_X1 U5436 ( .A1(n7006), .A2(n4796), .ZN(n4795) );
  AND2_X1 U5437 ( .A1(n7007), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U5438 ( .A1(n4795), .A2(n4794), .ZN(n4793) );
  INV_X1 U5439 ( .A(n7008), .ZN(n4794) );
  NOR2_X1 U5440 ( .A1(n7440), .A2(n7441), .ZN(n7688) );
  OR2_X1 U5441 ( .A1(n7688), .A2(n4788), .ZN(n4787) );
  AND2_X1 U5442 ( .A1(n7689), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4788) );
  AND2_X1 U5443 ( .A1(n4787), .A2(n4786), .ZN(n9374) );
  INV_X1 U5444 ( .A(n7690), .ZN(n4786) );
  NAND2_X1 U5445 ( .A1(n4801), .A2(n4479), .ZN(n4798) );
  OR2_X1 U5446 ( .A1(n9390), .A2(n4799), .ZN(n4797) );
  NAND2_X1 U5447 ( .A1(n4800), .A2(n4801), .ZN(n4799) );
  INV_X1 U5448 ( .A(n9389), .ZN(n4800) );
  NAND2_X1 U5449 ( .A1(n9519), .A2(n4395), .ZN(n8151) );
  AND2_X1 U5450 ( .A1(n9519), .A2(n5016), .ZN(n9480) );
  NAND2_X1 U5451 ( .A1(n9519), .A2(n9503), .ZN(n9498) );
  NAND2_X1 U5452 ( .A1(n4502), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U5453 ( .A1(n4998), .A2(n4557), .ZN(n4558) );
  OR2_X1 U5454 ( .A1(n9560), .A2(n9349), .ZN(n5045) );
  AND2_X1 U5455 ( .A1(n4561), .A2(n4415), .ZN(n9556) );
  NAND2_X1 U5456 ( .A1(n4562), .A2(n8021), .ZN(n4561) );
  INV_X1 U5457 ( .A(n9569), .ZN(n4562) );
  NAND2_X1 U5458 ( .A1(n9556), .A2(n9555), .ZN(n9554) );
  AND2_X1 U5459 ( .A1(n9135), .A2(n9129), .ZN(n9577) );
  INV_X1 U5460 ( .A(n4976), .ZN(n4975) );
  AND2_X1 U5461 ( .A1(n9603), .A2(n9602), .ZN(n9175) );
  NAND2_X1 U5462 ( .A1(n4539), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6417) );
  AND3_X1 U5463 ( .A1(n6375), .A2(n6374), .A3(n6373), .ZN(n9630) );
  NAND2_X1 U5464 ( .A1(n8034), .A2(n9650), .ZN(n9655) );
  NAND2_X1 U5465 ( .A1(n8011), .A2(n8012), .ZN(n4548) );
  AND2_X1 U5466 ( .A1(n4394), .A2(n9111), .ZN(n4672) );
  AND2_X1 U5467 ( .A1(n4673), .A2(n9111), .ZN(n5040) );
  AND2_X1 U5468 ( .A1(n9108), .A2(n7844), .ZN(n7845) );
  AND2_X1 U5469 ( .A1(n7842), .A2(n9100), .ZN(n9192) );
  AND2_X1 U5470 ( .A1(n9078), .A2(n9092), .ZN(n7507) );
  NAND2_X1 U5471 ( .A1(n5008), .A2(n7153), .ZN(n7503) );
  INV_X1 U5472 ( .A(n9656), .ZN(n9628) );
  NAND2_X1 U5473 ( .A1(n6580), .A2(n6579), .ZN(n9706) );
  NAND2_X1 U5474 ( .A1(n6565), .A2(n6564), .ZN(n9710) );
  NAND2_X1 U5475 ( .A1(n8902), .A2(n4377), .ZN(n6565) );
  NAND2_X1 U5476 ( .A1(n6416), .A2(n6415), .ZN(n9759) );
  INV_X1 U5477 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6055) );
  XNOR2_X1 U5478 ( .A(n5783), .B(n5782), .ZN(n9054) );
  NAND2_X1 U5479 ( .A1(n5805), .A2(n5804), .ZN(n5783) );
  NAND2_X1 U5480 ( .A1(n4935), .A2(n4933), .ZN(n5805) );
  NOR2_X1 U5481 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NOR2_X1 U5482 ( .A1(n6056), .A2(n6061), .ZN(n6062) );
  NAND2_X1 U5483 ( .A1(n6044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6040) );
  AND2_X1 U5484 ( .A1(n4959), .A2(n6021), .ZN(n4640) );
  XNOR2_X1 U5485 ( .A(n5544), .B(n5555), .ZN(n7992) );
  NOR2_X1 U5486 ( .A1(n5524), .A2(n4922), .ZN(n4921) );
  INV_X1 U5487 ( .A(n5504), .ZN(n4922) );
  OAI21_X1 U5488 ( .B1(n5506), .B2(n5505), .A(n5504), .ZN(n5525) );
  OR2_X1 U5489 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U5490 ( .A1(n4594), .A2(n4598), .ZN(n5451) );
  NAND2_X1 U5491 ( .A1(n5422), .A2(n4599), .ZN(n4594) );
  OAI21_X1 U5492 ( .B1(n6086), .B2(n6061), .A(n6087), .ZN(n6135) );
  NOR2_X1 U5493 ( .A1(n9854), .A2(n9853), .ZN(n9855) );
  NAND2_X1 U5494 ( .A1(n9858), .A2(n9859), .ZN(n9860) );
  NAND2_X1 U5495 ( .A1(n9864), .A2(n9865), .ZN(n9866) );
  INV_X1 U5496 ( .A(n8788), .ZN(n8207) );
  INV_X1 U5497 ( .A(n4875), .ZN(n4579) );
  NAND2_X1 U5498 ( .A1(n5532), .A2(n5531), .ZN(n8807) );
  NAND2_X1 U5499 ( .A1(n5460), .A2(n5459), .ZN(n8828) );
  AND2_X1 U5500 ( .A1(n7208), .A2(n7203), .ZN(n4885) );
  NAND2_X1 U5501 ( .A1(n7039), .A2(n4689), .ZN(n5409) );
  INV_X1 U5502 ( .A(n8420), .ZN(n8412) );
  AND4_X1 U5503 ( .A1(n5335), .A2(n5334), .A3(n5333), .A4(n5332), .ZN(n7969)
         );
  NAND2_X1 U5504 ( .A1(n6961), .A2(n10026), .ZN(n8386) );
  AND2_X1 U5505 ( .A1(n6976), .A2(n6972), .ZN(n8415) );
  INV_X1 U5506 ( .A(n8407), .ZN(n4543) );
  NAND2_X1 U5507 ( .A1(n8408), .A2(n8409), .ZN(n4542) );
  NAND2_X1 U5508 ( .A1(n4881), .A2(n4882), .ZN(n8408) );
  INV_X1 U5509 ( .A(n8386), .ZN(n8425) );
  OAI21_X1 U5510 ( .B1(n6001), .B2(n6000), .A(n4758), .ZN(n4642) );
  INV_X1 U5511 ( .A(n5999), .ZN(n4758) );
  XNOR2_X1 U5512 ( .A(n4923), .B(n5619), .ZN(n5992) );
  INV_X1 U5513 ( .A(n8282), .ZN(n8654) );
  INV_X1 U5514 ( .A(n8283), .ZN(n8686) );
  NAND2_X1 U5515 ( .A1(n7249), .A2(n4440), .ZN(n7236) );
  NAND2_X1 U5516 ( .A1(n7236), .A2(n7237), .ZN(n7235) );
  NOR2_X1 U5517 ( .A1(n5174), .A2(n4574), .ZN(n7234) );
  OAI21_X1 U5518 ( .B1(n5406), .B2(n4576), .A(n4575), .ZN(n4574) );
  NAND2_X1 U5519 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4576) );
  NAND2_X1 U5520 ( .A1(n8890), .A2(n5159), .ZN(n4575) );
  NAND2_X1 U5521 ( .A1(n7222), .A2(n4432), .ZN(n7062) );
  NAND2_X1 U5522 ( .A1(n8491), .A2(n8490), .ZN(n8489) );
  OAI21_X1 U5523 ( .B1(n8491), .B2(n4571), .A(n4569), .ZN(n4573) );
  INV_X1 U5524 ( .A(n4572), .ZN(n4571) );
  AOI21_X1 U5525 ( .B1(n4570), .B2(n4572), .A(n4455), .ZN(n4569) );
  NOR2_X1 U5526 ( .A1(n7363), .A2(n7364), .ZN(n7362) );
  NAND2_X1 U5527 ( .A1(n5816), .A2(n5815), .ZN(n5818) );
  NAND2_X1 U5528 ( .A1(n9049), .A2(n4689), .ZN(n5816) );
  INV_X1 U5529 ( .A(n8538), .ZN(n8539) );
  XNOR2_X1 U5530 ( .A(n4488), .B(n5950), .ZN(n8791) );
  NAND2_X1 U5531 ( .A1(n5027), .A2(n5714), .ZN(n4488) );
  INV_X1 U5532 ( .A(n8793), .ZN(n8565) );
  NAND2_X1 U5533 ( .A1(n8596), .A2(n5710), .ZN(n8580) );
  NAND2_X1 U5534 ( .A1(n5565), .A2(n5564), .ZN(n8799) );
  NAND2_X1 U5535 ( .A1(n7998), .A2(n4689), .ZN(n5565) );
  NAND2_X1 U5536 ( .A1(n8584), .A2(n8583), .ZN(n8797) );
  INV_X1 U5537 ( .A(n10026), .ZN(n10002) );
  NAND2_X1 U5538 ( .A1(n5680), .A2(n10026), .ZN(n10027) );
  AOI21_X1 U5539 ( .B1(n4774), .B2(n8911), .A(n8910), .ZN(n8912) );
  AND2_X1 U5540 ( .A1(n4774), .A2(n4393), .ZN(n6640) );
  NAND2_X1 U5541 ( .A1(n4549), .A2(n6253), .ZN(n7743) );
  NAND2_X1 U5542 ( .A1(n6249), .A2(n6578), .ZN(n4549) );
  NAND2_X1 U5543 ( .A1(n6470), .A2(n6469), .ZN(n9740) );
  INV_X1 U5544 ( .A(n4378), .ZN(n9340) );
  INV_X1 U5545 ( .A(n9208), .ZN(n9342) );
  NAND2_X1 U5546 ( .A1(n6573), .A2(n6572), .ZN(n9506) );
  OR2_X1 U5547 ( .A1(n9027), .A2(n6647), .ZN(n6573) );
  INV_X1 U5548 ( .A(n9517), .ZN(n9549) );
  AND2_X1 U5549 ( .A1(n6278), .A2(n6293), .ZN(n7097) );
  NAND2_X1 U5550 ( .A1(n9441), .A2(n9918), .ZN(n9444) );
  NOR2_X1 U5551 ( .A1(n9471), .A2(n9683), .ZN(n9450) );
  INV_X1 U5552 ( .A(n9477), .ZN(n4495) );
  OAI21_X1 U5553 ( .B1(n8154), .B2(n4684), .A(n4674), .ZN(n9469) );
  AOI21_X1 U5554 ( .B1(n8154), .B2(n4677), .A(n4675), .ZN(n4674) );
  INV_X1 U5555 ( .A(n8156), .ZN(n8157) );
  AOI21_X1 U5556 ( .B1(n9348), .B2(n9660), .A(n8155), .ZN(n8156) );
  INV_X1 U5557 ( .A(n4989), .ZN(n8149) );
  INV_X1 U5558 ( .A(n4996), .ZN(n4990) );
  AOI22_X1 U5559 ( .A1(n9489), .A2(n9660), .B1(n9659), .B2(n9488), .ZN(n9490)
         );
  INV_X1 U5560 ( .A(n9487), .ZN(n4566) );
  NAND2_X1 U5561 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5562 ( .A1(n9564), .A2(n9659), .ZN(n4537) );
  AND2_X1 U5563 ( .A1(n6525), .A2(n6524), .ZN(n9532) );
  INV_X1 U5564 ( .A(n9671), .ZN(n9635) );
  AND2_X1 U5565 ( .A1(n7131), .A2(n7118), .ZN(n9671) );
  AND2_X1 U5566 ( .A1(n7131), .A2(n7121), .ZN(n9600) );
  OR2_X1 U5567 ( .A1(n9724), .A2(n9962), .ZN(n4516) );
  XNOR2_X1 U5568 ( .A(n9866), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(n10476) );
  OAI21_X1 U5569 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10148), .ZN(n10472) );
  OAI22_X1 U5570 ( .A1(n5852), .A2(n5939), .B1(n5851), .B2(n5865), .ZN(n5860)
         );
  AOI21_X1 U5571 ( .B1(n5892), .B2(n5891), .A(n5883), .ZN(n4740) );
  AND3_X1 U5572 ( .A1(n4739), .A2(n5903), .A3(n4738), .ZN(n4737) );
  NAND2_X1 U5573 ( .A1(n9091), .A2(n9226), .ZN(n9096) );
  NOR2_X1 U5574 ( .A1(n4760), .A2(n5469), .ZN(n4759) );
  INV_X1 U5575 ( .A(n5913), .ZN(n4760) );
  AND2_X1 U5576 ( .A1(n9094), .A2(n9078), .ZN(n9089) );
  AND2_X1 U5577 ( .A1(n5926), .A2(n5925), .ZN(n4755) );
  INV_X1 U5578 ( .A(n5928), .ZN(n4754) );
  AND2_X1 U5579 ( .A1(n5831), .A2(n5044), .ZN(n5832) );
  NAND2_X1 U5580 ( .A1(n9119), .A2(n9175), .ZN(n4729) );
  AND2_X1 U5581 ( .A1(n9090), .A2(n9089), .ZN(n9226) );
  NOR2_X1 U5582 ( .A1(n10022), .A2(n4698), .ZN(n5980) );
  INV_X1 U5583 ( .A(n4921), .ZN(n4917) );
  INV_X1 U5584 ( .A(n5541), .ZN(n4916) );
  INV_X1 U5585 ( .A(n5172), .ZN(n4646) );
  INV_X1 U5586 ( .A(n5184), .ZN(n4648) );
  INV_X1 U5587 ( .A(n4734), .ZN(n4534) );
  AOI21_X1 U5588 ( .B1(n9140), .B2(n9157), .A(n9514), .ZN(n4734) );
  NOR2_X1 U5589 ( .A1(n9141), .A2(n4533), .ZN(n4532) );
  INV_X1 U5590 ( .A(n9142), .ZN(n4533) );
  NAND2_X1 U5591 ( .A1(n5558), .A2(n5557), .ZN(n5737) );
  AND2_X1 U5592 ( .A1(n4912), .A2(n5557), .ZN(n4585) );
  NOR2_X1 U5593 ( .A1(n4919), .A2(n4913), .ZN(n4912) );
  INV_X1 U5594 ( .A(n5053), .ZN(n4913) );
  INV_X1 U5595 ( .A(n4910), .ZN(n4909) );
  OAI21_X1 U5596 ( .B1(n4919), .B2(n4911), .A(n4915), .ZN(n4910) );
  NAND2_X1 U5597 ( .A1(n4414), .A2(n5053), .ZN(n4911) );
  AOI21_X1 U5598 ( .B1(n4917), .B2(n4918), .A(n4916), .ZN(n4915) );
  NAND2_X1 U5599 ( .A1(n5508), .A2(n5507), .ZN(n5523) );
  NAND2_X1 U5600 ( .A1(n4597), .A2(n5372), .ZN(n4590) );
  AOI21_X1 U5601 ( .B1(n4600), .B2(n4598), .A(n5450), .ZN(n4595) );
  NAND2_X1 U5602 ( .A1(n5373), .A2(n4592), .ZN(n4591) );
  NOR2_X1 U5603 ( .A1(n4596), .A2(n4593), .ZN(n4592) );
  INV_X1 U5604 ( .A(n5372), .ZN(n4593) );
  INV_X1 U5605 ( .A(n5338), .ZN(n4767) );
  NOR2_X1 U5606 ( .A1(n4771), .A2(n5338), .ZN(n4764) );
  NAND2_X1 U5607 ( .A1(n5342), .A2(n5341), .ZN(n5345) );
  INV_X1 U5608 ( .A(n4905), .ZN(n4904) );
  OAI21_X1 U5609 ( .B1(n4907), .B2(n4906), .A(n5055), .ZN(n4905) );
  XNOR2_X1 U5610 ( .A(n10070), .B(n7176), .ZN(n7189) );
  NOR2_X1 U5611 ( .A1(n8167), .A2(n4874), .ZN(n4873) );
  INV_X1 U5612 ( .A(n8070), .ZN(n4874) );
  NAND2_X1 U5613 ( .A1(n8197), .A2(n8189), .ZN(n8200) );
  OR2_X1 U5614 ( .A1(n8289), .A2(n8288), .ZN(n4883) );
  NOR2_X1 U5615 ( .A1(n5946), .A2(n5939), .ZN(n4745) );
  NOR2_X1 U5616 ( .A1(n4841), .A2(n4448), .ZN(n4742) );
  NAND2_X1 U5617 ( .A1(n5952), .A2(n5939), .ZN(n4606) );
  NAND2_X1 U5618 ( .A1(n5950), .A2(n5949), .ZN(n4743) );
  NOR2_X1 U5619 ( .A1(n8777), .A2(n4942), .ZN(n4941) );
  NOR2_X1 U5620 ( .A1(n8411), .A2(n4609), .ZN(n4608) );
  NAND2_X1 U5621 ( .A1(n8207), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U5622 ( .A1(n8543), .A2(n8258), .ZN(n5954) );
  INV_X1 U5623 ( .A(n5714), .ZN(n5030) );
  INV_X1 U5624 ( .A(n5029), .ZN(n5028) );
  OAI21_X1 U5625 ( .B1(n5988), .B2(n5030), .A(n5989), .ZN(n5029) );
  OR2_X1 U5626 ( .A1(n8793), .A2(n8196), .ZN(n5947) );
  AOI21_X1 U5627 ( .B1(n8599), .B2(n5710), .A(n4433), .ZN(n5033) );
  INV_X1 U5628 ( .A(n4848), .ZN(n4847) );
  INV_X1 U5629 ( .A(n5515), .ZN(n5514) );
  OR2_X1 U5630 ( .A1(n8807), .A2(n8639), .ZN(n5827) );
  OAI21_X1 U5631 ( .B1(n5470), .B2(n4838), .A(n5926), .ZN(n4837) );
  AND2_X1 U5632 ( .A1(n4717), .A2(n4722), .ZN(n4715) );
  INV_X1 U5633 ( .A(n4827), .ZN(n4826) );
  OAI21_X1 U5634 ( .B1(n5336), .B2(n4828), .A(n5891), .ZN(n4827) );
  OR2_X1 U5635 ( .A1(n4831), .A2(n4829), .ZN(n4828) );
  INV_X1 U5636 ( .A(n5881), .ZN(n4829) );
  NOR2_X1 U5637 ( .A1(n7696), .A2(n10095), .ZN(n4946) );
  NAND2_X1 U5638 ( .A1(n5255), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5276) );
  INV_X1 U5639 ( .A(n5257), .ZN(n5255) );
  INV_X1 U5640 ( .A(n10074), .ZN(n5217) );
  INV_X1 U5641 ( .A(n5195), .ZN(n4607) );
  XNOR2_X1 U5642 ( .A(n10074), .B(n8447), .ZN(n5216) );
  NAND2_X1 U5643 ( .A1(n5682), .A2(n10051), .ZN(n5853) );
  INV_X1 U5644 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4686) );
  INV_X1 U5645 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4685) );
  OR2_X1 U5646 ( .A1(n5347), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5358) );
  OR2_X1 U5647 ( .A1(n5324), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5248) );
  INV_X1 U5648 ( .A(n4635), .ZN(n4630) );
  NAND2_X1 U5649 ( .A1(n8975), .A2(n8971), .ZN(n4778) );
  AND3_X1 U5650 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U5651 ( .A1(n6510), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6110) );
  AND2_X1 U5652 ( .A1(n9375), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4785) );
  INV_X1 U5653 ( .A(n9414), .ZN(n4801) );
  NOR2_X1 U5654 ( .A1(n9710), .A2(n9715), .ZN(n5016) );
  NAND2_X1 U5655 ( .A1(n9504), .A2(n4412), .ZN(n4565) );
  AND2_X1 U5656 ( .A1(n4948), .A2(n4660), .ZN(n4659) );
  NOR2_X1 U5657 ( .A1(n4664), .A2(n4661), .ZN(n4660) );
  INV_X1 U5658 ( .A(n9247), .ZN(n4664) );
  INV_X1 U5659 ( .A(n9548), .ZN(n4661) );
  NAND2_X1 U5660 ( .A1(n9247), .A2(n4663), .ZN(n4662) );
  INV_X1 U5661 ( .A(n9137), .ZN(n4663) );
  NOR2_X1 U5662 ( .A1(n6508), .A2(n6052), .ZN(n4502) );
  AND2_X1 U5663 ( .A1(n4415), .A2(n4559), .ZN(n4557) );
  INV_X1 U5664 ( .A(n8021), .ZN(n4559) );
  AND2_X1 U5665 ( .A1(n4998), .A2(n4415), .ZN(n4560) );
  AOI21_X1 U5666 ( .B1(n4998), .B2(n5000), .A(n4443), .ZN(n4997) );
  INV_X1 U5667 ( .A(n4502), .ZN(n6526) );
  NAND2_X1 U5668 ( .A1(n9740), .A2(n9596), .ZN(n8021) );
  NAND2_X1 U5669 ( .A1(n6051), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6471) );
  INV_X1 U5670 ( .A(n6457), .ZN(n6051) );
  AND2_X1 U5671 ( .A1(n4973), .A2(n9174), .ZN(n4547) );
  AND2_X1 U5672 ( .A1(n4976), .A2(n9174), .ZN(n4972) );
  NAND2_X1 U5673 ( .A1(n4501), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6457) );
  NOR2_X1 U5674 ( .A1(n6417), .A2(n8989), .ZN(n4501) );
  INV_X1 U5675 ( .A(n9235), .ZN(n4966) );
  NOR2_X1 U5676 ( .A1(n6391), .A2(n6370), .ZN(n4539) );
  NAND2_X1 U5677 ( .A1(n4500), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6389) );
  INV_X1 U5678 ( .A(n6339), .ZN(n4500) );
  NOR2_X1 U5679 ( .A1(n9779), .A2(n7792), .ZN(n5012) );
  NAND2_X1 U5680 ( .A1(n4497), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6315) );
  INV_X1 U5681 ( .A(n6298), .ZN(n4497) );
  NAND2_X1 U5682 ( .A1(n4535), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6281) );
  INV_X1 U5683 ( .A(n6256), .ZN(n4535) );
  NAND2_X1 U5684 ( .A1(n6048), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6254) );
  INV_X1 U5685 ( .A(n6216), .ZN(n6048) );
  AND2_X1 U5686 ( .A1(n6084), .A2(n9281), .ZN(n6890) );
  INV_X1 U5687 ( .A(SI_14_), .ZN(n10337) );
  INV_X1 U5688 ( .A(SI_12_), .ZN(n10211) );
  NOR2_X1 U5689 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6064) );
  INV_X1 U5690 ( .A(n4961), .ZN(n4958) );
  INV_X1 U5691 ( .A(n6019), .ZN(n4957) );
  NAND2_X1 U5692 ( .A1(n4589), .A2(n4909), .ZN(n5558) );
  NAND2_X1 U5693 ( .A1(n5492), .A2(n4912), .ZN(n4589) );
  NAND2_X1 U5694 ( .A1(n6037), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U5695 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n4896) );
  NAND2_X1 U5696 ( .A1(n5375), .A2(n5374), .ZN(n5417) );
  AND3_X1 U5697 ( .A1(n4420), .A2(n4955), .A3(n4959), .ZN(n6364) );
  INV_X1 U5698 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U5699 ( .B1(n4380), .B2(n5156), .A(n4489), .ZN(n5171) );
  NAND2_X1 U5700 ( .A1(n4380), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4489) );
  INV_X1 U5701 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5095) );
  INV_X1 U5702 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5096) );
  INV_X1 U5703 ( .A(n8200), .ZN(n4876) );
  INV_X1 U5704 ( .A(n4883), .ZN(n4877) );
  NOR2_X1 U5705 ( .A1(n8409), .A2(n4880), .ZN(n4879) );
  INV_X1 U5706 ( .A(n4882), .ZN(n4880) );
  INV_X1 U5707 ( .A(n4879), .ZN(n4878) );
  AND2_X1 U5708 ( .A1(n8326), .A2(n8297), .ZN(n8300) );
  NAND2_X1 U5709 ( .A1(n5427), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5442) );
  CLKBUF_X1 U5710 ( .A(n8217), .Z(n8326) );
  AND2_X1 U5711 ( .A1(n4612), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5712 ( .A1(n5309), .A2(n4603), .ZN(n5363) );
  XNOR2_X1 U5713 ( .A(n8190), .B(n10051), .ZN(n7173) );
  NAND2_X1 U5714 ( .A1(n8289), .A2(n8288), .ZN(n4882) );
  AOI21_X1 U5715 ( .B1(n5757), .B2(n4425), .A(n4652), .ZN(n5819) );
  NAND2_X1 U5716 ( .A1(n4839), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U5717 ( .A1(n4930), .A2(n4924), .ZN(n4923) );
  INV_X1 U5718 ( .A(n5991), .ZN(n4930) );
  NOR2_X1 U5719 ( .A1(n5990), .A2(n4925), .ZN(n4924) );
  AND2_X1 U5720 ( .A1(n5554), .A2(n5553), .ZN(n8232) );
  AND2_X1 U5721 ( .A1(n5449), .A2(n5448), .ZN(n8331) );
  AND3_X1 U5722 ( .A1(n5414), .A2(n5413), .A3(n5412), .ZN(n8332) );
  NAND2_X1 U5723 ( .A1(n7229), .A2(n7230), .ZN(n7228) );
  NAND2_X1 U5724 ( .A1(n7257), .A2(n7258), .ZN(n7256) );
  NAND2_X1 U5725 ( .A1(n7056), .A2(n7057), .ZN(n7055) );
  INV_X1 U5726 ( .A(n8490), .ZN(n4570) );
  NOR2_X1 U5727 ( .A1(n7283), .A2(n4819), .ZN(n4572) );
  NAND2_X1 U5728 ( .A1(n7338), .A2(n6709), .ZN(n7368) );
  NOR2_X1 U5729 ( .A1(n7362), .A2(n4820), .ZN(n7482) );
  NOR2_X1 U5730 ( .A1(n6710), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4820) );
  OAI22_X1 U5731 ( .A1(n7482), .A2(n7481), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7483), .ZN(n6682) );
  XNOR2_X1 U5732 ( .A(n6713), .B(n7767), .ZN(n7764) );
  NAND2_X1 U5733 ( .A1(n4568), .A2(n6672), .ZN(n4817) );
  OAI21_X1 U5734 ( .B1(n8509), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8502), .ZN(
        n6716) );
  NOR2_X1 U5735 ( .A1(n8104), .A2(n4815), .ZN(n8105) );
  AND2_X1 U5736 ( .A1(n8109), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U5737 ( .A1(n5947), .A2(n5944), .ZN(n5988) );
  NAND2_X1 U5738 ( .A1(n8793), .A2(n8196), .ZN(n5944) );
  OR2_X1 U5739 ( .A1(n8799), .A2(n8592), .ZN(n8566) );
  AND2_X1 U5740 ( .A1(n5607), .A2(n5586), .ZN(n8574) );
  INV_X1 U5741 ( .A(n5988), .ZN(n8568) );
  NAND2_X1 U5742 ( .A1(n5514), .A2(n4601), .ZN(n5567) );
  AND2_X1 U5743 ( .A1(n4404), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n4601) );
  OR2_X1 U5744 ( .A1(n8620), .A2(n8639), .ZN(n5046) );
  NAND2_X1 U5745 ( .A1(n4688), .A2(n8591), .ZN(n8596) );
  INV_X1 U5746 ( .A(n8598), .ZN(n4688) );
  NAND2_X1 U5747 ( .A1(n5514), .A2(n5513), .ZN(n5533) );
  NAND2_X1 U5748 ( .A1(n5514), .A2(n4404), .ZN(n5547) );
  AOI21_X1 U5749 ( .B1(n4707), .B2(n4709), .A(n4446), .ZN(n4706) );
  INV_X1 U5750 ( .A(n8665), .ZN(n4707) );
  INV_X1 U5751 ( .A(n4709), .ZN(n4708) );
  CLKBUF_X1 U5752 ( .A(n8703), .Z(n8704) );
  AND3_X1 U5753 ( .A1(n5392), .A2(n5391), .A3(n5390), .ZN(n8731) );
  AND2_X1 U5754 ( .A1(n7985), .A2(n7989), .ZN(n8758) );
  NOR2_X1 U5755 ( .A1(n4604), .A2(n5362), .ZN(n4602) );
  NAND2_X1 U5756 ( .A1(n4825), .A2(n5881), .ZN(n7857) );
  NAND2_X1 U5757 ( .A1(n5296), .A2(n4831), .ZN(n4825) );
  AND2_X1 U5758 ( .A1(n7624), .A2(n4946), .ZN(n10007) );
  NAND2_X1 U5759 ( .A1(n10007), .A2(n10112), .ZN(n7866) );
  AND4_X1 U5760 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n7634)
         );
  NAND2_X1 U5761 ( .A1(n5888), .A2(n9993), .ZN(n7637) );
  AND4_X1 U5762 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n9997)
         );
  NAND2_X1 U5763 ( .A1(n4607), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5209) );
  AND4_X1 U5764 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n8391)
         );
  INV_X1 U5765 ( .A(n5216), .ZN(n7561) );
  NAND2_X1 U5766 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5195) );
  NOR2_X2 U5767 ( .A1(n7590), .A2(n7534), .ZN(n10023) );
  NAND2_X1 U5768 ( .A1(n7529), .A2(n5684), .ZN(n10021) );
  NAND2_X1 U5769 ( .A1(n10051), .A2(n10046), .ZN(n7590) );
  NAND2_X1 U5770 ( .A1(n7023), .A2(n4689), .ZN(n5383) );
  NAND2_X1 U5771 ( .A1(n5361), .A2(n5360), .ZN(n8858) );
  NAND2_X1 U5772 ( .A1(n6798), .A2(n4689), .ZN(n5361) );
  INV_X1 U5773 ( .A(n10096), .ZN(n10111) );
  INV_X1 U5774 ( .A(n6955), .ZN(n6002) );
  NOR2_X1 U5775 ( .A1(n5771), .A2(n5770), .ZN(n6003) );
  AND2_X1 U5776 ( .A1(n8904), .A2(n5663), .ZN(n10037) );
  XNOR2_X1 U5777 ( .A(n5088), .B(n5087), .ZN(n5090) );
  NAND2_X1 U5778 ( .A1(n5086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5779 ( .A1(n4746), .A2(n4439), .ZN(n5105) );
  NOR2_X1 U5780 ( .A1(n5648), .A2(n5647), .ZN(n5651) );
  OR2_X1 U5781 ( .A1(n5248), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5250) );
  NOR2_X1 U5782 ( .A1(n5041), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5783 ( .A1(n4629), .A2(n4628), .ZN(n4633) );
  INV_X1 U5784 ( .A(n7814), .ZN(n4638) );
  NAND2_X1 U5785 ( .A1(n4615), .A2(n9007), .ZN(n8094) );
  NAND2_X1 U5786 ( .A1(n9006), .A2(n9008), .ZN(n4615) );
  NAND2_X1 U5787 ( .A1(n4888), .A2(n7351), .ZN(n7717) );
  INV_X1 U5788 ( .A(n7457), .ZN(n7049) );
  OR2_X1 U5789 ( .A1(n6471), .A2(n10321), .ZN(n6508) );
  NAND2_X1 U5790 ( .A1(n6403), .A2(n6404), .ZN(n8975) );
  AND2_X1 U5791 ( .A1(n7015), .A2(n6131), .ZN(n4890) );
  AND2_X1 U5792 ( .A1(n7087), .A2(n6170), .ZN(n7571) );
  AND2_X1 U5793 ( .A1(n6184), .A2(n6183), .ZN(n7572) );
  NAND2_X1 U5794 ( .A1(n4726), .A2(n4473), .ZN(n4725) );
  INV_X1 U5795 ( .A(n9276), .ZN(n4726) );
  OAI21_X1 U5796 ( .B1(n6865), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6815), .ZN(
        n6862) );
  NAND2_X1 U5797 ( .A1(n4784), .A2(n4421), .ZN(n6989) );
  AOI21_X1 U5798 ( .B1(n4806), .B2(n4804), .A(n4803), .ZN(n4802) );
  AOI21_X1 U5799 ( .B1(n4810), .B2(n4808), .A(n4807), .ZN(n4806) );
  AND2_X1 U5800 ( .A1(n4793), .A2(n4792), .ZN(n7098) );
  NAND2_X1 U5801 ( .A1(n7097), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4792) );
  AND2_X1 U5802 ( .A1(n4797), .A2(n4485), .ZN(n9422) );
  NOR2_X1 U5803 ( .A1(n4438), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U5804 ( .A1(n4679), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5805 ( .A1(n4683), .A2(n4678), .ZN(n4676) );
  INV_X1 U5806 ( .A(n4680), .ZN(n4679) );
  AND2_X1 U5807 ( .A1(n6624), .A2(n6583), .ZN(n8914) );
  OR2_X1 U5808 ( .A1(n9710), .A2(n9506), .ZN(n9171) );
  NAND2_X1 U5809 ( .A1(n9172), .A2(n9171), .ZN(n9487) );
  NAND2_X1 U5810 ( .A1(n6053), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6542) );
  INV_X1 U5811 ( .A(n6540), .ZN(n6053) );
  AND2_X1 U5812 ( .A1(n6075), .A2(n6074), .ZN(n9518) );
  NAND2_X1 U5813 ( .A1(n8024), .A2(n9660), .ZN(n4538) );
  NOR2_X1 U5814 ( .A1(n9740), .A2(n9736), .ZN(n5014) );
  NAND2_X1 U5815 ( .A1(n5013), .A2(n9585), .ZN(n5056) );
  NOR2_X1 U5816 ( .A1(n9745), .A2(n9740), .ZN(n5013) );
  NAND2_X1 U5817 ( .A1(n9585), .A2(n9592), .ZN(n9586) );
  INV_X1 U5818 ( .A(n4501), .ZN(n6440) );
  INV_X1 U5819 ( .A(n4539), .ZN(n6372) );
  NOR2_X2 U5820 ( .A1(n9668), .A2(n9764), .ZN(n9634) );
  OAI21_X1 U5821 ( .B1(n7938), .B2(n4666), .A(n4665), .ZN(n9653) );
  INV_X1 U5822 ( .A(n4672), .ZN(n4666) );
  NAND2_X1 U5823 ( .A1(n7605), .A2(n5012), .ZN(n7850) );
  INV_X1 U5824 ( .A(n4554), .ZN(n4553) );
  OAI21_X1 U5825 ( .B1(n4555), .B2(n9176), .A(n7770), .ZN(n4554) );
  NAND2_X1 U5826 ( .A1(n7605), .A2(n9783), .ZN(n7776) );
  NOR2_X2 U5827 ( .A1(n5060), .A2(n9795), .ZN(n7523) );
  AND4_X1 U5828 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n7517)
         );
  AND4_X1 U5829 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n7788)
         );
  NAND2_X1 U5830 ( .A1(n7743), .A2(n7517), .ZN(n9087) );
  AND2_X1 U5831 ( .A1(n9090), .A2(n9087), .ZN(n9186) );
  AND2_X1 U5832 ( .A1(n5010), .A2(n9966), .ZN(n5009) );
  NAND2_X1 U5833 ( .A1(n7138), .A2(n9966), .ZN(n7428) );
  NAND2_X1 U5834 ( .A1(n6935), .A2(n7675), .ZN(n7676) );
  NAND2_X1 U5835 ( .A1(n6934), .A2(n6933), .ZN(n7670) );
  INV_X1 U5836 ( .A(n9179), .ZN(n6933) );
  CLKBUF_X1 U5837 ( .A(n7666), .Z(n9270) );
  AND2_X1 U5838 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  INV_X1 U5839 ( .A(n4986), .ZN(n9696) );
  NAND2_X1 U5840 ( .A1(n4988), .A2(n4397), .ZN(n4987) );
  OR2_X1 U5841 ( .A1(n7120), .A2(n9340), .ZN(n9944) );
  NAND2_X1 U5842 ( .A1(n6783), .A2(n4969), .ZN(n6160) );
  NOR2_X1 U5843 ( .A1(n5598), .A2(n4970), .ZN(n4969) );
  AND2_X1 U5844 ( .A1(n6804), .A2(n7119), .ZN(n9934) );
  OR2_X1 U5845 ( .A1(n9157), .A2(n9340), .ZN(n9939) );
  NOR2_X1 U5846 ( .A1(n7047), .A2(n9826), .ZN(n7113) );
  XNOR2_X1 U5847 ( .A(n5814), .B(n5813), .ZN(n9049) );
  XNOR2_X1 U5848 ( .A(n5796), .B(n5798), .ZN(n9063) );
  NAND2_X1 U5849 ( .A1(n4935), .A2(n5779), .ZN(n5796) );
  XNOR2_X1 U5850 ( .A(n5776), .B(n5775), .ZN(n8004) );
  XNOR2_X1 U5851 ( .A(n5604), .B(n5603), .ZN(n8899) );
  NAND2_X1 U5852 ( .A1(n5597), .A2(n5738), .ZN(n5604) );
  OR2_X1 U5853 ( .A1(n5592), .A2(n5733), .ZN(n5597) );
  XNOR2_X1 U5854 ( .A(n5581), .B(n5580), .ZN(n8902) );
  NAND2_X1 U5855 ( .A1(n5575), .A2(n5594), .ZN(n5581) );
  OR2_X1 U5856 ( .A1(n5592), .A2(n5591), .ZN(n5575) );
  XNOR2_X1 U5857 ( .A(n5592), .B(n5591), .ZN(n7998) );
  XNOR2_X1 U5858 ( .A(n5477), .B(n5476), .ZN(n7648) );
  INV_X1 U5859 ( .A(n6414), .ZN(n6033) );
  OAI21_X1 U5860 ( .B1(n5422), .B2(n5421), .A(n5058), .ZN(n5436) );
  XNOR2_X1 U5861 ( .A(n5339), .B(n5338), .ZN(n6794) );
  OAI21_X1 U5862 ( .B1(n5297), .B2(n4770), .A(n4768), .ZN(n5339) );
  NAND2_X1 U5863 ( .A1(n4773), .A2(n5298), .ZN(n5320) );
  NAND2_X1 U5864 ( .A1(n5297), .A2(n5054), .ZN(n4773) );
  XNOR2_X1 U5865 ( .A(n5297), .B(n5054), .ZN(n6768) );
  OAI21_X1 U5866 ( .B1(n4657), .B2(n4656), .A(n4654), .ZN(n5284) );
  INV_X1 U5867 ( .A(n4907), .ZN(n4656) );
  AOI21_X1 U5868 ( .B1(n4907), .B2(n4655), .A(n4906), .ZN(n4654) );
  OR2_X1 U5869 ( .A1(n6310), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U5870 ( .A1(n4647), .A2(n5184), .ZN(n5202) );
  NAND2_X1 U5871 ( .A1(n5182), .A2(n5181), .ZN(n4647) );
  AND2_X1 U5872 ( .A1(n6008), .A2(n6086), .ZN(n6154) );
  NOR2_X1 U5873 ( .A1(n10467), .A2(n9856), .ZN(n9857) );
  NAND2_X1 U5874 ( .A1(n9861), .A2(n9862), .ZN(n9863) );
  INV_X1 U5875 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10227) );
  AND2_X1 U5876 ( .A1(n8396), .A2(n7203), .ZN(n7209) );
  NAND2_X1 U5877 ( .A1(n6846), .A2(n4689), .ZN(n5350) );
  NAND2_X1 U5878 ( .A1(n8083), .A2(n8070), .ZN(n8168) );
  AND2_X1 U5879 ( .A1(n8548), .A2(n5630), .ZN(n8557) );
  NAND2_X1 U5880 ( .A1(n6249), .A2(n5272), .ZN(n5253) );
  AND2_X1 U5881 ( .A1(n8415), .A2(n10017), .ZN(n8421) );
  INV_X1 U5882 ( .A(n4865), .ZN(n4864) );
  OAI21_X1 U5883 ( .B1(n8366), .B2(n4866), .A(n8173), .ZN(n4865) );
  AND4_X1 U5884 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n9999)
         );
  AND2_X1 U5885 ( .A1(n7197), .A2(n7192), .ZN(n4884) );
  NAND2_X1 U5886 ( .A1(n8358), .A2(n7192), .ZN(n8316) );
  AND2_X1 U5887 ( .A1(n8065), .A2(n8059), .ZN(n8330) );
  NAND2_X1 U5888 ( .A1(n5546), .A2(n5545), .ZN(n8801) );
  NAND2_X1 U5889 ( .A1(n7824), .A2(n7822), .ZN(n7827) );
  OAI21_X1 U5890 ( .B1(n8066), .B2(n4872), .A(n4870), .ZN(n8367) );
  AND4_X1 U5891 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n8048)
         );
  INV_X1 U5892 ( .A(n8422), .ZN(n8383) );
  INV_X1 U5893 ( .A(n8421), .ZN(n8392) );
  NAND2_X1 U5894 ( .A1(n5512), .A2(n5511), .ZN(n8812) );
  NAND2_X1 U5895 ( .A1(n4859), .A2(n7805), .ZN(n4858) );
  NAND2_X1 U5896 ( .A1(n4860), .A2(n4863), .ZN(n4859) );
  AND2_X1 U5897 ( .A1(n8121), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8420) );
  NAND2_X1 U5898 ( .A1(n7235), .A2(n4436), .ZN(n7278) );
  NAND2_X1 U5899 ( .A1(n7278), .A2(n7279), .ZN(n7277) );
  NAND2_X1 U5900 ( .A1(n7264), .A2(n7265), .ZN(n7263) );
  NAND2_X1 U5901 ( .A1(n7263), .A2(n4567), .ZN(n7223) );
  NAND2_X1 U5902 ( .A1(n7262), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5903 ( .A1(n7223), .A2(n7224), .ZN(n7222) );
  NAND2_X1 U5904 ( .A1(n7061), .A2(n4437), .ZN(n8470) );
  NAND2_X1 U5905 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  NAND2_X1 U5906 ( .A1(n8484), .A2(n8485), .ZN(n8483) );
  NAND2_X1 U5907 ( .A1(n8489), .A2(n4818), .ZN(n7282) );
  NAND2_X1 U5908 ( .A1(n7290), .A2(n7289), .ZN(n7288) );
  NAND2_X1 U5909 ( .A1(n7342), .A2(n4474), .ZN(n7363) );
  INV_X1 U5910 ( .A(n4568), .ZN(n8511) );
  AND2_X1 U5911 ( .A1(n4817), .A2(n4816), .ZN(n8104) );
  INV_X1 U5912 ( .A(n6689), .ZN(n4816) );
  INV_X1 U5913 ( .A(n4817), .ZN(n6690) );
  INV_X1 U5914 ( .A(n9984), .ZN(n9978) );
  AND2_X1 U5915 ( .A1(n6721), .A2(n6720), .ZN(n8522) );
  INV_X1 U5916 ( .A(n5818), .ZN(n8161) );
  OR2_X1 U5917 ( .A1(n5629), .A2(n5628), .ZN(n8548) );
  XNOR2_X1 U5918 ( .A(n8542), .B(n8541), .ZN(n8556) );
  OR2_X1 U5919 ( .A1(n8610), .A2(n4848), .ZN(n8594) );
  CLKBUF_X1 U5920 ( .A(n8635), .Z(n8636) );
  INV_X1 U5921 ( .A(n8812), .ZN(n8634) );
  CLKBUF_X1 U5922 ( .A(n8651), .Z(n8652) );
  INV_X1 U5923 ( .A(n5721), .ZN(n8661) );
  AND2_X1 U5924 ( .A1(n4710), .A2(n4711), .ZN(n8646) );
  NAND2_X1 U5925 ( .A1(n8659), .A2(n8665), .ZN(n4710) );
  NAND2_X1 U5926 ( .A1(n8683), .A2(n5922), .ZN(n8666) );
  NAND2_X1 U5927 ( .A1(n4719), .A2(n4716), .ZN(n8691) );
  NAND2_X1 U5928 ( .A1(n8752), .A2(n4717), .ZN(n4716) );
  NAND2_X1 U5929 ( .A1(n5038), .A2(n4721), .ZN(n8710) );
  NAND2_X1 U5930 ( .A1(n4693), .A2(n4692), .ZN(n7926) );
  INV_X1 U5931 ( .A(n4694), .ZN(n4693) );
  INV_X1 U5932 ( .A(n10027), .ZN(n8766) );
  NAND2_X1 U5933 ( .A1(n5296), .A2(n5885), .ZN(n7746) );
  NAND2_X1 U5934 ( .A1(n7374), .A2(n5023), .ZN(n5022) );
  AND2_X1 U5935 ( .A1(n7557), .A2(n5063), .ZN(n5023) );
  NAND2_X1 U5936 ( .A1(n5158), .A2(n5272), .ZN(n5162) );
  NAND2_X1 U5937 ( .A1(n6717), .A2(n5679), .ZN(n10026) );
  INV_X1 U5938 ( .A(n10051), .ZN(n5123) );
  INV_X1 U5939 ( .A(n8763), .ZN(n10034) );
  AND2_X2 U5940 ( .A1(n6003), .A2(n6955), .ZN(n10142) );
  AOI21_X1 U5941 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(n8784) );
  NOR2_X1 U5942 ( .A1(n8787), .A2(n4508), .ZN(n8789) );
  AND2_X1 U5943 ( .A1(n8788), .A2(n10096), .ZN(n4508) );
  OAI21_X1 U5944 ( .B1(n8800), .B2(n10085), .A(n4451), .ZN(n8874) );
  NOR2_X1 U5945 ( .A1(n8798), .A2(n4854), .ZN(n4853) );
  INV_X1 U5946 ( .A(n8797), .ZN(n4855) );
  AND2_X1 U5947 ( .A1(n6964), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10044) );
  INV_X1 U5948 ( .A(n10039), .ZN(n10042) );
  INV_X1 U5949 ( .A(n5090), .ZN(n8897) );
  INV_X1 U5950 ( .A(n5674), .ZN(n8904) );
  INV_X1 U5951 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10176) );
  INV_X1 U5952 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6845) );
  INV_X1 U5953 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6797) );
  INV_X1 U5954 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6777) );
  INV_X1 U5955 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6765) );
  INV_X1 U5956 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6756) );
  INV_X1 U5957 ( .A(n4528), .ZN(n5189) );
  AND4_X1 U5958 ( .A1(n6178), .A2(n6177), .A3(n6176), .A4(n6175), .ZN(n7356)
         );
  NAND2_X1 U5959 ( .A1(n4889), .A2(n6270), .ZN(n7656) );
  AND2_X1 U5960 ( .A1(n7071), .A2(n6131), .ZN(n7017) );
  NAND2_X1 U5961 ( .A1(n4621), .A2(n4624), .ZN(n4617) );
  NAND2_X1 U5962 ( .A1(n8985), .A2(n4619), .ZN(n4618) );
  INV_X1 U5963 ( .A(n9354), .ZN(n7884) );
  AND3_X1 U5964 ( .A1(n6358), .A2(n6357), .A3(n6356), .ZN(n8991) );
  OR2_X1 U5965 ( .A1(n7361), .A2(n9965), .ZN(n8996) );
  AND4_X1 U5966 ( .A1(n6320), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(n7818)
         );
  INV_X1 U5967 ( .A(n5041), .ZN(n4634) );
  AND2_X1 U5968 ( .A1(n6533), .A2(n6532), .ZN(n9517) );
  AND2_X1 U5969 ( .A1(n6653), .A2(n8145), .ZN(n9040) );
  INV_X1 U5970 ( .A(n9040), .ZN(n9011) );
  NAND2_X1 U5971 ( .A1(n8985), .A2(n4625), .ZN(n9019) );
  NAND2_X1 U5972 ( .A1(n4620), .A2(n6452), .ZN(n9018) );
  NAND2_X1 U5973 ( .A1(n6438), .A2(n6437), .ZN(n9616) );
  OR2_X1 U5974 ( .A1(n6661), .A2(n6660), .ZN(n9039) );
  NAND2_X1 U5975 ( .A1(n9031), .A2(n9032), .ZN(n4900) );
  NOR2_X1 U5976 ( .A1(n9032), .A2(n4776), .ZN(n4775) );
  INV_X1 U5977 ( .A(n4777), .ZN(n4776) );
  AND2_X1 U5978 ( .A1(n9710), .A2(n9045), .ZN(n4898) );
  INV_X1 U5979 ( .A(n8996), .ZN(n9045) );
  INV_X1 U5980 ( .A(n8148), .ZN(n9467) );
  OR2_X1 U5981 ( .A1(n6395), .A2(n6394), .ZN(n9658) );
  AOI21_X1 U5982 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9882), .A(n9877), .ZN(
        n7029) );
  NAND2_X1 U5983 ( .A1(n6857), .A2(n6856), .ZN(n6855) );
  NAND2_X1 U5984 ( .A1(n6855), .A2(n4410), .ZN(n6819) );
  INV_X1 U5985 ( .A(n4795), .ZN(n7009) );
  INV_X1 U5986 ( .A(n4793), .ZN(n7096) );
  INV_X1 U5987 ( .A(n4787), .ZN(n7691) );
  NOR2_X1 U5988 ( .A1(n9387), .A2(n9386), .ZN(n9390) );
  NOR2_X1 U5989 ( .A1(n9390), .A2(n9389), .ZN(n9412) );
  INV_X1 U5990 ( .A(n9888), .ZN(n9910) );
  INV_X1 U5991 ( .A(n9901), .ZN(n9917) );
  INV_X1 U5992 ( .A(n9449), .ZN(n9682) );
  NAND2_X1 U5993 ( .A1(n9057), .A2(n9056), .ZN(n9683) );
  XNOR2_X1 U5994 ( .A(n9471), .B(n9683), .ZN(n9686) );
  NAND2_X1 U5995 ( .A1(n4964), .A2(n9215), .ZN(n8038) );
  INV_X1 U5996 ( .A(n4563), .ZN(n9497) );
  AOI21_X1 U5997 ( .B1(n9511), .B2(n8025), .A(n4412), .ZN(n4563) );
  NAND2_X1 U5998 ( .A1(n6538), .A2(n6537), .ZN(n9722) );
  NAND2_X1 U5999 ( .A1(n9554), .A2(n5045), .ZN(n9539) );
  NAND2_X1 U6000 ( .A1(n9562), .A2(n9563), .ZN(n9561) );
  NAND2_X1 U6001 ( .A1(n9576), .A2(n9129), .ZN(n9562) );
  NAND2_X1 U6002 ( .A1(n9619), .A2(n9174), .ZN(n9621) );
  NAND2_X1 U6003 ( .A1(n4977), .A2(n4975), .ZN(n9619) );
  INV_X1 U6004 ( .A(n8017), .ZN(n4978) );
  NAND2_X1 U6005 ( .A1(n9625), .A2(n9116), .ZN(n4980) );
  AND2_X1 U6006 ( .A1(n9655), .A2(n8035), .ZN(n9627) );
  NAND2_X1 U6007 ( .A1(n4673), .A2(n4672), .ZN(n8033) );
  NAND2_X1 U6008 ( .A1(n7596), .A2(n9176), .ZN(n4552) );
  NAND2_X1 U6009 ( .A1(n7503), .A2(n7502), .ZN(n7516) );
  AND2_X2 U6010 ( .A1(n7113), .A2(n6921), .ZN(n10175) );
  INV_X1 U6011 ( .A(n9926), .ZN(n9927) );
  AND2_X1 U6012 ( .A1(n6728), .A2(n6616), .ZN(n9925) );
  NAND2_X1 U6013 ( .A1(n6057), .A2(n4985), .ZN(n4984) );
  INV_X1 U6014 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4985) );
  CLKBUF_X1 U6015 ( .A(n6646), .Z(n8145) );
  NAND2_X1 U6016 ( .A1(n4914), .A2(n4918), .ZN(n5542) );
  NAND2_X1 U6017 ( .A1(n5506), .A2(n4921), .ZN(n4914) );
  INV_X1 U6018 ( .A(n6084), .ZN(n9328) );
  INV_X1 U6019 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6795) );
  XNOR2_X1 U6020 ( .A(n6294), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7439) );
  AND2_X1 U6021 ( .A1(n6252), .A2(n6272), .ZN(n9899) );
  XNOR2_X1 U6022 ( .A(n4901), .B(n4938), .ZN(n8046) );
  XNOR2_X1 U6023 ( .A(n5141), .B(n5151), .ZN(n4938) );
  OAI21_X1 U6024 ( .B1(n5598), .B2(n8045), .A(n4525), .ZN(n5141) );
  NAND2_X1 U6025 ( .A1(n5598), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U6026 ( .A1(n4790), .A2(n4789), .ZN(n4791) );
  NOR2_X1 U6027 ( .A1(n6087), .A2(n6061), .ZN(n4789) );
  XNOR2_X1 U6028 ( .A(n6098), .B(n6097), .ZN(n6823) );
  OAI21_X1 U6029 ( .B1(n10143), .B2(n9848), .A(n10145), .ZN(n10481) );
  AND2_X1 U6030 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9855), .ZN(n10468) );
  XNOR2_X1 U6031 ( .A(n9860), .B(n4522), .ZN(n10480) );
  INV_X1 U6032 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4522) );
  XNOR2_X1 U6033 ( .A(n9863), .B(n4523), .ZN(n10478) );
  NOR2_X1 U6034 ( .A1(n10475), .A2(n9867), .ZN(n10171) );
  NOR2_X1 U6035 ( .A1(n10171), .A2(n10170), .ZN(n10169) );
  AOI21_X1 U6036 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10169), .ZN(n10168) );
  AOI21_X1 U6037 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10166), .ZN(n10165) );
  OAI21_X1 U6038 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10163), .ZN(n10161) );
  NAND2_X1 U6039 ( .A1(n10161), .A2(n10162), .ZN(n10160) );
  NAND2_X1 U6040 ( .A1(n10160), .A2(n4519), .ZN(n10158) );
  NAND2_X1 U6041 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  INV_X1 U6042 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4521) );
  OAI21_X1 U6043 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10157), .ZN(n10155) );
  NAND2_X1 U6044 ( .A1(n10155), .A2(n10156), .ZN(n10154) );
  NAND2_X1 U6045 ( .A1(n10154), .A2(n4517), .ZN(n10152) );
  NAND2_X1 U6046 ( .A1(n7762), .A2(n4518), .ZN(n4517) );
  INV_X1 U6047 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4518) );
  INV_X1 U6048 ( .A(n4505), .ZN(n4504) );
  OAI21_X1 U6049 ( .B1(n8207), .B2(n8425), .A(n8206), .ZN(n4505) );
  NAND2_X1 U6050 ( .A1(n4541), .A2(n4540), .ZN(P2_U3242) );
  AND2_X1 U6051 ( .A1(n4477), .A2(n8416), .ZN(n4540) );
  NAND2_X1 U6052 ( .A1(n5994), .A2(n5974), .ZN(n4513) );
  INV_X1 U6053 ( .A(n4642), .ZN(n4512) );
  OAI21_X1 U6054 ( .B1(n8791), .B2(n8763), .A(n5730), .ZN(n5731) );
  NAND2_X1 U6055 ( .A1(n4713), .A2(n4712), .ZN(P2_U3545) );
  OR2_X1 U6056 ( .A1(n10142), .A2(n5571), .ZN(n4712) );
  NAND2_X1 U6057 ( .A1(n8874), .A2(n10142), .ZN(n4713) );
  NAND2_X1 U6058 ( .A1(n4852), .A2(n4851), .ZN(P2_U3513) );
  NAND2_X1 U6059 ( .A1(n10119), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U6060 ( .A1(n8874), .A2(n10121), .ZN(n4852) );
  OAI21_X1 U6061 ( .B1(n9030), .B2(n4899), .A(n4897), .ZN(P1_U3238) );
  NOR2_X1 U6062 ( .A1(n9033), .A2(n4898), .ZN(n4897) );
  INV_X1 U6063 ( .A(n4774), .ZN(n9030) );
  NAND2_X1 U6064 ( .A1(n4900), .A2(n8986), .ZN(n4899) );
  AND4_X1 U6065 ( .A1(n9338), .A2(n9337), .A3(n9336), .A4(n9335), .ZN(n9346)
         );
  INV_X1 U6066 ( .A(n9448), .ZN(n4812) );
  NAND2_X1 U6067 ( .A1(n9440), .A2(n9281), .ZN(n4813) );
  NAND2_X1 U6068 ( .A1(n9445), .A2(n9521), .ZN(n4814) );
  INV_X1 U6069 ( .A(n4494), .ZN(n4493) );
  OAI21_X1 U6070 ( .B1(n9478), .B2(n9645), .A(n4495), .ZN(n4494) );
  INV_X1 U6071 ( .A(n4529), .ZN(n8160) );
  OAI21_X1 U6072 ( .B1(n9703), .B2(n9679), .A(n4530), .ZN(n4529) );
  AOI21_X1 U6073 ( .B1(n9701), .B2(n9600), .A(n8159), .ZN(n4530) );
  NOR2_X1 U6074 ( .A1(n9713), .A2(n9679), .ZN(n9493) );
  NOR2_X1 U6075 ( .A1(n9728), .A2(n9679), .ZN(n9536) );
  NAND2_X1 U6076 ( .A1(n4515), .A2(n4514), .ZN(P1_U3547) );
  OR2_X1 U6077 ( .A1(n9977), .A2(n6545), .ZN(n4514) );
  OAI21_X1 U6078 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9871), .A(n10471), .ZN(
        n9874) );
  NOR2_X1 U6079 ( .A1(n8909), .A2(n8908), .ZN(n4392) );
  AND2_X1 U6080 ( .A1(n4392), .A2(n8986), .ZN(n4393) );
  AND2_X1 U6081 ( .A1(n9231), .A2(n9112), .ZN(n4394) );
  AND2_X1 U6082 ( .A1(n5016), .A2(n8919), .ZN(n4395) );
  AND2_X1 U6083 ( .A1(n8822), .A2(n8686), .ZN(n5709) );
  AND2_X1 U6084 ( .A1(n5933), .A2(n5937), .ZN(n8599) );
  INV_X1 U6085 ( .A(n9215), .ZN(n4963) );
  AND2_X1 U6086 ( .A1(n6270), .A2(n4434), .ZN(n4396) );
  INV_X1 U6087 ( .A(n9129), .ZN(n4952) );
  OR2_X1 U6088 ( .A1(n8258), .A2(n8543), .ZN(n5953) );
  INV_X1 U6089 ( .A(n5953), .ZN(n4841) );
  INV_X1 U6090 ( .A(n9231), .ZN(n4670) );
  AND2_X1 U6091 ( .A1(n9691), .A2(n4428), .ZN(n4397) );
  AND2_X1 U6092 ( .A1(n4595), .A2(n4444), .ZN(n4398) );
  NAND2_X1 U6093 ( .A1(n5885), .A2(n5880), .ZN(n4399) );
  INV_X1 U6094 ( .A(n4622), .ZN(n4621) );
  NAND2_X1 U6095 ( .A1(n4623), .A2(n9021), .ZN(n4622) );
  INV_X1 U6096 ( .A(n8637), .ZN(n4705) );
  AND2_X1 U6097 ( .A1(n5438), .A2(SI_17_), .ZN(n4400) );
  XNOR2_X1 U6098 ( .A(n5452), .B(SI_18_), .ZN(n5450) );
  NAND2_X1 U6099 ( .A1(n4722), .A2(n4456), .ZN(n4401) );
  AND2_X1 U6101 ( .A1(n5012), .A2(n5011), .ZN(n4402) );
  NAND2_X1 U6102 ( .A1(n6865), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6815) );
  NOR2_X1 U6103 ( .A1(n9412), .A2(n4479), .ZN(n4403) );
  INV_X1 U6104 ( .A(n8081), .ZN(n4871) );
  INV_X1 U6105 ( .A(n8426), .ZN(n8398) );
  AND2_X1 U6106 ( .A1(n5513), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4404) );
  AND2_X2 U6107 ( .A1(n6686), .A2(n4524), .ZN(n5272) );
  OR2_X1 U6108 ( .A1(n9706), .A2(n9489), .ZN(n4406) );
  INV_X1 U6109 ( .A(n6510), .ZN(n6647) );
  INV_X2 U6110 ( .A(n8190), .ZN(n7176) );
  XNOR2_X1 U6111 ( .A(n5371), .B(n10337), .ZN(n5370) );
  INV_X1 U6112 ( .A(n7813), .ZN(n4636) );
  AND2_X1 U6113 ( .A1(n5623), .A2(n5626), .ZN(n4407) );
  NAND2_X1 U6114 ( .A1(n5722), .A2(n4940), .ZN(n4408) );
  XNOR2_X1 U6115 ( .A(n5438), .B(n5423), .ZN(n5437) );
  AND2_X1 U6116 ( .A1(n4650), .A2(n4826), .ZN(n4409) );
  OR2_X1 U6117 ( .A1(n6860), .A2(n6818), .ZN(n4410) );
  OR2_X1 U6118 ( .A1(n10018), .A2(n10070), .ZN(n5842) );
  NAND2_X1 U6119 ( .A1(n7916), .A2(n8969), .ZN(n4411) );
  NAND2_X1 U6120 ( .A1(n6455), .A2(n6454), .ZN(n9745) );
  INV_X1 U6121 ( .A(n4919), .ZN(n4918) );
  OAI21_X1 U6122 ( .B1(n5524), .B2(n4920), .A(n5523), .ZN(n4919) );
  AND2_X1 U6123 ( .A1(n8103), .A2(n8963), .ZN(n4412) );
  NOR2_X1 U6124 ( .A1(n8650), .A2(n8638), .ZN(n4413) );
  OR2_X1 U6125 ( .A1(n5487), .A2(n5489), .ZN(n4414) );
  NAND2_X1 U6126 ( .A1(n5103), .A2(n5017), .ZN(n5086) );
  NAND2_X1 U6127 ( .A1(n7748), .A2(n5031), .ZN(n7862) );
  OR2_X1 U6128 ( .A1(n9596), .A2(n9740), .ZN(n4415) );
  AND2_X1 U6129 ( .A1(n5336), .A2(n5700), .ZN(n5031) );
  AND2_X1 U6130 ( .A1(n5325), .A2(n5405), .ZN(n4416) );
  OAI21_X1 U6131 ( .B1(n8659), .B2(n4708), .A(n4706), .ZN(n8627) );
  NAND2_X1 U6132 ( .A1(n9546), .A2(n9137), .ZN(n9533) );
  AND3_X1 U6133 ( .A1(n5987), .A2(n5975), .A3(n8599), .ZN(n4417) );
  NAND2_X1 U6134 ( .A1(n4633), .A2(n4632), .ZN(n7914) );
  INV_X1 U6135 ( .A(n9134), .ZN(n4951) );
  INV_X1 U6136 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5623) );
  INV_X1 U6137 ( .A(n8747), .ZN(n4718) );
  XNOR2_X1 U6138 ( .A(n5542), .B(n5541), .ZN(n6523) );
  AOI21_X1 U6139 ( .B1(n9563), .B2(n4952), .A(n4951), .ZN(n4950) );
  NAND2_X1 U6140 ( .A1(n6028), .A2(n6027), .ZN(n9715) );
  XNOR2_X1 U6141 ( .A(n4545), .B(n5266), .ZN(n6249) );
  AOI21_X1 U6142 ( .B1(n8752), .B2(n8747), .A(n5705), .ZN(n8726) );
  NAND2_X1 U6143 ( .A1(n5746), .A2(n5745), .ZN(n8258) );
  INV_X1 U6144 ( .A(n8258), .ZN(n4943) );
  XOR2_X1 U6145 ( .A(n4379), .B(n8799), .Z(n8289) );
  AND2_X1 U6146 ( .A1(n8113), .A2(n9979), .ZN(n4418) );
  INV_X1 U6147 ( .A(n8026), .ZN(n9489) );
  AND2_X1 U6148 ( .A1(n6589), .A2(n6588), .ZN(n8026) );
  AND2_X1 U6149 ( .A1(n9504), .A2(n8025), .ZN(n4419) );
  AND2_X1 U6150 ( .A1(n4641), .A2(n6008), .ZN(n4420) );
  AND2_X1 U6151 ( .A1(n6990), .A2(n6815), .ZN(n4421) );
  NAND2_X1 U6152 ( .A1(n5395), .A2(n5909), .ZN(n8728) );
  AND3_X1 U6153 ( .A1(n5432), .A2(n5431), .A3(n5430), .ZN(n8732) );
  NOR2_X1 U6154 ( .A1(n6084), .A2(n7119), .ZN(n4422) );
  OR2_X1 U6155 ( .A1(n8834), .A2(n8331), .ZN(n8681) );
  AND2_X1 U6156 ( .A1(n9759), .A2(n9607), .ZN(n4423) );
  AND2_X1 U6157 ( .A1(n9087), .A2(n7507), .ZN(n4424) );
  AND2_X1 U6158 ( .A1(n5756), .A2(n4842), .ZN(n4425) );
  NOR2_X1 U6159 ( .A1(n6271), .A2(n4887), .ZN(n4426) );
  AND2_X1 U6160 ( .A1(n4948), .A2(n9548), .ZN(n4427) );
  AND2_X1 U6161 ( .A1(n9690), .A2(n9958), .ZN(n4428) );
  OR2_X1 U6162 ( .A1(n8610), .A2(n5540), .ZN(n4429) );
  NOR2_X1 U6163 ( .A1(n9752), .A2(n8933), .ZN(n4430) );
  INV_X1 U6164 ( .A(n4771), .ZN(n4770) );
  NOR2_X1 U6165 ( .A1(n5319), .A2(n4772), .ZN(n4771) );
  AND2_X1 U6166 ( .A1(n8745), .A2(n5839), .ZN(n4431) );
  NAND2_X1 U6167 ( .A1(n5827), .A2(n5830), .ZN(n8615) );
  OR2_X1 U6168 ( .A1(n6741), .A2(n7564), .ZN(n4432) );
  AND2_X1 U6169 ( .A1(n8566), .A2(n5748), .ZN(n4433) );
  NAND2_X1 U6170 ( .A1(n7654), .A2(n6291), .ZN(n4434) );
  NAND2_X1 U6171 ( .A1(n5800), .A2(n5799), .ZN(n8777) );
  AND2_X1 U6172 ( .A1(n4735), .A2(n9164), .ZN(n4435) );
  INV_X1 U6173 ( .A(n9316), .ZN(n8027) );
  NAND2_X1 U6174 ( .A1(n9274), .A2(n9217), .ZN(n9316) );
  OR2_X1 U6175 ( .A1(n6732), .A2(n6674), .ZN(n4436) );
  OR2_X1 U6176 ( .A1(n7066), .A2(n7299), .ZN(n4437) );
  XNOR2_X1 U6177 ( .A(n5183), .B(SI_4_), .ZN(n5180) );
  OR2_X1 U6178 ( .A1(n9464), .A2(n9462), .ZN(n4438) );
  NAND2_X1 U6179 ( .A1(n9460), .A2(n9461), .ZN(n9205) );
  INV_X1 U6180 ( .A(n9205), .ZN(n4992) );
  AND2_X1 U6181 ( .A1(n4747), .A2(n4824), .ZN(n4439) );
  OR2_X1 U6182 ( .A1(n8047), .A2(n6673), .ZN(n4440) );
  INV_X1 U6183 ( .A(n8838), .ZN(n4936) );
  AND2_X1 U6184 ( .A1(n5696), .A2(n5695), .ZN(n4441) );
  OR2_X1 U6185 ( .A1(n7792), .A2(n9354), .ZN(n4442) );
  NOR2_X1 U6186 ( .A1(n9545), .A2(n8926), .ZN(n4443) );
  NAND2_X1 U6187 ( .A1(n5245), .A2(n5244), .ZN(n5265) );
  INV_X1 U6188 ( .A(n5265), .ZN(n4906) );
  OR2_X1 U6189 ( .A1(n4596), .A2(n4590), .ZN(n4444) );
  AND4_X1 U6190 ( .A1(n7588), .A2(n7532), .A3(n5978), .A4(n7541), .ZN(n4445)
         );
  AND2_X1 U6191 ( .A1(n8650), .A2(n8638), .ZN(n4446) );
  INV_X1 U6192 ( .A(n4819), .ZN(n4818) );
  NOR2_X1 U6193 ( .A1(n6770), .A2(n6679), .ZN(n4819) );
  INV_X1 U6194 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7003) );
  INV_X1 U6195 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7724) );
  AND2_X1 U6196 ( .A1(n7949), .A2(n9352), .ZN(n4447) );
  AND2_X1 U6197 ( .A1(n4606), .A2(n4605), .ZN(n4448) );
  AND2_X1 U6198 ( .A1(n8207), .A2(n8410), .ZN(n4449) );
  NAND2_X1 U6199 ( .A1(n8634), .A2(n8282), .ZN(n4450) );
  AND2_X1 U6200 ( .A1(n4855), .A2(n4853), .ZN(n4451) );
  INV_X1 U6201 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5101) );
  OR2_X1 U6202 ( .A1(n9715), .A2(n9488), .ZN(n4452) );
  AND2_X1 U6203 ( .A1(n6401), .A2(n4411), .ZN(n4453) );
  AND2_X1 U6204 ( .A1(n5421), .A2(n5437), .ZN(n4454) );
  AND2_X1 U6205 ( .A1(n6775), .A2(n6680), .ZN(n4455) );
  INV_X1 U6206 ( .A(n4684), .ZN(n4683) );
  NAND2_X1 U6207 ( .A1(n9464), .A2(n9461), .ZN(n4684) );
  AND2_X1 U6208 ( .A1(n8700), .A2(n8331), .ZN(n4456) );
  INV_X1 U6209 ( .A(n6452), .ZN(n4624) );
  AND2_X1 U6210 ( .A1(n5891), .A2(n5882), .ZN(n7864) );
  OR2_X1 U6211 ( .A1(n5216), .A2(n7551), .ZN(n4457) );
  AND2_X1 U6212 ( .A1(n5318), .A2(SI_11_), .ZN(n4458) );
  INV_X1 U6213 ( .A(n4600), .ZN(n4599) );
  NAND2_X1 U6214 ( .A1(n5058), .A2(n5437), .ZN(n4600) );
  AND2_X1 U6215 ( .A1(n9710), .A2(n9506), .ZN(n9170) );
  INV_X1 U6216 ( .A(n5707), .ZN(n4722) );
  AND2_X1 U6217 ( .A1(n4826), .A2(n4431), .ZN(n4459) );
  INV_X1 U6218 ( .A(n4626), .ZN(n4625) );
  OR2_X1 U6219 ( .A1(n6452), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U6220 ( .A1(n5960), .A2(n5961), .ZN(n8776) );
  INV_X1 U6221 ( .A(n8776), .ZN(n4929) );
  AND3_X1 U6222 ( .A1(n5162), .A2(n5161), .A3(n5160), .ZN(n10032) );
  INV_X1 U6223 ( .A(n10032), .ZN(n5163) );
  AND2_X1 U6224 ( .A1(n6204), .A2(n6170), .ZN(n4460) );
  INV_X1 U6225 ( .A(n8650), .ZN(n8817) );
  AND2_X1 U6226 ( .A1(n5494), .A2(n5493), .ZN(n8650) );
  OR2_X1 U6227 ( .A1(n9473), .A2(n6647), .ZN(n4461) );
  AND3_X1 U6228 ( .A1(n5178), .A2(n5177), .A3(n5176), .ZN(n10070) );
  INV_X1 U6229 ( .A(n5801), .ZN(n4842) );
  AND2_X1 U6230 ( .A1(n4997), .A2(n4558), .ZN(n4462) );
  AND2_X1 U6231 ( .A1(n6334), .A2(n4636), .ZN(n4463) );
  AND2_X1 U6232 ( .A1(n6504), .A2(n6518), .ZN(n4464) );
  AND2_X1 U6233 ( .A1(n8780), .A2(n8778), .ZN(n4465) );
  AND2_X1 U6234 ( .A1(n9069), .A2(n4662), .ZN(n4466) );
  AND2_X1 U6235 ( .A1(n4936), .A2(n8732), .ZN(n4467) );
  INV_X1 U6236 ( .A(n8773), .ZN(n8136) );
  AND2_X1 U6237 ( .A1(n5785), .A2(n5784), .ZN(n8773) );
  INV_X1 U6238 ( .A(n5005), .ZN(n5004) );
  NOR2_X1 U6239 ( .A1(n7504), .A2(n5006), .ZN(n5005) );
  AND2_X1 U6240 ( .A1(n5415), .A2(n5909), .ZN(n4468) );
  NAND2_X1 U6241 ( .A1(n5885), .A2(n5888), .ZN(n4469) );
  OR2_X1 U6242 ( .A1(n7743), .A2(n7517), .ZN(n9090) );
  AND2_X1 U6243 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n4470) );
  INV_X1 U6244 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5070) );
  INV_X1 U6245 ( .A(n5117), .ZN(n4823) );
  INV_X1 U6246 ( .A(n5763), .ZN(n5609) );
  NAND2_X1 U6247 ( .A1(n5692), .A2(n5691), .ZN(n7612) );
  NAND2_X1 U6248 ( .A1(n7827), .A2(n7710), .ZN(n7804) );
  AND2_X1 U6249 ( .A1(n7624), .A2(n5720), .ZN(n4471) );
  NAND2_X1 U6250 ( .A1(n9328), .A2(n9521), .ZN(n9157) );
  INV_X1 U6251 ( .A(n9196), .ZN(n4671) );
  NAND2_X1 U6252 ( .A1(n7840), .A2(n7839), .ZN(n7937) );
  NAND2_X1 U6253 ( .A1(n5003), .A2(n5001), .ZN(n7596) );
  NAND2_X1 U6254 ( .A1(n4552), .A2(n7597), .ZN(n7771) );
  NAND2_X1 U6255 ( .A1(n7506), .A2(n9087), .ZN(n7518) );
  NAND2_X1 U6256 ( .A1(n7750), .A2(n7749), .ZN(n7748) );
  AND2_X1 U6257 ( .A1(n8072), .A2(n8071), .ZN(n4472) );
  NAND2_X1 U6258 ( .A1(n7748), .A2(n5700), .ZN(n7863) );
  AND2_X1 U6259 ( .A1(n9169), .A2(n9157), .ZN(n4473) );
  NAND2_X1 U6260 ( .A1(n6621), .A2(n6620), .ZN(n9700) );
  INV_X1 U6261 ( .A(n9700), .ZN(n5015) );
  INV_X1 U6262 ( .A(n4507), .ZN(n8719) );
  AND2_X1 U6263 ( .A1(n5574), .A2(n5573), .ZN(n8592) );
  OR2_X1 U6264 ( .A1(n7345), .A2(n6681), .ZN(n4474) );
  INV_X1 U6265 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10241) );
  INV_X1 U6266 ( .A(n4604), .ZN(n4603) );
  NAND2_X1 U6267 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(n5308), .ZN(n4604) );
  AND2_X1 U6268 ( .A1(n4637), .A2(n4634), .ZN(n4475) );
  AND2_X1 U6269 ( .A1(n4980), .A2(n4978), .ZN(n4476) );
  OR2_X1 U6270 ( .A1(n8565), .A2(n8425), .ZN(n4477) );
  OR2_X1 U6271 ( .A1(n9503), .A2(n8996), .ZN(n4478) );
  INV_X1 U6272 ( .A(n5068), .ZN(n5024) );
  INV_X1 U6273 ( .A(n5557), .ZN(n4588) );
  AND2_X1 U6274 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  INV_X1 U6275 ( .A(n5709), .ZN(n4711) );
  INV_X1 U6276 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U6277 ( .A1(n4782), .A2(n4781), .ZN(n4784) );
  AND2_X2 U6278 ( .A1(n6003), .A2(n6002), .ZN(n10121) );
  AND2_X1 U6279 ( .A1(n9413), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U6280 ( .A1(n6338), .A2(n6337), .ZN(n7949) );
  INV_X1 U6281 ( .A(n7949), .ZN(n5011) );
  NAND2_X1 U6282 ( .A1(n6182), .A2(n6181), .ZN(n9943) );
  INV_X1 U6283 ( .A(n9943), .ZN(n5010) );
  INV_X1 U6284 ( .A(n7822), .ZN(n4862) );
  NAND2_X1 U6285 ( .A1(n5804), .A2(n5803), .ZN(n4480) );
  INV_X1 U6286 ( .A(n4809), .ZN(n9891) );
  NAND2_X1 U6287 ( .A1(n6855), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U6288 ( .A1(n5797), .A2(n10338), .ZN(n4481) );
  AND2_X1 U6289 ( .A1(n4608), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n4482) );
  AND2_X1 U6290 ( .A1(n7582), .A2(n5683), .ZN(n4483) );
  AND2_X1 U6291 ( .A1(n8489), .A2(n4572), .ZN(n4484) );
  AND2_X1 U6292 ( .A1(n4798), .A2(n9418), .ZN(n4485) );
  AND2_X1 U6293 ( .A1(n4784), .A2(n6815), .ZN(n4486) );
  INV_X1 U6294 ( .A(n4934), .ZN(n4933) );
  NAND2_X1 U6295 ( .A1(n4481), .A2(n5779), .ZN(n4934) );
  INV_X1 U6296 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6433) );
  INV_X1 U6297 ( .A(n9281), .ZN(n9521) );
  INV_X1 U6298 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6079) );
  INV_X1 U6299 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n4610) );
  INV_X1 U6300 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n4609) );
  INV_X1 U6301 ( .A(n5619), .ZN(n8575) );
  OR2_X1 U6302 ( .A1(n6910), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4487) );
  INV_X1 U6303 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4523) );
  INV_X1 U6304 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4583) );
  INV_X1 U6305 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4970) );
  INV_X1 U6306 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U6307 ( .A1(n4721), .A2(n5705), .ZN(n4720) );
  NAND2_X1 U6308 ( .A1(n4765), .A2(n4762), .ZN(n5357) );
  NAND2_X1 U6309 ( .A1(n7108), .A2(n4689), .ZN(n4490) );
  NOR2_X1 U6310 ( .A1(n8112), .A2(n4418), .ZN(n8117) );
  NAND2_X1 U6311 ( .A1(n8255), .A2(n8254), .ZN(n8263) );
  NOR2_X1 U6312 ( .A1(n8291), .A2(n4878), .ZN(n4578) );
  NAND2_X1 U6313 ( .A1(n7705), .A2(n7704), .ZN(n7823) );
  OAI21_X1 U6314 ( .B1(n4741), .B2(n4740), .A(n4737), .ZN(n5904) );
  AND2_X1 U6315 ( .A1(n5863), .A2(n7378), .ZN(n7549) );
  NAND2_X1 U6316 ( .A1(n4492), .A2(n5910), .ZN(n4531) );
  NAND3_X1 U6317 ( .A1(n5906), .A2(n4718), .A3(n5907), .ZN(n4492) );
  AOI21_X1 U6318 ( .B1(n5945), .B2(n5944), .A(n4745), .ZN(n4744) );
  AOI21_X1 U6319 ( .B1(n5927), .B2(n4755), .A(n4754), .ZN(n4753) );
  NAND3_X1 U6320 ( .A1(n6939), .A2(n6940), .A3(n9289), .ZN(n7666) );
  NAND2_X2 U6321 ( .A1(n9575), .A2(n9577), .ZN(n9576) );
  NAND2_X1 U6322 ( .A1(n4496), .A2(n4493), .ZN(P1_U3355) );
  NAND2_X1 U6323 ( .A1(n9687), .A2(n7131), .ZN(n4496) );
  NAND2_X1 U6324 ( .A1(n4506), .A2(n4504), .ZN(P2_U3216) );
  NAND2_X1 U6325 ( .A1(n8202), .A2(n8255), .ZN(n4506) );
  NAND2_X1 U6326 ( .A1(n7186), .A2(n8240), .ZN(n8242) );
  AOI21_X2 U6327 ( .B1(n8339), .B2(n8187), .A(n5050), .ZN(n8291) );
  NAND4_X1 U6328 ( .A1(n7932), .A2(n4937), .A3(n4936), .A4(n8741), .ZN(n4507)
         );
  XNOR2_X1 U6329 ( .A(n5111), .B(n5112), .ZN(n6762) );
  NAND2_X1 U6330 ( .A1(n5242), .A2(n4904), .ZN(n4723) );
  NAND3_X1 U6331 ( .A1(n4453), .A2(n4633), .A3(n4509), .ZN(n4631) );
  OR2_X2 U6332 ( .A1(n4630), .A2(n4510), .ZN(n4509) );
  AND2_X2 U6333 ( .A1(n7786), .A2(n6334), .ZN(n4510) );
  NAND2_X1 U6334 ( .A1(n4657), .A2(n5239), .ZN(n5242) );
  NAND3_X1 U6335 ( .A1(n4644), .A2(n4643), .A3(n5201), .ZN(n5235) );
  NAND4_X1 U6336 ( .A1(n4756), .A2(n4374), .A3(n4513), .A4(n4512), .ZN(
        P2_U3244) );
  NAND2_X1 U6337 ( .A1(n5754), .A2(n5753), .ZN(n5757) );
  NAND2_X1 U6338 ( .A1(n7617), .A2(n5264), .ZN(n7638) );
  NAND2_X1 U6339 ( .A1(n5795), .A2(n5953), .ZN(n8534) );
  INV_X1 U6340 ( .A(n7296), .ZN(n5232) );
  OAI21_X2 U6341 ( .B1(n7531), .B2(n7530), .A(n5855), .ZN(n10014) );
  NAND2_X1 U6342 ( .A1(n9808), .A2(n9977), .ZN(n4515) );
  NAND2_X1 U6343 ( .A1(n9723), .A2(n4516), .ZN(n9808) );
  AND4_X2 U6344 ( .A1(n4959), .A2(n6022), .A3(n6008), .A4(n6016), .ZN(n4956)
         );
  NAND2_X1 U6345 ( .A1(n4949), .A2(n4427), .ZN(n9546) );
  NAND2_X1 U6346 ( .A1(n9533), .A2(n9247), .ZN(n9513) );
  NAND2_X1 U6347 ( .A1(n7846), .A2(n7845), .ZN(n4947) );
  NOR2_X1 U6348 ( .A1(n10168), .A2(n10167), .ZN(n10166) );
  NOR2_X1 U6349 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10468), .ZN(n9856) );
  NAND3_X1 U6350 ( .A1(n8968), .A2(n8967), .A3(n4478), .ZN(P1_U3223) );
  NAND2_X2 U6351 ( .A1(n6428), .A2(n8982), .ZN(n8985) );
  NAND2_X1 U6352 ( .A1(n6402), .A2(n4778), .ZN(n6401) );
  NAND2_X1 U6353 ( .A1(n8779), .A2(n4465), .ZN(n8781) );
  NAND2_X1 U6354 ( .A1(n8550), .A2(n8549), .ZN(n8779) );
  NAND2_X1 U6355 ( .A1(n4527), .A2(n4526), .ZN(n5906) );
  NAND2_X1 U6356 ( .A1(n5904), .A2(n7924), .ZN(n4527) );
  AND2_X4 U6357 ( .A1(n5117), .A2(n5070), .ZN(n5406) );
  NAND2_X1 U6358 ( .A1(n4761), .A2(n4759), .ZN(n5919) );
  AOI21_X1 U6359 ( .B1(n5994), .B2(n4376), .A(n5993), .ZN(n4757) );
  NAND2_X1 U6360 ( .A1(n4949), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U6361 ( .A1(n4531), .A2(n5415), .ZN(n5911) );
  INV_X1 U6362 ( .A(n4757), .ZN(n4756) );
  AOI21_X1 U6363 ( .B1(n5850), .B2(n5844), .A(n5843), .ZN(n5852) );
  OAI21_X1 U6364 ( .B1(n4753), .B2(n4752), .A(n5937), .ZN(n5930) );
  OAI21_X1 U6365 ( .B1(n4744), .B2(n4743), .A(n4742), .ZN(n5957) );
  NAND2_X1 U6366 ( .A1(n9626), .A2(n9118), .ZN(n4731) );
  OAI21_X1 U6367 ( .B1(n4435), .B2(n4534), .A(n4532), .ZN(n9153) );
  NAND2_X1 U6368 ( .A1(n5919), .A2(n5918), .ZN(n5921) );
  OAI21_X1 U6369 ( .B1(n4730), .B2(n4729), .A(n9120), .ZN(n9124) );
  NOR2_X1 U6370 ( .A1(n9344), .A2(n9166), .ZN(n9213) );
  NAND3_X1 U6371 ( .A1(n4543), .A2(n4542), .A3(n8398), .ZN(n4541) );
  NAND2_X1 U6372 ( .A1(n4867), .A2(n4864), .ZN(n8279) );
  AOI21_X1 U6373 ( .B1(n7824), .B2(n4860), .A(n4858), .ZN(n4857) );
  NAND4_X1 U6374 ( .A1(n5406), .A2(n5325), .A3(n5405), .A4(n5079), .ZN(n5458)
         );
  NAND2_X1 U6375 ( .A1(n4901), .A2(n5153), .ZN(n4544) );
  NAND2_X1 U6376 ( .A1(n4544), .A2(n5155), .ZN(n5170) );
  NAND2_X1 U6377 ( .A1(n5173), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6378 ( .A1(n4550), .A2(n4553), .ZN(n7838) );
  NAND3_X1 U6379 ( .A1(n5003), .A2(n5001), .A3(n4551), .ZN(n4550) );
  NAND2_X1 U6380 ( .A1(n9569), .A2(n4560), .ZN(n4556) );
  NAND2_X1 U6381 ( .A1(n4556), .A2(n4462), .ZN(n9526) );
  XNOR2_X1 U6382 ( .A(n9479), .B(n4566), .ZN(n9714) );
  INV_X1 U6383 ( .A(n4573), .ZN(n7344) );
  OAI21_X2 U6384 ( .B1(n4579), .B2(n4578), .A(n8201), .ZN(n8255) );
  AND2_X4 U6385 ( .A1(n4581), .A2(n4580), .ZN(n5598) );
  NAND2_X1 U6386 ( .A1(n5492), .A2(n4585), .ZN(n4584) );
  NAND2_X1 U6387 ( .A1(n5309), .A2(n4602), .ZN(n5365) );
  NAND3_X1 U6388 ( .A1(n5951), .A2(n5959), .A3(n5954), .ZN(n4605) );
  NAND2_X1 U6389 ( .A1(n4607), .A2(n4470), .ZN(n5226) );
  NAND2_X1 U6390 ( .A1(n5566), .A2(n4482), .ZN(n5629) );
  NAND2_X1 U6391 ( .A1(n5566), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6392 ( .A1(n5427), .A2(n4611), .ZN(n5480) );
  INV_X1 U6393 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4614) );
  NOR2_X4 U6394 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6086) );
  NAND2_X1 U6395 ( .A1(n8948), .A2(n4464), .ZN(n9006) );
  NAND2_X1 U6396 ( .A1(n8948), .A2(n6504), .ZN(n4616) );
  NAND2_X1 U6397 ( .A1(n6500), .A2(n8946), .ZN(n8948) );
  NAND2_X2 U6398 ( .A1(n4618), .A2(n4617), .ZN(n8931) );
  NAND2_X1 U6399 ( .A1(n4637), .A2(n4635), .ZN(n4632) );
  NAND2_X1 U6400 ( .A1(n7786), .A2(n6334), .ZN(n4637) );
  AOI21_X1 U6401 ( .B1(n5041), .B2(n4636), .A(n4638), .ZN(n4628) );
  NAND2_X1 U6402 ( .A1(n7786), .A2(n4463), .ZN(n4629) );
  NAND2_X1 U6403 ( .A1(n4631), .A2(n6413), .ZN(n6428) );
  INV_X2 U6404 ( .A(n6090), .ZN(n6637) );
  NOR2_X2 U6405 ( .A1(n4422), .A2(n6090), .ZN(n6379) );
  NAND2_X2 U6406 ( .A1(n6728), .A2(n6889), .ZN(n6090) );
  NAND2_X2 U6407 ( .A1(n6047), .A2(n6611), .ZN(n6728) );
  NAND2_X1 U6408 ( .A1(n7087), .A2(n4460), .ZN(n4639) );
  NAND4_X1 U6409 ( .A1(n6039), .A2(n4420), .A3(n4955), .A4(n4640), .ZN(n6614)
         );
  AND2_X1 U6410 ( .A1(n4959), .A2(n6008), .ZN(n6196) );
  INV_X1 U6411 ( .A(n6015), .ZN(n4641) );
  NAND2_X1 U6412 ( .A1(n5180), .A2(n5184), .ZN(n4643) );
  NAND2_X1 U6413 ( .A1(n5283), .A2(n5282), .ZN(n7635) );
  INV_X1 U6414 ( .A(n7507), .ZN(n9188) );
  NAND2_X1 U6415 ( .A1(n4658), .A2(n4466), .ZN(n8037) );
  NAND2_X1 U6416 ( .A1(n8154), .A2(n9274), .ZN(n9463) );
  NAND3_X1 U6417 ( .A1(n5159), .A2(n4686), .A3(n4685), .ZN(n5403) );
  INV_X2 U6418 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6419 ( .A1(n4691), .A2(n4690), .ZN(n7984) );
  NAND3_X1 U6420 ( .A1(n4695), .A2(n5702), .A3(n5031), .ZN(n4691) );
  INV_X1 U6421 ( .A(n7750), .ZN(n4695) );
  NAND3_X1 U6422 ( .A1(n4445), .A2(n4700), .A3(n4699), .ZN(n4698) );
  NAND2_X1 U6423 ( .A1(n4715), .A2(n8752), .ZN(n4714) );
  NAND2_X1 U6424 ( .A1(n9163), .A2(n9276), .ZN(n4727) );
  AOI21_X1 U6425 ( .B1(n4733), .B2(n4732), .A(n4731), .ZN(n4730) );
  NAND2_X1 U6426 ( .A1(n5883), .A2(n4469), .ZN(n4738) );
  OR2_X1 U6427 ( .A1(n5879), .A2(n5878), .ZN(n4741) );
  NAND4_X1 U6428 ( .A1(n4748), .A2(n4750), .A3(n4749), .A4(n4416), .ZN(n4746)
         );
  AND2_X1 U6429 ( .A1(n5081), .A2(n5660), .ZN(n4751) );
  NAND3_X1 U6430 ( .A1(n5929), .A2(n5827), .A3(n5959), .ZN(n4752) );
  NAND3_X1 U6431 ( .A1(n5911), .A2(n5912), .A3(n8706), .ZN(n4761) );
  NAND2_X1 U6432 ( .A1(n5297), .A2(n4766), .ZN(n4765) );
  NAND2_X1 U6433 ( .A1(n8960), .A2(n4777), .ZN(n9031) );
  INV_X1 U6434 ( .A(n4784), .ZN(n6861) );
  INV_X1 U6435 ( .A(n6086), .ZN(n4790) );
  NAND2_X1 U6436 ( .A1(n6135), .A2(n4791), .ZN(n8044) );
  NAND2_X1 U6437 ( .A1(n4797), .A2(n4798), .ZN(n9419) );
  NAND2_X1 U6438 ( .A1(n6857), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U6439 ( .A1(n4805), .A2(n4802), .ZN(n9895) );
  NAND3_X1 U6440 ( .A1(n4814), .A2(n4813), .A3(n4812), .ZN(P1_U3260) );
  AOI22_X1 U6441 ( .A1(n6876), .A2(n6875), .B1(n6817), .B2(n6816), .ZN(n6857)
         );
  NOR2_X1 U6442 ( .A1(n9422), .A2(n9421), .ZN(n9435) );
  NOR2_X1 U6443 ( .A1(n7029), .A2(n7028), .ZN(n7027) );
  MUX2_X1 U6444 ( .A(n5840), .B(n7549), .S(n5959), .Z(n5850) );
  AOI21_X1 U6445 ( .B1(n5932), .B2(n5931), .A(n5930), .ZN(n5936) );
  NAND2_X1 U6446 ( .A1(n4822), .A2(n4821), .ZN(n5143) );
  NAND2_X1 U6447 ( .A1(n8890), .A2(n5070), .ZN(n4821) );
  NAND3_X1 U6448 ( .A1(n4823), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U6449 ( .A1(n5395), .A2(n4468), .ZN(n8703) );
  NAND2_X1 U6450 ( .A1(n8703), .A2(n5434), .ZN(n5435) );
  NAND2_X1 U6451 ( .A1(n8682), .A2(n4836), .ZN(n4833) );
  NAND2_X1 U6452 ( .A1(n4833), .A2(n4834), .ZN(n8651) );
  NAND2_X1 U6453 ( .A1(n5757), .A2(n5756), .ZN(n5795) );
  INV_X1 U6454 ( .A(n5960), .ZN(n4843) );
  XNOR2_X1 U6455 ( .A(n5163), .B(n8450), .ZN(n4850) );
  NAND2_X1 U6456 ( .A1(n10014), .A2(n4850), .ZN(n5164) );
  CLKBUF_X1 U6457 ( .A(n4850), .Z(n4849) );
  INV_X1 U6458 ( .A(n4849), .ZN(n10022) );
  OAI21_X1 U6459 ( .B1(n5849), .B2(n5848), .A(n4849), .ZN(n5851) );
  XNOR2_X1 U6460 ( .A(n10014), .B(n4849), .ZN(n10019) );
  NAND3_X1 U6461 ( .A1(n4457), .A2(n5869), .A3(n4856), .ZN(n7296) );
  NAND2_X1 U6462 ( .A1(n7550), .A2(n5215), .ZN(n4856) );
  NAND2_X1 U6463 ( .A1(n8066), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U6464 ( .A1(n8066), .A2(n8081), .ZN(n8083) );
  INV_X1 U6465 ( .A(n4873), .ZN(n4872) );
  AOI21_X1 U6466 ( .B1(n4877), .B2(n4879), .A(n4876), .ZN(n4875) );
  NAND2_X1 U6467 ( .A1(n8291), .A2(n4883), .ZN(n4881) );
  NAND2_X1 U6468 ( .A1(n4886), .A2(n7315), .ZN(n7705) );
  NAND2_X1 U6469 ( .A1(n7314), .A2(n7313), .ZN(n4886) );
  XNOR2_X2 U6470 ( .A(n5624), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5619) );
  NAND2_X2 U6471 ( .A1(n4889), .A2(n4396), .ZN(n7786) );
  NAND2_X2 U6472 ( .A1(n4888), .A2(n4426), .ZN(n4889) );
  NAND2_X1 U6473 ( .A1(n7071), .A2(n4890), .ZN(n4891) );
  NAND2_X1 U6474 ( .A1(n4891), .A2(n7014), .ZN(n7085) );
  OAI21_X1 U6475 ( .B1(n6078), .B2(n4895), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6035) );
  INV_X1 U6476 ( .A(n4892), .ZN(n6076) );
  NAND2_X1 U6477 ( .A1(n5140), .A2(n5139), .ZN(n4901) );
  NAND3_X1 U6478 ( .A1(n4929), .A2(n4927), .A3(n4926), .ZN(n4925) );
  NOR2_X1 U6479 ( .A1(n4928), .A2(n8541), .ZN(n4927) );
  OAI21_X1 U6480 ( .B1(n5776), .B2(n4934), .A(n4931), .ZN(n5810) );
  NAND2_X1 U6481 ( .A1(n5776), .A2(n5775), .ZN(n4935) );
  AND2_X2 U6482 ( .A1(n8719), .A2(n8700), .ZN(n8696) );
  NAND3_X1 U6483 ( .A1(n8741), .A2(n4937), .A3(n7985), .ZN(n8738) );
  INV_X1 U6484 ( .A(n8046), .ZN(n5142) );
  NAND2_X1 U6485 ( .A1(n5722), .A2(n4941), .ZN(n8549) );
  NAND2_X1 U6486 ( .A1(n5722), .A2(n8207), .ZN(n8135) );
  NAND3_X1 U6487 ( .A1(n4944), .A2(n10112), .A3(n7624), .ZN(n5042) );
  NAND2_X2 U6488 ( .A1(n4947), .A2(n9105), .ZN(n7938) );
  OAI21_X1 U6489 ( .B1(n9576), .B2(n9555), .A(n4950), .ZN(n9547) );
  NAND2_X1 U6490 ( .A1(n4950), .A2(n9555), .ZN(n4948) );
  NAND2_X1 U6491 ( .A1(n9576), .A2(n4950), .ZN(n4949) );
  NOR2_X1 U6492 ( .A1(n6015), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4954) );
  NAND3_X1 U6493 ( .A1(n4956), .A2(n4960), .A3(n6029), .ZN(n6024) );
  AND3_X2 U6494 ( .A1(n4956), .A2(n4960), .A3(n4953), .ZN(n6058) );
  INV_X1 U6495 ( .A(n6309), .ZN(n4955) );
  AND2_X2 U6496 ( .A1(n6086), .A2(n6009), .ZN(n4959) );
  NOR2_X2 U6497 ( .A1(n6019), .A2(n4961), .ZN(n4960) );
  NAND3_X1 U6498 ( .A1(n6079), .A2(n10416), .A3(n6037), .ZN(n4961) );
  NAND4_X1 U6499 ( .A1(n6012), .A2(n6011), .A3(n10441), .A4(n6010), .ZN(n6309)
         );
  NAND2_X1 U6500 ( .A1(n7519), .A2(n9078), .ZN(n7841) );
  NAND2_X1 U6501 ( .A1(n9485), .A2(n9312), .ZN(n4964) );
  NAND2_X2 U6502 ( .A1(n4964), .A2(n4962), .ZN(n8154) );
  NAND2_X2 U6503 ( .A1(n6783), .A2(n4524), .ZN(n9055) );
  NAND2_X4 U6504 ( .A1(n6646), .A2(n9835), .ZN(n6783) );
  INV_X1 U6505 ( .A(n9174), .ZN(n4974) );
  INV_X1 U6506 ( .A(n8018), .ZN(n4981) );
  NAND2_X1 U6507 ( .A1(n7840), .A2(n4982), .ZN(n8011) );
  OAI21_X1 U6508 ( .B1(n9479), .B2(n4993), .A(n4991), .ZN(n9689) );
  AOI21_X1 U6509 ( .B1(n9479), .B2(n4991), .A(n4987), .ZN(n4986) );
  AOI21_X1 U6510 ( .B1(n9479), .B2(n4990), .A(n4993), .ZN(n4989) );
  AOI21_X1 U6511 ( .B1(n9479), .B2(n9171), .A(n9170), .ZN(n8147) );
  NAND2_X1 U6512 ( .A1(n7154), .A2(n5005), .ZN(n5003) );
  INV_X1 U6513 ( .A(n7154), .ZN(n5008) );
  AND2_X2 U6514 ( .A1(n7605), .A2(n4402), .ZN(n7941) );
  NAND2_X1 U6515 ( .A1(n9557), .A2(n9545), .ZN(n9540) );
  AND3_X2 U6516 ( .A1(n5014), .A2(n9585), .A3(n9592), .ZN(n9557) );
  NAND2_X1 U6517 ( .A1(n7321), .A2(n5018), .ZN(n5021) );
  AND2_X1 U6518 ( .A1(n5690), .A2(n5687), .ZN(n5018) );
  AOI21_X1 U6519 ( .B1(n7321), .B2(n5687), .A(n5068), .ZN(n7374) );
  NAND3_X1 U6520 ( .A1(n5021), .A2(n5979), .A3(n5019), .ZN(n5692) );
  NAND2_X1 U6521 ( .A1(n5020), .A2(n5690), .ZN(n5019) );
  NAND3_X1 U6522 ( .A1(n7557), .A2(n5024), .A3(n5063), .ZN(n5020) );
  NAND2_X1 U6523 ( .A1(n5022), .A2(n5690), .ZN(n7294) );
  NAND2_X1 U6524 ( .A1(n8564), .A2(n5028), .ZN(n5026) );
  NAND2_X1 U6525 ( .A1(n8564), .A2(n5988), .ZN(n5027) );
  NAND2_X1 U6526 ( .A1(n5032), .A2(n5033), .ZN(n5713) );
  NAND2_X1 U6527 ( .A1(n8598), .A2(n5710), .ZN(n5032) );
  AOI21_X1 U6528 ( .B1(n5415), .B2(n4721), .A(n4467), .ZN(n5034) );
  NAND2_X1 U6529 ( .A1(n5036), .A2(n8711), .ZN(n5035) );
  NOR2_X1 U6530 ( .A1(n8725), .A2(n5706), .ZN(n8712) );
  NAND3_X1 U6531 ( .A1(n7582), .A2(n5683), .A3(n7530), .ZN(n7529) );
  NAND2_X1 U6532 ( .A1(n5976), .A2(n7583), .ZN(n7582) );
  NAND4_X2 U6533 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n6924)
         );
  NAND2_X1 U6534 ( .A1(n9059), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6112) );
  XNOR2_X1 U6535 ( .A(n8147), .B(n8027), .ZN(n9709) );
  AOI211_X2 U6536 ( .C1(n10036), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8578), .B(
        n8577), .ZN(n8579) );
  XNOR2_X1 U6537 ( .A(n6077), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6084) );
  CLKBUF_X1 U6538 ( .A(n8242), .Z(n8359) );
  NAND2_X1 U6539 ( .A1(n6004), .A2(n10142), .ZN(n5774) );
  NAND2_X2 U6540 ( .A1(n5763), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5091) );
  NAND4_X4 U6541 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n8451)
         );
  CLKBUF_X1 U6542 ( .A(n8660), .Z(n8674) );
  XNOR2_X1 U6543 ( .A(n5357), .B(n5052), .ZN(n6798) );
  NAND2_X1 U6544 ( .A1(n5719), .A2(n10070), .ZN(n7375) );
  INV_X1 U6545 ( .A(n7323), .ZN(n5719) );
  AND2_X1 U6546 ( .A1(n8451), .A2(n5681), .ZN(n7583) );
  NAND2_X1 U6547 ( .A1(n6076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6077) );
  CLKBUF_X1 U6548 ( .A(n7932), .Z(n7985) );
  OR2_X1 U6549 ( .A1(n8767), .A2(n10113), .ZN(n8769) );
  XNOR2_X1 U6550 ( .A(n8162), .B(n8161), .ZN(n8767) );
  NAND2_X1 U6551 ( .A1(n7166), .A2(n5821), .ZN(n10020) );
  NAND2_X1 U6552 ( .A1(n6191), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6093) );
  INV_X2 U6553 ( .A(n5681), .ZN(n10046) );
  NAND2_X1 U6554 ( .A1(n9832), .A2(n6068), .ZN(n6393) );
  INV_X2 U6555 ( .A(n5089), .ZN(n8894) );
  NAND2_X1 U6556 ( .A1(n7456), .A2(n7457), .ZN(n7455) );
  NAND2_X1 U6557 ( .A1(n5763), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5128) );
  XNOR2_X1 U6558 ( .A(n5284), .B(n5055), .ZN(n6759) );
  AOI21_X2 U6559 ( .B1(n8217), .B2(n8064), .A(n5048), .ZN(n8080) );
  NAND2_X2 U6560 ( .A1(n6026), .A2(n6063), .ZN(n9835) );
  OR2_X1 U6561 ( .A1(n10113), .A2(n8575), .ZN(n6962) );
  INV_X1 U6562 ( .A(n8610), .ZN(n8611) );
  OR2_X1 U6563 ( .A1(n8790), .A2(n10036), .ZN(n5039) );
  OR2_X1 U6564 ( .A1(n5937), .A2(n5959), .ZN(n5043) );
  INV_X1 U6565 ( .A(n9722), .ZN(n8103) );
  OR2_X1 U6566 ( .A1(n5830), .A2(n5939), .ZN(n5044) );
  AND2_X1 U6567 ( .A1(n4718), .A2(n5394), .ZN(n5047) );
  NOR2_X1 U6568 ( .A1(n8063), .A2(n8327), .ZN(n5048) );
  OR2_X1 U6569 ( .A1(n9592), .A2(n9001), .ZN(n5049) );
  AND2_X1 U6570 ( .A1(n8186), .A2(n8185), .ZN(n5050) );
  OR2_X1 U6571 ( .A1(n4524), .A2(n6735), .ZN(n5051) );
  AND2_X1 U6572 ( .A1(n5345), .A2(n5344), .ZN(n5052) );
  AND2_X1 U6573 ( .A1(n5491), .A2(n5490), .ZN(n5053) );
  INV_X1 U6574 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5156) );
  AND2_X1 U6575 ( .A1(n5298), .A2(n5288), .ZN(n5054) );
  INV_X1 U6576 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6810) );
  AND2_X1 U6577 ( .A1(n6897), .A2(n9327), .ZN(n9659) );
  INV_X1 U6578 ( .A(n9659), .ZN(n9631) );
  AND2_X1 U6579 ( .A1(n5285), .A2(n5271), .ZN(n5055) );
  INV_X1 U6580 ( .A(n8638), .ZN(n8668) );
  AND2_X1 U6581 ( .A1(n8768), .A2(n8771), .ZN(n5057) );
  AND2_X1 U6582 ( .A1(n5420), .A2(n5419), .ZN(n5058) );
  AND2_X1 U6583 ( .A1(n9076), .A2(n9123), .ZN(n5059) );
  INV_X1 U6584 ( .A(n9518), .ZN(n9488) );
  OR2_X2 U6585 ( .A1(n7156), .A2(n7743), .ZN(n5060) );
  INV_X1 U6586 ( .A(n7912), .ZN(n5822) );
  INV_X1 U6587 ( .A(n10095), .ZN(n5720) );
  NAND2_X1 U6588 ( .A1(n8176), .A2(n8380), .ZN(n5061) );
  AND2_X1 U6589 ( .A1(n5234), .A2(n5233), .ZN(n5062) );
  OR2_X1 U6590 ( .A1(n10074), .A2(n7210), .ZN(n5063) );
  INV_X1 U6591 ( .A(n9484), .ZN(n9071) );
  AND2_X1 U6592 ( .A1(n9692), .A2(n9934), .ZN(n5064) );
  NOR3_X1 U6593 ( .A1(n9691), .A2(n9962), .A3(n9690), .ZN(n5065) );
  INV_X1 U6594 ( .A(n9116), .ZN(n9626) );
  OR2_X1 U6595 ( .A1(n6929), .A2(n4388), .ZN(n5066) );
  OR2_X1 U6596 ( .A1(n10105), .A2(n7830), .ZN(n5067) );
  INV_X1 U6597 ( .A(n9584), .ZN(n8036) );
  NOR2_X1 U6598 ( .A1(n5686), .A2(n7328), .ZN(n5068) );
  NAND2_X1 U6599 ( .A1(n9117), .A2(n8035), .ZN(n9652) );
  OR2_X1 U6600 ( .A1(n6783), .A2(n6823), .ZN(n5069) );
  NAND2_X1 U6601 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  AND2_X1 U6602 ( .A1(n5947), .A2(n5941), .ZN(n5942) );
  NAND2_X1 U6603 ( .A1(n5943), .A2(n5942), .ZN(n5945) );
  INV_X1 U6604 ( .A(n9075), .ZN(n9141) );
  INV_X1 U6605 ( .A(n8729), .ZN(n5415) );
  AND2_X1 U6606 ( .A1(n9293), .A2(n9299), .ZN(n9264) );
  INV_X1 U6607 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6013) );
  OR2_X1 U6608 ( .A1(n5489), .A2(n5488), .ZN(n5491) );
  INV_X1 U6609 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5267) );
  INV_X1 U6610 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5618) );
  AND2_X1 U6611 ( .A1(n6556), .A2(n8956), .ZN(n6557) );
  INV_X1 U6612 ( .A(n6522), .ZN(n6518) );
  OR2_X1 U6613 ( .A1(n7046), .A2(n7042), .ZN(n6125) );
  INV_X1 U6614 ( .A(n8963), .ZN(n8024) );
  NOR2_X1 U6615 ( .A1(n8026), .A2(n9631), .ZN(n8155) );
  INV_X1 U6616 ( .A(n7138), .ZN(n7137) );
  OR2_X1 U6617 ( .A1(n5591), .A2(n5596), .ZN(n5733) );
  NAND2_X1 U6618 ( .A1(n5286), .A2(n10365), .ZN(n5298) );
  NOR2_X1 U6619 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6008) );
  INV_X1 U6620 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7828) );
  AND2_X1 U6621 ( .A1(n8834), .A2(n8708), .ZN(n5707) );
  NOR2_X2 U6622 ( .A1(n5042), .A2(n8858), .ZN(n7932) );
  XNOR2_X1 U6623 ( .A(n8788), .B(n8410), .ZN(n5989) );
  NAND2_X1 U6624 ( .A1(n5620), .A2(n5618), .ZN(n5648) );
  OAI21_X1 U6625 ( .B1(n6163), .B2(n7451), .A(n6118), .ZN(n6983) );
  NAND2_X1 U6626 ( .A1(n4391), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6109) );
  INV_X1 U6627 ( .A(n9637), .ZN(n9669) );
  AND2_X1 U6628 ( .A1(n6924), .A2(n7122), .ZN(n6926) );
  AND2_X1 U6629 ( .A1(n5556), .A2(n5530), .ZN(n5541) );
  NAND2_X1 U6630 ( .A1(n5321), .A2(n10211), .ZN(n5337) );
  INV_X1 U6631 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U6632 ( .A1(n7170), .A2(n7169), .ZN(n8271) );
  INV_X1 U6633 ( .A(n8315), .ZN(n7197) );
  OR2_X1 U6634 ( .A1(n8426), .A2(n8251), .ZN(n8402) );
  NAND2_X1 U6635 ( .A1(n5763), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5107) );
  INV_X1 U6636 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10379) );
  INV_X1 U6637 ( .A(n7624), .ZN(n7642) );
  AND2_X1 U6638 ( .A1(n5996), .A2(n5845), .ZN(n6974) );
  INV_X1 U6639 ( .A(n5989), .ZN(n5950) );
  INV_X1 U6640 ( .A(n10113), .ZN(n10097) );
  INV_X1 U6641 ( .A(n10015), .ZN(n9998) );
  AND2_X1 U6642 ( .A1(n6536), .A2(n6535), .ZN(n8921) );
  INV_X1 U6643 ( .A(n7084), .ZN(n6164) );
  INV_X1 U6644 ( .A(n9039), .ZN(n9013) );
  OR2_X1 U6645 ( .A1(n9934), .A2(n6897), .ZN(n6655) );
  INV_X1 U6646 ( .A(n9731), .ZN(n9545) );
  AND2_X1 U6647 ( .A1(n9106), .A2(n9111), .ZN(n9196) );
  OR2_X1 U6648 ( .A1(n9166), .A2(n9327), .ZN(n9633) );
  INV_X1 U6649 ( .A(n9490), .ZN(n9491) );
  INV_X1 U6650 ( .A(n9944), .ZN(n9935) );
  AND2_X1 U6651 ( .A1(n6893), .A2(n6892), .ZN(n9688) );
  NAND2_X1 U6652 ( .A1(n5417), .A2(n5377), .ZN(n5416) );
  INV_X1 U6653 ( .A(n7556), .ZN(n8321) );
  AND2_X1 U6654 ( .A1(n8415), .A2(n10015), .ZN(n8422) );
  AND4_X1 U6655 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n8208)
         );
  AND2_X1 U6656 ( .A1(n5667), .A2(n5666), .ZN(n6968) );
  INV_X1 U6657 ( .A(n9983), .ZN(n8510) );
  AND2_X1 U6658 ( .A1(n6692), .A2(n6688), .ZN(n9979) );
  INV_X1 U6659 ( .A(n8166), .ZN(n10029) );
  NAND2_X1 U6660 ( .A1(n5842), .A2(n7378), .ZN(n7328) );
  INV_X1 U6661 ( .A(n10031), .ZN(n8756) );
  AND2_X1 U6662 ( .A1(n5676), .A2(n5675), .ZN(n6955) );
  OR2_X1 U6663 ( .A1(n8783), .A2(n8774), .ZN(n8786) );
  AND2_X1 U6664 ( .A1(n8736), .A2(n10102), .ZN(n10085) );
  INV_X1 U6665 ( .A(n10085), .ZN(n10117) );
  XNOR2_X1 U6666 ( .A(n5650), .B(n5649), .ZN(n5674) );
  AND2_X1 U6667 ( .A1(n4461), .A2(n6652), .ZN(n9067) );
  AND2_X1 U6668 ( .A1(n6446), .A2(n6445), .ZN(n8933) );
  AND2_X1 U6669 ( .A1(n9133), .A2(n9137), .ZN(n9548) );
  INV_X1 U6670 ( .A(n7150), .ZN(n9185) );
  INV_X1 U6671 ( .A(n9688), .ZN(n9665) );
  INV_X1 U6672 ( .A(n9934), .ZN(n9965) );
  AND2_X1 U6673 ( .A1(n9688), .A2(n9939), .ZN(n9962) );
  AND2_X1 U6674 ( .A1(n6803), .A2(n6802), .ZN(n6921) );
  NAND2_X1 U6675 ( .A1(n6976), .A2(n6975), .ZN(n8426) );
  INV_X1 U6676 ( .A(n8592), .ZN(n8436) );
  INV_X1 U6677 ( .A(n8232), .ZN(n8613) );
  OR2_X1 U6678 ( .A1(n6714), .A2(n8900), .ZN(n9984) );
  INV_X1 U6679 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9872) );
  INV_X1 U6680 ( .A(n5731), .ZN(n5732) );
  OR2_X1 U6681 ( .A1(n8725), .A2(n8727), .ZN(n8845) );
  OR2_X1 U6682 ( .A1(n10036), .A2(n5718), .ZN(n8763) );
  INV_X2 U6683 ( .A(n10027), .ZN(n10036) );
  INV_X1 U6684 ( .A(n10142), .ZN(n10139) );
  OR2_X1 U6685 ( .A1(n10121), .A2(n6005), .ZN(n6006) );
  OR3_X1 U6686 ( .A1(n8868), .A2(n8867), .A3(n8866), .ZN(n8887) );
  INV_X1 U6687 ( .A(n10121), .ZN(n10119) );
  NOR2_X1 U6688 ( .A1(n10038), .A2(n10037), .ZN(n10039) );
  XNOR2_X1 U6689 ( .A(n5661), .B(n5660), .ZN(n7997) );
  INV_X1 U6690 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6772) );
  INV_X1 U6691 ( .A(n9706), .ZN(n8919) );
  INV_X1 U6692 ( .A(n9715), .ZN(n9503) );
  INV_X1 U6693 ( .A(n8986), .ZN(n9047) );
  INV_X1 U6694 ( .A(n9067), .ZN(n9348) );
  INV_X1 U6695 ( .A(n9630), .ZN(n9351) );
  OR2_X1 U6696 ( .A1(n6840), .A2(n8145), .ZN(n9893) );
  OR2_X1 U6697 ( .A1(P1_U3083), .A2(n6778), .ZN(n9923) );
  NAND2_X1 U6698 ( .A1(n7131), .A2(n7130), .ZN(n9645) );
  INV_X1 U6699 ( .A(n9977), .ZN(n9974) );
  AND2_X2 U6700 ( .A1(n6921), .A2(n6920), .ZN(n9977) );
  OR3_X1 U6701 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(n9822) );
  INV_X1 U6702 ( .A(n10175), .ZN(n10173) );
  AND2_X1 U6703 ( .A1(n9925), .A2(n9924), .ZN(n9926) );
  INV_X1 U6704 ( .A(n6618), .ZN(n9210) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7107) );
  INV_X1 U6706 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U6707 ( .A1(n6909), .A2(n10476), .ZN(n10475) );
  INV_X1 U6708 ( .A(n8449), .ZN(P2_U3966) );
  NAND2_X1 U6709 ( .A1(n5039), .A2(n5732), .ZN(P2_U3269) );
  NAND2_X1 U6710 ( .A1(n5072), .A2(n5071), .ZN(n5073) );
  NOR2_X2 U6711 ( .A1(n5403), .A2(n5073), .ZN(n5079) );
  NOR2_X2 U6712 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5076) );
  NOR2_X2 U6713 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5075) );
  NOR2_X2 U6714 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5074) );
  AND3_X2 U6715 ( .A1(n5076), .A2(n5075), .A3(n5074), .ZN(n5325) );
  NOR2_X1 U6716 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5078) );
  INV_X1 U6717 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5080) );
  INV_X2 U6718 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5668) );
  NOR2_X1 U6719 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5081) );
  INV_X2 U6720 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5660) );
  INV_X1 U6721 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5083) );
  OR2_X2 U6722 ( .A1(n8888), .A2(n8890), .ZN(n5085) );
  INV_X1 U6723 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5084) );
  XNOR2_X2 U6724 ( .A(n5085), .B(n5084), .ZN(n5089) );
  INV_X1 U6725 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5087) );
  AND2_X4 U6726 ( .A1(n5089), .A2(n8897), .ZN(n5787) );
  NAND2_X1 U6727 ( .A1(n5787), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6728 ( .A1(n5089), .A2(n5090), .ZN(n5254) );
  NAND2_X1 U6729 ( .A1(n5444), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5093) );
  AND2_X2 U6730 ( .A1(n8894), .A2(n5090), .ZN(n5193) );
  NAND2_X1 U6731 ( .A1(n5193), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5092) );
  AND2_X4 U6732 ( .A1(n8894), .A2(n8897), .ZN(n5763) );
  NAND2_X1 U6733 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  NAND2_X1 U6734 ( .A1(n5098), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6735 ( .A1(n4524), .A2(SI_0_), .ZN(n5100) );
  XNOR2_X1 U6736 ( .A(n5100), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8907) );
  XNOR2_X1 U6737 ( .A(n5102), .B(n5101), .ZN(n5114) );
  MUX2_X1 U6738 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8907), .S(n6686), .Z(n5681) );
  OR2_X2 U6739 ( .A1(n8451), .A2(n10046), .ZN(n7585) );
  NAND2_X1 U6740 ( .A1(n5787), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6741 ( .A1(n5444), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6742 ( .A1(n5193), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5106) );
  NAND4_X2 U6743 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5682)
         );
  INV_X1 U6744 ( .A(n5682), .ZN(n5124) );
  NAND2_X1 U6745 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5130) );
  AND2_X1 U6746 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6747 ( .A1(n5598), .A2(n5135), .ZN(n6115) );
  OAI21_X1 U6748 ( .B1(n5598), .B2(n5130), .A(n6115), .ZN(n5110) );
  INV_X1 U6749 ( .A(SI_1_), .ZN(n5134) );
  XNOR2_X1 U6750 ( .A(n5110), .B(n5134), .ZN(n5112) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4380), .Z(n5111) );
  INV_X1 U6752 ( .A(n6762), .ZN(n5113) );
  NAND2_X1 U6753 ( .A1(n5272), .A2(n5113), .ZN(n5122) );
  INV_X1 U6755 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6735) );
  AOI21_X1 U6756 ( .B1(n8138), .B2(n6691), .A(n5051), .ZN(n5115) );
  INV_X1 U6757 ( .A(n5115), .ZN(n5120) );
  NAND2_X1 U6758 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5116) );
  MUX2_X1 U6759 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5116), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5118) );
  NAND2_X1 U6760 ( .A1(n5118), .A2(n4823), .ZN(n6736) );
  INV_X1 U6761 ( .A(n6736), .ZN(n8452) );
  NAND3_X1 U6762 ( .A1(n8138), .A2(n6691), .A3(n8452), .ZN(n5119) );
  AND2_X1 U6763 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  AND2_X2 U6764 ( .A1(n5122), .A2(n5121), .ZN(n10051) );
  NAND2_X1 U6765 ( .A1(n7585), .A2(n5854), .ZN(n5125) );
  NAND2_X1 U6766 ( .A1(n5125), .A2(n5853), .ZN(n7531) );
  NAND2_X1 U6767 ( .A1(n5444), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6768 ( .A1(n5787), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6769 ( .A1(n5193), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5126) );
  NAND4_X4 U6770 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n10016)
         );
  AND3_X1 U6771 ( .A1(SI_1_), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5133) );
  AOI21_X1 U6772 ( .B1(n5134), .B2(n5130), .A(n6735), .ZN(n5132) );
  OAI21_X1 U6773 ( .B1(n5133), .B2(n5132), .A(n5131), .ZN(n5140) );
  INV_X1 U6774 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U6775 ( .A1(n6761), .A2(n5134), .ZN(n5136) );
  AOI22_X1 U6776 ( .A1(n5136), .A2(n5135), .B1(P2_DATAO_REG_1__SCAN_IN), .B2(
        SI_1_), .ZN(n5137) );
  INV_X1 U6777 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6778 ( .A1(n5138), .A2(n5598), .ZN(n5139) );
  INV_X1 U6779 ( .A(SI_2_), .ZN(n5151) );
  NAND2_X1 U6780 ( .A1(n5272), .A2(n5142), .ZN(n5146) );
  NAND2_X1 U6781 ( .A1(n5186), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5145) );
  INV_X1 U6782 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8890) );
  NOR2_X1 U6783 ( .A1(n5143), .A2(n5406), .ZN(n7248) );
  NAND2_X1 U6784 ( .A1(n6718), .A2(n7248), .ZN(n5144) );
  AND3_X2 U6785 ( .A1(n5146), .A2(n5145), .A3(n5144), .ZN(n10057) );
  NAND2_X2 U6786 ( .A1(n8239), .A2(n7534), .ZN(n5855) );
  NAND2_X1 U6787 ( .A1(n10016), .A2(n10057), .ZN(n5857) );
  NAND2_X2 U6788 ( .A1(n5855), .A2(n5857), .ZN(n7530) );
  NAND2_X1 U6789 ( .A1(n5444), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6790 ( .A1(n5193), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6791 ( .A1(n5787), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6792 ( .A1(n5763), .A2(n8246), .ZN(n5147) );
  NAND4_X1 U6793 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n8450)
         );
  INV_X1 U6794 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U6795 ( .A1(n4380), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5152) );
  OAI211_X1 U6796 ( .C1(n5598), .C2(n8045), .A(n5152), .B(n5151), .ZN(n5153)
         );
  INV_X1 U6797 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U6798 ( .A1(n4380), .A2(n10304), .ZN(n5154) );
  OAI211_X1 U6799 ( .C1(n5598), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5154), .B(
        SI_2_), .ZN(n5155) );
  INV_X1 U6800 ( .A(SI_3_), .ZN(n5157) );
  XNOR2_X1 U6801 ( .A(n5171), .B(n5157), .ZN(n5169) );
  XNOR2_X1 U6802 ( .A(n5170), .B(n5169), .ZN(n6749) );
  INV_X1 U6803 ( .A(n6749), .ZN(n5158) );
  NAND2_X1 U6804 ( .A1(n5582), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6805 ( .A1(n6718), .A2(n7234), .ZN(n5160) );
  OR2_X1 U6806 ( .A1(n8450), .A2(n10032), .ZN(n5841) );
  NAND2_X1 U6807 ( .A1(n5164), .A2(n5841), .ZN(n7327) );
  INV_X1 U6808 ( .A(n7327), .ZN(n5179) );
  OAI21_X1 U6809 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5195), .ZN(n7324) );
  INV_X1 U6810 ( .A(n7324), .ZN(n8356) );
  NAND2_X1 U6811 ( .A1(n5763), .A2(n8356), .ZN(n5168) );
  NAND2_X1 U6812 ( .A1(n5786), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6813 ( .A1(n5193), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6814 ( .A1(n5787), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6815 ( .A1(n5171), .A2(SI_3_), .ZN(n5172) );
  XNOR2_X1 U6816 ( .A(n5182), .B(n5180), .ZN(n6733) );
  NAND2_X1 U6817 ( .A1(n6733), .A2(n5272), .ZN(n5178) );
  NAND2_X1 U6818 ( .A1(n5582), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6819 ( .A1(n5187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5175) );
  XNOR2_X1 U6820 ( .A(n5175), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7276) );
  NAND2_X1 U6821 ( .A1(n6718), .A2(n7276), .ZN(n5176) );
  INV_X1 U6822 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6823 ( .A1(n5183), .A2(SI_4_), .ZN(n5184) );
  INV_X1 U6824 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6739) );
  INV_X1 U6825 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6744) );
  MUX2_X1 U6826 ( .A(n6739), .B(n6744), .S(n4380), .Z(n5203) );
  XNOR2_X1 U6827 ( .A(n5203), .B(SI_5_), .ZN(n5201) );
  INV_X1 U6828 ( .A(n5201), .ZN(n5185) );
  NAND2_X1 U6829 ( .A1(n6737), .A2(n5272), .ZN(n5192) );
  NAND2_X1 U6830 ( .A1(n5189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5188) );
  MUX2_X1 U6831 ( .A(n5188), .B(P2_IR_REG_31__SCAN_IN), .S(n10348), .Z(n5190)
         );
  NAND2_X1 U6832 ( .A1(n5190), .A2(n5324), .ZN(n6738) );
  INV_X1 U6833 ( .A(n6738), .ZN(n7262) );
  AOI22_X1 U6834 ( .A1(n5582), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6718), .B2(
        n7262), .ZN(n5191) );
  NAND2_X1 U6835 ( .A1(n5193), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6836 ( .A1(n5786), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5199) );
  INV_X1 U6837 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6838 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  AND2_X1 U6839 ( .A1(n5209), .A2(n5196), .ZN(n8320) );
  NAND2_X1 U6840 ( .A1(n5763), .A2(n8320), .ZN(n5198) );
  NAND2_X1 U6841 ( .A1(n5787), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6842 ( .A1(n7556), .A2(n8448), .ZN(n5863) );
  NAND2_X1 U6843 ( .A1(n10018), .A2(n10070), .ZN(n7378) );
  INV_X1 U6844 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6845 ( .A1(n5204), .A2(SI_5_), .ZN(n5234) );
  NAND2_X1 U6846 ( .A1(n5235), .A2(n5234), .ZN(n5220) );
  MUX2_X1 U6847 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4380), .Z(n5236) );
  XNOR2_X1 U6848 ( .A(n5236), .B(SI_6_), .ZN(n5218) );
  XNOR2_X1 U6849 ( .A(n5220), .B(n5218), .ZN(n6740) );
  NAND2_X1 U6850 ( .A1(n6740), .A2(n5272), .ZN(n5207) );
  NAND2_X1 U6851 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6852 ( .A(n5205), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7221) );
  AOI22_X1 U6853 ( .A1(n5582), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6718), .B2(
        n7221), .ZN(n5206) );
  NAND2_X1 U6854 ( .A1(n5791), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6855 ( .A1(n5786), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5213) );
  INV_X1 U6856 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6857 ( .A1(n5209), .A2(n5208), .ZN(n5210) );
  AND2_X1 U6858 ( .A1(n5226), .A2(n5210), .ZN(n8395) );
  NAND2_X1 U6859 ( .A1(n5763), .A2(n8395), .ZN(n5212) );
  NAND2_X1 U6860 ( .A1(n5787), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5211) );
  AND4_X2 U6861 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n7210)
         );
  AND2_X1 U6863 ( .A1(n7549), .A2(n7561), .ZN(n5215) );
  NAND2_X1 U6864 ( .A1(n5217), .A2(n7210), .ZN(n5869) );
  INV_X1 U6865 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U6866 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NAND2_X1 U6867 ( .A1(n5236), .A2(SI_6_), .ZN(n5233) );
  NAND2_X1 U6868 ( .A1(n5221), .A2(n5233), .ZN(n5222) );
  MUX2_X1 U6869 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5598), .Z(n5240) );
  XNOR2_X1 U6870 ( .A(n5240), .B(SI_7_), .ZN(n5238) );
  NAND2_X1 U6871 ( .A1(n6752), .A2(n5272), .ZN(n5225) );
  NAND2_X1 U6872 ( .A1(n5248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5223) );
  XNOR2_X1 U6873 ( .A(n5223), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6702) );
  AOI22_X1 U6874 ( .A1(n5582), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6718), .B2(
        n6702), .ZN(n5224) );
  NAND2_X1 U6875 ( .A1(n5225), .A2(n5224), .ZN(n10081) );
  NAND2_X1 U6876 ( .A1(n5791), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6877 ( .A1(n5786), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6878 ( .A1(n5226), .A2(n10227), .ZN(n5227) );
  AND2_X1 U6879 ( .A1(n5257), .A2(n5227), .ZN(n7303) );
  NAND2_X1 U6880 ( .A1(n5763), .A2(n7303), .ZN(n5229) );
  NAND2_X1 U6881 ( .A1(n5787), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6882 ( .A1(n10081), .A2(n8391), .ZN(n5871) );
  NAND2_X1 U6883 ( .A1(n5232), .A2(n5871), .ZN(n7617) );
  NOR2_X1 U6884 ( .A1(n5236), .A2(SI_6_), .ZN(n5237) );
  NOR2_X1 U6885 ( .A1(n5238), .A2(n5237), .ZN(n5239) );
  NAND2_X1 U6886 ( .A1(n5240), .A2(SI_7_), .ZN(n5241) );
  INV_X1 U6887 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5243) );
  MUX2_X1 U6888 ( .A(n6756), .B(n5243), .S(n4380), .Z(n5245) );
  INV_X1 U6889 ( .A(SI_8_), .ZN(n5244) );
  INV_X1 U6890 ( .A(n5245), .ZN(n5246) );
  NAND2_X1 U6891 ( .A1(n5246), .A2(SI_8_), .ZN(n5247) );
  NAND2_X1 U6892 ( .A1(n5250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5249) );
  MUX2_X1 U6893 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5249), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5251) );
  NAND2_X1 U6894 ( .A1(n5251), .A2(n5289), .ZN(n6754) );
  INV_X1 U6895 ( .A(n6754), .ZN(n8465) );
  AOI22_X1 U6896 ( .A1(n6718), .A2(n8465), .B1(n5582), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6897 ( .A1(n5791), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6898 ( .A1(n5786), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5262) );
  INV_X1 U6899 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6900 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6901 ( .A1(n5276), .A2(n5258), .ZN(n7626) );
  INV_X1 U6902 ( .A(n7626), .ZN(n5259) );
  NAND2_X1 U6903 ( .A1(n5763), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U6904 ( .A1(n5787), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6905 ( .A1(n10088), .A2(n7634), .ZN(n5876) );
  NAND2_X1 U6906 ( .A1(n10088), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U6907 ( .A1(n5876), .A2(n7636), .ZN(n5693) );
  OR2_X1 U6908 ( .A1(n10081), .A2(n8391), .ZN(n7616) );
  AND2_X1 U6909 ( .A1(n7619), .A2(n7616), .ZN(n5264) );
  NAND2_X1 U6910 ( .A1(n7638), .A2(n7636), .ZN(n5283) );
  MUX2_X1 U6911 ( .A(n6765), .B(n5267), .S(n5598), .Z(n5269) );
  INV_X1 U6912 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6913 ( .A1(n5270), .A2(SI_9_), .ZN(n5271) );
  NAND2_X1 U6914 ( .A1(n6759), .A2(n5272), .ZN(n5275) );
  NAND2_X1 U6915 ( .A1(n5289), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  AOI22_X1 U6916 ( .A1(n6718), .A2(n8482), .B1(n5582), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6917 ( .A1(n5791), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6918 ( .A1(n5444), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6919 ( .A1(n5276), .A2(n7828), .ZN(n5277) );
  AND2_X1 U6920 ( .A1(n5307), .A2(n5277), .ZN(n7829) );
  NAND2_X1 U6921 ( .A1(n5763), .A2(n7829), .ZN(n5279) );
  NAND2_X1 U6922 ( .A1(n5787), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6923 ( .A1(n10095), .A2(n9997), .ZN(n9993) );
  INV_X1 U6924 ( .A(n7637), .ZN(n5282) );
  MUX2_X1 U6925 ( .A(n6772), .B(n6769), .S(n4380), .Z(n5286) );
  INV_X1 U6926 ( .A(n5286), .ZN(n5287) );
  NAND2_X1 U6927 ( .A1(n5287), .A2(SI_10_), .ZN(n5288) );
  XNOR2_X1 U6928 ( .A(n5301), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8495) );
  AOI22_X1 U6929 ( .A1(n8495), .A2(n6718), .B1(n5582), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6930 ( .A1(n5786), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5295) );
  XNOR2_X1 U6931 ( .A(n5307), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U6932 ( .A1(n5763), .A2(n10003), .ZN(n5294) );
  NAND2_X1 U6933 ( .A1(n5787), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6934 ( .A1(n5791), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6935 ( .A1(n7696), .A2(n7830), .ZN(n5880) );
  AND2_X1 U6936 ( .A1(n5880), .A2(n9993), .ZN(n5884) );
  MUX2_X1 U6937 ( .A(n6777), .B(n5299), .S(n5598), .Z(n5317) );
  XNOR2_X1 U6938 ( .A(n5320), .B(n5316), .ZN(n6773) );
  INV_X1 U6939 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6940 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  NAND2_X1 U6941 ( .A1(n5791), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6942 ( .A1(n5786), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5313) );
  INV_X1 U6943 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5306) );
  INV_X1 U6944 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7284) );
  OAI21_X1 U6945 ( .B1(n5307), .B2(n5306), .A(n7284), .ZN(n5310) );
  AND2_X1 U6946 ( .A1(n5310), .A2(n5330), .ZN(n7810) );
  NAND2_X1 U6947 ( .A1(n5763), .A2(n7810), .ZN(n5312) );
  NAND2_X1 U6948 ( .A1(n5787), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5311) );
  INV_X1 U6949 ( .A(n5887), .ZN(n5315) );
  NAND2_X1 U6950 ( .A1(n7796), .A2(n9999), .ZN(n5881) );
  INV_X1 U6951 ( .A(n5317), .ZN(n5318) );
  MUX2_X1 U6952 ( .A(n6797), .B(n6795), .S(n4380), .Z(n5321) );
  INV_X1 U6953 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6954 ( .A1(n5322), .A2(SI_12_), .ZN(n5323) );
  INV_X1 U6955 ( .A(n5324), .ZN(n5326) );
  NAND2_X1 U6956 ( .A1(n5326), .A2(n5325), .ZN(n5347) );
  NAND2_X1 U6957 ( .A1(n5347), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5327) );
  XNOR2_X1 U6958 ( .A(n5327), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6708) );
  AOI22_X1 U6959 ( .A1(n5582), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6718), .B2(
        n6708), .ZN(n5328) );
  NAND2_X1 U6960 ( .A1(n5791), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6961 ( .A1(n5444), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6962 ( .A1(n5330), .A2(n10379), .ZN(n5331) );
  AND2_X1 U6963 ( .A1(n5363), .A2(n5331), .ZN(n7908) );
  NAND2_X1 U6964 ( .A1(n5763), .A2(n7908), .ZN(n5333) );
  NAND2_X1 U6965 ( .A1(n5787), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6966 ( .A1(n7893), .A2(n7969), .ZN(n5882) );
  INV_X1 U6967 ( .A(n7864), .ZN(n5336) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5340) );
  MUX2_X1 U6969 ( .A(n6845), .B(n5340), .S(n4380), .Z(n5342) );
  INV_X1 U6970 ( .A(SI_13_), .ZN(n5341) );
  INV_X1 U6971 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6972 ( .A1(n5343), .A2(SI_13_), .ZN(n5344) );
  NAND2_X1 U6973 ( .A1(n5357), .A2(n5052), .ZN(n5346) );
  MUX2_X1 U6974 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5598), .Z(n5371) );
  XNOR2_X1 U6975 ( .A(n5373), .B(n5370), .ZN(n6846) );
  NAND2_X1 U6976 ( .A1(n5348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5379) );
  XNOR2_X1 U6977 ( .A(n5379), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7483) );
  AOI22_X1 U6978 ( .A1(n6718), .A2(n7483), .B1(n5582), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6979 ( .A1(n5791), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5356) );
  INV_X1 U6980 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6981 ( .A1(n5365), .A2(n5351), .ZN(n5352) );
  AND2_X1 U6982 ( .A1(n5388), .A2(n5352), .ZN(n8212) );
  NAND2_X1 U6983 ( .A1(n5763), .A2(n8212), .ZN(n5355) );
  NAND2_X1 U6984 ( .A1(n5444), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6985 ( .A1(n5787), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6986 ( .A1(n5358), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5359) );
  XNOR2_X1 U6987 ( .A(n5359), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U6988 ( .A1(n5582), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6718), .B2(
        n6710), .ZN(n5360) );
  NAND2_X1 U6989 ( .A1(n5791), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6990 ( .A1(n5786), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5368) );
  INV_X1 U6991 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6992 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  AND2_X1 U6993 ( .A1(n5365), .A2(n5364), .ZN(n7972) );
  NAND2_X1 U6994 ( .A1(n5763), .A2(n7972), .ZN(n5367) );
  NAND2_X1 U6995 ( .A1(n5787), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6996 ( .A1(n5371), .A2(SI_14_), .ZN(n5372) );
  INV_X1 U6997 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7026) );
  MUX2_X1 U6998 ( .A(n10176), .B(n7026), .S(n5598), .Z(n5375) );
  INV_X1 U6999 ( .A(SI_15_), .ZN(n5374) );
  INV_X1 U7000 ( .A(n5375), .ZN(n5376) );
  NAND2_X1 U7001 ( .A1(n5376), .A2(SI_15_), .ZN(n5377) );
  INV_X1 U7002 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U7003 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  NAND2_X1 U7004 ( .A1(n5380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5381) );
  XNOR2_X1 U7005 ( .A(n5381), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7767) );
  AOI22_X1 U7006 ( .A1(n7767), .A2(n6718), .B1(n5582), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U7007 ( .A1(n5791), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U7008 ( .A1(n5786), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5384) );
  AND2_X1 U7009 ( .A1(n5385), .A2(n5384), .ZN(n5392) );
  INV_X1 U7010 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U7011 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U7012 ( .A1(n5410), .A2(n5389), .ZN(n8754) );
  OR2_X1 U7013 ( .A1(n8754), .A2(n5609), .ZN(n5391) );
  NAND2_X1 U7014 ( .A1(n5787), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U7015 ( .A1(n5704), .A2(n8731), .ZN(n5908) );
  NAND2_X1 U7016 ( .A1(n5909), .A2(n5908), .ZN(n8747) );
  NAND2_X1 U7017 ( .A1(n8854), .A2(n8048), .ZN(n5838) );
  NAND2_X1 U7018 ( .A1(n8858), .A2(n8208), .ZN(n7977) );
  NAND2_X1 U7019 ( .A1(n5838), .A2(n7977), .ZN(n5393) );
  NAND2_X1 U7020 ( .A1(n5393), .A2(n8745), .ZN(n5394) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5396) );
  MUX2_X1 U7022 ( .A(n5396), .B(n7107), .S(n5598), .Z(n5398) );
  INV_X1 U7023 ( .A(SI_16_), .ZN(n5397) );
  INV_X1 U7024 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U7025 ( .A1(n5399), .A2(SI_16_), .ZN(n5400) );
  INV_X1 U7026 ( .A(n5418), .ZN(n5401) );
  INV_X1 U7027 ( .A(n5403), .ZN(n5404) );
  NAND4_X1 U7028 ( .A1(n5325), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n5424)
         );
  NAND2_X1 U7029 ( .A1(n5424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U7030 ( .A(n5407), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8509) );
  AOI22_X1 U7031 ( .A1(n5582), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6718), .B2(
        n8509), .ZN(n5408) );
  INV_X1 U7032 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U7033 ( .A1(n5410), .A2(n10333), .ZN(n5411) );
  AND2_X1 U7034 ( .A1(n5428), .A2(n5411), .ZN(n8739) );
  NAND2_X1 U7035 ( .A1(n8739), .A2(n5763), .ZN(n5414) );
  AOI22_X1 U7036 ( .A1(n5791), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n5786), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7037 ( .A1(n5787), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5412) );
  OR2_X1 U7038 ( .A1(n8842), .A2(n8332), .ZN(n5837) );
  NAND2_X1 U7039 ( .A1(n8842), .A2(n8332), .ZN(n8705) );
  MUX2_X1 U7040 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5598), .Z(n5438) );
  INV_X1 U7041 ( .A(SI_17_), .ZN(n5423) );
  XNOR2_X1 U7042 ( .A(n5436), .B(n5437), .ZN(n7108) );
  OAI21_X1 U7043 ( .B1(n5424), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U7044 ( .A(n5425), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8109) );
  AOI22_X1 U7045 ( .A1(n5582), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6718), .B2(
        n8109), .ZN(n5426) );
  NAND2_X1 U7046 ( .A1(n5428), .A2(n4613), .ZN(n5429) );
  NAND2_X1 U7047 ( .A1(n5442), .A2(n5429), .ZN(n8715) );
  OR2_X1 U7048 ( .A1(n8715), .A2(n5609), .ZN(n5432) );
  AOI22_X1 U7049 ( .A1(n5791), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5786), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7050 ( .A1(n5787), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7051 ( .A1(n8838), .A2(n8732), .ZN(n5834) );
  INV_X1 U7052 ( .A(n8705), .ZN(n5433) );
  NOR2_X1 U7053 ( .A1(n8711), .A2(n5433), .ZN(n5434) );
  NAND2_X1 U7054 ( .A1(n5435), .A2(n5836), .ZN(n8693) );
  MUX2_X1 U7055 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5598), .Z(n5452) );
  XNOR2_X1 U7056 ( .A(n5451), .B(n5450), .ZN(n7332) );
  NAND2_X1 U7057 ( .A1(n7332), .A2(n4689), .ZN(n5441) );
  NAND2_X1 U7058 ( .A1(n5458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U7059 ( .A(n5439), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8110) );
  AOI22_X1 U7060 ( .A1(n5582), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6718), .B2(
        n8110), .ZN(n5440) );
  NAND2_X1 U7061 ( .A1(n5442), .A2(n4614), .ZN(n5443) );
  NAND2_X1 U7062 ( .A1(n5462), .A2(n5443), .ZN(n8086) );
  OR2_X1 U7063 ( .A1(n8086), .A2(n5609), .ZN(n5449) );
  INV_X1 U7064 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10256) );
  INV_X1 U7065 ( .A(n5787), .ZN(n5760) );
  NAND2_X1 U7066 ( .A1(n5791), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U7067 ( .A1(n5444), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5445) );
  OAI211_X1 U7068 ( .C1(n10256), .C2(n5760), .A(n5446), .B(n5445), .ZN(n5447)
         );
  INV_X1 U7069 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U7070 ( .A1(n8834), .A2(n8331), .ZN(n5918) );
  NAND2_X1 U7071 ( .A1(n5452), .A2(SI_18_), .ZN(n5453) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7492) );
  INV_X1 U7073 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7490) );
  MUX2_X1 U7074 ( .A(n7492), .B(n7490), .S(n4380), .Z(n5455) );
  INV_X1 U7075 ( .A(SI_19_), .ZN(n10331) );
  NAND2_X1 U7076 ( .A1(n5455), .A2(n10331), .ZN(n5488) );
  INV_X1 U7077 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U7078 ( .A1(n5456), .A2(SI_19_), .ZN(n5457) );
  NAND2_X1 U7079 ( .A1(n5488), .A2(n5457), .ZN(n5487) );
  XNOR2_X1 U7080 ( .A(n5492), .B(n5487), .ZN(n7489) );
  NAND2_X1 U7081 ( .A1(n7489), .A2(n4689), .ZN(n5460) );
  AOI22_X1 U7082 ( .A1(n5582), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5619), .B2(
        n6718), .ZN(n5459) );
  INV_X1 U7083 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7084 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  NAND2_X1 U7085 ( .A1(n5480), .A2(n5463), .ZN(n8677) );
  OR2_X1 U7086 ( .A1(n8677), .A2(n5609), .ZN(n5468) );
  INV_X1 U7087 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U7088 ( .A1(n5786), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7089 ( .A1(n5791), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5464) );
  OAI211_X1 U7090 ( .C1(n10422), .C2(n5760), .A(n5465), .B(n5464), .ZN(n5466)
         );
  INV_X1 U7091 ( .A(n5466), .ZN(n5467) );
  OR2_X1 U7092 ( .A1(n8828), .A2(n8695), .ZN(n5920) );
  NAND2_X1 U7093 ( .A1(n8828), .A2(n8695), .ZN(n5922) );
  NAND2_X1 U7094 ( .A1(n5920), .A2(n5922), .ZN(n5708) );
  INV_X1 U7095 ( .A(n8681), .ZN(n5469) );
  NOR2_X1 U7096 ( .A1(n5708), .A2(n5469), .ZN(n5470) );
  OR2_X1 U7097 ( .A1(n5492), .A2(n5487), .ZN(n5471) );
  NAND2_X1 U7098 ( .A1(n5471), .A2(n5488), .ZN(n5477) );
  INV_X1 U7099 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7650) );
  INV_X1 U7100 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7651) );
  MUX2_X1 U7101 ( .A(n7650), .B(n7651), .S(n5598), .Z(n5473) );
  INV_X1 U7102 ( .A(SI_20_), .ZN(n5472) );
  INV_X1 U7103 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U7104 ( .A1(n5474), .A2(SI_20_), .ZN(n5475) );
  INV_X1 U7105 ( .A(n5489), .ZN(n5476) );
  NAND2_X1 U7106 ( .A1(n7648), .A2(n4689), .ZN(n5479) );
  NAND2_X1 U7107 ( .A1(n5582), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5478) );
  INV_X1 U7108 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U7109 ( .A1(n5480), .A2(n8368), .ZN(n5481) );
  NAND2_X1 U7110 ( .A1(n5515), .A2(n5481), .ZN(n8369) );
  INV_X1 U7111 ( .A(n8369), .ZN(n8662) );
  NAND2_X1 U7112 ( .A1(n8662), .A2(n5763), .ZN(n5486) );
  INV_X1 U7113 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U7114 ( .A1(n5787), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7115 ( .A1(n5786), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U7116 ( .C1(n5790), .C2(n10205), .A(n5483), .B(n5482), .ZN(n5484)
         );
  INV_X1 U7117 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U7118 ( .A1(n8822), .A2(n8283), .ZN(n5923) );
  MUX2_X1 U7119 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4380), .Z(n5503) );
  INV_X1 U7120 ( .A(SI_21_), .ZN(n10259) );
  XNOR2_X1 U7121 ( .A(n5503), .B(n10259), .ZN(n5502) );
  XNOR2_X1 U7122 ( .A(n5506), .B(n5502), .ZN(n7728) );
  NAND2_X1 U7123 ( .A1(n7728), .A2(n4689), .ZN(n5494) );
  NAND2_X1 U7124 ( .A1(n5186), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5493) );
  XNOR2_X1 U7125 ( .A(n5515), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7126 ( .A1(n8648), .A2(n5763), .ZN(n5500) );
  INV_X1 U7127 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7128 ( .A1(n5786), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7129 ( .A1(n5791), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U7130 ( .C1(n5760), .C2(n5497), .A(n5496), .B(n5495), .ZN(n5498)
         );
  INV_X1 U7131 ( .A(n5498), .ZN(n5499) );
  XOR2_X1 U7132 ( .A(n8650), .B(n8638), .Z(n5986) );
  NAND2_X1 U7133 ( .A1(n8651), .A2(n8653), .ZN(n5501) );
  NAND2_X1 U7134 ( .A1(n8817), .A2(n8638), .ZN(n5928) );
  NAND2_X1 U7135 ( .A1(n5501), .A2(n5928), .ZN(n8635) );
  INV_X1 U7136 ( .A(n5502), .ZN(n5505) );
  NAND2_X1 U7137 ( .A1(n5503), .A2(SI_21_), .ZN(n5504) );
  INV_X1 U7138 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8092) );
  INV_X1 U7139 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7889) );
  MUX2_X1 U7140 ( .A(n8092), .B(n7889), .S(n4380), .Z(n5508) );
  INV_X1 U7141 ( .A(SI_22_), .ZN(n5507) );
  INV_X1 U7142 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7143 ( .A1(n5509), .A2(SI_22_), .ZN(n5510) );
  XNOR2_X1 U7144 ( .A(n5525), .B(n5524), .ZN(n7888) );
  NAND2_X1 U7145 ( .A1(n7888), .A2(n4689), .ZN(n5512) );
  NAND2_X1 U7146 ( .A1(n5582), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5511) );
  AND2_X1 U7147 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5513) );
  INV_X1 U7148 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8280) );
  INV_X1 U7149 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8382) );
  OAI21_X1 U7150 ( .B1(n5515), .B2(n8280), .A(n8382), .ZN(n5516) );
  NAND2_X1 U7151 ( .A1(n5533), .A2(n5516), .ZN(n8631) );
  OR2_X1 U7152 ( .A1(n8631), .A2(n5609), .ZN(n5522) );
  INV_X1 U7153 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7154 ( .A1(n5791), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7155 ( .A1(n5786), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5517) );
  OAI211_X1 U7156 ( .C1(n5519), .C2(n5760), .A(n5518), .B(n5517), .ZN(n5520)
         );
  INV_X1 U7157 ( .A(n5520), .ZN(n5521) );
  NAND2_X1 U7158 ( .A1(n8812), .A2(n8282), .ZN(n5828) );
  NAND2_X1 U7159 ( .A1(n5929), .A2(n5828), .ZN(n8637) );
  INV_X1 U7160 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10300) );
  INV_X1 U7161 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5526) );
  MUX2_X1 U7162 ( .A(n10300), .B(n5526), .S(n5598), .Z(n5528) );
  INV_X1 U7163 ( .A(SI_23_), .ZN(n5527) );
  NAND2_X1 U7164 ( .A1(n5528), .A2(n5527), .ZN(n5556) );
  INV_X1 U7165 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U7166 ( .A1(n5529), .A2(SI_23_), .ZN(n5530) );
  NAND2_X1 U7167 ( .A1(n6523), .A2(n4689), .ZN(n5532) );
  NAND2_X1 U7168 ( .A1(n5582), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5531) );
  INV_X1 U7169 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U7170 ( .A1(n5533), .A2(n8231), .ZN(n5534) );
  NAND2_X1 U7171 ( .A1(n5547), .A2(n5534), .ZN(n8621) );
  OR2_X1 U7172 ( .A1(n8621), .A2(n5609), .ZN(n5539) );
  INV_X1 U7173 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U7174 ( .A1(n5791), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U7175 ( .A1(n5787), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U7176 ( .C1(n5254), .C2(n10210), .A(n5536), .B(n5535), .ZN(n5537)
         );
  INV_X1 U7177 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U7178 ( .A1(n8807), .A2(n8639), .ZN(n5830) );
  INV_X1 U7179 ( .A(n5830), .ZN(n5540) );
  NAND2_X1 U7180 ( .A1(n5558), .A2(n5556), .ZN(n5544) );
  MUX2_X1 U7181 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4380), .Z(n5559) );
  INV_X1 U7182 ( .A(SI_24_), .ZN(n5543) );
  XNOR2_X1 U7183 ( .A(n5559), .B(n5543), .ZN(n5555) );
  NAND2_X1 U7184 ( .A1(n7992), .A2(n4689), .ZN(n5546) );
  NAND2_X1 U7185 ( .A1(n5582), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5545) );
  INV_X1 U7186 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U7187 ( .A1(n5547), .A2(n8345), .ZN(n5548) );
  AND2_X1 U7188 ( .A1(n5567), .A2(n5548), .ZN(n8602) );
  NAND2_X1 U7189 ( .A1(n8602), .A2(n5763), .ZN(n5554) );
  INV_X1 U7190 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7191 ( .A1(n5786), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7192 ( .A1(n5787), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5549) );
  OAI211_X1 U7193 ( .C1(n5790), .C2(n5551), .A(n5550), .B(n5549), .ZN(n5552)
         );
  INV_X1 U7194 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U7195 ( .A1(n8801), .A2(n8232), .ZN(n5937) );
  NAND2_X1 U7196 ( .A1(n5559), .A2(SI_24_), .ZN(n5735) );
  INV_X1 U7197 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8000) );
  INV_X1 U7198 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8003) );
  MUX2_X1 U7199 ( .A(n8000), .B(n8003), .S(n5598), .Z(n5561) );
  INV_X1 U7200 ( .A(SI_25_), .ZN(n5560) );
  NAND2_X1 U7201 ( .A1(n5561), .A2(n5560), .ZN(n5594) );
  INV_X1 U7202 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7203 ( .A1(n5562), .A2(SI_25_), .ZN(n5563) );
  NAND2_X1 U7204 ( .A1(n5594), .A2(n5563), .ZN(n5591) );
  NAND2_X1 U7205 ( .A1(n5582), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7206 ( .A1(n5567), .A2(n4609), .ZN(n5568) );
  NAND2_X1 U7207 ( .A1(n5585), .A2(n5568), .ZN(n8586) );
  INV_X1 U7208 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7209 ( .A1(n5791), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7210 ( .A1(n5786), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U7211 ( .C1(n5571), .C2(n5760), .A(n5570), .B(n5569), .ZN(n5572)
         );
  INV_X1 U7212 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7213 ( .A1(n8799), .A2(n8592), .ZN(n5748) );
  NAND2_X1 U7214 ( .A1(n8582), .A2(n4433), .ZN(n8581) );
  INV_X1 U7215 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5576) );
  INV_X1 U7216 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9838) );
  MUX2_X1 U7217 ( .A(n5576), .B(n9838), .S(n4380), .Z(n5578) );
  INV_X1 U7218 ( .A(SI_26_), .ZN(n5577) );
  NAND2_X1 U7219 ( .A1(n5578), .A2(n5577), .ZN(n5593) );
  INV_X1 U7220 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7221 ( .A1(n5579), .A2(SI_26_), .ZN(n5590) );
  AND2_X1 U7222 ( .A1(n5593), .A2(n5590), .ZN(n5580) );
  NAND2_X1 U7223 ( .A1(n8902), .A2(n4689), .ZN(n5584) );
  NAND2_X1 U7224 ( .A1(n5582), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5583) );
  INV_X1 U7225 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U7226 ( .A1(n5585), .A2(n8411), .ZN(n5586) );
  INV_X1 U7227 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U7228 ( .A1(n5791), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7229 ( .A1(n5786), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5587) );
  OAI211_X1 U7230 ( .C1(n10247), .C2(n5760), .A(n5588), .B(n5587), .ZN(n5589)
         );
  NAND3_X1 U7231 ( .A1(n8581), .A2(n8568), .A3(n8566), .ZN(n8567) );
  NAND2_X1 U7232 ( .A1(n8567), .A2(n5944), .ZN(n5616) );
  INV_X1 U7233 ( .A(n5590), .ZN(n5596) );
  AND2_X1 U7234 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  INV_X1 U7235 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5599) );
  INV_X1 U7236 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9836) );
  MUX2_X1 U7237 ( .A(n5599), .B(n9836), .S(n5598), .Z(n5600) );
  INV_X1 U7238 ( .A(SI_27_), .ZN(n10229) );
  NAND2_X1 U7239 ( .A1(n5600), .A2(n10229), .ZN(n5742) );
  INV_X1 U7240 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7241 ( .A1(n5601), .A2(SI_27_), .ZN(n5602) );
  NAND2_X1 U7242 ( .A1(n5742), .A2(n5602), .ZN(n5739) );
  INV_X1 U7243 ( .A(n5739), .ZN(n5603) );
  NAND2_X1 U7244 ( .A1(n5582), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7245 ( .A1(n5607), .A2(n4610), .ZN(n5608) );
  NAND2_X1 U7246 ( .A1(n5629), .A2(n5608), .ZN(n8203) );
  INV_X1 U7247 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7248 ( .A1(n5787), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7249 ( .A1(n5786), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5610) );
  OAI211_X1 U7250 ( .C1(n5790), .C2(n5612), .A(n5611), .B(n5610), .ZN(n5613)
         );
  INV_X1 U7251 ( .A(n5613), .ZN(n5614) );
  XNOR2_X1 U7252 ( .A(n5616), .B(n5950), .ZN(n5638) );
  XNOR2_X2 U7253 ( .A(n5657), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7254 ( .A1(n5678), .A2(n5619), .ZN(n7166) );
  INV_X1 U7255 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7256 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  NAND2_X1 U7257 ( .A1(n5625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7258 ( .A1(n5845), .A2(n5978), .ZN(n5821) );
  INV_X1 U7259 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7260 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  INV_X1 U7261 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7262 ( .A1(n5787), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7263 ( .A1(n5786), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5631) );
  OAI211_X1 U7264 ( .C1(n5790), .C2(n5633), .A(n5632), .B(n5631), .ZN(n5634)
         );
  INV_X1 U7265 ( .A(n6974), .ZN(n5715) );
  INV_X1 U7266 ( .A(n6691), .ZN(n5635) );
  OR2_X1 U7267 ( .A1(n8543), .A2(n10000), .ZN(n5637) );
  OR2_X1 U7268 ( .A1(n8196), .A2(n9998), .ZN(n5636) );
  NAND2_X1 U7269 ( .A1(n5637), .A2(n5636), .ZN(n8205) );
  AOI21_X2 U7270 ( .B1(n5638), .B2(n10020), .A(n8205), .ZN(n8790) );
  NOR4_X1 U7271 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5642) );
  NOR4_X1 U7272 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5641) );
  NOR4_X1 U7273 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5640) );
  NOR4_X1 U7274 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5639) );
  NAND4_X1 U7275 ( .A1(n5642), .A2(n5641), .A3(n5640), .A4(n5639), .ZN(n5665)
         );
  NOR2_X1 U7276 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5646) );
  NOR4_X1 U7277 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5645) );
  NOR4_X1 U7278 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5644) );
  NOR4_X1 U7279 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5643) );
  NAND4_X1 U7280 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(n5664)
         );
  NAND3_X1 U7281 ( .A1(n5660), .A2(n5656), .A3(n5668), .ZN(n5647) );
  INV_X1 U7282 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7283 ( .A1(n5651), .A2(n5652), .ZN(n5654) );
  NAND2_X1 U7284 ( .A1(n5654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5650) );
  INV_X1 U7285 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5649) );
  OR2_X1 U7286 ( .A1(n5651), .A2(n8890), .ZN(n5653) );
  MUX2_X1 U7287 ( .A(n5653), .B(P2_IR_REG_31__SCAN_IN), .S(n5652), .Z(n5655)
         );
  NAND2_X1 U7288 ( .A1(n5655), .A2(n5654), .ZN(n7999) );
  NAND2_X1 U7289 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U7290 ( .A1(n5658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7291 ( .A1(n5669), .A2(n5668), .ZN(n5659) );
  NAND2_X1 U7292 ( .A1(n5659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U7293 ( .A(n7997), .B(P2_B_REG_SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7294 ( .A1(n7999), .A2(n5662), .ZN(n5663) );
  OAI21_X1 U7295 ( .B1(n5665), .B2(n5664), .A(n10037), .ZN(n6958) );
  INV_X1 U7296 ( .A(n7997), .ZN(n5667) );
  NOR2_X1 U7297 ( .A1(n5674), .A2(n7999), .ZN(n5666) );
  XNOR2_X1 U7298 ( .A(n5669), .B(n5668), .ZN(n6964) );
  INV_X1 U7299 ( .A(n10044), .ZN(n5670) );
  NAND2_X1 U7300 ( .A1(n4376), .A2(n8575), .ZN(n6971) );
  AND2_X1 U7301 ( .A1(n6974), .A2(n6971), .ZN(n6966) );
  NOR2_X1 U7302 ( .A1(n10038), .A2(n6966), .ZN(n5671) );
  NAND2_X1 U7303 ( .A1(n6958), .A2(n5671), .ZN(n5771) );
  INV_X1 U7304 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U7305 ( .A1(n10037), .A2(n10289), .ZN(n5673) );
  AND2_X1 U7306 ( .A1(n5674), .A2(n7999), .ZN(n10043) );
  INV_X1 U7307 ( .A(n10043), .ZN(n5672) );
  NAND2_X1 U7308 ( .A1(n5673), .A2(n5672), .ZN(n6954) );
  NOR2_X1 U7309 ( .A1(n5771), .A2(n6954), .ZN(n5726) );
  INV_X1 U7310 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U7311 ( .A1(n10037), .A2(n10040), .ZN(n5676) );
  AND2_X1 U7312 ( .A1(n7997), .A2(n5674), .ZN(n10041) );
  INV_X1 U7313 ( .A(n10041), .ZN(n5675) );
  NAND2_X1 U7314 ( .A1(n5726), .A2(n6002), .ZN(n5680) );
  OR2_X4 U7315 ( .A1(n10045), .A2(n5978), .ZN(n10113) );
  INV_X1 U7316 ( .A(n6962), .ZN(n5679) );
  NAND2_X1 U7317 ( .A1(n5854), .A2(n5853), .ZN(n5976) );
  NAND2_X1 U7318 ( .A1(n5682), .A2(n5123), .ZN(n5683) );
  OR2_X1 U7319 ( .A1(n10016), .A2(n7534), .ZN(n5684) );
  OR2_X1 U7320 ( .A1(n8450), .A2(n5163), .ZN(n7320) );
  INV_X1 U7321 ( .A(n10070), .ZN(n8357) );
  OR2_X1 U7322 ( .A1(n10018), .A2(n8357), .ZN(n5685) );
  AND2_X1 U7323 ( .A1(n7320), .A2(n5685), .ZN(n5687) );
  INV_X1 U7324 ( .A(n5685), .ZN(n5686) );
  OAI21_X1 U7325 ( .B1(n8448), .B2(n8321), .A(n8447), .ZN(n5689) );
  NOR2_X1 U7326 ( .A1(n8448), .A2(n8447), .ZN(n5688) );
  AOI22_X1 U7327 ( .A1(n10074), .A2(n5689), .B1(n5688), .B2(n7556), .ZN(n5690)
         );
  NAND2_X1 U7328 ( .A1(n7616), .A2(n5871), .ZN(n5979) );
  INV_X1 U7329 ( .A(n8391), .ZN(n8446) );
  OR2_X1 U7330 ( .A1(n10081), .A2(n8446), .ZN(n5691) );
  INV_X1 U7331 ( .A(n7634), .ZN(n8445) );
  AND2_X1 U7332 ( .A1(n10088), .A2(n8445), .ZN(n7631) );
  NOR2_X1 U7333 ( .A1(n5693), .A2(n7631), .ZN(n5694) );
  NAND2_X1 U7334 ( .A1(n7637), .A2(n5694), .ZN(n5696) );
  INV_X1 U7335 ( .A(n9997), .ZN(n8444) );
  OR2_X1 U7336 ( .A1(n10095), .A2(n8444), .ZN(n5695) );
  NAND2_X1 U7337 ( .A1(n4441), .A2(n4399), .ZN(n5699) );
  INV_X1 U7338 ( .A(n7696), .ZN(n10105) );
  INV_X1 U7339 ( .A(n7631), .ZN(n5697) );
  NAND2_X1 U7340 ( .A1(n7637), .A2(n5697), .ZN(n9990) );
  NAND3_X1 U7341 ( .A1(n4441), .A2(n4399), .A3(n9990), .ZN(n5698) );
  NAND2_X1 U7342 ( .A1(n5887), .A2(n5881), .ZN(n7749) );
  INV_X1 U7343 ( .A(n9999), .ZN(n8442) );
  NAND2_X1 U7344 ( .A1(n7796), .A2(n8442), .ZN(n5700) );
  NAND2_X1 U7345 ( .A1(n5839), .A2(n7977), .ZN(n7927) );
  INV_X1 U7346 ( .A(n7969), .ZN(n8441) );
  OR2_X1 U7347 ( .A1(n7893), .A2(n8441), .ZN(n7925) );
  AND2_X1 U7348 ( .A1(n7927), .A2(n7925), .ZN(n5701) );
  INV_X1 U7349 ( .A(n8208), .ZN(n8440) );
  NAND2_X1 U7350 ( .A1(n8858), .A2(n8440), .ZN(n5702) );
  NAND2_X1 U7351 ( .A1(n8745), .A2(n5838), .ZN(n7983) );
  NAND2_X1 U7352 ( .A1(n7984), .A2(n7983), .ZN(n7982) );
  INV_X1 U7353 ( .A(n8048), .ZN(n8749) );
  OR2_X1 U7354 ( .A1(n8854), .A2(n8749), .ZN(n5703) );
  NAND2_X1 U7355 ( .A1(n7982), .A2(n5703), .ZN(n8752) );
  INV_X1 U7356 ( .A(n8731), .ZN(n8439) );
  NOR2_X1 U7357 ( .A1(n5704), .A2(n8439), .ZN(n5705) );
  INV_X1 U7358 ( .A(n8332), .ZN(n8750) );
  INV_X1 U7359 ( .A(n8732), .ZN(n8438) );
  INV_X1 U7360 ( .A(n8331), .ZN(n8708) );
  INV_X1 U7361 ( .A(n8828), .ZN(n8680) );
  NAND2_X1 U7362 ( .A1(n5926), .A2(n5923), .ZN(n8665) );
  NAND2_X1 U7363 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  INV_X1 U7364 ( .A(n8807), .ZN(n8620) );
  OR2_X1 U7365 ( .A1(n8801), .A2(n8613), .ZN(n5710) );
  NAND2_X1 U7366 ( .A1(n5711), .A2(n8592), .ZN(n5712) );
  NAND2_X1 U7367 ( .A1(n8565), .A2(n8196), .ZN(n5714) );
  OR2_X1 U7368 ( .A1(n5715), .A2(n5978), .ZN(n5995) );
  NAND2_X1 U7369 ( .A1(n5845), .A2(n4376), .ZN(n7167) );
  AOI21_X1 U7370 ( .B1(n5716), .B2(n7167), .A(n5619), .ZN(n5717) );
  NAND2_X1 U7371 ( .A1(n5995), .A2(n5717), .ZN(n8736) );
  OR2_X1 U7372 ( .A1(n7167), .A2(n8575), .ZN(n7614) );
  AND2_X1 U7373 ( .A1(n8736), .A2(n7614), .ZN(n5718) );
  NAND2_X1 U7374 ( .A1(n10023), .A2(n10032), .ZN(n7323) );
  NOR2_X2 U7375 ( .A1(n7375), .A2(n8321), .ZN(n7563) );
  INV_X1 U7376 ( .A(n10081), .ZN(n7305) );
  NAND2_X1 U7377 ( .A1(n7300), .A2(n7305), .ZN(n7301) );
  INV_X1 U7378 ( .A(n7796), .ZN(n10112) );
  INV_X1 U7379 ( .A(n8854), .ZN(n7989) );
  INV_X1 U7380 ( .A(n8842), .ZN(n8741) );
  INV_X1 U7381 ( .A(n5704), .ZN(n8757) );
  NAND2_X1 U7382 ( .A1(n8696), .A2(n8680), .ZN(n8660) );
  OR2_X2 U7383 ( .A1(n8628), .A2(n8807), .ZN(n8618) );
  NOR2_X2 U7384 ( .A1(n8799), .A2(n8601), .ZN(n8572) );
  AND2_X2 U7385 ( .A1(n8572), .A2(n8565), .ZN(n5722) );
  INV_X1 U7386 ( .A(n5722), .ZN(n5724) );
  INV_X1 U7387 ( .A(n8135), .ZN(n5723) );
  AOI211_X1 U7388 ( .C1(n8788), .C2(n5724), .A(n10113), .B(n5723), .ZN(n8787)
         );
  NOR2_X1 U7389 ( .A1(n6955), .A2(n5619), .ZN(n5725) );
  NAND2_X1 U7390 ( .A1(n5726), .A2(n5725), .ZN(n8551) );
  INV_X1 U7391 ( .A(n8551), .ZN(n8720) );
  OR2_X1 U7392 ( .A1(n10045), .A2(n4376), .ZN(n6959) );
  OR2_X2 U7393 ( .A1(n10036), .A2(n6959), .ZN(n10031) );
  INV_X1 U7394 ( .A(n8203), .ZN(n5727) );
  AOI22_X1 U7395 ( .A1(n5727), .A2(n10002), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8766), .ZN(n5728) );
  OAI21_X1 U7396 ( .B1(n8207), .B2(n10031), .A(n5728), .ZN(n5729) );
  AOI21_X1 U7397 ( .B1(n8787), .B2(n8720), .A(n5729), .ZN(n5730) );
  NOR2_X1 U7398 ( .A1(n5733), .A2(n5739), .ZN(n5734) );
  AND2_X1 U7399 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  NAND2_X1 U7400 ( .A1(n5737), .A2(n5736), .ZN(n5741) );
  INV_X1 U7401 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5744) );
  INV_X1 U7402 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8146) );
  MUX2_X1 U7403 ( .A(n5744), .B(n8146), .S(n4380), .Z(n5778) );
  XNOR2_X1 U7404 ( .A(n5778), .B(SI_28_), .ZN(n5775) );
  NAND2_X1 U7405 ( .A1(n8004), .A2(n5272), .ZN(n5746) );
  NAND2_X1 U7406 ( .A1(n5186), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5745) );
  AND2_X1 U7407 ( .A1(n4376), .A2(n5619), .ZN(n5747) );
  NAND2_X1 U7408 ( .A1(n5716), .A2(n5747), .ZN(n10102) );
  NAND2_X1 U7409 ( .A1(n8556), .A2(n10117), .ZN(n5769) );
  AND2_X1 U7410 ( .A1(n5944), .A2(n5748), .ZN(n5946) );
  NAND2_X1 U7411 ( .A1(n8788), .A2(n8410), .ZN(n5951) );
  NAND3_X1 U7412 ( .A1(n8582), .A2(n5946), .A3(n5951), .ZN(n5754) );
  INV_X1 U7413 ( .A(n8410), .ZN(n8434) );
  NAND2_X1 U7414 ( .A1(n5947), .A2(n8566), .ZN(n5749) );
  NAND3_X1 U7415 ( .A1(n5749), .A2(n8434), .A3(n5944), .ZN(n5750) );
  NAND2_X1 U7416 ( .A1(n5750), .A2(n8788), .ZN(n5752) );
  NAND3_X1 U7417 ( .A1(n5947), .A2(n8410), .A3(n8566), .ZN(n5751) );
  OAI211_X1 U7418 ( .C1(n5944), .C2(n8434), .A(n5752), .B(n5751), .ZN(n5753)
         );
  INV_X1 U7419 ( .A(n5757), .ZN(n5755) );
  AOI21_X1 U7420 ( .B1(n5755), .B2(n8541), .A(n9995), .ZN(n5766) );
  INV_X1 U7421 ( .A(n8541), .ZN(n5756) );
  INV_X1 U7422 ( .A(n8548), .ZN(n5764) );
  INV_X1 U7423 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7424 ( .A1(n5791), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7425 ( .A1(n5786), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5758) );
  OAI211_X1 U7426 ( .C1(n5761), .C2(n5760), .A(n5759), .B(n5758), .ZN(n5762)
         );
  AOI21_X1 U7427 ( .B1(n5764), .B2(n5763), .A(n5762), .ZN(n8265) );
  OAI22_X1 U7428 ( .A1(n8265), .A2(n10000), .B1(n8410), .B2(n9998), .ZN(n5765)
         );
  AOI21_X1 U7429 ( .B1(n5766), .B2(n5795), .A(n5765), .ZN(n8563) );
  XNOR2_X1 U7430 ( .A(n4943), .B(n8135), .ZN(n8560) );
  INV_X1 U7431 ( .A(n10045), .ZN(n5972) );
  AND2_X2 U7432 ( .A1(n5972), .A2(n6971), .ZN(n10096) );
  AOI22_X1 U7433 ( .A1(n8560), .A2(n10097), .B1(n10096), .B2(n8258), .ZN(n5767) );
  NAND2_X1 U7434 ( .A1(n6954), .A2(n6962), .ZN(n5770) );
  INV_X1 U7435 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5772) );
  OR2_X1 U7436 ( .A1(n10142), .A2(n5772), .ZN(n5773) );
  NAND2_X1 U7437 ( .A1(n5774), .A2(n5773), .ZN(P2_U3548) );
  INV_X1 U7438 ( .A(SI_28_), .ZN(n5777) );
  NAND2_X1 U7439 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  INV_X1 U7440 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5780) );
  INV_X1 U7441 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9833) );
  MUX2_X1 U7442 ( .A(n5780), .B(n9833), .S(n5598), .Z(n5797) );
  INV_X1 U7443 ( .A(SI_29_), .ZN(n10338) );
  INV_X1 U7444 ( .A(n5797), .ZN(n5781) );
  NAND2_X1 U7445 ( .A1(n5781), .A2(SI_29_), .ZN(n5804) );
  MUX2_X1 U7446 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4524), .Z(n5806) );
  XNOR2_X1 U7447 ( .A(n5806), .B(SI_30_), .ZN(n5782) );
  NAND2_X1 U7448 ( .A1(n9054), .A2(n5272), .ZN(n5785) );
  NAND2_X1 U7449 ( .A1(n5186), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5784) );
  INV_X1 U7450 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U7451 ( .A1(n5786), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7452 ( .A1(n5787), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5788) );
  OAI211_X1 U7453 ( .C1(n5790), .C2(n10330), .A(n5789), .B(n5788), .ZN(n8535)
         );
  INV_X1 U7454 ( .A(n8535), .ZN(n5817) );
  NOR2_X1 U7455 ( .A1(n8136), .A2(n5817), .ZN(n5824) );
  NAND2_X1 U7456 ( .A1(n5787), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7457 ( .A1(n5791), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7458 ( .A1(n5786), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5792) );
  AND3_X1 U7459 ( .A1(n5794), .A2(n5793), .A3(n5792), .ZN(n8141) );
  NAND2_X1 U7460 ( .A1(n8141), .A2(n5845), .ZN(n5802) );
  XNOR2_X1 U7461 ( .A(n5797), .B(SI_29_), .ZN(n5798) );
  NAND2_X1 U7462 ( .A1(n9063), .A2(n5272), .ZN(n5800) );
  NAND2_X1 U7463 ( .A1(n5186), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7464 ( .A1(n8777), .A2(n8265), .ZN(n5961) );
  OAI21_X1 U7465 ( .B1(n8773), .B2(n5802), .A(n5961), .ZN(n5801) );
  NAND2_X1 U7466 ( .A1(n5806), .A2(SI_30_), .ZN(n5803) );
  INV_X1 U7467 ( .A(n5806), .ZN(n5808) );
  INV_X1 U7468 ( .A(SI_30_), .ZN(n5807) );
  NAND2_X1 U7469 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  NAND2_X1 U7470 ( .A1(n5810), .A2(n5809), .ZN(n5814) );
  INV_X1 U7471 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9050) );
  INV_X1 U7472 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5811) );
  MUX2_X1 U7473 ( .A(n9050), .B(n5811), .S(n4524), .Z(n5812) );
  XNOR2_X1 U7474 ( .A(n5812), .B(SI_31_), .ZN(n5813) );
  NAND2_X1 U7475 ( .A1(n5582), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5815) );
  OR2_X1 U7476 ( .A1(n5818), .A2(n8141), .ZN(n5968) );
  NAND2_X1 U7477 ( .A1(n8136), .A2(n5817), .ZN(n5962) );
  NAND2_X1 U7478 ( .A1(n5818), .A2(n8141), .ZN(n5967) );
  XNOR2_X1 U7479 ( .A(n5820), .B(n8575), .ZN(n6001) );
  OR2_X4 U7480 ( .A1(n10113), .A2(n5619), .ZN(n8188) );
  NAND2_X1 U7481 ( .A1(n8188), .A2(n5821), .ZN(n5823) );
  OR2_X1 U7482 ( .A1(n6964), .A2(P2_U3152), .ZN(n7912) );
  NAND2_X1 U7483 ( .A1(n5823), .A2(n5822), .ZN(n6000) );
  OR3_X1 U7484 ( .A1(n7912), .A2(n5978), .A3(n7166), .ZN(n5971) );
  INV_X1 U7485 ( .A(n5824), .ZN(n5963) );
  NAND2_X1 U7486 ( .A1(n5967), .A2(n5963), .ZN(n5991) );
  NAND2_X1 U7487 ( .A1(n5845), .A2(n5619), .ZN(n5825) );
  MUX2_X1 U7488 ( .A(n5990), .B(n5991), .S(n5959), .Z(n5970) );
  INV_X1 U7489 ( .A(n8615), .ZN(n5975) );
  AND2_X1 U7490 ( .A1(n5828), .A2(n5939), .ZN(n5826) );
  NAND2_X1 U7491 ( .A1(n5975), .A2(n5826), .ZN(n5833) );
  NOR2_X1 U7492 ( .A1(n5828), .A2(n5939), .ZN(n5829) );
  NAND2_X1 U7493 ( .A1(n5827), .A2(n5829), .ZN(n5831) );
  NAND2_X1 U7494 ( .A1(n5833), .A2(n5832), .ZN(n5932) );
  AND2_X1 U7495 ( .A1(n5918), .A2(n5834), .ZN(n5835) );
  MUX2_X1 U7496 ( .A(n5836), .B(n5835), .S(n5939), .Z(n5913) );
  MUX2_X1 U7497 ( .A(n5837), .B(n8705), .S(n5959), .Z(n5912) );
  INV_X1 U7498 ( .A(n8711), .ZN(n8706) );
  MUX2_X1 U7499 ( .A(n5838), .B(n8745), .S(n5959), .Z(n5907) );
  INV_X1 U7500 ( .A(n7983), .ZN(n7976) );
  MUX2_X1 U7501 ( .A(n5839), .B(n7977), .S(n5959), .Z(n5905) );
  INV_X1 U7502 ( .A(n7927), .ZN(n7924) );
  AND2_X1 U7503 ( .A1(n5842), .A2(n7551), .ZN(n5840) );
  NAND2_X1 U7504 ( .A1(n5842), .A2(n5841), .ZN(n5844) );
  NAND2_X1 U7505 ( .A1(n5869), .A2(n7551), .ZN(n5843) );
  NAND2_X1 U7506 ( .A1(n8451), .A2(n10046), .ZN(n7541) );
  NAND3_X1 U7507 ( .A1(n5853), .A2(n7541), .A3(n5845), .ZN(n5847) );
  INV_X1 U7508 ( .A(n5857), .ZN(n5846) );
  AOI21_X1 U7509 ( .B1(n7531), .B2(n5847), .A(n5846), .ZN(n5849) );
  NAND2_X1 U7510 ( .A1(n5855), .A2(n5959), .ZN(n5848) );
  INV_X1 U7511 ( .A(n5850), .ZN(n5865) );
  NAND2_X1 U7512 ( .A1(n10074), .A2(n8447), .ZN(n5862) );
  NAND2_X1 U7513 ( .A1(n7541), .A2(n5853), .ZN(n5856) );
  NAND3_X1 U7514 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(n5858) );
  NAND3_X1 U7515 ( .A1(n5858), .A2(n5939), .A3(n5857), .ZN(n5859) );
  NAND3_X1 U7516 ( .A1(n5860), .A2(n5862), .A3(n5859), .ZN(n5868) );
  NAND2_X1 U7517 ( .A1(n8450), .A2(n10032), .ZN(n5861) );
  AND2_X1 U7518 ( .A1(n7378), .A2(n5861), .ZN(n5864) );
  OAI211_X1 U7519 ( .C1(n5865), .C2(n5864), .A(n5863), .B(n5862), .ZN(n5866)
         );
  NAND2_X1 U7520 ( .A1(n5866), .A2(n5939), .ZN(n5867) );
  NAND2_X1 U7521 ( .A1(n5868), .A2(n5867), .ZN(n5875) );
  NOR2_X1 U7522 ( .A1(n5869), .A2(n5959), .ZN(n5870) );
  NOR2_X1 U7523 ( .A1(n5979), .A2(n5870), .ZN(n5874) );
  MUX2_X1 U7524 ( .A(n7616), .B(n5871), .S(n5959), .Z(n5872) );
  NAND2_X1 U7525 ( .A1(n7619), .A2(n5872), .ZN(n5873) );
  AOI21_X1 U7526 ( .B1(n5875), .B2(n5874), .A(n5873), .ZN(n5879) );
  MUX2_X1 U7527 ( .A(n5876), .B(n7636), .S(n5939), .Z(n5877) );
  NAND2_X1 U7528 ( .A1(n5877), .A2(n9993), .ZN(n5878) );
  INV_X1 U7529 ( .A(n5884), .ZN(n5889) );
  AND2_X1 U7530 ( .A1(n5885), .A2(n5959), .ZN(n5886) );
  OAI211_X1 U7531 ( .C1(n5889), .C2(n5888), .A(n5887), .B(n5886), .ZN(n5890)
         );
  INV_X1 U7532 ( .A(n5890), .ZN(n5892) );
  INV_X1 U7533 ( .A(n7893), .ZN(n8864) );
  NAND2_X1 U7534 ( .A1(n9999), .A2(n5959), .ZN(n5896) );
  INV_X1 U7535 ( .A(n5896), .ZN(n5893) );
  AOI22_X1 U7536 ( .A1(n7796), .A2(n5893), .B1(n7969), .B2(n5959), .ZN(n5901)
         );
  OR2_X1 U7537 ( .A1(n9999), .A2(n5959), .ZN(n5895) );
  OAI22_X1 U7538 ( .A1(n7796), .A2(n5895), .B1(n7969), .B2(n5959), .ZN(n5894)
         );
  NAND2_X1 U7539 ( .A1(n8864), .A2(n5894), .ZN(n5900) );
  NOR2_X1 U7540 ( .A1(n5895), .A2(n7969), .ZN(n5898) );
  OAI21_X1 U7541 ( .B1(n8441), .B2(n5896), .A(n7796), .ZN(n5897) );
  OAI21_X1 U7542 ( .B1(n5898), .B2(n7796), .A(n5897), .ZN(n5899) );
  OAI211_X1 U7543 ( .C1(n8864), .C2(n5901), .A(n5900), .B(n5899), .ZN(n5902)
         );
  INV_X1 U7544 ( .A(n5902), .ZN(n5903) );
  MUX2_X1 U7545 ( .A(n5909), .B(n5908), .S(n5959), .Z(n5910) );
  NAND2_X1 U7546 ( .A1(n5919), .A2(n8681), .ZN(n5914) );
  NAND2_X1 U7547 ( .A1(n5914), .A2(n5922), .ZN(n5915) );
  NAND3_X1 U7548 ( .A1(n5915), .A2(n5926), .A3(n5920), .ZN(n5916) );
  NAND3_X1 U7549 ( .A1(n5916), .A2(n5923), .A3(n5928), .ZN(n5917) );
  NAND2_X1 U7550 ( .A1(n8650), .A2(n8668), .ZN(n5925) );
  NAND4_X1 U7551 ( .A1(n5929), .A2(n5939), .A3(n5917), .A4(n5925), .ZN(n5931)
         );
  NAND2_X1 U7552 ( .A1(n5921), .A2(n5920), .ZN(n5924) );
  NAND3_X1 U7553 ( .A1(n5924), .A2(n5923), .A3(n5922), .ZN(n5927) );
  INV_X1 U7554 ( .A(n5933), .ZN(n5935) );
  AND2_X1 U7555 ( .A1(n5933), .A2(n5827), .ZN(n5934) );
  OAI22_X1 U7556 ( .A1(n5936), .A2(n5935), .B1(n5934), .B2(n5959), .ZN(n5938)
         );
  NAND3_X1 U7557 ( .A1(n5938), .A2(n4433), .A3(n5043), .ZN(n5943) );
  INV_X1 U7558 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U7559 ( .A1(n5948), .A2(n5959), .ZN(n5949) );
  OR2_X1 U7560 ( .A1(n8788), .A2(n8410), .ZN(n5952) );
  INV_X1 U7561 ( .A(n8543), .ZN(n8537) );
  OAI21_X1 U7562 ( .B1(n5939), .B2(n8258), .A(n5954), .ZN(n5955) );
  OAI21_X1 U7563 ( .B1(n5939), .B2(n8537), .A(n5955), .ZN(n5956) );
  NAND2_X1 U7564 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  NAND2_X1 U7565 ( .A1(n5958), .A2(n4929), .ZN(n5966) );
  MUX2_X1 U7566 ( .A(n5961), .B(n5960), .S(n5959), .Z(n5965) );
  NAND2_X1 U7567 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  MUX2_X1 U7568 ( .A(n5968), .B(n5967), .S(n5939), .Z(n5969) );
  INV_X1 U7569 ( .A(n7166), .ZN(n5973) );
  NOR4_X1 U7570 ( .A1(n5973), .A2(n7912), .A3(n5972), .A4(n5978), .ZN(n5974)
         );
  INV_X1 U7571 ( .A(n7585), .ZN(n5977) );
  NOR2_X1 U7572 ( .A1(n5976), .A2(n5977), .ZN(n7588) );
  INV_X1 U7573 ( .A(n7530), .ZN(n7532) );
  INV_X1 U7574 ( .A(n5979), .ZN(n7295) );
  NAND4_X1 U7575 ( .A1(n5980), .A2(n7295), .A3(n7619), .A4(n7561), .ZN(n5981)
         );
  NOR4_X1 U7576 ( .A1(n7749), .A2(n4399), .A3(n7637), .A4(n5981), .ZN(n5982)
         );
  NAND4_X1 U7577 ( .A1(n7976), .A2(n7924), .A3(n7864), .A4(n5982), .ZN(n5983)
         );
  NOR4_X1 U7578 ( .A1(n8711), .A2(n8729), .A3(n8747), .A4(n5983), .ZN(n5984)
         );
  NAND3_X1 U7579 ( .A1(n8684), .A2(n8692), .A3(n5984), .ZN(n5985) );
  NOR4_X1 U7580 ( .A1(n8637), .A2(n5986), .A3(n8665), .A4(n5985), .ZN(n5987)
         );
  NAND3_X1 U7581 ( .A1(n5992), .A2(n5822), .A3(n7729), .ZN(n5993) );
  NOR4_X1 U7582 ( .A1(n5995), .A2(n5619), .A3(n6691), .A4(n8138), .ZN(n5998)
         );
  OAI21_X1 U7583 ( .B1(n7912), .B2(n5996), .A(P2_B_REG_SCAN_IN), .ZN(n5997) );
  AOI21_X1 U7584 ( .B1(n6717), .B2(n5998), .A(n5997), .ZN(n5999) );
  NAND2_X1 U7585 ( .A1(n6004), .A2(n10121), .ZN(n6007) );
  INV_X1 U7586 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7587 ( .A1(n6007), .A2(n6006), .ZN(P2_U3516) );
  NOR2_X1 U7588 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6012) );
  NAND3_X1 U7589 ( .A1(n6014), .A2(n6013), .A3(n6179), .ZN(n6015) );
  NOR2_X1 U7590 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6016) );
  INV_X1 U7591 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6018) );
  INV_X1 U7592 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6017) );
  NAND4_X1 U7593 ( .A1(n6365), .A2(n6433), .A3(n6018), .A4(n6017), .ZN(n6019)
         );
  INV_X1 U7594 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6021) );
  INV_X1 U7595 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6020) );
  XNOR2_X2 U7596 ( .A(n6023), .B(n6055), .ZN(n6646) );
  NAND2_X1 U7597 ( .A1(n6024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  INV_X1 U7598 ( .A(n6058), .ZN(n6063) );
  NAND2_X1 U7599 ( .A1(n6783), .A2(n5598), .ZN(n6139) );
  NAND2_X1 U7600 ( .A1(n7998), .A2(n6578), .ZN(n6028) );
  NAND2_X1 U7601 ( .A1(n9064), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6027) );
  NOR2_X1 U7602 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6030) );
  NOR2_X1 U7603 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6032) );
  INV_X1 U7604 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6034) );
  INV_X2 U7605 ( .A(n6889), .ZN(n6641) );
  NAND2_X1 U7606 ( .A1(n6042), .A2(n6041), .ZN(n6044) );
  OR2_X1 U7607 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND2_X1 U7608 ( .A1(n6044), .A2(n6043), .ZN(n8001) );
  NAND2_X1 U7609 ( .A1(n6614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  XNOR2_X1 U7610 ( .A(n6046), .B(n6045), .ZN(n7994) );
  NOR2_X1 U7611 ( .A1(n8001), .A2(n7994), .ZN(n6047) );
  INV_X1 U7612 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6370) );
  INV_X1 U7613 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8989) );
  INV_X1 U7614 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U7615 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6052) );
  INV_X1 U7616 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10432) );
  NAND2_X1 U7617 ( .A1(n6542), .A2(n10432), .ZN(n6054) );
  AND2_X1 U7618 ( .A1(n6567), .A2(n6054), .ZN(n9501) );
  INV_X1 U7619 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6056) );
  AND2_X1 U7620 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  INV_X1 U7621 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6059) );
  AND2_X2 U7622 ( .A1(n6067), .A2(n6066), .ZN(n6069) );
  AND2_X4 U7623 ( .A1(n6068), .A2(n6069), .ZN(n6510) );
  NAND2_X1 U7624 ( .A1(n9501), .A2(n6510), .ZN(n6075) );
  AND2_X4 U7625 ( .A1(n4386), .A2(n6069), .ZN(n9059) );
  INV_X1 U7626 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10310) );
  INV_X2 U7627 ( .A(n6069), .ZN(n9832) );
  NAND2_X1 U7628 ( .A1(n4391), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6072) );
  INV_X2 U7629 ( .A(n4383), .ZN(n9058) );
  NAND2_X1 U7630 ( .A1(n9058), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6071) );
  OAI211_X1 U7631 ( .C1(n6650), .C2(n10310), .A(n6072), .B(n6071), .ZN(n6073)
         );
  INV_X1 U7632 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7633 ( .A1(n6078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6080) );
  INV_X1 U7634 ( .A(n6891), .ZN(n7119) );
  NOR2_X1 U7635 ( .A1(n9518), .A2(n6163), .ZN(n6081) );
  AOI21_X1 U7636 ( .B1(n9715), .B2(n6465), .A(n6081), .ZN(n6560) );
  INV_X1 U7637 ( .A(n6560), .ZN(n6563) );
  NAND2_X1 U7638 ( .A1(n9715), .A2(n6637), .ZN(n6083) );
  NAND2_X1 U7639 ( .A1(n9488), .A2(n6622), .ZN(n6082) );
  NAND2_X1 U7640 ( .A1(n6083), .A2(n6082), .ZN(n6085) );
  XNOR2_X1 U7641 ( .A(n6085), .B(n7129), .ZN(n6562) );
  NAND2_X1 U7642 ( .A1(n9059), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7643 ( .A1(n6510), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6094) );
  INV_X1 U7644 ( .A(n6393), .ZN(n6191) );
  NAND2_X1 U7645 ( .A1(n4390), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6092) );
  INV_X1 U7646 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6087) );
  OR2_X1 U7647 ( .A1(n6139), .A2(n8046), .ZN(n6089) );
  OR2_X1 U7648 ( .A1(n9055), .A2(n10304), .ZN(n6088) );
  OAI211_X1 U7649 ( .C1(n6783), .C2(n8044), .A(n6089), .B(n6088), .ZN(n6096)
         );
  INV_X1 U7650 ( .A(n6096), .ZN(n7473) );
  OAI22_X1 U7651 ( .A1(n6132), .A2(n4388), .B1(n7473), .B2(n6090), .ZN(n6091)
         );
  XNOR2_X1 U7652 ( .A(n6091), .B(n7129), .ZN(n6128) );
  AOI22_X1 U7653 ( .A1(n6379), .A2(n9364), .B1(n6121), .B2(n7076), .ZN(n6129)
         );
  XNOR2_X1 U7654 ( .A(n6128), .B(n6129), .ZN(n7069) );
  NAND2_X1 U7655 ( .A1(n9059), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6104) );
  AND2_X1 U7656 ( .A1(n6068), .A2(n9832), .ZN(n6134) );
  NAND2_X1 U7657 ( .A1(n6134), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7658 ( .A1(n6510), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7659 ( .A1(n4389), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7660 ( .A1(n6379), .A2(n9365), .ZN(n6102) );
  OR2_X1 U7661 ( .A1(n6139), .A2(n6762), .ZN(n6100) );
  OR2_X1 U7662 ( .A1(n9055), .A2(n6761), .ZN(n6099) );
  NAND2_X1 U7663 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6098) );
  INV_X1 U7664 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6097) );
  AND3_X4 U7665 ( .A1(n6100), .A2(n6099), .A3(n5069), .ZN(n7457) );
  NAND2_X1 U7666 ( .A1(n6465), .A2(n7049), .ZN(n6101) );
  NAND2_X1 U7667 ( .A1(n6102), .A2(n6101), .ZN(n7046) );
  OAI22_X1 U7668 ( .A1(n6132), .A2(n7080), .B1(n7457), .B2(n6090), .ZN(n6107)
         );
  XNOR2_X1 U7669 ( .A(n6107), .B(n7129), .ZN(n7042) );
  NAND2_X1 U7670 ( .A1(n7046), .A2(n7042), .ZN(n6108) );
  NAND2_X1 U7671 ( .A1(n6134), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6111) );
  INV_X1 U7672 ( .A(n7052), .ZN(n7451) );
  INV_X1 U7673 ( .A(SI_0_), .ZN(n6114) );
  INV_X1 U7674 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7675 ( .B1(n4524), .B2(n6114), .A(n6113), .ZN(n6116) );
  AND2_X1 U7676 ( .A1(n6116), .A2(n6115), .ZN(n9842) );
  MUX2_X1 U7677 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9842), .S(n6783), .Z(n7122) );
  INV_X1 U7678 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6986) );
  NOR2_X1 U7679 ( .A1(n6728), .A2(n6986), .ZN(n6117) );
  AOI21_X1 U7680 ( .B1(n6121), .B2(n7122), .A(n6117), .ZN(n6118) );
  INV_X1 U7681 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6119) );
  NOR2_X1 U7682 ( .A1(n6728), .A2(n6119), .ZN(n6120) );
  AOI21_X1 U7683 ( .B1(n6637), .B2(n7122), .A(n6120), .ZN(n6123) );
  NAND2_X1 U7684 ( .A1(n6121), .A2(n7052), .ZN(n6122) );
  AND2_X1 U7685 ( .A1(n6123), .A2(n6122), .ZN(n6984) );
  OR2_X1 U7686 ( .A1(n6983), .A2(n6984), .ZN(n6981) );
  NAND2_X1 U7687 ( .A1(n6984), .A2(n7129), .ZN(n6124) );
  AND2_X1 U7688 ( .A1(n6981), .A2(n6124), .ZN(n7041) );
  NAND2_X1 U7689 ( .A1(n7041), .A2(n6125), .ZN(n6126) );
  INV_X1 U7690 ( .A(n6128), .ZN(n6130) );
  NAND2_X1 U7691 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  NAND2_X1 U7692 ( .A1(n9059), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6144) );
  INV_X1 U7693 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7694 ( .A1(n6510), .A2(n6133), .ZN(n6143) );
  NAND2_X1 U7695 ( .A1(n6134), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7696 ( .A1(n4389), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6141) );
  AND4_X1 U7697 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n7074)
         );
  NAND2_X1 U7698 ( .A1(n6135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6136) );
  XNOR2_X2 U7699 ( .A(n6136), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U7700 ( .A1(n6453), .A2(n6865), .ZN(n6138) );
  INV_X1 U7701 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6750) );
  OR2_X1 U7702 ( .A1(n9055), .A2(n6750), .ZN(n6137) );
  OAI211_X1 U7703 ( .C1(n6139), .C2(n6749), .A(n6138), .B(n6137), .ZN(n9933)
         );
  OAI22_X1 U7704 ( .A1(n6132), .A2(n7074), .B1(n6935), .B2(n6090), .ZN(n6140)
         );
  XNOR2_X1 U7705 ( .A(n6634), .B(n6140), .ZN(n6145) );
  NAND4_X1 U7706 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n9363)
         );
  INV_X1 U7707 ( .A(n6935), .ZN(n7679) );
  AOI22_X1 U7708 ( .A1(n6201), .A2(n9363), .B1(n6121), .B2(n7679), .ZN(n6146)
         );
  NAND2_X1 U7709 ( .A1(n6145), .A2(n6146), .ZN(n7015) );
  INV_X1 U7710 ( .A(n6145), .ZN(n6148) );
  INV_X1 U7711 ( .A(n6146), .ZN(n6147) );
  NAND2_X1 U7712 ( .A1(n6148), .A2(n6147), .ZN(n7014) );
  INV_X1 U7713 ( .A(n7085), .ZN(n6165) );
  NAND2_X1 U7714 ( .A1(n9059), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6153) );
  INV_X1 U7715 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6149) );
  XNOR2_X1 U7716 ( .A(n6149), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U7717 ( .A1(n6510), .A2(n7493), .ZN(n6152) );
  NAND2_X1 U7718 ( .A1(n6191), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7719 ( .A1(n4391), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6150) );
  NOR2_X1 U7720 ( .A1(n6154), .A2(n6061), .ZN(n6155) );
  MUX2_X1 U7721 ( .A(n6061), .B(n6155), .S(P1_IR_REG_4__SCAN_IN), .Z(n6156) );
  INV_X1 U7722 ( .A(n6156), .ZN(n6158) );
  INV_X1 U7723 ( .A(n6196), .ZN(n6157) );
  NAND2_X1 U7724 ( .A1(n6158), .A2(n6157), .ZN(n6830) );
  NAND2_X1 U7725 ( .A1(n6733), .A2(n4377), .ZN(n6161) );
  OAI211_X1 U7726 ( .C1(n6783), .C2(n6830), .A(n6161), .B(n6160), .ZN(n6946)
         );
  OAI22_X1 U7727 ( .A1(n6132), .A2(n7667), .B1(n7497), .B2(n6090), .ZN(n6162)
         );
  XNOR2_X1 U7728 ( .A(n6162), .B(n7129), .ZN(n6166) );
  OAI22_X1 U7729 ( .A1(n6163), .A2(n7667), .B1(n6132), .B2(n7497), .ZN(n6167)
         );
  XNOR2_X1 U7730 ( .A(n6166), .B(n6167), .ZN(n7084) );
  INV_X1 U7731 ( .A(n6166), .ZN(n6169) );
  INV_X1 U7732 ( .A(n6167), .ZN(n6168) );
  NAND2_X1 U7733 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7734 ( .A1(n9059), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6178) );
  INV_X1 U7735 ( .A(n6171), .ZN(n6190) );
  INV_X1 U7736 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7737 ( .A1(n6190), .A2(n6172), .ZN(n6173) );
  AND2_X1 U7738 ( .A1(n6216), .A2(n6173), .ZN(n7576) );
  NAND2_X1 U7739 ( .A1(n6510), .A2(n7576), .ZN(n6177) );
  NAND2_X1 U7740 ( .A1(n9058), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7741 ( .A1(n4391), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6175) );
  INV_X1 U7742 ( .A(n7356), .ZN(n9359) );
  NAND2_X1 U7743 ( .A1(n6201), .A2(n9359), .ZN(n6184) );
  NAND2_X1 U7744 ( .A1(n6740), .A2(n6578), .ZN(n6182) );
  NAND2_X1 U7745 ( .A1(n6196), .A2(n6179), .ZN(n6310) );
  NAND2_X1 U7746 ( .A1(n6310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U7747 ( .A(n6180), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7748 ( .A1(n9064), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6453), .B2(
        n6833), .ZN(n6181) );
  NAND2_X1 U7749 ( .A1(n6465), .A2(n9943), .ZN(n6183) );
  NAND2_X1 U7750 ( .A1(n9943), .A2(n6637), .ZN(n6185) );
  OAI21_X1 U7751 ( .B1(n6132), .B2(n7356), .A(n6185), .ZN(n6186) );
  XNOR2_X1 U7752 ( .A(n6634), .B(n6186), .ZN(n7573) );
  NAND2_X1 U7753 ( .A1(n9059), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6195) );
  INV_X1 U7754 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7755 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6187) );
  NAND2_X1 U7756 ( .A1(n6188), .A2(n6187), .ZN(n6189) );
  AND2_X1 U7757 ( .A1(n6190), .A2(n6189), .ZN(n7465) );
  NAND2_X1 U7758 ( .A1(n6510), .A2(n7465), .ZN(n6194) );
  NAND2_X1 U7759 ( .A1(n6191), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7760 ( .A1(n4390), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6192) );
  NAND4_X1 U7761 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n9360)
         );
  INV_X1 U7762 ( .A(n9360), .ZN(n7423) );
  NAND2_X1 U7763 ( .A1(n6737), .A2(n6578), .ZN(n6199) );
  OR2_X1 U7764 ( .A1(n6196), .A2(n6061), .ZN(n6197) );
  XNOR2_X1 U7765 ( .A(n6197), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6877) );
  AOI22_X1 U7766 ( .A1(n9064), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6453), .B2(
        n6877), .ZN(n6198) );
  OAI22_X1 U7767 ( .A1(n6132), .A2(n7423), .B1(n9966), .B2(n6090), .ZN(n6200)
         );
  XNOR2_X1 U7768 ( .A(n6634), .B(n6200), .ZN(n7461) );
  NAND2_X1 U7769 ( .A1(n6201), .A2(n9360), .ZN(n6203) );
  NAND2_X1 U7770 ( .A1(n6465), .A2(n7144), .ZN(n6202) );
  AND2_X1 U7771 ( .A1(n6203), .A2(n6202), .ZN(n7463) );
  AOI22_X1 U7772 ( .A1(n7572), .A2(n7573), .B1(n7461), .B2(n7463), .ZN(n6204)
         );
  INV_X1 U7773 ( .A(n7573), .ZN(n6210) );
  INV_X1 U7774 ( .A(n7461), .ZN(n7570) );
  INV_X1 U7775 ( .A(n7463), .ZN(n6205) );
  NAND2_X1 U7776 ( .A1(n7570), .A2(n6205), .ZN(n6206) );
  NAND2_X1 U7777 ( .A1(n6206), .A2(n7572), .ZN(n6209) );
  INV_X1 U7778 ( .A(n6206), .ZN(n6208) );
  INV_X1 U7779 ( .A(n7572), .ZN(n6207) );
  AOI22_X1 U7780 ( .A1(n6210), .A2(n6209), .B1(n6208), .B2(n6207), .ZN(n6211)
         );
  NAND2_X1 U7781 ( .A1(n6752), .A2(n6578), .ZN(n6214) );
  NAND2_X1 U7782 ( .A1(n6231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6212) );
  AOI22_X1 U7783 ( .A1(n9064), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6453), .B2(
        n6910), .ZN(n6213) );
  NAND2_X1 U7784 ( .A1(n6214), .A2(n6213), .ZN(n7404) );
  NAND2_X1 U7785 ( .A1(n7404), .A2(n6637), .ZN(n6223) );
  NAND2_X1 U7786 ( .A1(n9059), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6221) );
  INV_X1 U7787 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7788 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  AND2_X1 U7789 ( .A1(n6254), .A2(n6217), .ZN(n7355) );
  NAND2_X1 U7790 ( .A1(n6510), .A2(n7355), .ZN(n6220) );
  NAND2_X1 U7791 ( .A1(n9058), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7792 ( .A1(n4391), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7793 ( .A1(n7741), .A2(n6132), .ZN(n6222) );
  NAND2_X1 U7794 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  XNOR2_X1 U7795 ( .A(n6224), .B(n6634), .ZN(n6227) );
  NAND2_X1 U7796 ( .A1(n7404), .A2(n6622), .ZN(n6226) );
  INV_X1 U7797 ( .A(n7741), .ZN(n9358) );
  NAND2_X1 U7798 ( .A1(n6379), .A2(n9358), .ZN(n6225) );
  AND2_X1 U7799 ( .A1(n6226), .A2(n6225), .ZN(n6228) );
  NAND2_X1 U7800 ( .A1(n6227), .A2(n6228), .ZN(n7350) );
  INV_X1 U7801 ( .A(n6227), .ZN(n6230) );
  INV_X1 U7802 ( .A(n6228), .ZN(n6229) );
  NAND2_X1 U7803 ( .A1(n6230), .A2(n6229), .ZN(n7351) );
  NAND2_X1 U7804 ( .A1(n6759), .A2(n6578), .ZN(n6238) );
  INV_X1 U7805 ( .A(n6231), .ZN(n6233) );
  INV_X1 U7806 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7807 ( .A1(n6233), .A2(n6232), .ZN(n6250) );
  INV_X1 U7808 ( .A(n6250), .ZN(n6235) );
  INV_X1 U7809 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7810 ( .A1(n6235), .A2(n6234), .ZN(n6272) );
  NAND2_X1 U7811 ( .A1(n6272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6236) );
  XNOR2_X1 U7812 ( .A(n6236), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U7813 ( .A1(n9064), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7007), .B2(
        n6453), .ZN(n6237) );
  NAND2_X1 U7814 ( .A1(n9795), .A2(n6637), .ZN(n6245) );
  NAND2_X1 U7815 ( .A1(n9059), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7816 ( .A1(n6256), .A2(n7724), .ZN(n6239) );
  AND2_X1 U7817 ( .A1(n6281), .A2(n6239), .ZN(n7721) );
  NAND2_X1 U7818 ( .A1(n6510), .A2(n7721), .ZN(n6242) );
  NAND2_X1 U7819 ( .A1(n9058), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7820 ( .A1(n4390), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6240) );
  NAND4_X1 U7821 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(n9356)
         );
  NAND2_X1 U7822 ( .A1(n6465), .A2(n9356), .ZN(n6244) );
  NAND2_X1 U7823 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  XNOR2_X1 U7824 ( .A(n6246), .B(n6634), .ZN(n7719) );
  NAND2_X1 U7825 ( .A1(n9795), .A2(n6622), .ZN(n6248) );
  NAND2_X1 U7826 ( .A1(n6201), .A2(n9356), .ZN(n6247) );
  NAND2_X1 U7827 ( .A1(n6248), .A2(n6247), .ZN(n7718) );
  INV_X1 U7828 ( .A(n7718), .ZN(n6267) );
  NAND2_X1 U7829 ( .A1(n6250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6251) );
  MUX2_X1 U7830 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6251), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6252) );
  AOI22_X1 U7831 ( .A1(n9064), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9899), .B2(
        n6453), .ZN(n6253) );
  NAND2_X1 U7832 ( .A1(n7743), .A2(n6622), .ZN(n6262) );
  NAND2_X1 U7833 ( .A1(n9059), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6260) );
  INV_X1 U7834 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U7835 ( .A1(n6254), .A2(n10204), .ZN(n6255) );
  AND2_X1 U7836 ( .A1(n6256), .A2(n6255), .ZN(n7739) );
  NAND2_X1 U7837 ( .A1(n6510), .A2(n7739), .ZN(n6259) );
  NAND2_X1 U7838 ( .A1(n9058), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7839 ( .A1(n4390), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6257) );
  INV_X1 U7840 ( .A(n7517), .ZN(n9357) );
  NAND2_X1 U7841 ( .A1(n6201), .A2(n9357), .ZN(n6261) );
  NAND2_X1 U7842 ( .A1(n6262), .A2(n6261), .ZN(n7716) );
  INV_X1 U7843 ( .A(n7716), .ZN(n6266) );
  NAND2_X1 U7844 ( .A1(n7743), .A2(n6637), .ZN(n6264) );
  OR2_X1 U7845 ( .A1(n7517), .A2(n6132), .ZN(n6263) );
  NAND2_X1 U7846 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  XNOR2_X1 U7847 ( .A(n6265), .B(n7129), .ZN(n7715) );
  INV_X1 U7848 ( .A(n7715), .ZN(n7733) );
  OAI22_X1 U7849 ( .A1(n7719), .A2(n6267), .B1(n6266), .B2(n7733), .ZN(n6271)
         );
  OAI21_X1 U7850 ( .B1(n7715), .B2(n7716), .A(n7718), .ZN(n6269) );
  NOR2_X1 U7851 ( .A1(n7718), .A2(n7716), .ZN(n6268) );
  AOI22_X1 U7852 ( .A1(n7719), .A2(n6269), .B1(n6268), .B2(n7733), .ZN(n6270)
         );
  NAND2_X1 U7853 ( .A1(n6768), .A2(n6578), .ZN(n6280) );
  INV_X1 U7854 ( .A(n6272), .ZN(n6274) );
  INV_X1 U7855 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6273) );
  AOI21_X1 U7856 ( .B1(n6274), .B2(n6273), .A(n6061), .ZN(n6275) );
  NAND2_X1 U7857 ( .A1(n6275), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6278) );
  INV_X1 U7858 ( .A(n6275), .ZN(n6277) );
  INV_X1 U7859 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7860 ( .A1(n6277), .A2(n6276), .ZN(n6293) );
  AOI22_X1 U7861 ( .A1(n7097), .A2(n6453), .B1(n9064), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7862 ( .A1(n9790), .A2(n6637), .ZN(n6288) );
  NAND2_X1 U7863 ( .A1(n9059), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7864 ( .A1(n6281), .A2(n7003), .ZN(n6282) );
  AND2_X1 U7865 ( .A1(n6298), .A2(n6282), .ZN(n7658) );
  NAND2_X1 U7866 ( .A1(n6510), .A2(n7658), .ZN(n6285) );
  NAND2_X1 U7867 ( .A1(n9058), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7868 ( .A1(n4390), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6283) );
  OR2_X1 U7869 ( .A1(n7788), .A2(n6132), .ZN(n6287) );
  NAND2_X1 U7870 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  XNOR2_X1 U7871 ( .A(n6289), .B(n6634), .ZN(n7654) );
  NOR2_X1 U7872 ( .A1(n6163), .A2(n7788), .ZN(n6290) );
  AOI21_X1 U7873 ( .B1(n9790), .B2(n6465), .A(n6290), .ZN(n6291) );
  INV_X1 U7874 ( .A(n7654), .ZN(n6292) );
  INV_X1 U7875 ( .A(n6291), .ZN(n7653) );
  NAND2_X1 U7876 ( .A1(n6292), .A2(n7653), .ZN(n7785) );
  NAND2_X1 U7877 ( .A1(n6773), .A2(n6578), .ZN(n6296) );
  NAND2_X1 U7878 ( .A1(n6293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6294) );
  AOI22_X1 U7879 ( .A1(n7439), .A2(n6453), .B1(n9064), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7880 ( .A1(n7792), .A2(n6637), .ZN(n6305) );
  NAND2_X1 U7881 ( .A1(n9059), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6303) );
  INV_X1 U7882 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7883 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  AND2_X1 U7884 ( .A1(n6315), .A2(n6299), .ZN(n7787) );
  NAND2_X1 U7885 ( .A1(n6510), .A2(n7787), .ZN(n6302) );
  NAND2_X1 U7886 ( .A1(n4391), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7887 ( .A1(n9058), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6300) );
  NAND4_X1 U7888 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n9354)
         );
  NAND2_X1 U7889 ( .A1(n6465), .A2(n9354), .ZN(n6304) );
  NAND2_X1 U7890 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  XNOR2_X1 U7891 ( .A(n6306), .B(n7129), .ZN(n6329) );
  NOR2_X1 U7892 ( .A1(n6163), .A2(n7884), .ZN(n6307) );
  AOI21_X1 U7893 ( .B1(n7792), .B2(n6465), .A(n6307), .ZN(n6328) );
  INV_X1 U7894 ( .A(n6328), .ZN(n6308) );
  NAND2_X1 U7895 ( .A1(n6329), .A2(n6308), .ZN(n7877) );
  NAND2_X1 U7896 ( .A1(n6794), .A2(n6578), .ZN(n6313) );
  OR2_X1 U7897 ( .A1(n6310), .A2(n6309), .ZN(n6335) );
  NAND2_X1 U7898 ( .A1(n6335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6311) );
  XNOR2_X1 U7899 ( .A(n6311), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7689) );
  AOI22_X1 U7900 ( .A1(n9064), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6453), .B2(
        n7689), .ZN(n6312) );
  NAND2_X1 U7901 ( .A1(n9779), .A2(n6637), .ZN(n6322) );
  NAND2_X1 U7902 ( .A1(n9059), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6320) );
  INV_X1 U7903 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7904 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  AND2_X1 U7905 ( .A1(n6339), .A2(n6316), .ZN(n7881) );
  NAND2_X1 U7906 ( .A1(n6510), .A2(n7881), .ZN(n6319) );
  NAND2_X1 U7907 ( .A1(n9058), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7908 ( .A1(n4390), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6317) );
  OR2_X1 U7909 ( .A1(n7818), .A2(n6132), .ZN(n6321) );
  NAND2_X1 U7910 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  XNOR2_X1 U7911 ( .A(n6323), .B(n6634), .ZN(n6332) );
  INV_X1 U7912 ( .A(n6332), .ZN(n6326) );
  NOR2_X1 U7913 ( .A1(n6163), .A2(n7818), .ZN(n6324) );
  AOI21_X1 U7914 ( .B1(n9779), .B2(n6465), .A(n6324), .ZN(n6331) );
  INV_X1 U7915 ( .A(n6331), .ZN(n6325) );
  NAND2_X1 U7916 ( .A1(n6326), .A2(n6325), .ZN(n7874) );
  AND2_X1 U7917 ( .A1(n7785), .A2(n6327), .ZN(n6334) );
  INV_X1 U7918 ( .A(n6327), .ZN(n6330) );
  XNOR2_X1 U7919 ( .A(n6329), .B(n6328), .ZN(n7875) );
  OR2_X1 U7920 ( .A1(n6330), .A2(n7875), .ZN(n6333) );
  NAND2_X1 U7921 ( .A1(n6332), .A2(n6331), .ZN(n7873) );
  NAND2_X1 U7922 ( .A1(n6798), .A2(n4377), .ZN(n6338) );
  OAI21_X1 U7923 ( .B1(n6335), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6336) );
  XNOR2_X1 U7924 ( .A(n6336), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9375) );
  AOI22_X1 U7925 ( .A1(n9064), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6453), .B2(
        n9375), .ZN(n6337) );
  NAND2_X1 U7926 ( .A1(n7949), .A2(n6637), .ZN(n6346) );
  NAND2_X1 U7927 ( .A1(n9059), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7928 ( .A1(n6339), .A2(n10241), .ZN(n6340) );
  AND2_X1 U7929 ( .A1(n6389), .A2(n6340), .ZN(n7852) );
  NAND2_X1 U7930 ( .A1(n6510), .A2(n7852), .ZN(n6343) );
  NAND2_X1 U7931 ( .A1(n9058), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7932 ( .A1(n4391), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6341) );
  NAND4_X1 U7933 ( .A1(n6344), .A2(n6343), .A3(n6342), .A4(n6341), .ZN(n9352)
         );
  NAND2_X1 U7934 ( .A1(n6465), .A2(n9352), .ZN(n6345) );
  NAND2_X1 U7935 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U7936 ( .A(n6347), .B(n7129), .ZN(n7813) );
  NAND2_X1 U7937 ( .A1(n7949), .A2(n6622), .ZN(n6349) );
  NAND2_X1 U7938 ( .A1(n6201), .A2(n9352), .ZN(n6348) );
  NAND2_X1 U7939 ( .A1(n6349), .A2(n6348), .ZN(n7814) );
  NAND2_X1 U7940 ( .A1(n7039), .A2(n4377), .ZN(n6353) );
  OR2_X1 U7941 ( .A1(n6350), .A2(n6061), .ZN(n6351) );
  XNOR2_X1 U7942 ( .A(n6351), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9413) );
  AOI22_X1 U7943 ( .A1(n9064), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6453), .B2(
        n9413), .ZN(n6352) );
  NAND2_X1 U7944 ( .A1(n9764), .A2(n6637), .ZN(n6360) );
  INV_X1 U7945 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7946 ( .A1(n6372), .A2(n6354), .ZN(n6355) );
  NAND2_X1 U7947 ( .A1(n6417), .A2(n6355), .ZN(n9638) );
  OR2_X1 U7948 ( .A1(n9638), .A2(n6647), .ZN(n6358) );
  AOI22_X1 U7949 ( .A1(n9059), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9058), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7950 ( .A1(n4391), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6356) );
  INV_X1 U7951 ( .A(n8991), .ZN(n9661) );
  NAND2_X1 U7952 ( .A1(n9661), .A2(n6622), .ZN(n6359) );
  NAND2_X1 U7953 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  NAND2_X1 U7954 ( .A1(n9764), .A2(n6622), .ZN(n6363) );
  NAND2_X1 U7955 ( .A1(n9661), .A2(n6201), .ZN(n6362) );
  NAND2_X1 U7956 ( .A1(n6363), .A2(n6362), .ZN(n6404) );
  NAND2_X1 U7957 ( .A1(n7023), .A2(n4377), .ZN(n6369) );
  OR2_X1 U7958 ( .A1(n6364), .A2(n6061), .ZN(n6385) );
  NAND2_X1 U7959 ( .A1(n6385), .A2(n6365), .ZN(n6366) );
  NAND2_X1 U7960 ( .A1(n6366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6367) );
  XNOR2_X1 U7961 ( .A(n6367), .B(n10416), .ZN(n9392) );
  INV_X1 U7962 ( .A(n9392), .ZN(n9382) );
  AOI22_X1 U7963 ( .A1(n9064), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9382), .B2(
        n6453), .ZN(n6368) );
  NAND2_X1 U7964 ( .A1(n9672), .A2(n6637), .ZN(n6377) );
  NAND2_X1 U7965 ( .A1(n6391), .A2(n6370), .ZN(n6371) );
  AND2_X1 U7966 ( .A1(n6372), .A2(n6371), .ZN(n9670) );
  NAND2_X1 U7967 ( .A1(n9670), .A2(n6510), .ZN(n6375) );
  AOI22_X1 U7968 ( .A1(n9059), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9058), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7969 ( .A1(n4390), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7970 ( .A1(n9351), .A2(n6622), .ZN(n6376) );
  NAND2_X1 U7971 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  XNOR2_X1 U7972 ( .A(n6378), .B(n6634), .ZN(n8971) );
  NAND2_X1 U7973 ( .A1(n9672), .A2(n6622), .ZN(n6381) );
  NAND2_X1 U7974 ( .A1(n9351), .A2(n6201), .ZN(n6380) );
  NAND2_X1 U7975 ( .A1(n6381), .A2(n6380), .ZN(n9037) );
  OR2_X1 U7976 ( .A1(n6404), .A2(n9037), .ZN(n6382) );
  NAND2_X1 U7977 ( .A1(n6403), .A2(n6382), .ZN(n6384) );
  NAND2_X1 U7978 ( .A1(n6404), .A2(n9037), .ZN(n6383) );
  NAND2_X1 U7979 ( .A1(n6384), .A2(n6383), .ZN(n6402) );
  NAND2_X1 U7980 ( .A1(n6846), .A2(n6578), .ZN(n6387) );
  XNOR2_X1 U7981 ( .A(n6385), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U7982 ( .A1(n9064), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6453), .B2(
        n9909), .ZN(n6386) );
  NAND2_X1 U7983 ( .A1(n9774), .A2(n6637), .ZN(n6397) );
  INV_X1 U7984 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U7985 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U7986 ( .A1(n6391), .A2(n6390), .ZN(n7918) );
  INV_X1 U7987 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10374) );
  OAI22_X1 U7988 ( .A1(n7918), .A2(n6647), .B1(n6586), .B2(n10374), .ZN(n6395)
         );
  INV_X1 U7989 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9369) );
  INV_X1 U7990 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6392) );
  OAI22_X1 U7991 ( .A1(n6650), .A2(n9369), .B1(n4383), .B2(n6392), .ZN(n6394)
         );
  NAND2_X1 U7992 ( .A1(n6465), .A2(n9658), .ZN(n6396) );
  NAND2_X1 U7993 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  XNOR2_X1 U7994 ( .A(n6398), .B(n7129), .ZN(n7916) );
  NAND2_X1 U7995 ( .A1(n9774), .A2(n6622), .ZN(n6400) );
  NAND2_X1 U7996 ( .A1(n6201), .A2(n9658), .ZN(n6399) );
  NAND2_X1 U7997 ( .A1(n6400), .A2(n6399), .ZN(n8969) );
  INV_X1 U7998 ( .A(n6402), .ZN(n6412) );
  INV_X1 U7999 ( .A(n6403), .ZN(n6406) );
  INV_X1 U8000 ( .A(n6404), .ZN(n6405) );
  NAND2_X1 U8001 ( .A1(n6406), .A2(n6405), .ZN(n8981) );
  INV_X1 U8002 ( .A(n8971), .ZN(n6407) );
  INV_X1 U8003 ( .A(n7916), .ZN(n8973) );
  INV_X1 U8004 ( .A(n8969), .ZN(n7915) );
  NAND2_X1 U8005 ( .A1(n8973), .A2(n7915), .ZN(n6408) );
  NAND3_X1 U8006 ( .A1(n8981), .A2(n6407), .A3(n6408), .ZN(n6411) );
  INV_X1 U8007 ( .A(n6408), .ZN(n6409) );
  AND2_X1 U8008 ( .A1(n8971), .A2(n6409), .ZN(n6410) );
  AOI22_X1 U8009 ( .A1(n6412), .A2(n6411), .B1(n6410), .B2(n8975), .ZN(n6413)
         );
  NAND2_X1 U8010 ( .A1(n7108), .A2(n4377), .ZN(n6416) );
  NAND2_X1 U8011 ( .A1(n6414), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6434) );
  XNOR2_X1 U8012 ( .A(n6434), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9426) );
  AOI22_X1 U8013 ( .A1(n9064), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9426), .B2(
        n6453), .ZN(n6415) );
  NAND2_X1 U8014 ( .A1(n9759), .A2(n6637), .ZN(n6425) );
  NAND2_X1 U8015 ( .A1(n6417), .A2(n8989), .ZN(n6418) );
  AND2_X1 U8016 ( .A1(n6440), .A2(n6418), .ZN(n8990) );
  NAND2_X1 U8017 ( .A1(n8990), .A2(n6510), .ZN(n6423) );
  INV_X1 U8018 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U8019 ( .A1(n9058), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8020 ( .A1(n4391), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6419) );
  OAI211_X1 U8021 ( .C1(n6650), .C2(n10249), .A(n6420), .B(n6419), .ZN(n6421)
         );
  INV_X1 U8022 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8023 ( .A1(n6423), .A2(n6422), .ZN(n9607) );
  NAND2_X1 U8024 ( .A1(n9607), .A2(n6622), .ZN(n6424) );
  NAND2_X1 U8025 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  XNOR2_X1 U8026 ( .A(n6426), .B(n7129), .ZN(n6429) );
  AND2_X1 U8027 ( .A1(n9607), .A2(n6201), .ZN(n6427) );
  AOI21_X1 U8028 ( .B1(n9759), .B2(n6622), .A(n6427), .ZN(n6430) );
  XNOR2_X1 U8029 ( .A(n6429), .B(n6430), .ZN(n8982) );
  INV_X1 U8030 ( .A(n6429), .ZN(n6431) );
  NAND2_X1 U8031 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  NAND2_X1 U8032 ( .A1(n7332), .A2(n4377), .ZN(n6438) );
  NAND2_X1 U8033 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  NAND2_X1 U8034 ( .A1(n6435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6436) );
  XNOR2_X1 U8035 ( .A(n6436), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9437) );
  AOI22_X1 U8036 ( .A1(n9437), .A2(n6453), .B1(n9064), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8037 ( .A1(n9616), .A2(n6637), .ZN(n6448) );
  INV_X1 U8038 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8039 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U8040 ( .A1(n6457), .A2(n6441), .ZN(n9613) );
  OR2_X1 U8041 ( .A1(n9613), .A2(n6647), .ZN(n6446) );
  INV_X1 U8042 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10287) );
  INV_X1 U8043 ( .A(n4391), .ZN(n6586) );
  NAND2_X1 U8044 ( .A1(n9059), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8045 ( .A1(n9058), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6442) );
  OAI211_X1 U8046 ( .C1(n10287), .C2(n6586), .A(n6443), .B(n6442), .ZN(n6444)
         );
  INV_X1 U8047 ( .A(n6444), .ZN(n6445) );
  INV_X1 U8048 ( .A(n8933), .ZN(n9595) );
  NAND2_X1 U8049 ( .A1(n9595), .A2(n6622), .ZN(n6447) );
  NAND2_X1 U8050 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  XNOR2_X1 U8051 ( .A(n6449), .B(n6634), .ZN(n6452) );
  NAND2_X1 U8052 ( .A1(n9616), .A2(n6622), .ZN(n6451) );
  NAND2_X1 U8053 ( .A1(n9595), .A2(n6201), .ZN(n6450) );
  NAND2_X1 U8054 ( .A1(n6451), .A2(n6450), .ZN(n9021) );
  NAND2_X1 U8055 ( .A1(n7489), .A2(n4377), .ZN(n6455) );
  AOI22_X1 U8056 ( .A1(n6453), .A2(n9521), .B1(n9064), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6454) );
  INV_X1 U8057 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8058 ( .A1(n6457), .A2(n6456), .ZN(n6458) );
  NAND2_X1 U8059 ( .A1(n6471), .A2(n6458), .ZN(n9589) );
  OR2_X1 U8060 ( .A1(n9589), .A2(n6647), .ZN(n6463) );
  INV_X1 U8061 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U8062 ( .A1(n9058), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8063 ( .A1(n4390), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6459) );
  OAI211_X1 U8064 ( .C1(n6650), .C2(n9438), .A(n6460), .B(n6459), .ZN(n6461)
         );
  INV_X1 U8065 ( .A(n6461), .ZN(n6462) );
  NAND2_X1 U8066 ( .A1(n6463), .A2(n6462), .ZN(n9608) );
  AND2_X1 U8067 ( .A1(n9608), .A2(n6201), .ZN(n6464) );
  AOI21_X1 U8068 ( .B1(n9745), .B2(n6465), .A(n6464), .ZN(n8942) );
  NAND2_X1 U8069 ( .A1(n9745), .A2(n6637), .ZN(n6467) );
  NAND2_X1 U8070 ( .A1(n9608), .A2(n6622), .ZN(n6466) );
  NAND2_X1 U8071 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  XNOR2_X1 U8072 ( .A(n6468), .B(n6634), .ZN(n8940) );
  NAND2_X1 U8073 ( .A1(n7648), .A2(n4377), .ZN(n6470) );
  NAND2_X1 U8074 ( .A1(n9064), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U8075 ( .A1(n9740), .A2(n6637), .ZN(n6480) );
  NAND2_X1 U8076 ( .A1(n6471), .A2(n10321), .ZN(n6472) );
  NAND2_X1 U8077 ( .A1(n6508), .A2(n6472), .ZN(n9571) );
  OR2_X1 U8078 ( .A1(n9571), .A2(n6647), .ZN(n6478) );
  INV_X1 U8079 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U8080 ( .A1(n9058), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8081 ( .A1(n4391), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6473) );
  OAI211_X1 U8082 ( .C1(n6650), .C2(n6475), .A(n6474), .B(n6473), .ZN(n6476)
         );
  INV_X1 U8083 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U8084 ( .A1(n6478), .A2(n6477), .ZN(n9596) );
  NAND2_X1 U8085 ( .A1(n9596), .A2(n6622), .ZN(n6479) );
  NAND2_X1 U8086 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  XNOR2_X1 U8087 ( .A(n6481), .B(n7129), .ZN(n6484) );
  NAND2_X1 U8088 ( .A1(n9740), .A2(n6622), .ZN(n6483) );
  NAND2_X1 U8089 ( .A1(n9596), .A2(n6201), .ZN(n6482) );
  NAND2_X1 U8090 ( .A1(n6483), .A2(n6482), .ZN(n6485) );
  NAND2_X1 U8091 ( .A1(n6484), .A2(n6485), .ZN(n8944) );
  OAI21_X1 U8092 ( .B1(n8942), .B2(n8940), .A(n8944), .ZN(n6489) );
  INV_X1 U8093 ( .A(n6484), .ZN(n6487) );
  INV_X1 U8094 ( .A(n6485), .ZN(n6486) );
  NAND2_X1 U8095 ( .A1(n6487), .A2(n6486), .ZN(n8945) );
  NAND3_X1 U8096 ( .A1(n8944), .A2(n8942), .A3(n8940), .ZN(n6488) );
  OAI211_X1 U8097 ( .C1(n8931), .C2(n6489), .A(n8945), .B(n6488), .ZN(n6500)
         );
  NAND2_X1 U8098 ( .A1(n7728), .A2(n4377), .ZN(n6491) );
  NAND2_X1 U8099 ( .A1(n9064), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8100 ( .A1(n9736), .A2(n6637), .ZN(n6497) );
  XNOR2_X1 U8101 ( .A(n6508), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9558) );
  INV_X1 U8102 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8103 ( .A1(n4390), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8104 ( .A1(n9058), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6492) );
  OAI211_X1 U8105 ( .C1(n6650), .C2(n6494), .A(n6493), .B(n6492), .ZN(n6495)
         );
  OR2_X1 U8106 ( .A1(n9349), .A2(n6132), .ZN(n6496) );
  NAND2_X1 U8107 ( .A1(n6497), .A2(n6496), .ZN(n6498) );
  XNOR2_X1 U8108 ( .A(n6498), .B(n7129), .ZN(n6501) );
  NOR2_X1 U8109 ( .A1(n9349), .A2(n6163), .ZN(n6499) );
  AOI21_X1 U8110 ( .B1(n9736), .B2(n6622), .A(n6499), .ZN(n6502) );
  XNOR2_X1 U8111 ( .A(n6501), .B(n6502), .ZN(n8946) );
  INV_X1 U8112 ( .A(n6501), .ZN(n6503) );
  NAND2_X1 U8113 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  NAND2_X1 U8114 ( .A1(n7888), .A2(n4377), .ZN(n6506) );
  NAND2_X1 U8115 ( .A1(n9064), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6505) );
  INV_X1 U8116 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6507) );
  INV_X1 U8117 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9010) );
  OAI21_X1 U8118 ( .B1(n6508), .B2(n6507), .A(n9010), .ZN(n6509) );
  AND2_X1 U8119 ( .A1(n6526), .A2(n6509), .ZN(n9543) );
  NAND2_X1 U8120 ( .A1(n9543), .A2(n6510), .ZN(n6516) );
  INV_X1 U8121 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8122 ( .A1(n9058), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U8123 ( .A1(n4390), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6511) );
  OAI211_X1 U8124 ( .C1(n6650), .C2(n6513), .A(n6512), .B(n6511), .ZN(n6514)
         );
  INV_X1 U8125 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U8126 ( .A1(n6516), .A2(n6515), .ZN(n9564) );
  AND2_X1 U8127 ( .A1(n9564), .A2(n6201), .ZN(n6517) );
  AOI21_X1 U8128 ( .B1(n9731), .B2(n6622), .A(n6517), .ZN(n6522) );
  NAND2_X1 U8129 ( .A1(n9731), .A2(n6637), .ZN(n6520) );
  NAND2_X1 U8130 ( .A1(n9564), .A2(n6622), .ZN(n6519) );
  NAND2_X1 U8131 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  XNOR2_X1 U8132 ( .A(n6521), .B(n6634), .ZN(n9008) );
  INV_X1 U8133 ( .A(n8094), .ZN(n6559) );
  NAND2_X1 U8134 ( .A1(n6523), .A2(n6578), .ZN(n6525) );
  NAND2_X1 U8135 ( .A1(n9064), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6524) );
  INV_X1 U8136 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U8137 ( .A1(n6526), .A2(n10261), .ZN(n6527) );
  NAND2_X1 U8138 ( .A1(n6540), .A2(n6527), .ZN(n9529) );
  OR2_X1 U8139 ( .A1(n9529), .A2(n6647), .ZN(n6533) );
  INV_X1 U8140 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8141 ( .A1(n9058), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8142 ( .A1(n4391), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6528) );
  OAI211_X1 U8143 ( .C1(n6650), .C2(n6530), .A(n6529), .B(n6528), .ZN(n6531)
         );
  INV_X1 U8144 ( .A(n6531), .ZN(n6532) );
  OAI22_X1 U8145 ( .A1(n9532), .A2(n6090), .B1(n9517), .B2(n6132), .ZN(n6534)
         );
  XNOR2_X1 U8146 ( .A(n6534), .B(n6634), .ZN(n8095) );
  OR2_X1 U8147 ( .A1(n9532), .A2(n6132), .ZN(n6536) );
  NAND2_X1 U8148 ( .A1(n9549), .A2(n6379), .ZN(n6535) );
  NAND2_X1 U8149 ( .A1(n7992), .A2(n4377), .ZN(n6538) );
  NAND2_X1 U8150 ( .A1(n9064), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6537) );
  INV_X1 U8151 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8152 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NAND2_X1 U8153 ( .A1(n6542), .A2(n6541), .ZN(n9520) );
  OR2_X1 U8154 ( .A1(n9520), .A2(n6647), .ZN(n6548) );
  INV_X1 U8155 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8156 ( .A1(n9058), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8157 ( .A1(n4390), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6543) );
  OAI211_X1 U8158 ( .C1(n6650), .C2(n6545), .A(n6544), .B(n6543), .ZN(n6546)
         );
  INV_X1 U8159 ( .A(n6546), .ZN(n6547) );
  OAI22_X1 U8160 ( .A1(n8103), .A2(n6090), .B1(n8963), .B2(n6132), .ZN(n6549)
         );
  XNOR2_X1 U8161 ( .A(n6549), .B(n7129), .ZN(n6552) );
  OR2_X1 U8162 ( .A1(n8103), .A2(n6132), .ZN(n6551) );
  NAND2_X1 U8163 ( .A1(n8024), .A2(n6201), .ZN(n6550) );
  NAND2_X1 U8164 ( .A1(n6551), .A2(n6550), .ZN(n6553) );
  NAND2_X1 U8165 ( .A1(n6552), .A2(n6553), .ZN(n8096) );
  OAI21_X1 U8166 ( .B1(n8095), .B2(n8921), .A(n8096), .ZN(n6558) );
  NAND3_X1 U8167 ( .A1(n8096), .A2(n8095), .A3(n8921), .ZN(n6556) );
  INV_X1 U8168 ( .A(n6552), .ZN(n6555) );
  INV_X1 U8169 ( .A(n6553), .ZN(n6554) );
  NAND2_X1 U8170 ( .A1(n6555), .A2(n6554), .ZN(n8956) );
  OAI21_X1 U8171 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6561) );
  XNOR2_X1 U8172 ( .A(n6562), .B(n6560), .ZN(n8957) );
  NAND2_X1 U8173 ( .A1(n6561), .A2(n8957), .ZN(n8960) );
  NAND2_X1 U8174 ( .A1(n9064), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6564) );
  INV_X1 U8175 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U8176 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  NAND2_X1 U8177 ( .A1(n6582), .A2(n6568), .ZN(n9027) );
  INV_X1 U8178 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U8179 ( .A1(n9058), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8180 ( .A1(n4390), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6569) );
  OAI211_X1 U8181 ( .C1(n6650), .C2(n10318), .A(n6570), .B(n6569), .ZN(n6571)
         );
  INV_X1 U8182 ( .A(n6571), .ZN(n6572) );
  AND2_X1 U8183 ( .A1(n9506), .A2(n6201), .ZN(n6574) );
  AOI21_X1 U8184 ( .B1(n9710), .B2(n6622), .A(n6574), .ZN(n6593) );
  NAND2_X1 U8185 ( .A1(n9710), .A2(n6637), .ZN(n6576) );
  NAND2_X1 U8186 ( .A1(n9506), .A2(n6622), .ZN(n6575) );
  NAND2_X1 U8187 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  XNOR2_X1 U8188 ( .A(n6577), .B(n7129), .ZN(n6595) );
  XOR2_X1 U8189 ( .A(n6593), .B(n6595), .Z(n9032) );
  NAND2_X1 U8190 ( .A1(n8899), .A2(n6578), .ZN(n6580) );
  NAND2_X1 U8191 ( .A1(n9064), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6579) );
  INV_X1 U8192 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U8193 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND2_X1 U8194 ( .A1(n8914), .A2(n6510), .ZN(n6589) );
  INV_X1 U8195 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U8196 ( .A1(n9059), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U8197 ( .A1(n9058), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6584) );
  OAI211_X1 U8198 ( .C1(n6586), .C2(n10320), .A(n6585), .B(n6584), .ZN(n6587)
         );
  INV_X1 U8199 ( .A(n6587), .ZN(n6588) );
  OAI22_X1 U8200 ( .A1(n8919), .A2(n6090), .B1(n8026), .B2(n6132), .ZN(n6590)
         );
  XOR2_X1 U8201 ( .A(n7129), .B(n6590), .Z(n6592) );
  AOI22_X1 U8202 ( .A1(n9706), .A2(n6622), .B1(n6201), .B2(n9489), .ZN(n6591)
         );
  NAND2_X1 U8203 ( .A1(n6592), .A2(n6591), .ZN(n6665) );
  OAI21_X1 U8204 ( .B1(n6592), .B2(n6591), .A(n6665), .ZN(n8909) );
  INV_X1 U8205 ( .A(n6593), .ZN(n6594) );
  AND2_X1 U8206 ( .A1(n6595), .A2(n6594), .ZN(n8908) );
  INV_X1 U8207 ( .A(n8913), .ZN(n6619) );
  NAND2_X1 U8208 ( .A1(n8001), .A2(P1_B_REG_SCAN_IN), .ZN(n6596) );
  INV_X1 U8209 ( .A(n7994), .ZN(n6610) );
  MUX2_X1 U8210 ( .A(n6596), .B(P1_B_REG_SCAN_IN), .S(n6610), .Z(n6597) );
  NAND2_X1 U8211 ( .A1(n6597), .A2(n6611), .ZN(n9924) );
  INV_X1 U8212 ( .A(n6611), .ZN(n9841) );
  NAND2_X1 U8213 ( .A1(n9841), .A2(n8001), .ZN(n6598) );
  OAI21_X1 U8214 ( .B1(n9924), .B2(P1_D_REG_1__SCAN_IN), .A(n6598), .ZN(n6801)
         );
  INV_X1 U8215 ( .A(n6801), .ZN(n9825) );
  NOR4_X1 U8216 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6602) );
  NOR4_X1 U8217 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6601) );
  NOR4_X1 U8218 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6600) );
  NOR4_X1 U8219 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6599) );
  NAND4_X1 U8220 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n6609)
         );
  NOR2_X1 U8221 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .ZN(
        n6606) );
  NOR4_X1 U8222 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6605) );
  NOR4_X1 U8223 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6604) );
  NOR4_X1 U8224 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6603) );
  NAND4_X1 U8225 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6608)
         );
  INV_X1 U8226 ( .A(n9924), .ZN(n6607) );
  OAI21_X1 U8227 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(n6800) );
  AND2_X1 U8228 ( .A1(n9825), .A2(n6800), .ZN(n7112) );
  OAI22_X1 U8229 ( .A1(n9924), .A2(P1_D_REG_0__SCAN_IN), .B1(n6611), .B2(n6610), .ZN(n6919) );
  INV_X1 U8230 ( .A(n6919), .ZN(n9826) );
  NAND2_X1 U8231 ( .A1(n7112), .A2(n9826), .ZN(n7048) );
  NAND2_X1 U8232 ( .A1(n6612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6613) );
  MUX2_X1 U8233 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6613), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6615) );
  NAND2_X1 U8234 ( .A1(n6615), .A2(n6614), .ZN(n6729) );
  AND2_X1 U8235 ( .A1(n6729), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6616) );
  INV_X1 U8236 ( .A(n9925), .ZN(n6617) );
  NAND2_X1 U8237 ( .A1(n9328), .A2(n9210), .ZN(n7120) );
  INV_X1 U8238 ( .A(n7120), .ZN(n6804) );
  NAND2_X1 U8239 ( .A1(n6084), .A2(n6618), .ZN(n9166) );
  INV_X1 U8240 ( .A(n9166), .ZN(n6897) );
  NOR2_X2 U8241 ( .A1(n6645), .A2(n6655), .ZN(n8986) );
  NAND3_X1 U8242 ( .A1(n6619), .A2(n8986), .A3(n6665), .ZN(n6671) );
  NAND2_X1 U8243 ( .A1(n8004), .A2(n4377), .ZN(n6621) );
  NAND2_X1 U8244 ( .A1(n9064), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8245 ( .A1(n9700), .A2(n6622), .ZN(n6633) );
  INV_X1 U8246 ( .A(n6624), .ZN(n6623) );
  NAND2_X1 U8247 ( .A1(n6623), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9473) );
  INV_X1 U8248 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U8249 ( .A1(n6624), .A2(n10245), .ZN(n6625) );
  NAND2_X1 U8250 ( .A1(n9473), .A2(n6625), .ZN(n6654) );
  INV_X1 U8251 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U8252 ( .A1(n9058), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8253 ( .A1(n4391), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6626) );
  OAI211_X1 U8254 ( .C1(n6650), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6629)
         );
  INV_X1 U8255 ( .A(n6629), .ZN(n6630) );
  NAND2_X1 U8256 ( .A1(n9467), .A2(n6379), .ZN(n6632) );
  NAND2_X1 U8257 ( .A1(n6633), .A2(n6632), .ZN(n6635) );
  XNOR2_X1 U8258 ( .A(n6635), .B(n6634), .ZN(n6639) );
  NOR2_X1 U8259 ( .A1(n8148), .A2(n6132), .ZN(n6636) );
  AOI21_X1 U8260 ( .B1(n9700), .B2(n6637), .A(n6636), .ZN(n6638) );
  XNOR2_X1 U8261 ( .A(n6639), .B(n6638), .ZN(n6664) );
  INV_X1 U8262 ( .A(n6664), .ZN(n6670) );
  NAND2_X1 U8263 ( .A1(n6640), .A2(n6670), .ZN(n6669) );
  NAND2_X1 U8264 ( .A1(n6890), .A2(n6641), .ZN(n9331) );
  INV_X1 U8265 ( .A(n9331), .ZN(n6805) );
  NOR2_X1 U8266 ( .A1(n7120), .A2(n4378), .ZN(n7118) );
  OR2_X1 U8267 ( .A1(n6805), .A2(n7118), .ZN(n6642) );
  AND3_X1 U8268 ( .A1(n7048), .A2(n6642), .A3(n9925), .ZN(n6660) );
  INV_X1 U8269 ( .A(n6660), .ZN(n6644) );
  OR2_X1 U8270 ( .A1(n9166), .A2(n6891), .ZN(n6657) );
  NAND2_X1 U8271 ( .A1(n6657), .A2(n9925), .ZN(n7047) );
  INV_X1 U8272 ( .A(n7047), .ZN(n6643) );
  NAND2_X1 U8273 ( .A1(n6644), .A2(n6643), .ZN(n7361) );
  NOR2_X1 U8274 ( .A1(n6645), .A2(n9331), .ZN(n6653) );
  INV_X1 U8275 ( .A(n8145), .ZN(n9327) );
  NAND2_X1 U8276 ( .A1(n6653), .A2(n9327), .ZN(n9042) );
  INV_X1 U8277 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U8278 ( .A1(n9058), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8279 ( .A1(n4390), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6648) );
  OAI211_X1 U8280 ( .C1(n6650), .C2(n10273), .A(n6649), .B(n6648), .ZN(n6651)
         );
  INV_X1 U8281 ( .A(n6651), .ZN(n6652) );
  NAND2_X1 U8282 ( .A1(n9348), .A2(n9040), .ZN(n6663) );
  INV_X1 U8283 ( .A(n6654), .ZN(n8152) );
  INV_X1 U8284 ( .A(n6655), .ZN(n6656) );
  NAND2_X1 U8285 ( .A1(n6656), .A2(n7048), .ZN(n6659) );
  AND3_X1 U8286 ( .A1(n6657), .A2(n6729), .A3(n6728), .ZN(n6658) );
  AOI21_X1 U8287 ( .B1(n6659), .B2(n6658), .A(P1_U3084), .ZN(n6661) );
  AOI22_X1 U8288 ( .A1(n8152), .A2(n9039), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6662) );
  OAI211_X1 U8289 ( .C1(n8026), .C2(n9042), .A(n6663), .B(n6662), .ZN(n6667)
         );
  NOR3_X1 U8290 ( .A1(n6665), .A2(n6664), .A3(n9047), .ZN(n6666) );
  AOI211_X1 U8291 ( .C1(n9045), .C2(n9700), .A(n6667), .B(n6666), .ZN(n6668)
         );
  OAI211_X1 U8292 ( .C1(n6671), .C2(n6670), .A(n6669), .B(n6668), .ZN(P1_U3218) );
  INV_X1 U8293 ( .A(n6729), .ZN(n7890) );
  NOR2_X1 U8294 ( .A1(n6728), .A2(n7890), .ZN(n6778) );
  NAND2_X2 U8295 ( .A1(n6968), .A2(n10044), .ZN(n8449) );
  NAND2_X1 U8296 ( .A1(n8509), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U8297 ( .B1(n8509), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6672), .ZN(
        n8513) );
  INV_X1 U8298 ( .A(n7767), .ZN(n7024) );
  INV_X1 U8299 ( .A(n6710), .ZN(n7365) );
  INV_X1 U8300 ( .A(n6708), .ZN(n7345) );
  INV_X1 U8301 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6681) );
  INV_X1 U8302 ( .A(n7287), .ZN(n6775) );
  INV_X1 U8303 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6680) );
  INV_X1 U8304 ( .A(n8495), .ZN(n6770) );
  INV_X1 U8305 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6679) );
  INV_X1 U8306 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6678) );
  INV_X1 U8307 ( .A(n8482), .ZN(n6763) );
  INV_X1 U8308 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6677) );
  INV_X1 U8309 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7299) );
  INV_X1 U8310 ( .A(n6702), .ZN(n7066) );
  INV_X1 U8311 ( .A(n7221), .ZN(n6741) );
  INV_X1 U8312 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7564) );
  INV_X1 U8313 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6676) );
  INV_X1 U8314 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6675) );
  INV_X1 U8315 ( .A(n7276), .ZN(n6734) );
  INV_X1 U8316 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6674) );
  INV_X1 U8317 ( .A(n7234), .ZN(n6732) );
  INV_X1 U8318 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6673) );
  INV_X1 U8319 ( .A(n7248), .ZN(n8047) );
  MUX2_X1 U8320 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6673), .S(n7248), .Z(n7251)
         );
  INV_X1 U8321 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7595) );
  XNOR2_X1 U8322 ( .A(n6736), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n8455) );
  AND2_X1 U8323 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8454) );
  NAND2_X1 U8324 ( .A1(n8455), .A2(n8454), .ZN(n8453) );
  OAI21_X1 U8325 ( .B1(n6736), .B2(n7595), .A(n8453), .ZN(n7250) );
  NAND2_X1 U8326 ( .A1(n7251), .A2(n7250), .ZN(n7249) );
  MUX2_X1 U8327 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6674), .S(n7234), .Z(n7237)
         );
  XOR2_X1 U8328 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7276), .Z(n7279) );
  OAI21_X1 U8329 ( .B1(n6675), .B2(n6734), .A(n7277), .ZN(n7264) );
  XNOR2_X1 U8330 ( .A(n6738), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7265) );
  XOR2_X1 U8331 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7221), .Z(n7224) );
  MUX2_X1 U8332 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7299), .S(n6702), .Z(n7063)
         );
  MUX2_X1 U8333 ( .A(n6677), .B(P2_REG2_REG_8__SCAN_IN), .S(n6754), .Z(n8471)
         );
  OAI21_X1 U8334 ( .B1(n6677), .B2(n6754), .A(n8469), .ZN(n8477) );
  XOR2_X1 U8335 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8482), .Z(n8476) );
  NAND2_X1 U8336 ( .A1(n8477), .A2(n8476), .ZN(n8475) );
  OAI21_X1 U8337 ( .B1(n6678), .B2(n6763), .A(n8475), .ZN(n8491) );
  XOR2_X1 U8338 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8495), .Z(n8490) );
  XNOR2_X1 U8339 ( .A(n7287), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n7283) );
  XOR2_X1 U8340 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6708), .Z(n7343) );
  NAND2_X1 U8341 ( .A1(n7344), .A2(n7343), .ZN(n7342) );
  XNOR2_X1 U8342 ( .A(n6710), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n7364) );
  XNOR2_X1 U8343 ( .A(n7483), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U8344 ( .A1(n7024), .A2(n6682), .ZN(n6683) );
  XNOR2_X1 U8345 ( .A(n6682), .B(n7767), .ZN(n7759) );
  INV_X1 U8346 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U8347 ( .A1(n7759), .A2(n7758), .ZN(n7757) );
  NAND2_X1 U8348 ( .A1(n6683), .A2(n7757), .ZN(n8512) );
  NAND2_X1 U8349 ( .A1(n8109), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6684) );
  OAI21_X1 U8350 ( .B1(n8109), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6684), .ZN(
        n6689) );
  NOR2_X1 U8351 ( .A1(n6691), .A2(P2_U3152), .ZN(n8005) );
  AOI21_X1 U8352 ( .B1(n6968), .B2(n8005), .A(n5822), .ZN(n6685) );
  OAI21_X1 U8353 ( .B1(n10038), .B2(n6974), .A(n6685), .ZN(n6687) );
  NAND2_X1 U8354 ( .A1(n6687), .A2(n6686), .ZN(n6714) );
  NAND2_X1 U8355 ( .A1(n6714), .A2(n8449), .ZN(n6692) );
  NOR2_X1 U8356 ( .A1(n6691), .A2(n8138), .ZN(n6688) );
  INV_X1 U8357 ( .A(n9979), .ZN(n9982) );
  AOI211_X1 U8358 ( .C1(n6690), .C2(n6689), .A(n8104), .B(n9982), .ZN(n6727)
         );
  NAND2_X1 U8359 ( .A1(n6692), .A2(n6691), .ZN(n9983) );
  INV_X1 U8360 ( .A(n8109), .ZN(n6693) );
  NOR2_X1 U8361 ( .A1(n9983), .A2(n6693), .ZN(n6726) );
  XOR2_X1 U8362 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8509), .Z(n8503) );
  INV_X1 U8363 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10126) );
  MUX2_X1 U8364 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10126), .S(n7248), .Z(n7244)
         );
  XNOR2_X1 U8365 ( .A(n6736), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n8458) );
  AND2_X1 U8366 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8457) );
  NAND2_X1 U8367 ( .A1(n8458), .A2(n8457), .ZN(n8456) );
  NAND2_X1 U8368 ( .A1(n8452), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U8369 ( .A1(n8456), .A2(n6694), .ZN(n7243) );
  NAND2_X1 U8370 ( .A1(n7244), .A2(n7243), .ZN(n7242) );
  NAND2_X1 U8371 ( .A1(n7248), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8372 ( .A1(n7242), .A2(n6695), .ZN(n7229) );
  INV_X1 U8373 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U8374 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10128), .S(n7234), .Z(n7230)
         );
  NAND2_X1 U8375 ( .A1(n7234), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U8376 ( .A1(n7228), .A2(n6696), .ZN(n7271) );
  INV_X1 U8377 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6697) );
  XNOR2_X1 U8378 ( .A(n7276), .B(n6697), .ZN(n7272) );
  NAND2_X1 U8379 ( .A1(n7271), .A2(n7272), .ZN(n7270) );
  NAND2_X1 U8380 ( .A1(n7276), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8381 ( .A1(n7270), .A2(n6698), .ZN(n7257) );
  XNOR2_X1 U8382 ( .A(n6738), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7258) );
  NAND2_X1 U8383 ( .A1(n7262), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8384 ( .A1(n7256), .A2(n6699), .ZN(n7216) );
  INV_X1 U8385 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6700) );
  XNOR2_X1 U8386 ( .A(n7221), .B(n6700), .ZN(n7217) );
  NAND2_X1 U8387 ( .A1(n7216), .A2(n7217), .ZN(n7215) );
  NAND2_X1 U8388 ( .A1(n7221), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U8389 ( .A1(n7215), .A2(n6701), .ZN(n7056) );
  INV_X1 U8390 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10132) );
  MUX2_X1 U8391 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10132), .S(n6702), .Z(n7057)
         );
  NAND2_X1 U8392 ( .A1(n6702), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8393 ( .A1(n7055), .A2(n6703), .ZN(n8467) );
  INV_X1 U8394 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10134) );
  MUX2_X1 U8395 ( .A(n10134), .B(P2_REG1_REG_8__SCAN_IN), .S(n6754), .Z(n8468)
         );
  NAND2_X1 U8396 ( .A1(n8467), .A2(n8468), .ZN(n8466) );
  NAND2_X1 U8397 ( .A1(n8465), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8398 ( .A1(n8466), .A2(n6704), .ZN(n8484) );
  INV_X1 U8399 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10136) );
  MUX2_X1 U8400 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10136), .S(n8482), .Z(n8485)
         );
  NAND2_X1 U8401 ( .A1(n8482), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8402 ( .A1(n8483), .A2(n6705), .ZN(n8498) );
  INV_X1 U8403 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10335) );
  MUX2_X1 U8404 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10335), .S(n8495), .Z(n8497) );
  NAND2_X1 U8405 ( .A1(n8498), .A2(n8497), .ZN(n8496) );
  NAND2_X1 U8406 ( .A1(n8495), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U8407 ( .A1(n8496), .A2(n6706), .ZN(n7290) );
  INV_X1 U8408 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10140) );
  MUX2_X1 U8409 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10140), .S(n7287), .Z(n7289) );
  NAND2_X1 U8410 ( .A1(n7287), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U8411 ( .A1(n7288), .A2(n6707), .ZN(n7340) );
  XNOR2_X1 U8412 ( .A(n6708), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7341) );
  OR2_X1 U8413 ( .A1(n6708), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6709) );
  INV_X1 U8414 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10262) );
  XNOR2_X1 U8415 ( .A(n6710), .B(n10262), .ZN(n7369) );
  NAND2_X1 U8416 ( .A1(n7368), .A2(n7369), .ZN(n7367) );
  OR2_X1 U8417 ( .A1(n6710), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U8418 ( .A1(n7367), .A2(n6711), .ZN(n7479) );
  INV_X1 U8419 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10366) );
  XNOR2_X1 U8420 ( .A(n7483), .B(n10366), .ZN(n7480) );
  NOR2_X1 U8421 ( .A1(n7483), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6712) );
  AOI21_X1 U8422 ( .B1(n7479), .B2(n7480), .A(n6712), .ZN(n6713) );
  INV_X1 U8423 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10352) );
  NOR2_X1 U8424 ( .A1(n7764), .A2(n10352), .ZN(n7763) );
  AOI21_X1 U8425 ( .B1(n6713), .B2(n7767), .A(n7763), .ZN(n8504) );
  NAND2_X1 U8426 ( .A1(n8503), .A2(n8504), .ZN(n8502) );
  XNOR2_X1 U8427 ( .A(n8109), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U8428 ( .A1(n6715), .A2(n6716), .ZN(n8108) );
  INV_X1 U8429 ( .A(n8138), .ZN(n8900) );
  AOI211_X1 U8430 ( .C1(n6716), .C2(n6715), .A(n8108), .B(n9984), .ZN(n6725)
         );
  NAND2_X1 U8431 ( .A1(n6717), .A2(n6974), .ZN(n6721) );
  NAND2_X1 U8432 ( .A1(n10038), .A2(n7912), .ZN(n6719) );
  NAND2_X1 U8433 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  INV_X1 U8434 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U8435 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n6722) );
  OAI21_X1 U8436 ( .B1(n8522), .B2(n6723), .A(n6722), .ZN(n6724) );
  OR4_X1 U8437 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(P2_U3262)
         );
  NAND2_X1 U8438 ( .A1(n9166), .A2(n6728), .ZN(n6730) );
  NAND2_X1 U8439 ( .A1(n6730), .A2(n6729), .ZN(n6785) );
  NAND2_X1 U8440 ( .A1(n6785), .A2(n6783), .ZN(n6731) );
  NAND2_X1 U8441 ( .A1(n6731), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U8442 ( .A1(n4524), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8903) );
  INV_X1 U8443 ( .A(n8903), .ZN(n8093) );
  AND2_X1 U8444 ( .A1(n4524), .A2(P2_U3152), .ZN(n7911) );
  INV_X2 U8445 ( .A(n7911), .ZN(n8906) );
  OAI222_X1 U8446 ( .A1(n8093), .A2(n5156), .B1(n8906), .B2(n6749), .C1(
        P2_U3152), .C2(n6732), .ZN(P2_U3355) );
  INV_X1 U8447 ( .A(n6733), .ZN(n6747) );
  OAI222_X1 U8448 ( .A1(n8093), .A2(n4583), .B1(n8906), .B2(n6747), .C1(
        P2_U3152), .C2(n6734), .ZN(P2_U3354) );
  OAI222_X1 U8449 ( .A1(n6736), .A2(P2_U3152), .B1(n8906), .B2(n6762), .C1(
        n6735), .C2(n8093), .ZN(P2_U3357) );
  INV_X1 U8450 ( .A(n6737), .ZN(n6743) );
  OAI222_X1 U8451 ( .A1(n8093), .A2(n6739), .B1(n8906), .B2(n6743), .C1(
        P2_U3152), .C2(n6738), .ZN(P2_U3353) );
  INV_X1 U8452 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6742) );
  INV_X1 U8453 ( .A(n6740), .ZN(n6745) );
  OAI222_X1 U8454 ( .A1(n8093), .A2(n6742), .B1(n8906), .B2(n6745), .C1(
        P2_U3152), .C2(n6741), .ZN(P2_U3352) );
  NAND2_X1 U8455 ( .A1(n4524), .A2(P1_U3084), .ZN(n9837) );
  INV_X1 U8456 ( .A(n6877), .ZN(n6816) );
  OAI222_X1 U8457 ( .A1(n9837), .A2(n6744), .B1(n9840), .B2(n6743), .C1(
        P1_U3084), .C2(n6816), .ZN(P1_U3348) );
  INV_X1 U8458 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6746) );
  INV_X1 U8459 ( .A(n6833), .ZN(n6860) );
  OAI222_X1 U8460 ( .A1(n9837), .A2(n6746), .B1(n9840), .B2(n6745), .C1(
        P1_U3084), .C2(n6860), .ZN(P1_U3347) );
  OAI222_X1 U8461 ( .A1(n9837), .A2(n4970), .B1(n9840), .B2(n6747), .C1(
        P1_U3084), .C2(n6830), .ZN(P1_U3349) );
  INV_X1 U8462 ( .A(n6865), .ZN(n6748) );
  OAI222_X1 U8463 ( .A1(n9837), .A2(n6750), .B1(n9840), .B2(n6749), .C1(
        P1_U3084), .C2(n6748), .ZN(P1_U3350) );
  INV_X1 U8464 ( .A(n6249), .ZN(n6755) );
  INV_X1 U8465 ( .A(n9837), .ZN(n9828) );
  AOI22_X1 U8466 ( .A1(n9899), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9828), .ZN(n6751) );
  OAI21_X1 U8467 ( .B1(n6755), .B2(n9840), .A(n6751), .ZN(P1_U3345) );
  INV_X1 U8468 ( .A(n6752), .ZN(n6757) );
  AOI22_X1 U8469 ( .A1(n6910), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9828), .ZN(n6753) );
  OAI21_X1 U8470 ( .B1(n6757), .B2(n9840), .A(n6753), .ZN(P1_U3346) );
  OAI222_X1 U8471 ( .A1(n8093), .A2(n6756), .B1(n8906), .B2(n6755), .C1(
        P2_U3152), .C2(n6754), .ZN(P2_U3350) );
  INV_X1 U8472 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6758) );
  OAI222_X1 U8473 ( .A1(n8093), .A2(n6758), .B1(n8906), .B2(n6757), .C1(
        P2_U3152), .C2(n7066), .ZN(P2_U3351) );
  INV_X1 U8474 ( .A(n6759), .ZN(n6764) );
  AOI22_X1 U8475 ( .A1(n7007), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9828), .ZN(n6760) );
  OAI21_X1 U8476 ( .B1(n6764), .B2(n9840), .A(n6760), .ZN(P1_U3344) );
  OAI222_X1 U8477 ( .A1(n6823), .A2(P1_U3084), .B1(n9840), .B2(n6762), .C1(
        n6761), .C2(n9837), .ZN(P1_U3352) );
  OAI222_X1 U8478 ( .A1(n8093), .A2(n6765), .B1(n8906), .B2(n6764), .C1(n6763), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8479 ( .A(n8141), .ZN(n6766) );
  NAND2_X1 U8480 ( .A1(n6766), .A2(P2_U3966), .ZN(n6767) );
  OAI21_X1 U8481 ( .B1(n9050), .B2(P2_U3966), .A(n6767), .ZN(P2_U3583) );
  INV_X1 U8482 ( .A(n8522), .ZN(n9981) );
  NOR2_X1 U8483 ( .A1(n9981), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8484 ( .A(n6768), .ZN(n6771) );
  INV_X1 U8485 ( .A(n7097), .ZN(n7093) );
  OAI222_X1 U8486 ( .A1(n9837), .A2(n6769), .B1(n9840), .B2(n6771), .C1(n7093), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  OAI222_X1 U8487 ( .A1(n8093), .A2(n6772), .B1(n8906), .B2(n6771), .C1(n6770), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8488 ( .A(n6773), .ZN(n6776) );
  AOI22_X1 U8489 ( .A1(n7439), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9828), .ZN(n6774) );
  OAI21_X1 U8490 ( .B1(n6776), .B2(n9840), .A(n6774), .ZN(P1_U3342) );
  OAI222_X1 U8491 ( .A1(n8093), .A2(n6777), .B1(n8906), .B2(n6776), .C1(n6775), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8492 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6788) );
  AOI21_X1 U8493 ( .B1(n9835), .B2(n6119), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6781) );
  INV_X1 U8494 ( .A(n9835), .ZN(n9326) );
  INV_X1 U8495 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8496 ( .A1(n9326), .A2(n6779), .ZN(n6780) );
  NAND2_X1 U8497 ( .A1(n9327), .A2(n6780), .ZN(n6985) );
  MUX2_X1 U8498 ( .A(n6781), .B(P1_IR_REG_0__SCAN_IN), .S(n6985), .Z(n6782) );
  AND4_X1 U8499 ( .A1(n6785), .A2(P1_STATE_REG_SCAN_IN), .A3(n6783), .A4(n6782), .ZN(n6784) );
  AOI21_X1 U8500 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n6784), .ZN(
        n6787) );
  NAND2_X1 U8501 ( .A1(n6785), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6821) );
  OR3_X1 U8502 ( .A1(n6821), .A2(n9326), .A3(n8145), .ZN(n9901) );
  NAND3_X1 U8503 ( .A1(n9917), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6119), .ZN(
        n6786) );
  OAI211_X1 U8504 ( .C1(n6788), .C2(n9923), .A(n6787), .B(n6786), .ZN(P1_U3241) );
  NAND2_X1 U8505 ( .A1(n9059), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8506 ( .A1(n9058), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8507 ( .A1(n4390), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6789) );
  AND3_X1 U8508 ( .A1(n6791), .A2(n6790), .A3(n6789), .ZN(n9053) );
  INV_X1 U8509 ( .A(n9053), .ZN(n9452) );
  NAND2_X1 U8510 ( .A1(P1_U4006), .A2(n9452), .ZN(n6792) );
  OAI21_X1 U8511 ( .B1(P1_U4006), .B2(n5811), .A(n6792), .ZN(P1_U3586) );
  INV_X1 U8512 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U8513 ( .A1(P1_U4006), .A2(n7052), .ZN(n6793) );
  OAI21_X1 U8514 ( .B1(P1_U4006), .B2(n10430), .A(n6793), .ZN(P1_U3555) );
  INV_X1 U8515 ( .A(n6794), .ZN(n6796) );
  INV_X1 U8516 ( .A(n7689), .ZN(n7685) );
  OAI222_X1 U8517 ( .A1(n9837), .A2(n6795), .B1(n9840), .B2(n6796), .C1(
        P1_U3084), .C2(n7685), .ZN(P1_U3341) );
  OAI222_X1 U8518 ( .A1(n8093), .A2(n6797), .B1(n8906), .B2(n6796), .C1(
        P2_U3152), .C2(n7345), .ZN(P2_U3346) );
  INV_X1 U8519 ( .A(n6798), .ZN(n6844) );
  AOI22_X1 U8520 ( .A1(n9375), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9828), .ZN(n6799) );
  OAI21_X1 U8521 ( .B1(n6844), .B2(n9840), .A(n6799), .ZN(P1_U3340) );
  OR2_X1 U8522 ( .A1(n9939), .A2(n6618), .ZN(n6803) );
  AND2_X1 U8523 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  INV_X1 U8524 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6808) );
  NOR2_X2 U8525 ( .A1(n6924), .A2(n7456), .ZN(n7450) );
  AND2_X1 U8526 ( .A1(n7052), .A2(n7456), .ZN(n9286) );
  NOR2_X1 U8527 ( .A1(n7450), .A2(n9286), .ZN(n9180) );
  NOR3_X1 U8528 ( .A1(n9180), .A2(n6805), .A3(n6804), .ZN(n6806) );
  AOI21_X1 U8529 ( .B1(n9660), .B2(n9365), .A(n6806), .ZN(n7115) );
  OAI21_X1 U8530 ( .B1(n7456), .B2(n7120), .A(n7115), .ZN(n6922) );
  NAND2_X1 U8531 ( .A1(n6922), .A2(n10175), .ZN(n6807) );
  OAI21_X1 U8532 ( .B1(n10175), .B2(n6808), .A(n6807), .ZN(P1_U3454) );
  INV_X1 U8533 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6809) );
  MUX2_X1 U8534 ( .A(n6809), .B(P1_REG2_REG_7__SCAN_IN), .S(n6910), .Z(n6820)
         );
  INV_X1 U8535 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6818) );
  INV_X1 U8536 ( .A(n6830), .ZN(n6992) );
  INV_X1 U8537 ( .A(n8044), .ZN(n6813) );
  INV_X1 U8538 ( .A(n6823), .ZN(n9882) );
  NAND2_X1 U8539 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9879) );
  NOR2_X1 U8540 ( .A1(n9878), .A2(n9879), .ZN(n9877) );
  INV_X1 U8541 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8542 ( .A(n6811), .B(P1_REG2_REG_2__SCAN_IN), .S(n8044), .Z(n6812)
         );
  INV_X1 U8543 ( .A(n6812), .ZN(n7028) );
  INV_X1 U8544 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6814) );
  XNOR2_X1 U8545 ( .A(n6830), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6990) );
  INV_X1 U8546 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6817) );
  XNOR2_X1 U8547 ( .A(n6877), .B(n6817), .ZN(n6875) );
  XOR2_X1 U8548 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6833), .Z(n6856) );
  AOI21_X1 U8549 ( .B1(n6820), .B2(n6819), .A(n9891), .ZN(n6843) );
  OR2_X1 U8550 ( .A1(n6821), .A2(n9835), .ZN(n6840) );
  INV_X1 U8551 ( .A(n9923), .ZN(n9397) );
  AND2_X1 U8552 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7358) );
  INV_X1 U8553 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6822) );
  MUX2_X1 U8554 ( .A(n6822), .B(P1_REG1_REG_2__SCAN_IN), .S(n8044), .Z(n7031)
         );
  INV_X1 U8555 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6824) );
  MUX2_X1 U8556 ( .A(n6824), .B(P1_REG1_REG_1__SCAN_IN), .S(n6823), .Z(n9884)
         );
  AND2_X1 U8557 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9885) );
  NAND2_X1 U8558 ( .A1(n9884), .A2(n9885), .ZN(n9883) );
  NAND2_X1 U8559 ( .A1(n9882), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8560 ( .A1(n9883), .A2(n6825), .ZN(n7032) );
  NAND2_X1 U8561 ( .A1(n7031), .A2(n7032), .ZN(n7030) );
  OR2_X1 U8562 ( .A1(n8044), .A2(n6822), .ZN(n6866) );
  NAND2_X1 U8563 ( .A1(n7030), .A2(n6866), .ZN(n6828) );
  INV_X1 U8564 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6826) );
  MUX2_X1 U8565 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6826), .S(n6865), .Z(n6827)
         );
  NAND2_X1 U8566 ( .A1(n6828), .A2(n6827), .ZN(n6869) );
  NAND2_X1 U8567 ( .A1(n6865), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6829) );
  AND2_X1 U8568 ( .A1(n6869), .A2(n6829), .ZN(n6995) );
  INV_X1 U8569 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6953) );
  MUX2_X1 U8570 ( .A(n6953), .B(P1_REG1_REG_4__SCAN_IN), .S(n6830), .Z(n6994)
         );
  NAND2_X1 U8571 ( .A1(n6995), .A2(n6994), .ZN(n6993) );
  NAND2_X1 U8572 ( .A1(n6830), .A2(n6953), .ZN(n6831) );
  NAND2_X1 U8573 ( .A1(n6993), .A2(n6831), .ZN(n6882) );
  INV_X1 U8574 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9971) );
  MUX2_X1 U8575 ( .A(n9971), .B(P1_REG1_REG_5__SCAN_IN), .S(n6877), .Z(n6881)
         );
  OR2_X1 U8576 ( .A1(n6882), .A2(n6881), .ZN(n6879) );
  NAND2_X1 U8577 ( .A1(n6877), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6832) );
  AND2_X1 U8578 ( .A1(n6879), .A2(n6832), .ZN(n6850) );
  INV_X1 U8579 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U8580 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9972), .S(n6833), .Z(n6849)
         );
  NAND2_X1 U8581 ( .A1(n6850), .A2(n6849), .ZN(n6848) );
  OR2_X1 U8582 ( .A1(n6833), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8583 ( .A1(n6848), .A2(n6836), .ZN(n6834) );
  INV_X1 U8584 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9975) );
  MUX2_X1 U8585 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9975), .S(n6910), .Z(n6835)
         );
  NAND2_X1 U8586 ( .A1(n6834), .A2(n6835), .ZN(n6906) );
  INV_X1 U8587 ( .A(n6835), .ZN(n6837) );
  NAND3_X1 U8588 ( .A1(n6848), .A2(n6837), .A3(n6836), .ZN(n6838) );
  AOI21_X1 U8589 ( .B1(n6906), .B2(n6838), .A(n9901), .ZN(n6839) );
  AOI211_X1 U8590 ( .C1(n9397), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7358), .B(
        n6839), .ZN(n6842) );
  OR2_X1 U8591 ( .A1(n6840), .A2(n9327), .ZN(n9888) );
  NAND2_X1 U8592 ( .A1(n9910), .A2(n6910), .ZN(n6841) );
  OAI211_X1 U8593 ( .C1(n6843), .C2(n9893), .A(n6842), .B(n6841), .ZN(P1_U3248) );
  OAI222_X1 U8594 ( .A1(n8093), .A2(n6845), .B1(n8906), .B2(n6844), .C1(n7365), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8595 ( .A(n6846), .ZN(n6886) );
  AOI22_X1 U8596 ( .A1(n7483), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n8903), .ZN(n6847) );
  OAI21_X1 U8597 ( .B1(n6886), .B2(n8906), .A(n6847), .ZN(P2_U3344) );
  OAI21_X1 U8598 ( .B1(n6850), .B2(n6849), .A(n6848), .ZN(n6854) );
  NAND2_X1 U8599 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7577) );
  INV_X1 U8600 ( .A(n7577), .ZN(n6853) );
  INV_X1 U8601 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U8602 ( .A1(n9923), .A2(n6851), .ZN(n6852) );
  AOI211_X1 U8603 ( .C1(n9917), .C2(n6854), .A(n6853), .B(n6852), .ZN(n6859)
         );
  INV_X1 U8604 ( .A(n9893), .ZN(n9918) );
  OAI211_X1 U8605 ( .C1(n6857), .C2(n6856), .A(n6855), .B(n9918), .ZN(n6858)
         );
  OAI211_X1 U8606 ( .C1(n9888), .C2(n6860), .A(n6859), .B(n6858), .ZN(P1_U3247) );
  INV_X1 U8607 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6874) );
  AOI211_X1 U8608 ( .C1(n6863), .C2(n6862), .A(n6861), .B(n9893), .ZN(n6864)
         );
  AOI21_X1 U8609 ( .B1(n9910), .B2(n6865), .A(n6864), .ZN(n6873) );
  MUX2_X1 U8610 ( .A(n6826), .B(P1_REG1_REG_3__SCAN_IN), .S(n6865), .Z(n6867)
         );
  NAND3_X1 U8611 ( .A1(n6867), .A2(n7030), .A3(n6866), .ZN(n6868) );
  AND3_X1 U8612 ( .A1(n9917), .A2(n6869), .A3(n6868), .ZN(n6871) );
  NOR2_X1 U8613 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6133), .ZN(n6870) );
  NOR2_X1 U8614 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  OAI211_X1 U8615 ( .C1(n6874), .C2(n9923), .A(n6873), .B(n6872), .ZN(P1_U3244) );
  INV_X1 U8616 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10469) );
  XNOR2_X1 U8617 ( .A(n6876), .B(n6875), .ZN(n6878) );
  AOI22_X1 U8618 ( .A1(n6878), .A2(n9918), .B1(n6877), .B2(n9910), .ZN(n6885)
         );
  INV_X1 U8619 ( .A(n6879), .ZN(n6880) );
  AOI211_X1 U8620 ( .C1(n6882), .C2(n6881), .A(n6880), .B(n9901), .ZN(n6883)
         );
  AND2_X1 U8621 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7464) );
  NOR2_X1 U8622 ( .A1(n6883), .A2(n7464), .ZN(n6884) );
  OAI211_X1 U8623 ( .C1(n10469), .C2(n9923), .A(n6885), .B(n6884), .ZN(
        P1_U3246) );
  INV_X1 U8624 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6887) );
  INV_X1 U8625 ( .A(n9909), .ZN(n9376) );
  OAI222_X1 U8626 ( .A1(n9837), .A2(n6887), .B1(n9840), .B2(n6886), .C1(n9376), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8627 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6904) );
  XNOR2_X1 U8628 ( .A(n4388), .B(n7473), .ZN(n9178) );
  XNOR2_X1 U8629 ( .A(n7080), .B(n7457), .ZN(n9177) );
  NOR2_X1 U8630 ( .A1(n9177), .A2(n6925), .ZN(n7447) );
  AOI21_X1 U8631 ( .B1(n7049), .B2(n9365), .A(n7447), .ZN(n6888) );
  XOR2_X1 U8632 ( .A(n9178), .B(n6888), .Z(n6901) );
  INV_X1 U8633 ( .A(n6901), .ZN(n7478) );
  NAND2_X1 U8634 ( .A1(n6890), .A2(n6889), .ZN(n6893) );
  NAND3_X1 U8635 ( .A1(n9328), .A2(n6618), .A3(n6891), .ZN(n6892) );
  NAND2_X1 U8636 ( .A1(n9177), .A2(n7450), .ZN(n7449) );
  INV_X1 U8637 ( .A(n6938), .ZN(n6894) );
  NAND2_X1 U8638 ( .A1(n7449), .A2(n6894), .ZN(n9292) );
  XOR2_X1 U8639 ( .A(n9178), .B(n9292), .Z(n6899) );
  NAND2_X1 U8640 ( .A1(n6084), .A2(n9521), .ZN(n6896) );
  NAND2_X1 U8641 ( .A1(n6618), .A2(n9340), .ZN(n6895) );
  AOI22_X1 U8642 ( .A1(n9660), .A2(n9363), .B1(n9659), .B2(n9365), .ZN(n6898)
         );
  OAI21_X1 U8643 ( .B1(n6899), .B2(n9628), .A(n6898), .ZN(n6900) );
  AOI21_X1 U8644 ( .B1(n6901), .B2(n9665), .A(n6900), .ZN(n7471) );
  NOR2_X2 U8645 ( .A1(n7455), .A2(n7076), .ZN(n7675) );
  AOI21_X1 U8646 ( .B1(n7076), .B2(n7455), .A(n7675), .ZN(n7475) );
  AOI22_X1 U8647 ( .A1(n7475), .A2(n9935), .B1(n9934), .B2(n7076), .ZN(n6902)
         );
  OAI211_X1 U8648 ( .C1(n7478), .C2(n9939), .A(n7471), .B(n6902), .ZN(n9800)
         );
  NAND2_X1 U8649 ( .A1(n9800), .A2(n10175), .ZN(n6903) );
  OAI21_X1 U8650 ( .B1(n10175), .B2(n6904), .A(n6903), .ZN(P1_U3460) );
  XNOR2_X1 U8651 ( .A(n7007), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7002) );
  OR2_X1 U8652 ( .A1(n6910), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8653 ( .A1(n6906), .A2(n6905), .ZN(n9902) );
  NAND2_X1 U8654 ( .A1(n9899), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6907) );
  NOR2_X1 U8655 ( .A1(n9899), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9903) );
  AOI21_X1 U8656 ( .B1(n9902), .B2(n6907), .A(n9903), .ZN(n9900) );
  XOR2_X1 U8657 ( .A(n7002), .B(n9900), .Z(n6918) );
  INV_X1 U8658 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8659 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n6908) );
  OAI21_X1 U8660 ( .B1(n9923), .B2(n6909), .A(n6908), .ZN(n6916) );
  XNOR2_X1 U8661 ( .A(n7007), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6914) );
  INV_X1 U8662 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6911) );
  MUX2_X1 U8663 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6911), .S(n9899), .Z(n6912)
         );
  OAI21_X1 U8664 ( .B1(n9899), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9895), .ZN(
        n6913) );
  AOI211_X1 U8665 ( .C1(n6914), .C2(n6913), .A(n9893), .B(n7006), .ZN(n6915)
         );
  AOI211_X1 U8666 ( .C1(n9910), .C2(n7007), .A(n6916), .B(n6915), .ZN(n6917)
         );
  OAI21_X1 U8667 ( .B1(n9901), .B2(n6918), .A(n6917), .ZN(P1_U3250) );
  NOR2_X1 U8668 ( .A1(n7047), .A2(n6919), .ZN(n6920) );
  NAND2_X1 U8669 ( .A1(n6922), .A2(n9977), .ZN(n6923) );
  OAI21_X1 U8670 ( .B1(n9977), .B2(n6119), .A(n6923), .ZN(P1_U3523) );
  INV_X1 U8671 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6950) );
  NAND2_X1 U8672 ( .A1(n6924), .A2(n7122), .ZN(n6925) );
  NAND2_X1 U8673 ( .A1(n6925), .A2(n7080), .ZN(n6930) );
  NAND2_X1 U8674 ( .A1(n6930), .A2(n7049), .ZN(n6927) );
  NAND2_X1 U8675 ( .A1(n6926), .A2(n9365), .ZN(n6929) );
  NAND3_X1 U8676 ( .A1(n6927), .A2(n6929), .A3(n4388), .ZN(n6928) );
  NAND2_X1 U8677 ( .A1(n6928), .A2(n7076), .ZN(n6932) );
  NAND3_X1 U8678 ( .A1(n6930), .A2(n9364), .A3(n7049), .ZN(n6931) );
  NAND3_X1 U8679 ( .A1(n6932), .A2(n5066), .A3(n6931), .ZN(n7669) );
  INV_X1 U8680 ( .A(n7669), .ZN(n6934) );
  NAND2_X1 U8681 ( .A1(n9363), .A2(n6935), .ZN(n9259) );
  AND2_X2 U8682 ( .A1(n9293), .A2(n9259), .ZN(n9179) );
  NAND2_X1 U8683 ( .A1(n7074), .A2(n6935), .ZN(n6936) );
  NAND2_X1 U8684 ( .A1(n7670), .A2(n6936), .ZN(n6937) );
  NAND2_X1 U8685 ( .A1(n7667), .A2(n6946), .ZN(n9299) );
  INV_X1 U8686 ( .A(n7667), .ZN(n9361) );
  NAND2_X1 U8687 ( .A1(n9361), .A2(n7497), .ZN(n9265) );
  NAND2_X1 U8688 ( .A1(n9299), .A2(n9265), .ZN(n9181) );
  NAND2_X1 U8689 ( .A1(n6937), .A2(n9181), .ZN(n7126) );
  OAI21_X1 U8690 ( .B1(n6937), .B2(n9181), .A(n7126), .ZN(n7499) );
  INV_X1 U8691 ( .A(n7499), .ZN(n6948) );
  NAND2_X1 U8692 ( .A1(n9365), .A2(n7457), .ZN(n9287) );
  NAND3_X1 U8693 ( .A1(n9287), .A2(n9295), .A3(n7450), .ZN(n6940) );
  NAND2_X1 U8694 ( .A1(n6938), .A2(n9295), .ZN(n6939) );
  NAND2_X1 U8695 ( .A1(n7666), .A2(n9179), .ZN(n7132) );
  NAND2_X1 U8696 ( .A1(n7132), .A2(n9293), .ZN(n6941) );
  XNOR2_X1 U8697 ( .A(n6941), .B(n9181), .ZN(n6943) );
  AOI22_X1 U8698 ( .A1(n9660), .A2(n9360), .B1(n9659), .B2(n9363), .ZN(n6942)
         );
  OAI21_X1 U8699 ( .B1(n6943), .B2(n9628), .A(n6942), .ZN(n6944) );
  AOI21_X1 U8700 ( .B1(n7499), .B2(n9665), .A(n6944), .ZN(n7501) );
  NAND2_X1 U8701 ( .A1(n7676), .A2(n6946), .ZN(n6945) );
  AND2_X1 U8702 ( .A1(n7137), .A2(n6945), .ZN(n7494) );
  AOI22_X1 U8703 ( .A1(n7494), .A2(n9935), .B1(n9934), .B2(n6946), .ZN(n6947)
         );
  OAI211_X1 U8704 ( .C1(n6948), .C2(n9939), .A(n7501), .B(n6947), .ZN(n6951)
         );
  NAND2_X1 U8705 ( .A1(n6951), .A2(n10175), .ZN(n6949) );
  OAI21_X1 U8706 ( .B1(n10175), .B2(n6950), .A(n6949), .ZN(P1_U3466) );
  NAND2_X1 U8707 ( .A1(n6951), .A2(n9977), .ZN(n6952) );
  OAI21_X1 U8708 ( .B1(n9977), .B2(n6953), .A(n6952), .ZN(P1_U3527) );
  INV_X1 U8709 ( .A(n6954), .ZN(n6956) );
  AND2_X1 U8710 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  NAND2_X1 U8711 ( .A1(n6958), .A2(n6957), .ZN(n6963) );
  INV_X1 U8712 ( .A(n6959), .ZN(n6960) );
  NAND2_X1 U8713 ( .A1(n6976), .A2(n6960), .ZN(n6961) );
  NAND2_X1 U8714 ( .A1(n6963), .A2(n6962), .ZN(n6970) );
  INV_X1 U8715 ( .A(n6964), .ZN(n6965) );
  OR2_X1 U8716 ( .A1(n6966), .A2(n6965), .ZN(n6967) );
  NOR2_X1 U8717 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  NAND2_X1 U8718 ( .A1(n6970), .A2(n6969), .ZN(n8121) );
  AND2_X1 U8719 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9980) );
  INV_X1 U8720 ( .A(n6971), .ZN(n6972) );
  INV_X1 U8721 ( .A(n8415), .ZN(n8292) );
  NAND2_X1 U8722 ( .A1(n5682), .A2(n10017), .ZN(n7542) );
  NOR2_X1 U8723 ( .A1(n8292), .A2(n7542), .ZN(n6973) );
  AOI211_X1 U8724 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n8121), .A(n9980), .B(
        n6973), .ZN(n6980) );
  NOR2_X1 U8725 ( .A1(n10096), .A2(n6974), .ZN(n6975) );
  INV_X2 U8726 ( .A(n8188), .ZN(n8251) );
  INV_X1 U8727 ( .A(n8451), .ZN(n6977) );
  OAI22_X1 U8728 ( .A1(n8402), .A2(n6977), .B1(n10046), .B2(n8426), .ZN(n6978)
         );
  NAND2_X1 U8729 ( .A1(n7583), .A2(n8188), .ZN(n7170) );
  NAND2_X1 U8730 ( .A1(n6978), .A2(n7170), .ZN(n6979) );
  OAI211_X1 U8731 ( .C1(n8425), .C2(n10046), .A(n6980), .B(n6979), .ZN(
        P2_U3234) );
  INV_X1 U8732 ( .A(n6981), .ZN(n6982) );
  AOI21_X1 U8733 ( .B1(n6984), .B2(n6983), .A(n6982), .ZN(n7079) );
  MUX2_X1 U8734 ( .A(n7079), .B(P1_IR_REG_0__SCAN_IN), .S(n9326), .Z(n6987) );
  MUX2_X1 U8735 ( .A(n6987), .B(n6986), .S(n6985), .Z(n6988) );
  INV_X1 U8736 ( .A(P1_U4006), .ZN(n9350) );
  NOR2_X1 U8737 ( .A1(n6988), .A2(n9350), .ZN(n7038) );
  OAI21_X1 U8738 ( .B1(n6990), .B2(n4486), .A(n6989), .ZN(n6991) );
  AOI22_X1 U8739 ( .A1(n6992), .A2(n9910), .B1(n9918), .B2(n6991), .ZN(n7000)
         );
  NAND2_X1 U8740 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6999) );
  NAND2_X1 U8741 ( .A1(n9397), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U8742 ( .B1(n6995), .B2(n6994), .A(n6993), .ZN(n6996) );
  NAND2_X1 U8743 ( .A1(n9917), .A2(n6996), .ZN(n6997) );
  NAND4_X1 U8744 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7001)
         );
  OR2_X1 U8745 ( .A1(n7038), .A2(n7001), .ZN(P1_U3245) );
  XOR2_X1 U8746 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7097), .Z(n7094) );
  OAI22_X1 U8747 ( .A1(n9900), .A2(n7002), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n7007), .ZN(n7095) );
  XOR2_X1 U8748 ( .A(n7094), .B(n7095), .Z(n7013) );
  INV_X1 U8749 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U8750 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7003), .ZN(n7662) );
  INV_X1 U8751 ( .A(n7662), .ZN(n7004) );
  OAI21_X1 U8752 ( .B1(n9923), .B2(n7005), .A(n7004), .ZN(n7011) );
  XNOR2_X1 U8753 ( .A(n7097), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7008) );
  AOI211_X1 U8754 ( .C1(n7009), .C2(n7008), .A(n9893), .B(n7096), .ZN(n7010)
         );
  AOI211_X1 U8755 ( .C1(n9910), .C2(n7097), .A(n7011), .B(n7010), .ZN(n7012)
         );
  OAI21_X1 U8756 ( .B1(n9901), .B2(n7013), .A(n7012), .ZN(P1_U3251) );
  NAND2_X1 U8757 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  XNOR2_X1 U8758 ( .A(n7017), .B(n7016), .ZN(n7021) );
  INV_X1 U8759 ( .A(n9042), .ZN(n8951) );
  AOI22_X1 U8760 ( .A1(n8951), .A2(n9364), .B1(n6133), .B2(n9039), .ZN(n7019)
         );
  AOI22_X1 U8761 ( .A1(n9040), .A2(n9361), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n7018) );
  OAI211_X1 U8762 ( .C1(n6935), .C2(n8996), .A(n7019), .B(n7018), .ZN(n7020)
         );
  AOI21_X1 U8763 ( .B1(n8986), .B2(n7021), .A(n7020), .ZN(n7022) );
  INV_X1 U8764 ( .A(n7022), .ZN(P1_U3216) );
  INV_X1 U8765 ( .A(n7023), .ZN(n7025) );
  OAI222_X1 U8766 ( .A1(n8093), .A2(n10176), .B1(n8906), .B2(n7025), .C1(
        P2_U3152), .C2(n7024), .ZN(P2_U3343) );
  OAI222_X1 U8767 ( .A1(n9837), .A2(n7026), .B1(n9840), .B2(n7025), .C1(
        P1_U3084), .C2(n9392), .ZN(P1_U3338) );
  AOI211_X1 U8768 ( .C1(n7029), .C2(n7028), .A(n7027), .B(n9893), .ZN(n7037)
         );
  INV_X1 U8769 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10274) );
  OAI211_X1 U8770 ( .C1(n7032), .C2(n7031), .A(n9917), .B(n7030), .ZN(n7033)
         );
  OAI21_X1 U8771 ( .B1(n10274), .B2(n9923), .A(n7033), .ZN(n7034) );
  AOI21_X1 U8772 ( .B1(P1_U3084), .B2(P1_REG3_REG_2__SCAN_IN), .A(n7034), .ZN(
        n7035) );
  OAI21_X1 U8773 ( .B1(n9888), .B2(n8044), .A(n7035), .ZN(n7036) );
  OR3_X1 U8774 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(P1_U3243) );
  INV_X1 U8775 ( .A(n7039), .ZN(n7106) );
  AOI22_X1 U8776 ( .A1(n8509), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8903), .ZN(n7040) );
  OAI21_X1 U8777 ( .B1(n7106), .B2(n8906), .A(n7040), .ZN(P2_U3342) );
  INV_X1 U8778 ( .A(n7041), .ZN(n7044) );
  INV_X1 U8779 ( .A(n7042), .ZN(n7043) );
  NAND2_X1 U8780 ( .A1(n7044), .A2(n7043), .ZN(n7067) );
  OAI21_X1 U8781 ( .B1(n7044), .B2(n7043), .A(n7067), .ZN(n7045) );
  NOR2_X1 U8782 ( .A1(n7045), .A2(n7046), .ZN(n7070) );
  AOI21_X1 U8783 ( .B1(n7046), .B2(n7045), .A(n7070), .ZN(n7054) );
  OAI21_X1 U8784 ( .B1(n7048), .B2(n7047), .A(n8996), .ZN(n7083) );
  INV_X1 U8785 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9875) );
  NOR2_X1 U8786 ( .A1(n7083), .A2(n9875), .ZN(n7051) );
  NAND2_X1 U8787 ( .A1(n9934), .A2(n7049), .ZN(n9929) );
  OAI22_X1 U8788 ( .A1(n9011), .A2(n4388), .B1(n9929), .B2(n7361), .ZN(n7050)
         );
  AOI211_X1 U8789 ( .C1(n8951), .C2(n7052), .A(n7051), .B(n7050), .ZN(n7053)
         );
  OAI21_X1 U8790 ( .B1(n7054), .B2(n9047), .A(n7053), .ZN(P1_U3220) );
  INV_X1 U8791 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10479) );
  OAI211_X1 U8792 ( .C1(n7057), .C2(n7056), .A(n9978), .B(n7055), .ZN(n7059)
         );
  NAND2_X1 U8793 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n7058) );
  OAI211_X1 U8794 ( .C1(n8522), .C2(n10479), .A(n7059), .B(n7058), .ZN(n7060)
         );
  INV_X1 U8795 ( .A(n7060), .ZN(n7065) );
  OAI211_X1 U8796 ( .C1(n7063), .C2(n7062), .A(n9979), .B(n7061), .ZN(n7064)
         );
  OAI211_X1 U8797 ( .C1(n9983), .C2(n7066), .A(n7065), .B(n7064), .ZN(P2_U3252) );
  INV_X1 U8798 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7472) );
  INV_X1 U8799 ( .A(n7067), .ZN(n7068) );
  NOR3_X1 U8800 ( .A1(n7070), .A2(n7069), .A3(n7068), .ZN(n7073) );
  INV_X1 U8801 ( .A(n7071), .ZN(n7072) );
  OAI21_X1 U8802 ( .B1(n7073), .B2(n7072), .A(n8986), .ZN(n7078) );
  OAI22_X1 U8803 ( .A1(n9011), .A2(n7074), .B1(n7080), .B2(n9042), .ZN(n7075)
         );
  AOI21_X1 U8804 ( .B1(n9045), .B2(n7076), .A(n7075), .ZN(n7077) );
  OAI211_X1 U8805 ( .C1(n7472), .C2(n7083), .A(n7078), .B(n7077), .ZN(P1_U3235) );
  INV_X1 U8806 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7116) );
  OAI22_X1 U8807 ( .A1(n9011), .A2(n7080), .B1(n7079), .B2(n9047), .ZN(n7081)
         );
  AOI21_X1 U8808 ( .B1(n7122), .B2(n9045), .A(n7081), .ZN(n7082) );
  OAI21_X1 U8809 ( .B1(n7116), .B2(n7083), .A(n7082), .ZN(P1_U3230) );
  NAND2_X1 U8810 ( .A1(n7085), .A2(n7084), .ZN(n7086) );
  AOI21_X1 U8811 ( .B1(n7087), .B2(n7086), .A(n9047), .ZN(n7091) );
  AOI22_X1 U8812 ( .A1(n8951), .A2(n9363), .B1(n7493), .B2(n9039), .ZN(n7089)
         );
  AOI22_X1 U8813 ( .A1(n9040), .A2(n9360), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3084), .ZN(n7088) );
  OAI211_X1 U8814 ( .C1(n7497), .C2(n8996), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OR2_X1 U8815 ( .A1(n7091), .A2(n7090), .ZN(P1_U3228) );
  XNOR2_X1 U8816 ( .A(n7439), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7435) );
  INV_X1 U8817 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7092) );
  AOI22_X1 U8818 ( .A1(n7095), .A2(n7094), .B1(n7093), .B2(n7092), .ZN(n7436)
         );
  XOR2_X1 U8819 ( .A(n7435), .B(n7436), .Z(n7105) );
  XOR2_X1 U8820 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7439), .Z(n7099) );
  NAND2_X1 U8821 ( .A1(n7098), .A2(n7099), .ZN(n7438) );
  OAI21_X1 U8822 ( .B1(n7099), .B2(n7098), .A(n7438), .ZN(n7100) );
  NAND2_X1 U8823 ( .A1(n7100), .A2(n9918), .ZN(n7104) );
  AND2_X1 U8824 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7791) );
  INV_X1 U8825 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7101) );
  NOR2_X1 U8826 ( .A1(n9923), .A2(n7101), .ZN(n7102) );
  AOI211_X1 U8827 ( .C1(n9910), .C2(n7439), .A(n7791), .B(n7102), .ZN(n7103)
         );
  OAI211_X1 U8828 ( .C1(n7105), .C2(n9901), .A(n7104), .B(n7103), .ZN(P1_U3252) );
  INV_X1 U8829 ( .A(n9413), .ZN(n9400) );
  OAI222_X1 U8830 ( .A1(n9837), .A2(n7107), .B1(n9840), .B2(n7106), .C1(n9400), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8831 ( .A(n7108), .ZN(n7111) );
  AOI22_X1 U8832 ( .A1(n8109), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n8903), .ZN(n7109) );
  OAI21_X1 U8833 ( .B1(n7111), .B2(n8906), .A(n7109), .ZN(P2_U3341) );
  AOI22_X1 U8834 ( .A1(n9426), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9828), .ZN(n7110) );
  OAI21_X1 U8835 ( .B1(n7111), .B2(n9840), .A(n7110), .ZN(P1_U3336) );
  NAND2_X1 U8836 ( .A1(n7113), .A2(n7112), .ZN(n7405) );
  NAND2_X1 U8837 ( .A1(n9925), .A2(n9210), .ZN(n7114) );
  OAI21_X1 U8838 ( .B1(n7116), .B2(n9637), .A(n7115), .ZN(n7117) );
  NAND2_X1 U8839 ( .A1(n7117), .A2(n7131), .ZN(n7124) );
  NOR2_X1 U8840 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  OAI21_X1 U8841 ( .B1(n9671), .B2(n9600), .A(n7122), .ZN(n7123) );
  OAI211_X1 U8842 ( .C1(n6779), .C2(n7131), .A(n7124), .B(n7123), .ZN(P1_U3291) );
  NAND2_X1 U8843 ( .A1(n7667), .A2(n7497), .ZN(n7125) );
  NAND2_X1 U8844 ( .A1(n7126), .A2(n7125), .ZN(n7146) );
  INV_X1 U8845 ( .A(n7146), .ZN(n7127) );
  NAND2_X1 U8846 ( .A1(n7423), .A2(n7144), .ZN(n9300) );
  NAND2_X1 U8847 ( .A1(n9966), .A2(n9360), .ZN(n9266) );
  AND2_X1 U8848 ( .A1(n9266), .A2(n9300), .ZN(n7147) );
  INV_X1 U8849 ( .A(n7147), .ZN(n9182) );
  NAND2_X1 U8850 ( .A1(n7127), .A2(n9182), .ZN(n7420) );
  NAND2_X1 U8851 ( .A1(n7146), .A2(n7147), .ZN(n7128) );
  NAND2_X1 U8852 ( .A1(n7420), .A2(n7128), .ZN(n9963) );
  AND2_X1 U8853 ( .A1(n7129), .A2(n9331), .ZN(n7130) );
  AOI22_X1 U8854 ( .A1(n9671), .A2(n7144), .B1(n9679), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7143) );
  NAND2_X1 U8855 ( .A1(n7132), .A2(n9264), .ZN(n7133) );
  XNOR2_X1 U8856 ( .A(n4381), .B(n9182), .ZN(n7134) );
  NAND2_X1 U8857 ( .A1(n7134), .A2(n9656), .ZN(n7136) );
  AOI22_X1 U8858 ( .A1(n9660), .A2(n9359), .B1(n9659), .B2(n9361), .ZN(n7135)
         );
  NAND2_X1 U8859 ( .A1(n7136), .A2(n7135), .ZN(n9968) );
  AOI21_X1 U8860 ( .B1(n7137), .B2(n7144), .A(n9944), .ZN(n7139) );
  NAND2_X1 U8861 ( .A1(n7139), .A2(n7428), .ZN(n9964) );
  INV_X1 U8862 ( .A(n7465), .ZN(n7140) );
  OAI22_X1 U8863 ( .A1(n9964), .A2(n9521), .B1(n9637), .B2(n7140), .ZN(n7141)
         );
  OAI21_X1 U8864 ( .B1(n9968), .B2(n7141), .A(n7131), .ZN(n7142) );
  OAI211_X1 U8865 ( .C1(n9963), .C2(n9645), .A(n7143), .B(n7142), .ZN(P1_U3286) );
  INV_X1 U8866 ( .A(n9939), .ZN(n9949) );
  OR2_X1 U8867 ( .A1(n7356), .A2(n9943), .ZN(n9260) );
  NAND2_X1 U8868 ( .A1(n9943), .A2(n7356), .ZN(n9301) );
  NAND2_X1 U8869 ( .A1(n9260), .A2(n9301), .ZN(n9085) );
  NAND2_X1 U8870 ( .A1(n9360), .A2(n7144), .ZN(n7419) );
  AND2_X1 U8871 ( .A1(n9085), .A2(n7419), .ZN(n7145) );
  NAND2_X1 U8872 ( .A1(n7146), .A2(n7145), .ZN(n7396) );
  OR2_X1 U8873 ( .A1(n7404), .A2(n7741), .ZN(n9262) );
  NAND2_X1 U8874 ( .A1(n7404), .A2(n7741), .ZN(n9086) );
  NAND2_X1 U8875 ( .A1(n9262), .A2(n9086), .ZN(n7150) );
  NAND3_X1 U8876 ( .A1(n9085), .A2(n7147), .A3(n7419), .ZN(n7149) );
  OR2_X1 U8877 ( .A1(n9359), .A2(n9943), .ZN(n7148) );
  NAND2_X1 U8878 ( .A1(n7149), .A2(n7148), .ZN(n7394) );
  NAND2_X1 U8879 ( .A1(n7394), .A2(n7150), .ZN(n7152) );
  OR2_X1 U8880 ( .A1(n7404), .A2(n9358), .ZN(n7151) );
  OAI211_X1 U8881 ( .C1(n7396), .C2(n9185), .A(n7152), .B(n7151), .ZN(n7154)
         );
  NAND2_X1 U8882 ( .A1(n7154), .A2(n9186), .ZN(n7155) );
  NAND2_X1 U8883 ( .A1(n7503), .A2(n7155), .ZN(n7163) );
  INV_X1 U8884 ( .A(n7163), .ZN(n7392) );
  INV_X1 U8885 ( .A(n7404), .ZN(n7407) );
  NAND2_X1 U8886 ( .A1(n7401), .A2(n7407), .ZN(n7156) );
  INV_X1 U8887 ( .A(n7156), .ZN(n7402) );
  INV_X1 U8888 ( .A(n7743), .ZN(n7157) );
  OAI21_X1 U8889 ( .B1(n7402), .B2(n7157), .A(n5060), .ZN(n7388) );
  OAI22_X1 U8890 ( .A1(n7388), .A2(n9944), .B1(n7157), .B2(n9965), .ZN(n7164)
         );
  AOI22_X1 U8891 ( .A1(n9660), .A2(n9356), .B1(n9659), .B2(n9358), .ZN(n7162)
         );
  INV_X1 U8892 ( .A(n9266), .ZN(n9261) );
  NAND2_X1 U8893 ( .A1(n7422), .A2(n9260), .ZN(n7159) );
  NAND2_X1 U8894 ( .A1(n7159), .A2(n9301), .ZN(n7399) );
  NAND2_X1 U8895 ( .A1(n7399), .A2(n9185), .ZN(n7398) );
  NAND2_X1 U8896 ( .A1(n7398), .A2(n9086), .ZN(n7505) );
  XNOR2_X1 U8897 ( .A(n7505), .B(n9186), .ZN(n7160) );
  NAND2_X1 U8898 ( .A1(n7160), .A2(n9656), .ZN(n7161) );
  OAI211_X1 U8899 ( .C1(n7163), .C2(n9688), .A(n7162), .B(n7161), .ZN(n7389)
         );
  AOI211_X1 U8900 ( .C1(n9949), .C2(n7392), .A(n7164), .B(n7389), .ZN(n7335)
         );
  NAND2_X1 U8901 ( .A1(n9974), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7165) );
  OAI21_X1 U8902 ( .B1(n7335), .B2(n9974), .A(n7165), .ZN(P1_U3531) );
  NAND2_X1 U8903 ( .A1(n5682), .A2(n8188), .ZN(n7174) );
  XNOR2_X1 U8904 ( .A(n7173), .B(n7174), .ZN(n8272) );
  INV_X1 U8905 ( .A(n8272), .ZN(n7172) );
  NAND2_X1 U8906 ( .A1(n10046), .A2(n7176), .ZN(n7169) );
  INV_X1 U8907 ( .A(n8271), .ZN(n7171) );
  NAND2_X1 U8908 ( .A1(n7172), .A2(n7171), .ZN(n8270) );
  NAND2_X1 U8909 ( .A1(n7174), .A2(n7173), .ZN(n7175) );
  XNOR2_X1 U8910 ( .A(n10057), .B(n7176), .ZN(n7177) );
  AND2_X1 U8911 ( .A1(n10016), .A2(n8188), .ZN(n7178) );
  NAND2_X1 U8912 ( .A1(n7177), .A2(n7178), .ZN(n7181) );
  INV_X1 U8913 ( .A(n7177), .ZN(n8238) );
  INV_X1 U8914 ( .A(n7178), .ZN(n7179) );
  NAND2_X1 U8915 ( .A1(n8238), .A2(n7179), .ZN(n7180) );
  AND2_X1 U8916 ( .A1(n7181), .A2(n7180), .ZN(n8124) );
  NAND2_X1 U8917 ( .A1(n8123), .A2(n7181), .ZN(n7186) );
  XNOR2_X1 U8918 ( .A(n10032), .B(n7176), .ZN(n8352) );
  AND2_X1 U8919 ( .A1(n8450), .A2(n8188), .ZN(n7182) );
  NAND2_X1 U8920 ( .A1(n8352), .A2(n7182), .ZN(n7187) );
  INV_X1 U8921 ( .A(n8352), .ZN(n7184) );
  INV_X1 U8922 ( .A(n7182), .ZN(n7183) );
  NAND2_X1 U8923 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  AND2_X1 U8924 ( .A1(n7187), .A2(n7185), .ZN(n8240) );
  NAND2_X1 U8925 ( .A1(n10018), .A2(n8188), .ZN(n7190) );
  AND2_X1 U8926 ( .A1(n8360), .A2(n7187), .ZN(n7188) );
  INV_X1 U8927 ( .A(n7189), .ZN(n7191) );
  NAND2_X1 U8928 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  XNOR2_X1 U8929 ( .A(n7556), .B(n7176), .ZN(n7193) );
  AND2_X1 U8930 ( .A1(n8448), .A2(n8188), .ZN(n7194) );
  NAND2_X1 U8931 ( .A1(n7193), .A2(n7194), .ZN(n7198) );
  INV_X1 U8932 ( .A(n7193), .ZN(n8401) );
  INV_X1 U8933 ( .A(n7194), .ZN(n7195) );
  NAND2_X1 U8934 ( .A1(n8401), .A2(n7195), .ZN(n7196) );
  NAND2_X1 U8935 ( .A1(n7198), .A2(n7196), .ZN(n8315) );
  XNOR2_X1 U8936 ( .A(n10074), .B(n4379), .ZN(n7202) );
  NOR2_X1 U8937 ( .A1(n7210), .A2(n8251), .ZN(n7200) );
  XNOR2_X1 U8938 ( .A(n7202), .B(n7200), .ZN(n8400) );
  AND2_X1 U8939 ( .A1(n8400), .A2(n7198), .ZN(n7199) );
  INV_X1 U8940 ( .A(n7200), .ZN(n7201) );
  NAND2_X1 U8941 ( .A1(n7202), .A2(n7201), .ZN(n7203) );
  XNOR2_X1 U8942 ( .A(n10081), .B(n4379), .ZN(n7204) );
  NOR2_X1 U8943 ( .A1(n8391), .A2(n8251), .ZN(n7205) );
  NAND2_X1 U8944 ( .A1(n7204), .A2(n7205), .ZN(n7313) );
  INV_X1 U8945 ( .A(n7204), .ZN(n7312) );
  INV_X1 U8946 ( .A(n7205), .ZN(n7206) );
  NAND2_X1 U8947 ( .A1(n7312), .A2(n7206), .ZN(n7207) );
  AND2_X1 U8948 ( .A1(n7313), .A2(n7207), .ZN(n7208) );
  OAI211_X1 U8949 ( .C1(n7209), .C2(n7208), .A(n7314), .B(n8398), .ZN(n7214)
         );
  OAI22_X1 U8950 ( .A1(n7210), .A2(n9998), .B1(n7634), .B2(n10000), .ZN(n7297)
         );
  INV_X1 U8951 ( .A(n7297), .ZN(n7211) );
  OAI22_X1 U8952 ( .A1(n8292), .A2(n7211), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10227), .ZN(n7212) );
  AOI21_X1 U8953 ( .B1(n7303), .B2(n8420), .A(n7212), .ZN(n7213) );
  OAI211_X1 U8954 ( .C1(n7305), .C2(n8425), .A(n7214), .B(n7213), .ZN(P2_U3215) );
  INV_X1 U8955 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U8956 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8390) );
  OAI21_X1 U8957 ( .B1(n8522), .B2(n10465), .A(n8390), .ZN(n7220) );
  OAI21_X1 U8958 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(n7218) );
  NOR2_X1 U8959 ( .A1(n9984), .A2(n7218), .ZN(n7219) );
  AOI211_X1 U8960 ( .C1(n8510), .C2(n7221), .A(n7220), .B(n7219), .ZN(n7226)
         );
  OAI211_X1 U8961 ( .C1(n7224), .C2(n7223), .A(n9979), .B(n7222), .ZN(n7225)
         );
  NAND2_X1 U8962 ( .A1(n7226), .A2(n7225), .ZN(P2_U3251) );
  INV_X1 U8963 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U8964 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n7227) );
  OAI21_X1 U8965 ( .B1(n8522), .B2(n10315), .A(n7227), .ZN(n7233) );
  OAI21_X1 U8966 ( .B1(n7230), .B2(n7229), .A(n7228), .ZN(n7231) );
  NOR2_X1 U8967 ( .A1(n9984), .A2(n7231), .ZN(n7232) );
  AOI211_X1 U8968 ( .C1(n8510), .C2(n7234), .A(n7233), .B(n7232), .ZN(n7239)
         );
  OAI211_X1 U8969 ( .C1(n7237), .C2(n7236), .A(n9979), .B(n7235), .ZN(n7238)
         );
  NAND2_X1 U8970 ( .A1(n7239), .A2(n7238), .ZN(P2_U3248) );
  INV_X1 U8971 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7241) );
  INV_X1 U8972 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7240) );
  OAI22_X1 U8973 ( .A1(n8522), .A2(n7241), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7240), .ZN(n7247) );
  OAI21_X1 U8974 ( .B1(n7244), .B2(n7243), .A(n7242), .ZN(n7245) );
  NOR2_X1 U8975 ( .A1(n9984), .A2(n7245), .ZN(n7246) );
  AOI211_X1 U8976 ( .C1(n8510), .C2(n7248), .A(n7247), .B(n7246), .ZN(n7253)
         );
  OAI211_X1 U8977 ( .C1(n7251), .C2(n7250), .A(n9979), .B(n7249), .ZN(n7252)
         );
  NAND2_X1 U8978 ( .A1(n7253), .A2(n7252), .ZN(P2_U3247) );
  INV_X1 U8979 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7255) );
  NAND2_X1 U8980 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7254) );
  OAI21_X1 U8981 ( .B1(n8522), .B2(n7255), .A(n7254), .ZN(n7261) );
  OAI21_X1 U8982 ( .B1(n7258), .B2(n7257), .A(n7256), .ZN(n7259) );
  NOR2_X1 U8983 ( .A1(n9984), .A2(n7259), .ZN(n7260) );
  AOI211_X1 U8984 ( .C1(n8510), .C2(n7262), .A(n7261), .B(n7260), .ZN(n7267)
         );
  OAI211_X1 U8985 ( .C1(n7265), .C2(n7264), .A(n9979), .B(n7263), .ZN(n7266)
         );
  NAND2_X1 U8986 ( .A1(n7267), .A2(n7266), .ZN(P2_U3250) );
  INV_X1 U8987 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U8988 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7268) );
  OAI21_X1 U8989 ( .B1(n8522), .B2(n7269), .A(n7268), .ZN(n7275) );
  OAI21_X1 U8990 ( .B1(n7272), .B2(n7271), .A(n7270), .ZN(n7273) );
  NOR2_X1 U8991 ( .A1(n9984), .A2(n7273), .ZN(n7274) );
  AOI211_X1 U8992 ( .C1(n8510), .C2(n7276), .A(n7275), .B(n7274), .ZN(n7281)
         );
  OAI211_X1 U8993 ( .C1(n7279), .C2(n7278), .A(n9979), .B(n7277), .ZN(n7280)
         );
  NAND2_X1 U8994 ( .A1(n7281), .A2(n7280), .ZN(P2_U3249) );
  AOI21_X1 U8995 ( .B1(n7283), .B2(n7282), .A(n4484), .ZN(n7293) );
  INV_X1 U8996 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7285) );
  OAI22_X1 U8997 ( .A1(n8522), .A2(n7285), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7284), .ZN(n7286) );
  AOI21_X1 U8998 ( .B1(n8510), .B2(n7287), .A(n7286), .ZN(n7292) );
  OAI211_X1 U8999 ( .C1(n7290), .C2(n7289), .A(n7288), .B(n9978), .ZN(n7291)
         );
  OAI211_X1 U9000 ( .C1(n7293), .C2(n9982), .A(n7292), .B(n7291), .ZN(P2_U3256) );
  XNOR2_X1 U9001 ( .A(n7294), .B(n7295), .ZN(n10084) );
  XNOR2_X1 U9002 ( .A(n7296), .B(n7295), .ZN(n7298) );
  AOI21_X1 U9003 ( .B1(n7298), .B2(n10020), .A(n7297), .ZN(n10082) );
  MUX2_X1 U9004 ( .A(n7299), .B(n10082), .S(n10027), .Z(n7308) );
  INV_X1 U9005 ( .A(n7300), .ZN(n7562) );
  INV_X1 U9006 ( .A(n7301), .ZN(n7302) );
  AOI211_X1 U9007 ( .C1(n10081), .C2(n7562), .A(n10113), .B(n7302), .ZN(n10080) );
  INV_X1 U9008 ( .A(n7303), .ZN(n7304) );
  OAI22_X1 U9009 ( .A1(n10031), .A2(n7305), .B1(n10026), .B2(n7304), .ZN(n7306) );
  AOI21_X1 U9010 ( .B1(n10080), .B2(n8720), .A(n7306), .ZN(n7307) );
  OAI211_X1 U9011 ( .C1(n10084), .C2(n8763), .A(n7308), .B(n7307), .ZN(
        P2_U3289) );
  NAND2_X1 U9012 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8463) );
  OAI21_X1 U9013 ( .B1(n8412), .B2(n7626), .A(n8463), .ZN(n7310) );
  OAI22_X1 U9014 ( .A1(n8391), .A2(n8383), .B1(n8392), .B2(n9997), .ZN(n7309)
         );
  AOI211_X1 U9015 ( .C1(n10088), .C2(n8386), .A(n7310), .B(n7309), .ZN(n7319)
         );
  XNOR2_X1 U9016 ( .A(n10088), .B(n7176), .ZN(n7701) );
  NOR2_X1 U9017 ( .A1(n7634), .A2(n8251), .ZN(n7702) );
  XNOR2_X1 U9018 ( .A(n7701), .B(n7702), .ZN(n7315) );
  INV_X1 U9019 ( .A(n7315), .ZN(n7311) );
  AOI21_X1 U9020 ( .B1(n7314), .B2(n7311), .A(n8426), .ZN(n7317) );
  NOR3_X1 U9021 ( .A1(n8402), .A2(n8391), .A3(n7312), .ZN(n7316) );
  OAI21_X1 U9022 ( .B1(n7317), .B2(n7316), .A(n7705), .ZN(n7318) );
  NAND2_X1 U9023 ( .A1(n7319), .A2(n7318), .ZN(P2_U3223) );
  NAND2_X1 U9024 ( .A1(n7321), .A2(n7320), .ZN(n7322) );
  XOR2_X1 U9025 ( .A(n7328), .B(n7322), .Z(n10068) );
  INV_X1 U9026 ( .A(n7323), .ZN(n10024) );
  OAI211_X1 U9027 ( .C1(n10024), .C2(n10070), .A(n10097), .B(n7375), .ZN(
        n10069) );
  OAI22_X1 U9028 ( .A1(n8551), .A2(n10069), .B1(n7324), .B2(n10026), .ZN(n7326) );
  NOR2_X1 U9029 ( .A1(n10027), .A2(n6675), .ZN(n7325) );
  AOI211_X1 U9030 ( .C1(n8756), .C2(n8357), .A(n7326), .B(n7325), .ZN(n7331)
         );
  XNOR2_X1 U9031 ( .A(n7328), .B(n7327), .ZN(n7329) );
  AOI22_X1 U9032 ( .A1(n10017), .A2(n8448), .B1(n8450), .B2(n10015), .ZN(n8354) );
  OAI21_X1 U9033 ( .B1(n7329), .B2(n9995), .A(n8354), .ZN(n10072) );
  NAND2_X1 U9034 ( .A1(n10027), .A2(n10072), .ZN(n7330) );
  OAI211_X1 U9035 ( .C1(n10068), .C2(n8763), .A(n7331), .B(n7330), .ZN(
        P2_U3292) );
  INV_X1 U9036 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7333) );
  INV_X1 U9037 ( .A(n7332), .ZN(n7334) );
  INV_X1 U9038 ( .A(n8110), .ZN(n8530) );
  OAI222_X1 U9039 ( .A1(n8093), .A2(n7333), .B1(n8906), .B2(n7334), .C1(
        P2_U3152), .C2(n8530), .ZN(P2_U3340) );
  INV_X1 U9040 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10302) );
  INV_X1 U9041 ( .A(n9437), .ZN(n9424) );
  OAI222_X1 U9042 ( .A1(n9837), .A2(n10302), .B1(n9840), .B2(n7334), .C1(
        P1_U3084), .C2(n9424), .ZN(P1_U3335) );
  INV_X1 U9043 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7337) );
  OR2_X1 U9044 ( .A1(n7335), .A2(n10173), .ZN(n7336) );
  OAI21_X1 U9045 ( .B1(n10175), .B2(n7337), .A(n7336), .ZN(P1_U3478) );
  INV_X1 U9046 ( .A(n7338), .ZN(n7339) );
  AOI21_X1 U9047 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(n7349) );
  OAI211_X1 U9048 ( .C1(n7344), .C2(n7343), .A(n7342), .B(n9979), .ZN(n7348)
         );
  NOR2_X1 U9049 ( .A1(n10379), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7907) );
  NOR2_X1 U9050 ( .A1(n9983), .A2(n7345), .ZN(n7346) );
  AOI211_X1 U9051 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n9981), .A(n7907), .B(
        n7346), .ZN(n7347) );
  OAI211_X1 U9052 ( .C1(n7349), .C2(n9984), .A(n7348), .B(n7347), .ZN(P2_U3257) );
  NAND2_X1 U9053 ( .A1(n9934), .A2(n7404), .ZN(n9954) );
  NAND2_X1 U9054 ( .A1(n7351), .A2(n7350), .ZN(n7352) );
  XNOR2_X1 U9055 ( .A(n7353), .B(n7352), .ZN(n7354) );
  NAND2_X1 U9056 ( .A1(n7354), .A2(n8986), .ZN(n7360) );
  INV_X1 U9057 ( .A(n7355), .ZN(n7406) );
  OAI22_X1 U9058 ( .A1(n9013), .A2(n7406), .B1(n9042), .B2(n7356), .ZN(n7357)
         );
  AOI211_X1 U9059 ( .C1(n9040), .C2(n9357), .A(n7358), .B(n7357), .ZN(n7359)
         );
  OAI211_X1 U9060 ( .C1(n7361), .C2(n9954), .A(n7360), .B(n7359), .ZN(P1_U3211) );
  AOI21_X1 U9061 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(n7373) );
  AND2_X1 U9062 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7971) );
  NOR2_X1 U9063 ( .A1(n9983), .A2(n7365), .ZN(n7366) );
  AOI211_X1 U9064 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9981), .A(n7971), .B(
        n7366), .ZN(n7372) );
  OAI21_X1 U9065 ( .B1(n7369), .B2(n7368), .A(n7367), .ZN(n7370) );
  NAND2_X1 U9066 ( .A1(n7370), .A2(n9978), .ZN(n7371) );
  OAI211_X1 U9067 ( .C1(n7373), .C2(n9982), .A(n7372), .B(n7371), .ZN(P2_U3258) );
  INV_X1 U9068 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7383) );
  INV_X1 U9069 ( .A(n7374), .ZN(n7559) );
  XNOR2_X1 U9070 ( .A(n7559), .B(n7557), .ZN(n7414) );
  NAND2_X1 U9071 ( .A1(n7375), .A2(n8321), .ZN(n7376) );
  NAND2_X1 U9072 ( .A1(n7376), .A2(n10097), .ZN(n7377) );
  NOR2_X1 U9073 ( .A1(n7563), .A2(n7377), .ZN(n7411) );
  NAND2_X1 U9074 ( .A1(n7550), .A2(n7378), .ZN(n7379) );
  XOR2_X1 U9075 ( .A(n7557), .B(n7379), .Z(n7380) );
  AOI22_X1 U9076 ( .A1(n8447), .A2(n10017), .B1(n10015), .B2(n10018), .ZN(
        n8318) );
  OAI21_X1 U9077 ( .B1(n7380), .B2(n9995), .A(n8318), .ZN(n7417) );
  AOI211_X1 U9078 ( .C1(n10096), .C2(n8321), .A(n7411), .B(n7417), .ZN(n7381)
         );
  OAI21_X1 U9079 ( .B1(n10085), .B2(n7414), .A(n7381), .ZN(n7384) );
  NAND2_X1 U9080 ( .A1(n7384), .A2(n10142), .ZN(n7382) );
  OAI21_X1 U9081 ( .B1(n10142), .B2(n7383), .A(n7382), .ZN(P2_U3525) );
  INV_X1 U9082 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9083 ( .A1(n7384), .A2(n10121), .ZN(n7385) );
  OAI21_X1 U9084 ( .B1(n10121), .B2(n7386), .A(n7385), .ZN(P2_U3466) );
  NOR3_X2 U9085 ( .A1(n9679), .A2(n6889), .A3(n9281), .ZN(n9677) );
  INV_X1 U9086 ( .A(n9600), .ZN(n9675) );
  AOI22_X1 U9087 ( .A1(n9671), .A2(n7743), .B1(n9669), .B2(n7739), .ZN(n7387)
         );
  OAI21_X1 U9088 ( .B1(n7388), .B2(n9675), .A(n7387), .ZN(n7391) );
  MUX2_X1 U9089 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7389), .S(n7131), .Z(n7390)
         );
  AOI211_X1 U9090 ( .C1(n7392), .C2(n9677), .A(n7391), .B(n7390), .ZN(n7393)
         );
  INV_X1 U9091 ( .A(n7393), .ZN(P1_U3283) );
  INV_X1 U9092 ( .A(n7394), .ZN(n7395) );
  NAND2_X1 U9093 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  XNOR2_X1 U9094 ( .A(n7397), .B(n9185), .ZN(n9951) );
  OAI21_X1 U9095 ( .B1(n9185), .B2(n7399), .A(n7398), .ZN(n7400) );
  AOI222_X1 U9096 ( .A1(n9656), .A2(n7400), .B1(n9357), .B2(n9660), .C1(n9359), 
        .C2(n9659), .ZN(n9955) );
  MUX2_X1 U9097 ( .A(n6809), .B(n9955), .S(n7131), .Z(n7410) );
  INV_X1 U9098 ( .A(n7401), .ZN(n7403) );
  AOI211_X1 U9099 ( .C1(n7404), .C2(n7403), .A(n9944), .B(n7402), .ZN(n9952)
         );
  NOR2_X1 U9100 ( .A1(n7405), .A2(n9521), .ZN(n9642) );
  OAI22_X1 U9101 ( .A1(n9635), .A2(n7407), .B1(n7406), .B2(n9637), .ZN(n7408)
         );
  AOI21_X1 U9102 ( .B1(n9952), .B2(n9642), .A(n7408), .ZN(n7409) );
  OAI211_X1 U9103 ( .C1(n9951), .C2(n9645), .A(n7410), .B(n7409), .ZN(P1_U3284) );
  NAND2_X1 U9104 ( .A1(n8720), .A2(n7411), .ZN(n7413) );
  AOI22_X1 U9105 ( .A1(n8766), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8320), .B2(
        n10002), .ZN(n7412) );
  OAI211_X1 U9106 ( .C1(n7556), .C2(n10031), .A(n7413), .B(n7412), .ZN(n7416)
         );
  NOR2_X1 U9107 ( .A1(n7414), .A2(n8763), .ZN(n7415) );
  AOI211_X1 U9108 ( .C1(n10027), .C2(n7417), .A(n7416), .B(n7415), .ZN(n7418)
         );
  INV_X1 U9109 ( .A(n7418), .ZN(P2_U3291) );
  NAND2_X1 U9110 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  XNOR2_X1 U9111 ( .A(n7421), .B(n9085), .ZN(n7427) );
  INV_X1 U9112 ( .A(n9085), .ZN(n9184) );
  XNOR2_X1 U9113 ( .A(n4385), .B(n9184), .ZN(n7425) );
  OAI22_X1 U9114 ( .A1(n9631), .A2(n7423), .B1(n7741), .B2(n9633), .ZN(n7424)
         );
  AOI21_X1 U9115 ( .B1(n7425), .B2(n9656), .A(n7424), .ZN(n7426) );
  OAI21_X1 U9116 ( .B1(n7427), .B2(n9688), .A(n7426), .ZN(n9946) );
  INV_X1 U9117 ( .A(n9946), .ZN(n7434) );
  INV_X1 U9118 ( .A(n7427), .ZN(n9948) );
  AND2_X1 U9119 ( .A1(n7428), .A2(n9943), .ZN(n7429) );
  OR2_X1 U9120 ( .A1(n7429), .A2(n7401), .ZN(n9945) );
  AOI22_X1 U9121 ( .A1(n9679), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7576), .B2(
        n9669), .ZN(n7431) );
  NAND2_X1 U9122 ( .A1(n9671), .A2(n9943), .ZN(n7430) );
  OAI211_X1 U9123 ( .C1(n9675), .C2(n9945), .A(n7431), .B(n7430), .ZN(n7432)
         );
  AOI21_X1 U9124 ( .B1(n9948), .B2(n9677), .A(n7432), .ZN(n7433) );
  OAI21_X1 U9125 ( .B1(n7434), .B2(n9679), .A(n7433), .ZN(P1_U3285) );
  XOR2_X1 U9126 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7689), .Z(n7686) );
  OAI22_X1 U9127 ( .A1(n7436), .A2(n7435), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7439), .ZN(n7687) );
  XOR2_X1 U9128 ( .A(n7686), .B(n7687), .Z(n7445) );
  INV_X1 U9129 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9130 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7882) );
  OAI21_X1 U9131 ( .B1(n9923), .B2(n7437), .A(n7882), .ZN(n7443) );
  XNOR2_X1 U9132 ( .A(n7689), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7441) );
  OAI21_X1 U9133 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7439), .A(n7438), .ZN(
        n7440) );
  AOI211_X1 U9134 ( .C1(n7441), .C2(n7440), .A(n9893), .B(n7688), .ZN(n7442)
         );
  AOI211_X1 U9135 ( .C1(n9910), .C2(n7689), .A(n7443), .B(n7442), .ZN(n7444)
         );
  OAI21_X1 U9136 ( .B1(n9901), .B2(n7445), .A(n7444), .ZN(P1_U3253) );
  INV_X1 U9137 ( .A(n9677), .ZN(n7680) );
  AND2_X1 U9138 ( .A1(n9177), .A2(n6925), .ZN(n7446) );
  OR2_X1 U9139 ( .A1(n7447), .A2(n7446), .ZN(n9930) );
  OAI22_X1 U9140 ( .A1(n9635), .A2(n7457), .B1(n6810), .B2(n7131), .ZN(n7448)
         );
  INV_X1 U9141 ( .A(n7448), .ZN(n7460) );
  OAI21_X1 U9142 ( .B1(n7450), .B2(n9177), .A(n7449), .ZN(n7453) );
  OAI22_X1 U9143 ( .A1(n9631), .A2(n7451), .B1(n4388), .B2(n9633), .ZN(n7452)
         );
  AOI21_X1 U9144 ( .B1(n9656), .B2(n7453), .A(n7452), .ZN(n7454) );
  OAI21_X1 U9145 ( .B1(n9688), .B2(n9930), .A(n7454), .ZN(n9932) );
  OAI211_X1 U9146 ( .C1(n7457), .C2(n7456), .A(n9935), .B(n7455), .ZN(n9928)
         );
  OAI22_X1 U9147 ( .A1(n9928), .A2(n9521), .B1(n9637), .B2(n9875), .ZN(n7458)
         );
  OAI21_X1 U9148 ( .B1(n9932), .B2(n7458), .A(n7131), .ZN(n7459) );
  OAI211_X1 U9149 ( .C1(n7680), .C2(n9930), .A(n7460), .B(n7459), .ZN(P1_U3290) );
  XNOR2_X1 U9150 ( .A(n7571), .B(n7461), .ZN(n7462) );
  NAND2_X1 U9151 ( .A1(n7462), .A2(n7463), .ZN(n7569) );
  OAI21_X1 U9152 ( .B1(n7463), .B2(n7462), .A(n7569), .ZN(n7469) );
  AOI21_X1 U9153 ( .B1(n8951), .B2(n9361), .A(n7464), .ZN(n7467) );
  AOI22_X1 U9154 ( .A1(n9040), .A2(n9359), .B1(n9039), .B2(n7465), .ZN(n7466)
         );
  OAI211_X1 U9155 ( .C1(n9966), .C2(n8996), .A(n7467), .B(n7466), .ZN(n7468)
         );
  AOI21_X1 U9156 ( .B1(n7469), .B2(n8986), .A(n7468), .ZN(n7470) );
  INV_X1 U9157 ( .A(n7470), .ZN(P1_U3225) );
  MUX2_X1 U9158 ( .A(n6811), .B(n7471), .S(n7131), .Z(n7477) );
  OAI22_X1 U9159 ( .A1(n9635), .A2(n7473), .B1(n9637), .B2(n7472), .ZN(n7474)
         );
  AOI21_X1 U9160 ( .B1(n9600), .B2(n7475), .A(n7474), .ZN(n7476) );
  OAI211_X1 U9161 ( .C1(n7478), .C2(n7680), .A(n7477), .B(n7476), .ZN(P1_U3289) );
  XOR2_X1 U9162 ( .A(n7480), .B(n7479), .Z(n7488) );
  XNOR2_X1 U9163 ( .A(n7482), .B(n7481), .ZN(n7486) );
  INV_X1 U9164 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U9165 ( .A1(n8510), .A2(n7483), .ZN(n7484) );
  NAND2_X1 U9166 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U9167 ( .C1(n8522), .C2(n10392), .A(n7484), .B(n8215), .ZN(n7485)
         );
  AOI21_X1 U9168 ( .B1(n7486), .B2(n9979), .A(n7485), .ZN(n7487) );
  OAI21_X1 U9169 ( .B1(n9984), .B2(n7488), .A(n7487), .ZN(P2_U3259) );
  INV_X1 U9170 ( .A(n7489), .ZN(n7491) );
  OAI222_X1 U9171 ( .A1(n9837), .A2(n7490), .B1(n9840), .B2(n7491), .C1(
        P1_U3084), .C2(n9281), .ZN(P1_U3334) );
  OAI222_X1 U9172 ( .A1(n8093), .A2(n7492), .B1(n8906), .B2(n7491), .C1(
        P2_U3152), .C2(n8575), .ZN(P2_U3339) );
  AOI22_X1 U9173 ( .A1(n9679), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7493), .B2(
        n9669), .ZN(n7496) );
  NAND2_X1 U9174 ( .A1(n9600), .A2(n7494), .ZN(n7495) );
  OAI211_X1 U9175 ( .C1(n9635), .C2(n7497), .A(n7496), .B(n7495), .ZN(n7498)
         );
  AOI21_X1 U9176 ( .B1(n9677), .B2(n7499), .A(n7498), .ZN(n7500) );
  OAI21_X1 U9177 ( .B1(n9679), .B2(n7501), .A(n7500), .ZN(P1_U3287) );
  NAND2_X1 U9178 ( .A1(n7743), .A2(n9357), .ZN(n7502) );
  AND2_X1 U9179 ( .A1(n9795), .A2(n9356), .ZN(n7504) );
  OR2_X1 U9180 ( .A1(n9790), .A2(n7788), .ZN(n9094) );
  NAND2_X1 U9181 ( .A1(n9790), .A2(n7788), .ZN(n9093) );
  NAND2_X1 U9182 ( .A1(n9094), .A2(n9093), .ZN(n9176) );
  XNOR2_X1 U9183 ( .A(n7596), .B(n9176), .ZN(n9788) );
  INV_X1 U9184 ( .A(n9356), .ZN(n7659) );
  OAI22_X1 U9185 ( .A1(n9631), .A2(n7659), .B1(n7884), .B2(n9633), .ZN(n7510)
         );
  NAND2_X1 U9186 ( .A1(n7505), .A2(n9090), .ZN(n7506) );
  NAND2_X1 U9187 ( .A1(n9795), .A2(n7659), .ZN(n9092) );
  OR2_X1 U9188 ( .A1(n7841), .A2(n9176), .ZN(n7599) );
  NAND2_X1 U9189 ( .A1(n7841), .A2(n9176), .ZN(n7508) );
  AOI21_X1 U9190 ( .B1(n7599), .B2(n7508), .A(n9628), .ZN(n7509) );
  AOI211_X1 U9191 ( .C1(n9665), .C2(n9788), .A(n7510), .B(n7509), .ZN(n9792)
         );
  INV_X1 U9192 ( .A(n9790), .ZN(n7665) );
  INV_X1 U9193 ( .A(n7523), .ZN(n7511) );
  AND2_X2 U9194 ( .A1(n7523), .A2(n7665), .ZN(n7605) );
  AOI211_X1 U9195 ( .C1(n9790), .C2(n7511), .A(n9944), .B(n7605), .ZN(n9789)
         );
  NAND2_X1 U9196 ( .A1(n9789), .A2(n9642), .ZN(n7513) );
  AOI22_X1 U9197 ( .A1(n9679), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7658), .B2(
        n9669), .ZN(n7512) );
  OAI211_X1 U9198 ( .C1(n7665), .C2(n9635), .A(n7513), .B(n7512), .ZN(n7514)
         );
  AOI21_X1 U9199 ( .B1(n9788), .B2(n9677), .A(n7514), .ZN(n7515) );
  OAI21_X1 U9200 ( .B1(n9792), .B2(n9679), .A(n7515), .ZN(P1_U3281) );
  XNOR2_X1 U9201 ( .A(n7516), .B(n7507), .ZN(n9794) );
  OAI22_X1 U9202 ( .A1(n9631), .A2(n7517), .B1(n7788), .B2(n9633), .ZN(n7522)
         );
  INV_X1 U9203 ( .A(n7519), .ZN(n7520) );
  AOI211_X1 U9204 ( .C1(n9188), .C2(n7518), .A(n9628), .B(n7520), .ZN(n7521)
         );
  AOI211_X1 U9205 ( .C1(n9794), .C2(n9665), .A(n7522), .B(n7521), .ZN(n9798)
         );
  INV_X1 U9206 ( .A(n9795), .ZN(n7526) );
  AOI21_X1 U9207 ( .B1(n9795), .B2(n5060), .A(n7523), .ZN(n9796) );
  NAND2_X1 U9208 ( .A1(n9796), .A2(n9600), .ZN(n7525) );
  AOI22_X1 U9209 ( .A1(n9679), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7721), .B2(
        n9669), .ZN(n7524) );
  OAI211_X1 U9210 ( .C1(n7526), .C2(n9635), .A(n7525), .B(n7524), .ZN(n7527)
         );
  AOI21_X1 U9211 ( .B1(n9794), .B2(n9677), .A(n7527), .ZN(n7528) );
  OAI21_X1 U9212 ( .B1(n9798), .B2(n9679), .A(n7528), .ZN(P1_U3282) );
  OAI21_X1 U9213 ( .B1(n4483), .B2(n7530), .A(n7529), .ZN(n10056) );
  XNOR2_X1 U9214 ( .A(n7532), .B(n7531), .ZN(n7533) );
  AOI22_X1 U9215 ( .A1(n10015), .A2(n5682), .B1(n8450), .B2(n10017), .ZN(n8120) );
  OAI21_X1 U9216 ( .B1(n7533), .B2(n9995), .A(n8120), .ZN(n10060) );
  MUX2_X1 U9217 ( .A(n10060), .B(P2_REG2_REG_2__SCAN_IN), .S(n10036), .Z(n7539) );
  NAND2_X1 U9218 ( .A1(n7534), .A2(n7590), .ZN(n7535) );
  NAND2_X1 U9219 ( .A1(n7535), .A2(n10097), .ZN(n7536) );
  NOR2_X1 U9220 ( .A1(n10023), .A2(n7536), .ZN(n10059) );
  AOI22_X1 U9221 ( .A1(n8720), .A2(n10059), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n10002), .ZN(n7537) );
  OAI21_X1 U9222 ( .B1(n10031), .B2(n10057), .A(n7537), .ZN(n7538) );
  AOI211_X1 U9223 ( .C1(n10034), .C2(n10056), .A(n7539), .B(n7538), .ZN(n7540)
         );
  INV_X1 U9224 ( .A(n7540), .ZN(P2_U3294) );
  NAND2_X1 U9225 ( .A1(n7585), .A2(n7541), .ZN(n10049) );
  NAND2_X1 U9226 ( .A1(n10049), .A2(n10020), .ZN(n7543) );
  NAND2_X1 U9227 ( .A1(n7543), .A2(n7542), .ZN(n10047) );
  AOI21_X1 U9228 ( .B1(n10002), .B2(P2_REG3_REG_0__SCAN_IN), .A(n10047), .ZN(
        n7545) );
  NAND2_X1 U9229 ( .A1(n10036), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7544) );
  OAI21_X1 U9230 ( .B1(n10036), .B2(n7545), .A(n7544), .ZN(n7547) );
  OR2_X1 U9231 ( .A1(n8551), .A2(n10113), .ZN(n8166) );
  AOI21_X1 U9232 ( .B1(n10031), .B2(n8166), .A(n10046), .ZN(n7546) );
  AOI211_X1 U9233 ( .C1(n10034), .C2(n10049), .A(n7547), .B(n7546), .ZN(n7548)
         );
  INV_X1 U9234 ( .A(n7548), .ZN(P2_U3296) );
  INV_X1 U9235 ( .A(n8448), .ZN(n7555) );
  NAND2_X1 U9236 ( .A1(n7550), .A2(n7549), .ZN(n7552) );
  NAND2_X1 U9237 ( .A1(n7552), .A2(n7551), .ZN(n7553) );
  XOR2_X1 U9238 ( .A(n7561), .B(n7553), .Z(n7554) );
  OAI222_X1 U9239 ( .A1(n10000), .A2(n8391), .B1(n9998), .B2(n7555), .C1(n9995), .C2(n7554), .ZN(n10076) );
  AOI21_X1 U9240 ( .B1(n8395), .B2(n10002), .A(n10076), .ZN(n7568) );
  AOI21_X1 U9241 ( .B1(n7374), .B2(n7557), .A(n7556), .ZN(n7558) );
  AOI21_X1 U9242 ( .B1(n7559), .B2(n8448), .A(n7558), .ZN(n7560) );
  XOR2_X1 U9243 ( .A(n7561), .B(n7560), .Z(n10078) );
  NOR2_X1 U9244 ( .A1(n10031), .A2(n10074), .ZN(n7566) );
  OAI21_X1 U9245 ( .B1(n10074), .B2(n7563), .A(n7562), .ZN(n10075) );
  OAI22_X1 U9246 ( .A1(n10027), .A2(n7564), .B1(n8166), .B2(n10075), .ZN(n7565) );
  AOI211_X1 U9247 ( .C1(n10078), .C2(n10034), .A(n7566), .B(n7565), .ZN(n7567)
         );
  OAI21_X1 U9248 ( .B1(n10036), .B2(n7568), .A(n7567), .ZN(P2_U3290) );
  OAI21_X1 U9249 ( .B1(n7571), .B2(n7570), .A(n7569), .ZN(n7575) );
  XNOR2_X1 U9250 ( .A(n7573), .B(n7572), .ZN(n7574) );
  XNOR2_X1 U9251 ( .A(n7575), .B(n7574), .ZN(n7581) );
  AOI22_X1 U9252 ( .A1(n8951), .A2(n9360), .B1(n7576), .B2(n9039), .ZN(n7580)
         );
  OAI21_X1 U9253 ( .B1(n9011), .B2(n7741), .A(n7577), .ZN(n7578) );
  AOI21_X1 U9254 ( .B1(n9045), .B2(n9943), .A(n7578), .ZN(n7579) );
  OAI211_X1 U9255 ( .C1(n7581), .C2(n9047), .A(n7580), .B(n7579), .ZN(P1_U3237) );
  OAI21_X1 U9256 ( .B1(n5976), .B2(n7583), .A(n7582), .ZN(n7584) );
  INV_X1 U9257 ( .A(n7584), .ZN(n10054) );
  AOI22_X1 U9258 ( .A1(n10054), .A2(n10034), .B1(n8756), .B2(n5123), .ZN(n7594) );
  INV_X1 U9259 ( .A(n5976), .ZN(n7586) );
  OAI21_X1 U9260 ( .B1(n7586), .B2(n7585), .A(n10020), .ZN(n7589) );
  AOI22_X1 U9261 ( .A1(n10015), .A2(n8451), .B1(n10016), .B2(n10017), .ZN(
        n7587) );
  OAI21_X1 U9262 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n10052) );
  OAI211_X1 U9263 ( .C1(n10046), .C2(n10051), .A(n10097), .B(n7590), .ZN(
        n10050) );
  INV_X1 U9264 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7591) );
  OAI22_X1 U9265 ( .A1(n8551), .A2(n10050), .B1(n7591), .B2(n10026), .ZN(n7592) );
  AOI21_X1 U9266 ( .B1(n10027), .B2(n10052), .A(n7592), .ZN(n7593) );
  OAI211_X1 U9267 ( .C1(n7595), .C2(n10027), .A(n7594), .B(n7593), .ZN(
        P2_U3295) );
  INV_X1 U9268 ( .A(n7788), .ZN(n9355) );
  OR2_X1 U9269 ( .A1(n9790), .A2(n9355), .ZN(n7597) );
  OR2_X1 U9270 ( .A1(n7792), .A2(n7884), .ZN(n7842) );
  NAND2_X1 U9271 ( .A1(n7792), .A2(n7884), .ZN(n9100) );
  INV_X1 U9272 ( .A(n9192), .ZN(n7598) );
  XNOR2_X1 U9273 ( .A(n7771), .B(n7598), .ZN(n9782) );
  NAND2_X1 U9274 ( .A1(n9782), .A2(n9665), .ZN(n7604) );
  NAND2_X1 U9275 ( .A1(n7599), .A2(n9093), .ZN(n7773) );
  XNOR2_X1 U9276 ( .A(n7773), .B(n9192), .ZN(n7602) );
  NAND2_X1 U9277 ( .A1(n9659), .A2(n9355), .ZN(n7600) );
  OAI21_X1 U9278 ( .B1(n7818), .B2(n9633), .A(n7600), .ZN(n7601) );
  AOI21_X1 U9279 ( .B1(n7602), .B2(n9656), .A(n7601), .ZN(n7603) );
  NAND2_X1 U9280 ( .A1(n7604), .A2(n7603), .ZN(n9787) );
  INV_X1 U9281 ( .A(n9787), .ZN(n7611) );
  INV_X1 U9282 ( .A(n7792), .ZN(n9783) );
  OR2_X1 U9283 ( .A1(n7605), .A2(n9783), .ZN(n7606) );
  NAND2_X1 U9284 ( .A1(n7776), .A2(n7606), .ZN(n9784) );
  AOI22_X1 U9285 ( .A1(n9679), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7787), .B2(
        n9669), .ZN(n7608) );
  NAND2_X1 U9286 ( .A1(n9671), .A2(n7792), .ZN(n7607) );
  OAI211_X1 U9287 ( .C1(n9784), .C2(n9675), .A(n7608), .B(n7607), .ZN(n7609)
         );
  AOI21_X1 U9288 ( .B1(n9782), .B2(n9677), .A(n7609), .ZN(n7610) );
  OAI21_X1 U9289 ( .B1(n7611), .B2(n9679), .A(n7610), .ZN(P1_U3280) );
  NOR2_X1 U9290 ( .A1(n7612), .A2(n7619), .ZN(n7632) );
  AND2_X1 U9291 ( .A1(n7612), .A2(n7619), .ZN(n7613) );
  OR2_X1 U9292 ( .A1(n7632), .A2(n7613), .ZN(n10091) );
  OR2_X1 U9293 ( .A1(n10036), .A2(n7614), .ZN(n10006) );
  OAI22_X1 U9294 ( .A1(n8391), .A2(n9998), .B1(n9997), .B2(n10000), .ZN(n7615)
         );
  INV_X1 U9295 ( .A(n7615), .ZN(n7622) );
  AND2_X1 U9296 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  OAI21_X1 U9297 ( .B1(n7619), .B2(n7618), .A(n7638), .ZN(n7620) );
  NAND2_X1 U9298 ( .A1(n7620), .A2(n10020), .ZN(n7621) );
  OAI211_X1 U9299 ( .C1(n10091), .C2(n8736), .A(n7622), .B(n7621), .ZN(n10093)
         );
  MUX2_X1 U9300 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10093), .S(n10027), .Z(n7623) );
  INV_X1 U9301 ( .A(n7623), .ZN(n7630) );
  NAND2_X1 U9302 ( .A1(n7301), .A2(n10088), .ZN(n7625) );
  AND2_X1 U9303 ( .A1(n7642), .A2(n7625), .ZN(n10089) );
  INV_X1 U9304 ( .A(n10088), .ZN(n7627) );
  OAI22_X1 U9305 ( .A1(n10031), .A2(n7627), .B1(n10026), .B2(n7626), .ZN(n7628) );
  AOI21_X1 U9306 ( .B1(n10029), .B2(n10089), .A(n7628), .ZN(n7629) );
  OAI211_X1 U9307 ( .C1(n10091), .C2(n10006), .A(n7630), .B(n7629), .ZN(
        P2_U3288) );
  NOR2_X1 U9308 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  XNOR2_X1 U9309 ( .A(n7633), .B(n7637), .ZN(n7644) );
  INV_X1 U9310 ( .A(n8736), .ZN(n10001) );
  OAI22_X1 U9311 ( .A1(n7830), .A2(n10000), .B1(n7634), .B2(n9998), .ZN(n7641)
         );
  NAND3_X1 U9312 ( .A1(n7638), .A2(n7637), .A3(n7636), .ZN(n7639) );
  AOI21_X1 U9313 ( .B1(n7635), .B2(n7639), .A(n9995), .ZN(n7640) );
  AOI211_X1 U9314 ( .C1(n7644), .C2(n10001), .A(n7641), .B(n7640), .ZN(n10100)
         );
  AOI21_X1 U9315 ( .B1(n10095), .B2(n7642), .A(n4471), .ZN(n10098) );
  AOI22_X1 U9316 ( .A1(n8766), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7829), .B2(
        n10002), .ZN(n7643) );
  OAI21_X1 U9317 ( .B1(n10031), .B2(n5720), .A(n7643), .ZN(n7646) );
  INV_X1 U9318 ( .A(n7644), .ZN(n10101) );
  NOR2_X1 U9319 ( .A1(n10101), .A2(n10006), .ZN(n7645) );
  AOI211_X1 U9320 ( .C1(n10029), .C2(n10098), .A(n7646), .B(n7645), .ZN(n7647)
         );
  OAI21_X1 U9321 ( .B1(n10036), .B2(n10100), .A(n7647), .ZN(P2_U3287) );
  INV_X1 U9322 ( .A(n7648), .ZN(n7652) );
  OAI222_X1 U9323 ( .A1(n8093), .A2(n7650), .B1(n8906), .B2(n7652), .C1(n4376), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U9324 ( .A1(P1_U3084), .A2(n4378), .B1(n9840), .B2(n7652), .C1(
        n7651), .C2(n9837), .ZN(P1_U3333) );
  XNOR2_X1 U9325 ( .A(n7654), .B(n7653), .ZN(n7655) );
  XNOR2_X1 U9326 ( .A(n7656), .B(n7655), .ZN(n7657) );
  NAND2_X1 U9327 ( .A1(n7657), .A2(n8986), .ZN(n7664) );
  INV_X1 U9328 ( .A(n7658), .ZN(n7660) );
  OAI22_X1 U9329 ( .A1(n9013), .A2(n7660), .B1(n9042), .B2(n7659), .ZN(n7661)
         );
  AOI211_X1 U9330 ( .C1(n9040), .C2(n9354), .A(n7662), .B(n7661), .ZN(n7663)
         );
  OAI211_X1 U9331 ( .C1(n7665), .C2(n8996), .A(n7664), .B(n7663), .ZN(P1_U3215) );
  OAI21_X1 U9332 ( .B1(n9179), .B2(n9270), .A(n7132), .ZN(n7674) );
  OAI22_X1 U9333 ( .A1(n9631), .A2(n4388), .B1(n7667), .B2(n9633), .ZN(n7673)
         );
  INV_X1 U9334 ( .A(n7670), .ZN(n7671) );
  AOI21_X1 U9335 ( .B1(n9179), .B2(n7669), .A(n7671), .ZN(n9940) );
  NOR2_X1 U9336 ( .A1(n9940), .A2(n9688), .ZN(n7672) );
  AOI211_X1 U9337 ( .C1(n9656), .C2(n7674), .A(n7673), .B(n7672), .ZN(n9938)
         );
  INV_X1 U9338 ( .A(n7675), .ZN(n7678) );
  INV_X1 U9339 ( .A(n7676), .ZN(n7677) );
  AOI21_X1 U9340 ( .B1(n7679), .B2(n7678), .A(n7677), .ZN(n9936) );
  OAI22_X1 U9341 ( .A1(n7131), .A2(n6814), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9637), .ZN(n7682) );
  OAI22_X1 U9342 ( .A1(n7680), .A2(n9940), .B1(n6935), .B2(n9635), .ZN(n7681)
         );
  AOI211_X1 U9343 ( .C1(n9600), .C2(n9936), .A(n7682), .B(n7681), .ZN(n7683)
         );
  OAI21_X1 U9344 ( .B1(n9679), .B2(n9938), .A(n7683), .ZN(P1_U3288) );
  XNOR2_X1 U9345 ( .A(n9375), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9367) );
  INV_X1 U9346 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7684) );
  AOI22_X1 U9347 ( .A1(n7687), .A2(n7686), .B1(n7685), .B2(n7684), .ZN(n9368)
         );
  XOR2_X1 U9348 ( .A(n9367), .B(n9368), .Z(n7695) );
  NAND2_X1 U9349 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7816) );
  OAI21_X1 U9350 ( .B1(n9923), .B2(n4520), .A(n7816), .ZN(n7693) );
  XNOR2_X1 U9351 ( .A(n9375), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7690) );
  AOI211_X1 U9352 ( .C1(n7691), .C2(n7690), .A(n9893), .B(n9374), .ZN(n7692)
         );
  AOI211_X1 U9353 ( .C1(n9910), .C2(n9375), .A(n7693), .B(n7692), .ZN(n7694)
         );
  OAI21_X1 U9354 ( .B1(n9901), .B2(n7695), .A(n7694), .ZN(P1_U3254) );
  XNOR2_X1 U9355 ( .A(n7696), .B(n4379), .ZN(n7697) );
  NOR2_X1 U9356 ( .A1(n7830), .A2(n8251), .ZN(n7698) );
  NAND2_X1 U9357 ( .A1(n7697), .A2(n7698), .ZN(n7803) );
  INV_X1 U9358 ( .A(n7697), .ZN(n7802) );
  INV_X1 U9359 ( .A(n7698), .ZN(n7699) );
  NAND2_X1 U9360 ( .A1(n7802), .A2(n7699), .ZN(n7700) );
  AND2_X1 U9361 ( .A1(n7803), .A2(n7700), .ZN(n7710) );
  INV_X1 U9362 ( .A(n7701), .ZN(n7703) );
  NAND2_X1 U9363 ( .A1(n7703), .A2(n7702), .ZN(n7704) );
  XNOR2_X1 U9364 ( .A(n10095), .B(n7176), .ZN(n7826) );
  OR2_X1 U9365 ( .A1(n9997), .A2(n8251), .ZN(n7707) );
  NAND2_X1 U9366 ( .A1(n7826), .A2(n7707), .ZN(n7706) );
  INV_X1 U9367 ( .A(n7826), .ZN(n7709) );
  INV_X1 U9368 ( .A(n7707), .ZN(n7708) );
  NAND2_X1 U9369 ( .A1(n7709), .A2(n7708), .ZN(n7822) );
  OAI211_X1 U9370 ( .C1(n7710), .C2(n7827), .A(n7804), .B(n8398), .ZN(n7714)
         );
  NAND2_X1 U9371 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8492) );
  INV_X1 U9372 ( .A(n8492), .ZN(n7712) );
  OAI22_X1 U9373 ( .A1(n9997), .A2(n8383), .B1(n8392), .B2(n9999), .ZN(n7711)
         );
  AOI211_X1 U9374 ( .C1(n10003), .C2(n8420), .A(n7712), .B(n7711), .ZN(n7713)
         );
  OAI211_X1 U9375 ( .C1(n10105), .C2(n8425), .A(n7714), .B(n7713), .ZN(
        P2_U3219) );
  OR2_X1 U9376 ( .A1(n7717), .A2(n7716), .ZN(n7737) );
  NAND2_X1 U9377 ( .A1(n7737), .A2(n7715), .ZN(n7732) );
  NAND2_X1 U9378 ( .A1(n7717), .A2(n7716), .ZN(n7734) );
  NAND2_X1 U9379 ( .A1(n7732), .A2(n7734), .ZN(n7731) );
  XNOR2_X1 U9380 ( .A(n7719), .B(n7718), .ZN(n7720) );
  XNOR2_X1 U9381 ( .A(n7731), .B(n7720), .ZN(n7727) );
  AOI22_X1 U9382 ( .A1(n8951), .A2(n9357), .B1(n7721), .B2(n9039), .ZN(n7723)
         );
  NAND2_X1 U9383 ( .A1(n9040), .A2(n9355), .ZN(n7722) );
  OAI211_X1 U9384 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7724), .A(n7723), .B(n7722), .ZN(n7725) );
  AOI21_X1 U9385 ( .B1(n9045), .B2(n9795), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9386 ( .B1(n7727), .B2(n9047), .A(n7726), .ZN(P1_U3229) );
  INV_X1 U9387 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7730) );
  INV_X1 U9388 ( .A(n7728), .ZN(n7783) );
  OAI222_X1 U9389 ( .A1(n8093), .A2(n7730), .B1(n8906), .B2(n7783), .C1(n7729), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U9390 ( .A(n7731), .ZN(n7738) );
  INV_X1 U9391 ( .A(n7732), .ZN(n7735) );
  AOI21_X1 U9392 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7736) );
  AOI21_X1 U9393 ( .B1(n7738), .B2(n7737), .A(n7736), .ZN(n7745) );
  AOI22_X1 U9394 ( .A1(n9040), .A2(n9356), .B1(n9039), .B2(n7739), .ZN(n7740)
         );
  NAND2_X1 U9395 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9890) );
  OAI211_X1 U9396 ( .C1(n7741), .C2(n9042), .A(n7740), .B(n9890), .ZN(n7742)
         );
  AOI21_X1 U9397 ( .B1(n9045), .B2(n7743), .A(n7742), .ZN(n7744) );
  OAI21_X1 U9398 ( .B1(n7745), .B2(n9047), .A(n7744), .ZN(P1_U3219) );
  XOR2_X1 U9399 ( .A(n7749), .B(n7746), .Z(n7747) );
  OAI222_X1 U9400 ( .A1(n10000), .A2(n7969), .B1(n9998), .B2(n7830), .C1(n9995), .C2(n7747), .ZN(n10115) );
  INV_X1 U9401 ( .A(n10115), .ZN(n7756) );
  OAI21_X1 U9402 ( .B1(n7750), .B2(n7749), .A(n7748), .ZN(n7751) );
  INV_X1 U9403 ( .A(n7751), .ZN(n10118) );
  OAI21_X1 U9404 ( .B1(n10007), .B2(n10112), .A(n7866), .ZN(n10114) );
  AOI22_X1 U9405 ( .A1(n10036), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7810), .B2(
        n10002), .ZN(n7753) );
  NAND2_X1 U9406 ( .A1(n8756), .A2(n7796), .ZN(n7752) );
  OAI211_X1 U9407 ( .C1(n10114), .C2(n8166), .A(n7753), .B(n7752), .ZN(n7754)
         );
  AOI21_X1 U9408 ( .B1(n10118), .B2(n10034), .A(n7754), .ZN(n7755) );
  OAI21_X1 U9409 ( .B1(n7756), .B2(n8766), .A(n7755), .ZN(P2_U3285) );
  OAI21_X1 U9410 ( .B1(n7759), .B2(n7758), .A(n7757), .ZN(n7760) );
  NAND2_X1 U9411 ( .A1(n7760), .A2(n9979), .ZN(n7769) );
  INV_X1 U9412 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U9413 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7761) );
  OAI21_X1 U9414 ( .B1(n8522), .B2(n7762), .A(n7761), .ZN(n7766) );
  AOI211_X1 U9415 ( .C1(n10352), .C2(n7764), .A(n9984), .B(n7763), .ZN(n7765)
         );
  AOI211_X1 U9416 ( .C1(n8510), .C2(n7767), .A(n7766), .B(n7765), .ZN(n7768)
         );
  NAND2_X1 U9417 ( .A1(n7769), .A2(n7768), .ZN(P2_U3260) );
  NAND2_X1 U9418 ( .A1(n7792), .A2(n9354), .ZN(n7770) );
  OR2_X1 U9419 ( .A1(n9779), .A2(n7818), .ZN(n9101) );
  NAND2_X1 U9420 ( .A1(n9779), .A2(n7818), .ZN(n9105) );
  NAND2_X1 U9421 ( .A1(n9101), .A2(n9105), .ZN(n9194) );
  XNOR2_X1 U9422 ( .A(n7838), .B(n9194), .ZN(n9781) );
  INV_X1 U9423 ( .A(n9352), .ZN(n7920) );
  INV_X1 U9424 ( .A(n9100), .ZN(n7772) );
  OAI21_X1 U9425 ( .B1(n7773), .B2(n7772), .A(n7842), .ZN(n7774) );
  INV_X1 U9426 ( .A(n9194), .ZN(n9099) );
  XNOR2_X1 U9427 ( .A(n7774), .B(n9099), .ZN(n7775) );
  OAI222_X1 U9428 ( .A1(n9633), .A2(n7920), .B1(n9631), .B2(n7884), .C1(n9628), 
        .C2(n7775), .ZN(n9777) );
  NAND2_X1 U9429 ( .A1(n9777), .A2(n7131), .ZN(n7782) );
  AOI21_X1 U9430 ( .B1(n7776), .B2(n9779), .A(n9944), .ZN(n7777) );
  AND2_X1 U9431 ( .A1(n7777), .A2(n7850), .ZN(n9778) );
  NAND2_X1 U9432 ( .A1(n9779), .A2(n9671), .ZN(n7779) );
  AOI22_X1 U9433 ( .A1(n9679), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7881), .B2(
        n9669), .ZN(n7778) );
  NAND2_X1 U9434 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  AOI21_X1 U9435 ( .B1(n9778), .B2(n9642), .A(n7780), .ZN(n7781) );
  OAI211_X1 U9436 ( .C1(n9645), .C2(n9781), .A(n7782), .B(n7781), .ZN(P1_U3279) );
  INV_X1 U9437 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7784) );
  OAI222_X1 U9438 ( .A1(n9837), .A2(n7784), .B1(P1_U3084), .B2(n9210), .C1(
        n9840), .C2(n7783), .ZN(P1_U3332) );
  NAND2_X1 U9439 ( .A1(n7786), .A2(n7785), .ZN(n7876) );
  XNOR2_X1 U9440 ( .A(n7876), .B(n7875), .ZN(n7795) );
  INV_X1 U9441 ( .A(n7818), .ZN(n9353) );
  INV_X1 U9442 ( .A(n7787), .ZN(n7789) );
  OAI22_X1 U9443 ( .A1(n9013), .A2(n7789), .B1(n9042), .B2(n7788), .ZN(n7790)
         );
  AOI211_X1 U9444 ( .C1(n9040), .C2(n9353), .A(n7791), .B(n7790), .ZN(n7794)
         );
  NAND2_X1 U9445 ( .A1(n9045), .A2(n7792), .ZN(n7793) );
  OAI211_X1 U9446 ( .C1(n7795), .C2(n9047), .A(n7794), .B(n7793), .ZN(P1_U3234) );
  XNOR2_X1 U9447 ( .A(n7796), .B(n4379), .ZN(n7797) );
  NOR2_X1 U9448 ( .A1(n9999), .A2(n8251), .ZN(n7798) );
  NAND2_X1 U9449 ( .A1(n7797), .A2(n7798), .ZN(n7900) );
  INV_X1 U9450 ( .A(n7797), .ZN(n7899) );
  INV_X1 U9451 ( .A(n7798), .ZN(n7799) );
  NAND2_X1 U9452 ( .A1(n7899), .A2(n7799), .ZN(n7800) );
  AND2_X1 U9453 ( .A1(n7900), .A2(n7800), .ZN(n7805) );
  INV_X1 U9454 ( .A(n7805), .ZN(n7801) );
  AOI21_X1 U9455 ( .B1(n7804), .B2(n7801), .A(n8426), .ZN(n7807) );
  NOR3_X1 U9456 ( .A1(n8402), .A2(n7802), .A3(n7830), .ZN(n7806) );
  OAI21_X1 U9457 ( .B1(n7807), .B2(n7806), .A(n7901), .ZN(n7812) );
  NOR2_X1 U9458 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7284), .ZN(n7809) );
  OAI22_X1 U9459 ( .A1(n7830), .A2(n8383), .B1(n8392), .B2(n7969), .ZN(n7808)
         );
  AOI211_X1 U9460 ( .C1(n8420), .C2(n7810), .A(n7809), .B(n7808), .ZN(n7811)
         );
  OAI211_X1 U9461 ( .C1(n10112), .C2(n8425), .A(n7812), .B(n7811), .ZN(
        P2_U3238) );
  XOR2_X1 U9462 ( .A(n7814), .B(n7813), .Z(n7815) );
  XNOR2_X1 U9463 ( .A(n4475), .B(n7815), .ZN(n7821) );
  AOI22_X1 U9464 ( .A1(n9040), .A2(n9658), .B1(n9039), .B2(n7852), .ZN(n7817)
         );
  OAI211_X1 U9465 ( .C1(n7818), .C2(n9042), .A(n7817), .B(n7816), .ZN(n7819)
         );
  AOI21_X1 U9466 ( .B1(n7949), .B2(n9045), .A(n7819), .ZN(n7820) );
  OAI21_X1 U9467 ( .B1(n7821), .B2(n9047), .A(n7820), .ZN(P1_U3232) );
  OAI21_X1 U9468 ( .B1(n7824), .B2(n4862), .A(n7823), .ZN(n7825) );
  OAI21_X1 U9469 ( .B1(n7827), .B2(n7826), .A(n7825), .ZN(n7836) );
  OR3_X1 U9470 ( .A1(n7827), .A2(n9997), .A3(n8402), .ZN(n7834) );
  NOR2_X1 U9471 ( .A1(n7828), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8478) );
  AOI21_X1 U9472 ( .B1(n8420), .B2(n7829), .A(n8478), .ZN(n7833) );
  INV_X1 U9473 ( .A(n7830), .ZN(n8443) );
  AOI22_X1 U9474 ( .A1(n8421), .A2(n8443), .B1(n8422), .B2(n8445), .ZN(n7832)
         );
  NAND2_X1 U9475 ( .A1(n8386), .A2(n10095), .ZN(n7831) );
  NAND4_X1 U9476 ( .A1(n7834), .A2(n7833), .A3(n7832), .A4(n7831), .ZN(n7835)
         );
  AOI21_X1 U9477 ( .B1(n8398), .B2(n7836), .A(n7835), .ZN(n7837) );
  INV_X1 U9478 ( .A(n7837), .ZN(P2_U3233) );
  NAND2_X1 U9479 ( .A1(n7838), .A2(n9194), .ZN(n7840) );
  NAND2_X1 U9480 ( .A1(n9779), .A2(n9353), .ZN(n7839) );
  OR2_X1 U9481 ( .A1(n7949), .A2(n7920), .ZN(n9106) );
  NAND2_X1 U9482 ( .A1(n7949), .A2(n7920), .ZN(n9111) );
  XNOR2_X1 U9483 ( .A(n7937), .B(n9196), .ZN(n7952) );
  NAND3_X1 U9484 ( .A1(n7841), .A2(n9100), .A3(n9093), .ZN(n7846) );
  AND2_X1 U9485 ( .A1(n9101), .A2(n7842), .ZN(n9108) );
  INV_X1 U9486 ( .A(n9094), .ZN(n7843) );
  NAND2_X1 U9487 ( .A1(n9100), .A2(n7843), .ZN(n7844) );
  XNOR2_X1 U9488 ( .A(n7938), .B(n4671), .ZN(n7848) );
  AOI22_X1 U9489 ( .A1(n9660), .A2(n9658), .B1(n9659), .B2(n9353), .ZN(n7847)
         );
  OAI21_X1 U9490 ( .B1(n7848), .B2(n9628), .A(n7847), .ZN(n7849) );
  AOI21_X1 U9491 ( .B1(n7952), .B2(n9665), .A(n7849), .ZN(n7954) );
  AND2_X1 U9492 ( .A1(n7850), .A2(n7949), .ZN(n7851) );
  OR2_X1 U9493 ( .A1(n7851), .A2(n7941), .ZN(n7950) );
  AOI22_X1 U9494 ( .A1(n9679), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7852), .B2(
        n9669), .ZN(n7854) );
  NAND2_X1 U9495 ( .A1(n7949), .A2(n9671), .ZN(n7853) );
  OAI211_X1 U9496 ( .C1(n7950), .C2(n9675), .A(n7854), .B(n7853), .ZN(n7855)
         );
  AOI21_X1 U9497 ( .B1(n7952), .B2(n9677), .A(n7855), .ZN(n7856) );
  OAI21_X1 U9498 ( .B1(n7954), .B2(n9679), .A(n7856), .ZN(P1_U3278) );
  XNOR2_X1 U9499 ( .A(n7857), .B(n7864), .ZN(n7858) );
  NAND2_X1 U9500 ( .A1(n7858), .A2(n10020), .ZN(n7861) );
  OAI22_X1 U9501 ( .A1(n9999), .A2(n9998), .B1(n8208), .B2(n10000), .ZN(n7859)
         );
  INV_X1 U9502 ( .A(n7859), .ZN(n7860) );
  NAND2_X1 U9503 ( .A1(n7861), .A2(n7860), .ZN(n8868) );
  INV_X1 U9504 ( .A(n8868), .ZN(n7872) );
  NAND2_X1 U9505 ( .A1(n7863), .A2(n7864), .ZN(n7865) );
  NAND2_X1 U9506 ( .A1(n7862), .A2(n7865), .ZN(n8863) );
  NAND2_X1 U9507 ( .A1(n7866), .A2(n7893), .ZN(n7867) );
  NAND2_X1 U9508 ( .A1(n5042), .A2(n7867), .ZN(n8865) );
  NOR2_X1 U9509 ( .A1(n8865), .A2(n8166), .ZN(n7870) );
  AOI22_X1 U9510 ( .A1(n8766), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7908), .B2(
        n10002), .ZN(n7868) );
  OAI21_X1 U9511 ( .B1(n10031), .B2(n8864), .A(n7868), .ZN(n7869) );
  AOI211_X1 U9512 ( .C1(n8863), .C2(n10034), .A(n7870), .B(n7869), .ZN(n7871)
         );
  OAI21_X1 U9513 ( .B1(n7872), .B2(n8766), .A(n7871), .ZN(P2_U3284) );
  NAND2_X1 U9514 ( .A1(n7874), .A2(n7873), .ZN(n7880) );
  NAND2_X1 U9515 ( .A1(n7876), .A2(n7875), .ZN(n7878) );
  NAND2_X1 U9516 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  XOR2_X1 U9517 ( .A(n7880), .B(n7879), .Z(n7887) );
  AOI22_X1 U9518 ( .A1(n9040), .A2(n9352), .B1(n9039), .B2(n7881), .ZN(n7883)
         );
  OAI211_X1 U9519 ( .C1(n7884), .C2(n9042), .A(n7883), .B(n7882), .ZN(n7885)
         );
  AOI21_X1 U9520 ( .B1(n9045), .B2(n9779), .A(n7885), .ZN(n7886) );
  OAI21_X1 U9521 ( .B1(n7887), .B2(n9047), .A(n7886), .ZN(P1_U3222) );
  INV_X1 U9522 ( .A(n7888), .ZN(n8091) );
  OAI222_X1 U9523 ( .A1(n9837), .A2(n7889), .B1(n9840), .B2(n8091), .C1(
        P1_U3084), .C2(n9328), .ZN(P1_U3331) );
  INV_X1 U9524 ( .A(n6523), .ZN(n7892) );
  NAND2_X1 U9525 ( .A1(n7890), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9212) );
  INV_X1 U9526 ( .A(n9212), .ZN(n9339) );
  AOI21_X1 U9527 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9828), .A(n9339), .ZN(
        n7891) );
  OAI21_X1 U9528 ( .B1(n7892), .B2(n9840), .A(n7891), .ZN(P1_U3330) );
  XNOR2_X1 U9529 ( .A(n7893), .B(n4379), .ZN(n7894) );
  NOR2_X1 U9530 ( .A1(n7969), .A2(n8251), .ZN(n7895) );
  NAND2_X1 U9531 ( .A1(n7894), .A2(n7895), .ZN(n7963) );
  INV_X1 U9532 ( .A(n7894), .ZN(n7962) );
  INV_X1 U9533 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9534 ( .A1(n7962), .A2(n7896), .ZN(n7897) );
  AND2_X1 U9535 ( .A1(n7963), .A2(n7897), .ZN(n7902) );
  INV_X1 U9536 ( .A(n7902), .ZN(n7898) );
  AOI21_X1 U9537 ( .B1(n7901), .B2(n7898), .A(n8426), .ZN(n7905) );
  NOR3_X1 U9538 ( .A1(n7899), .A2(n9999), .A3(n8402), .ZN(n7904) );
  NAND2_X1 U9539 ( .A1(n7901), .A2(n7900), .ZN(n7903) );
  OAI21_X1 U9540 ( .B1(n7905), .B2(n7904), .A(n7964), .ZN(n7910) );
  OAI22_X1 U9541 ( .A1(n9999), .A2(n8383), .B1(n8392), .B2(n8208), .ZN(n7906)
         );
  AOI211_X1 U9542 ( .C1(n8420), .C2(n7908), .A(n7907), .B(n7906), .ZN(n7909)
         );
  OAI211_X1 U9543 ( .C1(n8864), .C2(n8425), .A(n7910), .B(n7909), .ZN(P2_U3226) );
  NAND2_X1 U9544 ( .A1(n6523), .A2(n7911), .ZN(n7913) );
  OAI211_X1 U9545 ( .C1(n10300), .C2(n8093), .A(n7913), .B(n7912), .ZN(
        P2_U3335) );
  XNOR2_X1 U9546 ( .A(n7916), .B(n7915), .ZN(n7917) );
  XNOR2_X1 U9547 ( .A(n7914), .B(n7917), .ZN(n7923) );
  INV_X1 U9548 ( .A(n7918), .ZN(n7943) );
  AOI22_X1 U9549 ( .A1(n9040), .A2(n9351), .B1(n9039), .B2(n7943), .ZN(n7919)
         );
  NAND2_X1 U9550 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U9551 ( .C1(n7920), .C2(n9042), .A(n7919), .B(n9907), .ZN(n7921)
         );
  AOI21_X1 U9552 ( .B1(n9774), .B2(n9045), .A(n7921), .ZN(n7922) );
  OAI21_X1 U9553 ( .B1(n7923), .B2(n9047), .A(n7922), .ZN(P1_U3213) );
  NAND2_X1 U9554 ( .A1(n4409), .A2(n7924), .ZN(n7978) );
  OAI21_X1 U9555 ( .B1(n7924), .B2(n4409), .A(n7978), .ZN(n7931) );
  OAI22_X1 U9556 ( .A1(n7969), .A2(n9998), .B1(n8048), .B2(n10000), .ZN(n7930)
         );
  AND2_X1 U9557 ( .A1(n7862), .A2(n7925), .ZN(n7928) );
  OAI21_X1 U9558 ( .B1(n7928), .B2(n7927), .A(n7926), .ZN(n8862) );
  NOR2_X1 U9559 ( .A1(n8862), .A2(n8736), .ZN(n7929) );
  AOI211_X1 U9560 ( .C1(n7931), .C2(n10020), .A(n7930), .B(n7929), .ZN(n8861)
         );
  AOI21_X1 U9561 ( .B1(n8858), .B2(n5042), .A(n7985), .ZN(n8859) );
  INV_X1 U9562 ( .A(n8858), .ZN(n7975) );
  AOI22_X1 U9563 ( .A1(n8766), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7972), .B2(
        n10002), .ZN(n7933) );
  OAI21_X1 U9564 ( .B1(n7975), .B2(n10031), .A(n7933), .ZN(n7935) );
  NOR2_X1 U9565 ( .A1(n8862), .A2(n10006), .ZN(n7934) );
  AOI211_X1 U9566 ( .C1(n8859), .C2(n10029), .A(n7935), .B(n7934), .ZN(n7936)
         );
  OAI21_X1 U9567 ( .B1(n8861), .B2(n8766), .A(n7936), .ZN(P2_U3283) );
  OR2_X1 U9568 ( .A1(n7949), .A2(n9352), .ZN(n8008) );
  NAND2_X1 U9569 ( .A1(n8011), .A2(n8008), .ZN(n9647) );
  INV_X1 U9570 ( .A(n9658), .ZN(n9043) );
  NAND2_X1 U9571 ( .A1(n9774), .A2(n9043), .ZN(n9112) );
  XNOR2_X1 U9572 ( .A(n9647), .B(n4394), .ZN(n9776) );
  OAI211_X1 U9573 ( .C1(n5040), .C2(n4394), .A(n8033), .B(n9656), .ZN(n7940)
         );
  AOI22_X1 U9574 ( .A1(n9660), .A2(n9351), .B1(n9659), .B2(n9352), .ZN(n7939)
         );
  NAND2_X1 U9575 ( .A1(n7940), .A2(n7939), .ZN(n9772) );
  INV_X1 U9576 ( .A(n9774), .ZN(n7946) );
  INV_X1 U9577 ( .A(n7941), .ZN(n7942) );
  AND2_X2 U9578 ( .A1(n7941), .A2(n7946), .ZN(n9666) );
  AOI211_X1 U9579 ( .C1(n9774), .C2(n7942), .A(n9944), .B(n9666), .ZN(n9773)
         );
  NAND2_X1 U9580 ( .A1(n9773), .A2(n9642), .ZN(n7945) );
  AOI22_X1 U9581 ( .A1(n9679), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7943), .B2(
        n9669), .ZN(n7944) );
  OAI211_X1 U9582 ( .C1(n7946), .C2(n9635), .A(n7945), .B(n7944), .ZN(n7947)
         );
  AOI21_X1 U9583 ( .B1(n7131), .B2(n9772), .A(n7947), .ZN(n7948) );
  OAI21_X1 U9584 ( .B1(n9776), .B2(n9645), .A(n7948), .ZN(P1_U3277) );
  INV_X1 U9585 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7955) );
  OAI22_X1 U9586 ( .A1(n7950), .A2(n9944), .B1(n5011), .B2(n9965), .ZN(n7951)
         );
  AOI21_X1 U9587 ( .B1(n7952), .B2(n9949), .A(n7951), .ZN(n7953) );
  AND2_X1 U9588 ( .A1(n7954), .A2(n7953), .ZN(n9819) );
  MUX2_X1 U9589 ( .A(n7955), .B(n9819), .S(n9977), .Z(n7956) );
  INV_X1 U9590 ( .A(n7956), .ZN(P1_U3536) );
  XNOR2_X1 U9591 ( .A(n8858), .B(n4379), .ZN(n7957) );
  NOR2_X1 U9592 ( .A1(n8208), .A2(n8251), .ZN(n7958) );
  NAND2_X1 U9593 ( .A1(n7957), .A2(n7958), .ZN(n8049) );
  INV_X1 U9594 ( .A(n7957), .ZN(n8209) );
  INV_X1 U9595 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9596 ( .A1(n8209), .A2(n7959), .ZN(n7960) );
  AND2_X1 U9597 ( .A1(n8049), .A2(n7960), .ZN(n7965) );
  INV_X1 U9598 ( .A(n7965), .ZN(n7961) );
  AOI21_X1 U9599 ( .B1(n7964), .B2(n7961), .A(n8426), .ZN(n7968) );
  NOR3_X1 U9600 ( .A1(n7962), .A2(n7969), .A3(n8402), .ZN(n7967) );
  NAND2_X1 U9601 ( .A1(n7964), .A2(n7963), .ZN(n7966) );
  OAI21_X1 U9602 ( .B1(n7968), .B2(n7967), .A(n8051), .ZN(n7974) );
  OAI22_X1 U9603 ( .A1(n7969), .A2(n8383), .B1(n8392), .B2(n8048), .ZN(n7970)
         );
  AOI211_X1 U9604 ( .C1(n8420), .C2(n7972), .A(n7971), .B(n7970), .ZN(n7973)
         );
  OAI211_X1 U9605 ( .C1(n7975), .C2(n8425), .A(n7974), .B(n7973), .ZN(P2_U3236) );
  NAND3_X1 U9606 ( .A1(n7978), .A2(n7976), .A3(n7977), .ZN(n8746) );
  INV_X1 U9607 ( .A(n8746), .ZN(n7980) );
  AOI21_X1 U9608 ( .B1(n7978), .B2(n7977), .A(n7976), .ZN(n7979) );
  NOR3_X1 U9609 ( .A1(n7980), .A2(n7979), .A3(n9995), .ZN(n7981) );
  OAI22_X1 U9610 ( .A1(n8731), .A2(n10000), .B1(n8208), .B2(n9998), .ZN(n8213)
         );
  NOR2_X1 U9611 ( .A1(n7981), .A2(n8213), .ZN(n8856) );
  OAI21_X1 U9612 ( .B1(n7984), .B2(n7983), .A(n7982), .ZN(n8852) );
  INV_X1 U9613 ( .A(n7985), .ZN(n7986) );
  AOI211_X1 U9614 ( .C1(n8854), .C2(n7986), .A(n10113), .B(n8758), .ZN(n8853)
         );
  NAND2_X1 U9615 ( .A1(n8853), .A2(n8720), .ZN(n7988) );
  AOI22_X1 U9616 ( .A1(n10036), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8212), .B2(
        n10002), .ZN(n7987) );
  OAI211_X1 U9617 ( .C1(n7989), .C2(n10031), .A(n7988), .B(n7987), .ZN(n7990)
         );
  AOI21_X1 U9618 ( .B1(n10034), .B2(n8852), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9619 ( .B1(n8856), .B2(n8766), .A(n7991), .ZN(P2_U3282) );
  INV_X1 U9620 ( .A(n7992), .ZN(n7996) );
  INV_X1 U9621 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7993) );
  OAI222_X1 U9622 ( .A1(n7994), .A2(P1_U3084), .B1(n9840), .B2(n7996), .C1(
        n7993), .C2(n9837), .ZN(P1_U3329) );
  INV_X1 U9623 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7995) );
  OAI222_X1 U9624 ( .A1(P2_U3152), .A2(n7997), .B1(n8906), .B2(n7996), .C1(
        n7995), .C2(n8093), .ZN(P2_U3334) );
  INV_X1 U9625 ( .A(n7998), .ZN(n8002) );
  OAI222_X1 U9626 ( .A1(n8093), .A2(n8000), .B1(n8906), .B2(n8002), .C1(
        P2_U3152), .C2(n7999), .ZN(P2_U3333) );
  OAI222_X1 U9627 ( .A1(n9837), .A2(n8003), .B1(n9840), .B2(n8002), .C1(n8001), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9628 ( .A(n8004), .ZN(n8144) );
  AOI21_X1 U9629 ( .B1(n8903), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8005), .ZN(
        n8006) );
  OAI21_X1 U9630 ( .B1(n8144), .B2(n8906), .A(n8006), .ZN(P2_U3330) );
  NAND2_X1 U9631 ( .A1(n9672), .A2(n9351), .ZN(n8013) );
  INV_X1 U9632 ( .A(n8013), .ZN(n8007) );
  INV_X1 U9633 ( .A(n9672), .ZN(n8028) );
  NAND2_X1 U9634 ( .A1(n8028), .A2(n9351), .ZN(n9117) );
  NAND2_X1 U9635 ( .A1(n9672), .A2(n9630), .ZN(n8035) );
  NOR2_X1 U9636 ( .A1(n8007), .A2(n9652), .ZN(n8015) );
  NOR2_X1 U9637 ( .A1(n9774), .A2(n9658), .ZN(n9646) );
  INV_X1 U9638 ( .A(n8008), .ZN(n8009) );
  OR2_X1 U9639 ( .A1(n9646), .A2(n8009), .ZN(n8010) );
  NOR2_X1 U9640 ( .A1(n8015), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U9641 ( .A1(n9774), .A2(n9658), .ZN(n9648) );
  AND2_X1 U9642 ( .A1(n9648), .A2(n8013), .ZN(n8014) );
  OR2_X1 U9643 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U9644 ( .A1(n9764), .A2(n8991), .ZN(n9221) );
  NAND2_X1 U9645 ( .A1(n9235), .A2(n9221), .ZN(n9116) );
  AND2_X1 U9646 ( .A1(n9764), .A2(n9661), .ZN(n8017) );
  NOR2_X1 U9647 ( .A1(n9759), .A2(n9607), .ZN(n8018) );
  OR2_X1 U9648 ( .A1(n9616), .A2(n8933), .ZN(n9121) );
  NAND2_X1 U9649 ( .A1(n9616), .A2(n8933), .ZN(n9123) );
  NAND2_X1 U9650 ( .A1(n9121), .A2(n9123), .ZN(n9174) );
  INV_X1 U9651 ( .A(n9616), .ZN(n9752) );
  OR2_X1 U9652 ( .A1(n9745), .A2(n9608), .ZN(n8019) );
  NAND2_X1 U9653 ( .A1(n9583), .A2(n8019), .ZN(n8020) );
  INV_X1 U9654 ( .A(n9745), .ZN(n9592) );
  INV_X1 U9655 ( .A(n9608), .ZN(n9001) );
  NAND2_X1 U9656 ( .A1(n8020), .A2(n5049), .ZN(n9569) );
  INV_X1 U9657 ( .A(n9596), .ZN(n8934) );
  INV_X1 U9658 ( .A(n9740), .ZN(n9574) );
  OR2_X1 U9659 ( .A1(n9736), .A2(n9349), .ZN(n9130) );
  NAND2_X1 U9660 ( .A1(n9736), .A2(n9349), .ZN(n9134) );
  NAND2_X1 U9661 ( .A1(n9130), .A2(n9134), .ZN(n9555) );
  INV_X1 U9662 ( .A(n9736), .ZN(n9560) );
  INV_X1 U9663 ( .A(n9564), .ZN(n8926) );
  NAND2_X1 U9664 ( .A1(n9532), .A2(n9517), .ZN(n8023) );
  AOI22_X1 U9665 ( .A1(n9526), .A2(n8023), .B1(n9549), .B2(n9725), .ZN(n9511)
         );
  NAND2_X1 U9666 ( .A1(n9722), .A2(n8024), .ZN(n8025) );
  NAND2_X1 U9667 ( .A1(n9715), .A2(n9518), .ZN(n9143) );
  NAND2_X1 U9668 ( .A1(n9484), .A2(n9143), .ZN(n9504) );
  NAND2_X1 U9669 ( .A1(n9706), .A2(n8026), .ZN(n9217) );
  NAND2_X1 U9670 ( .A1(n9666), .A2(n8028), .ZN(n9668) );
  INV_X1 U9671 ( .A(n9759), .ZN(n8997) );
  AND2_X1 U9672 ( .A1(n9752), .A2(n8997), .ZN(n8029) );
  AND2_X2 U9673 ( .A1(n9634), .A2(n8029), .ZN(n9585) );
  OR2_X2 U9674 ( .A1(n9540), .A2(n9725), .ZN(n9527) );
  NOR2_X4 U9675 ( .A1(n9722), .A2(n9527), .ZN(n9519) );
  INV_X1 U9676 ( .A(n9480), .ZN(n8031) );
  INV_X1 U9677 ( .A(n8151), .ZN(n8030) );
  AOI211_X1 U9678 ( .C1(n9706), .C2(n8031), .A(n9944), .B(n8030), .ZN(n9705)
         );
  AOI22_X1 U9679 ( .A1(n8914), .A2(n9669), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9679), .ZN(n8032) );
  OAI21_X1 U9680 ( .B1(n8919), .B2(n9635), .A(n8032), .ZN(n8042) );
  INV_X1 U9681 ( .A(n9607), .ZN(n9632) );
  NAND2_X1 U9682 ( .A1(n9759), .A2(n9632), .ZN(n9602) );
  AND2_X1 U9683 ( .A1(n9123), .A2(n9602), .ZN(n9222) );
  OR2_X1 U9684 ( .A1(n9759), .A2(n9632), .ZN(n9603) );
  NAND2_X1 U9685 ( .A1(n9121), .A2(n9603), .ZN(n9076) );
  OR2_X1 U9686 ( .A1(n9745), .A2(n9001), .ZN(n9125) );
  NAND2_X1 U9687 ( .A1(n9745), .A2(n9001), .ZN(n9223) );
  NAND2_X1 U9688 ( .A1(n9125), .A2(n9223), .ZN(n9584) );
  NAND2_X1 U9689 ( .A1(n9594), .A2(n8036), .ZN(n9593) );
  OR2_X1 U9690 ( .A1(n9740), .A2(n8934), .ZN(n9135) );
  NAND2_X1 U9691 ( .A1(n9740), .A2(n8934), .ZN(n9129) );
  INV_X1 U9692 ( .A(n9555), .ZN(n9563) );
  OR2_X1 U9693 ( .A1(n9731), .A2(n8926), .ZN(n9133) );
  NAND2_X1 U9694 ( .A1(n9731), .A2(n8926), .ZN(n9137) );
  NAND2_X1 U9695 ( .A1(n9722), .A2(n8963), .ZN(n9070) );
  NAND2_X1 U9696 ( .A1(n9725), .A2(n9517), .ZN(n9512) );
  AND2_X1 U9697 ( .A1(n9070), .A2(n9512), .ZN(n9069) );
  NAND2_X1 U9698 ( .A1(n8037), .A2(n9249), .ZN(n9505) );
  INV_X1 U9699 ( .A(n9506), .ZN(n8964) );
  OR2_X1 U9700 ( .A1(n9710), .A2(n8964), .ZN(n9074) );
  NAND2_X1 U9701 ( .A1(n9710), .A2(n8964), .ZN(n9215) );
  AOI21_X1 U9702 ( .B1(n8038), .B2(n9316), .A(n9628), .ZN(n8040) );
  OAI22_X1 U9703 ( .A1(n8148), .A2(n9633), .B1(n8964), .B2(n9631), .ZN(n8039)
         );
  AOI21_X1 U9704 ( .B1(n8040), .B2(n8154), .A(n8039), .ZN(n9708) );
  NOR2_X1 U9705 ( .A1(n9708), .A2(n9679), .ZN(n8041) );
  AOI211_X1 U9706 ( .C1(n9642), .C2(n9705), .A(n8042), .B(n8041), .ZN(n8043)
         );
  OAI21_X1 U9707 ( .B1(n9709), .B2(n9645), .A(n8043), .ZN(P1_U3264) );
  OAI222_X1 U9708 ( .A1(n8044), .A2(P1_U3084), .B1(n9840), .B2(n8046), .C1(
        n10304), .C2(n9837), .ZN(P1_U3351) );
  OAI222_X1 U9709 ( .A1(n8047), .A2(P2_U3152), .B1(n8906), .B2(n8046), .C1(
        n8045), .C2(n8093), .ZN(P2_U3356) );
  INV_X1 U9710 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10272) );
  INV_X1 U9711 ( .A(n9054), .ZN(n8896) );
  OAI222_X1 U9712 ( .A1(n9837), .A2(n10272), .B1(n9840), .B2(n8896), .C1(n6070), .C2(P1_U3084), .ZN(P1_U3323) );
  XNOR2_X1 U9713 ( .A(n8854), .B(n7176), .ZN(n8054) );
  NOR2_X1 U9714 ( .A1(n8048), .A2(n8251), .ZN(n8052) );
  XNOR2_X1 U9715 ( .A(n8054), .B(n8052), .ZN(n8221) );
  AND2_X1 U9716 ( .A1(n8221), .A2(n8049), .ZN(n8050) );
  XNOR2_X1 U9717 ( .A(n8842), .B(n7176), .ZN(n8304) );
  OR2_X1 U9718 ( .A1(n8332), .A2(n8251), .ZN(n8303) );
  XNOR2_X1 U9719 ( .A(n5704), .B(n4379), .ZN(n8298) );
  NOR2_X1 U9720 ( .A1(n8731), .A2(n8251), .ZN(n8427) );
  INV_X1 U9721 ( .A(n8052), .ZN(n8053) );
  NAND2_X1 U9722 ( .A1(n8054), .A2(n8053), .ZN(n8297) );
  OAI21_X1 U9723 ( .B1(n8298), .B2(n8427), .A(n8297), .ZN(n8055) );
  AOI21_X1 U9724 ( .B1(n8304), .B2(n8303), .A(n8055), .ZN(n8325) );
  XNOR2_X1 U9725 ( .A(n8838), .B(n4379), .ZN(n8056) );
  NOR2_X1 U9726 ( .A1(n8732), .A2(n8251), .ZN(n8057) );
  NAND2_X1 U9727 ( .A1(n8056), .A2(n8057), .ZN(n8065) );
  INV_X1 U9728 ( .A(n8056), .ZN(n8082) );
  INV_X1 U9729 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U9730 ( .A1(n8082), .A2(n8058), .ZN(n8059) );
  AND2_X1 U9731 ( .A1(n8325), .A2(n8330), .ZN(n8064) );
  INV_X1 U9732 ( .A(n8330), .ZN(n8063) );
  INV_X1 U9733 ( .A(n8304), .ZN(n8062) );
  INV_X1 U9734 ( .A(n8298), .ZN(n8301) );
  INV_X1 U9735 ( .A(n8427), .ZN(n8307) );
  OAI21_X1 U9736 ( .B1(n8301), .B2(n8307), .A(n8303), .ZN(n8061) );
  NOR2_X1 U9737 ( .A1(n8303), .A2(n8307), .ZN(n8060) );
  AOI22_X1 U9738 ( .A1(n8062), .A2(n8061), .B1(n8060), .B2(n8298), .ZN(n8327)
         );
  XNOR2_X1 U9739 ( .A(n8700), .B(n4379), .ZN(n8067) );
  NOR2_X1 U9740 ( .A1(n8331), .A2(n8251), .ZN(n8068) );
  XNOR2_X1 U9741 ( .A(n8067), .B(n8068), .ZN(n8081) );
  INV_X1 U9742 ( .A(n8067), .ZN(n8069) );
  NAND2_X1 U9743 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  XNOR2_X1 U9744 ( .A(n8828), .B(n4379), .ZN(n8074) );
  INV_X1 U9745 ( .A(n8074), .ZN(n8072) );
  NOR2_X1 U9746 ( .A1(n8695), .A2(n8251), .ZN(n8073) );
  INV_X1 U9747 ( .A(n8073), .ZN(n8071) );
  AND2_X1 U9748 ( .A1(n8074), .A2(n8073), .ZN(n8167) );
  NOR2_X1 U9749 ( .A1(n4472), .A2(n8167), .ZN(n8075) );
  XNOR2_X1 U9750 ( .A(n8168), .B(n8075), .ZN(n8079) );
  AOI22_X1 U9751 ( .A1(n8422), .A2(n8708), .B1(n8421), .B2(n8686), .ZN(n8076)
         );
  NAND2_X1 U9752 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8118) );
  OAI211_X1 U9753 ( .C1(n8412), .C2(n8677), .A(n8076), .B(n8118), .ZN(n8077)
         );
  AOI21_X1 U9754 ( .B1(n8828), .B2(n8386), .A(n8077), .ZN(n8078) );
  OAI21_X1 U9755 ( .B1(n8079), .B2(n8426), .A(n8078), .ZN(P2_U3221) );
  AOI21_X1 U9756 ( .B1(n8080), .B2(n4871), .A(n8426), .ZN(n8085) );
  NOR3_X1 U9757 ( .A1(n8082), .A2(n8732), .A3(n8402), .ZN(n8084) );
  OAI21_X1 U9758 ( .B1(n8085), .B2(n8084), .A(n8083), .ZN(n8090) );
  INV_X1 U9759 ( .A(n8086), .ZN(n8697) );
  NAND2_X1 U9760 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8521) );
  INV_X1 U9761 ( .A(n8521), .ZN(n8088) );
  OAI22_X1 U9762 ( .A1(n8732), .A2(n8383), .B1(n8392), .B2(n8695), .ZN(n8087)
         );
  AOI211_X1 U9763 ( .C1(n8420), .C2(n8697), .A(n8088), .B(n8087), .ZN(n8089)
         );
  OAI211_X1 U9764 ( .C1(n8700), .C2(n8425), .A(n8090), .B(n8089), .ZN(P2_U3240) );
  OAI222_X1 U9765 ( .A1(n8093), .A2(n8092), .B1(n8906), .B2(n8091), .C1(
        P2_U3152), .C2(n5716), .ZN(P2_U3336) );
  NAND2_X1 U9766 ( .A1(n8922), .A2(n8921), .ZN(n8920) );
  NAND2_X1 U9767 ( .A1(n8094), .A2(n8095), .ZN(n8924) );
  NAND2_X1 U9768 ( .A1(n8096), .A2(n8956), .ZN(n8097) );
  AOI21_X1 U9769 ( .B1(n8920), .B2(n8924), .A(n8097), .ZN(n8959) );
  AND3_X1 U9770 ( .A1(n8920), .A2(n8924), .A3(n8097), .ZN(n8098) );
  OAI21_X1 U9771 ( .B1(n8959), .B2(n8098), .A(n8986), .ZN(n8102) );
  AOI22_X1 U9772 ( .A1(n9549), .A2(n8951), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8099) );
  OAI21_X1 U9773 ( .B1(n9013), .B2(n9520), .A(n8099), .ZN(n8100) );
  AOI21_X1 U9774 ( .B1(n9040), .B2(n9488), .A(n8100), .ZN(n8101) );
  OAI211_X1 U9775 ( .C1(n8103), .C2(n8996), .A(n8102), .B(n8101), .ZN(P1_U3227) );
  XNOR2_X1 U9776 ( .A(n8110), .B(n8105), .ZN(n8520) );
  INV_X1 U9777 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U9778 ( .A1(n8520), .A2(n8519), .ZN(n8518) );
  NAND2_X1 U9779 ( .A1(n8105), .A2(n8530), .ZN(n8106) );
  NAND2_X1 U9780 ( .A1(n8518), .A2(n8106), .ZN(n8107) );
  XNOR2_X1 U9781 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8107), .ZN(n8115) );
  INV_X1 U9782 ( .A(n8115), .ZN(n8113) );
  AOI21_X1 U9783 ( .B1(n8109), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8108), .ZN(
        n8526) );
  XNOR2_X1 U9784 ( .A(n8110), .B(n10256), .ZN(n8525) );
  NAND2_X1 U9785 ( .A1(n8526), .A2(n8525), .ZN(n8524) );
  OAI21_X1 U9786 ( .B1(n8110), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8524), .ZN(
        n8111) );
  XNOR2_X1 U9787 ( .A(n8111), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8114) );
  OAI21_X1 U9788 ( .B1(n8114), .B2(n9984), .A(n9983), .ZN(n8112) );
  AOI22_X1 U9789 ( .A1(n8115), .A2(n9979), .B1(n9978), .B2(n8114), .ZN(n8116)
         );
  MUX2_X1 U9790 ( .A(n8117), .B(n8116), .S(n8575), .Z(n8119) );
  OAI211_X1 U9791 ( .C1(n8522), .C2(n9872), .A(n8119), .B(n8118), .ZN(P2_U3264) );
  INV_X1 U9792 ( .A(n8120), .ZN(n8122) );
  OR2_X1 U9793 ( .A1(n8121), .A2(P2_U3152), .ZN(n8269) );
  AOI22_X1 U9794 ( .A1(n8415), .A2(n8122), .B1(n8269), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8127) );
  OAI211_X1 U9795 ( .C1(n8125), .C2(n8124), .A(n8398), .B(n8123), .ZN(n8126)
         );
  OAI211_X1 U9796 ( .C1(n8425), .C2(n10057), .A(n8127), .B(n8126), .ZN(
        P2_U3239) );
  XNOR2_X1 U9797 ( .A(n4476), .B(n9175), .ZN(n9761) );
  XNOR2_X1 U9798 ( .A(n4384), .B(n9175), .ZN(n8129) );
  OAI222_X1 U9799 ( .A1(n9633), .A2(n8933), .B1(n9631), .B2(n8991), .C1(n9628), 
        .C2(n8129), .ZN(n9757) );
  INV_X1 U9800 ( .A(n9634), .ZN(n8130) );
  AND2_X1 U9801 ( .A1(n9634), .A2(n8997), .ZN(n9611) );
  AOI211_X1 U9802 ( .C1(n9759), .C2(n8130), .A(n9944), .B(n9611), .ZN(n9758)
         );
  NAND2_X1 U9803 ( .A1(n9758), .A2(n9642), .ZN(n8132) );
  AOI22_X1 U9804 ( .A1(n9679), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8990), .B2(
        n9669), .ZN(n8131) );
  OAI211_X1 U9805 ( .C1(n8997), .C2(n9635), .A(n8132), .B(n8131), .ZN(n8133)
         );
  AOI21_X1 U9806 ( .B1(n9757), .B2(n7131), .A(n8133), .ZN(n8134) );
  OAI21_X1 U9807 ( .B1(n9645), .B2(n9761), .A(n8134), .ZN(P1_U3274) );
  AOI21_X1 U9808 ( .B1(n8136), .B2(n8549), .A(n8162), .ZN(n8770) );
  NAND2_X1 U9809 ( .A1(n8770), .A2(n10029), .ZN(n8143) );
  INV_X1 U9810 ( .A(P2_B_REG_SCAN_IN), .ZN(n8137) );
  NOR2_X1 U9811 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  NOR2_X1 U9812 ( .A1(n10000), .A2(n8139), .ZN(n8536) );
  INV_X1 U9813 ( .A(n8536), .ZN(n8140) );
  OR2_X1 U9814 ( .A1(n8141), .A2(n8140), .ZN(n8771) );
  NOR2_X1 U9815 ( .A1(n8766), .A2(n8771), .ZN(n8163) );
  AOI21_X1 U9816 ( .B1(n8766), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8163), .ZN(
        n8142) );
  OAI211_X1 U9817 ( .C1(n8773), .C2(n10031), .A(n8143), .B(n8142), .ZN(
        P2_U3266) );
  OAI222_X1 U9818 ( .A1(n9837), .A2(n8146), .B1(P1_U3084), .B2(n8145), .C1(
        n9840), .C2(n8144), .ZN(P1_U3325) );
  OAI21_X1 U9819 ( .B1(n8149), .B2(n9205), .A(n9689), .ZN(n9704) );
  INV_X1 U9820 ( .A(n9470), .ZN(n8150) );
  AOI21_X1 U9821 ( .B1(n9700), .B2(n8151), .A(n8150), .ZN(n9701) );
  AOI22_X1 U9822 ( .A1(n8152), .A2(n9669), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9679), .ZN(n8153) );
  OAI21_X1 U9823 ( .B1(n5015), .B2(n9635), .A(n8153), .ZN(n8159) );
  XNOR2_X1 U9824 ( .A(n9463), .B(n9205), .ZN(n8158) );
  AOI21_X2 U9825 ( .B1(n8158), .B2(n9656), .A(n8157), .ZN(n9703) );
  OAI21_X1 U9826 ( .B1(n9704), .B2(n9645), .A(n8160), .ZN(P1_U3263) );
  AOI21_X1 U9827 ( .B1(n10036), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8163), .ZN(
        n8165) );
  NAND2_X1 U9828 ( .A1(n5818), .A2(n8756), .ZN(n8164) );
  OAI211_X1 U9829 ( .C1(n8767), .C2(n8166), .A(n8165), .B(n8164), .ZN(P2_U3265) );
  XNOR2_X1 U9830 ( .A(n8822), .B(n7176), .ZN(n8169) );
  NAND2_X1 U9831 ( .A1(n8686), .A2(n8188), .ZN(n8170) );
  XNOR2_X1 U9832 ( .A(n8169), .B(n8170), .ZN(n8366) );
  INV_X1 U9833 ( .A(n8169), .ZN(n8172) );
  INV_X1 U9834 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U9835 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  XNOR2_X1 U9836 ( .A(n8650), .B(n7176), .ZN(n8179) );
  NAND2_X1 U9837 ( .A1(n8668), .A2(n8188), .ZN(n8175) );
  XNOR2_X1 U9838 ( .A(n8179), .B(n8175), .ZN(n8278) );
  NAND2_X1 U9839 ( .A1(n8279), .A2(n8278), .ZN(n8375) );
  INV_X1 U9840 ( .A(n8375), .ZN(n8174) );
  XNOR2_X1 U9841 ( .A(n8812), .B(n7176), .ZN(n8176) );
  NAND2_X1 U9842 ( .A1(n8654), .A2(n8188), .ZN(n8380) );
  NOR2_X1 U9843 ( .A1(n8639), .A2(n8251), .ZN(n8184) );
  XNOR2_X1 U9844 ( .A(n8807), .B(n4379), .ZN(n8183) );
  INV_X1 U9845 ( .A(n8175), .ZN(n8178) );
  NAND2_X1 U9846 ( .A1(n8179), .A2(n8178), .ZN(n8374) );
  NAND2_X1 U9847 ( .A1(n8374), .A2(n8380), .ZN(n8177) );
  INV_X1 U9848 ( .A(n8176), .ZN(n8376) );
  NAND2_X1 U9849 ( .A1(n8177), .A2(n8376), .ZN(n8181) );
  NAND3_X1 U9850 ( .A1(n8179), .A2(n8178), .A3(n8654), .ZN(n8180) );
  NAND2_X1 U9851 ( .A1(n8181), .A2(n8180), .ZN(n8223) );
  AOI21_X1 U9852 ( .B1(n8184), .B2(n8183), .A(n8223), .ZN(n8182) );
  XNOR2_X1 U9853 ( .A(n8801), .B(n7176), .ZN(n8340) );
  NAND2_X1 U9854 ( .A1(n8613), .A2(n8188), .ZN(n8343) );
  INV_X1 U9855 ( .A(n8183), .ZN(n8226) );
  INV_X1 U9856 ( .A(n8184), .ZN(n8228) );
  AND2_X1 U9857 ( .A1(n8226), .A2(n8228), .ZN(n8337) );
  AOI21_X1 U9858 ( .B1(n8340), .B2(n8343), .A(n8337), .ZN(n8187) );
  INV_X1 U9859 ( .A(n8340), .ZN(n8186) );
  INV_X1 U9860 ( .A(n8343), .ZN(n8185) );
  NAND2_X1 U9861 ( .A1(n8436), .A2(n8188), .ZN(n8288) );
  XNOR2_X1 U9862 ( .A(n8793), .B(n4379), .ZN(n8197) );
  NOR2_X1 U9863 ( .A1(n8196), .A2(n8251), .ZN(n8189) );
  OAI21_X1 U9864 ( .B1(n8197), .B2(n8189), .A(n8200), .ZN(n8409) );
  XNOR2_X1 U9865 ( .A(n8788), .B(n4379), .ZN(n8191) );
  NOR2_X1 U9866 ( .A1(n8410), .A2(n8251), .ZN(n8192) );
  NAND2_X1 U9867 ( .A1(n8191), .A2(n8192), .ZN(n8254) );
  INV_X1 U9868 ( .A(n8191), .ZN(n8194) );
  INV_X1 U9869 ( .A(n8192), .ZN(n8193) );
  NAND2_X1 U9870 ( .A1(n8194), .A2(n8193), .ZN(n8195) );
  AND2_X1 U9871 ( .A1(n8254), .A2(n8195), .ZN(n8201) );
  INV_X1 U9872 ( .A(n8402), .ZN(n8378) );
  INV_X1 U9873 ( .A(n8196), .ZN(n8435) );
  NAND3_X1 U9874 ( .A1(n8197), .A2(n8378), .A3(n8435), .ZN(n8198) );
  OAI21_X1 U9875 ( .B1(n8199), .B2(n8426), .A(n8198), .ZN(n8202) );
  OAI22_X1 U9876 ( .A1(n8203), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4610), .ZN(n8204) );
  AOI21_X1 U9877 ( .B1(n8205), .B2(n8415), .A(n8204), .ZN(n8206) );
  INV_X1 U9878 ( .A(n8051), .ZN(n8211) );
  NOR3_X1 U9879 ( .A1(n8209), .A2(n8208), .A3(n8402), .ZN(n8210) );
  AOI21_X1 U9880 ( .B1(n8211), .B2(n8398), .A(n8210), .ZN(n8222) );
  INV_X1 U9881 ( .A(n8212), .ZN(n8216) );
  NAND2_X1 U9882 ( .A1(n8415), .A2(n8213), .ZN(n8214) );
  OAI211_X1 U9883 ( .C1(n8412), .C2(n8216), .A(n8215), .B(n8214), .ZN(n8219)
         );
  NOR2_X1 U9884 ( .A1(n8326), .A2(n8426), .ZN(n8218) );
  AOI211_X1 U9885 ( .C1(n8854), .C2(n8386), .A(n8219), .B(n8218), .ZN(n8220)
         );
  OAI21_X1 U9886 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(P2_U3217) );
  INV_X1 U9887 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U9888 ( .A1(n8225), .A2(n8224), .ZN(n8227) );
  XNOR2_X1 U9889 ( .A(n8227), .B(n8226), .ZN(n8229) );
  NAND3_X1 U9890 ( .A1(n8229), .A2(n8398), .A3(n8228), .ZN(n8237) );
  INV_X1 U9891 ( .A(n8229), .ZN(n8230) );
  INV_X1 U9892 ( .A(n8639), .ZN(n8437) );
  NAND3_X1 U9893 ( .A1(n8230), .A2(n8378), .A3(n8437), .ZN(n8236) );
  OAI22_X1 U9894 ( .A1(n8412), .A2(n8621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8231), .ZN(n8234) );
  OAI22_X1 U9895 ( .A1(n8232), .A2(n8392), .B1(n8383), .B2(n8282), .ZN(n8233)
         );
  AOI211_X1 U9896 ( .C1(n8807), .C2(n8386), .A(n8234), .B(n8233), .ZN(n8235)
         );
  NAND3_X1 U9897 ( .A1(n8237), .A2(n8236), .A3(n8235), .ZN(P2_U3218) );
  NOR3_X1 U9898 ( .A1(n8402), .A2(n8239), .A3(n8238), .ZN(n8244) );
  INV_X1 U9899 ( .A(n8240), .ZN(n8241) );
  AOI21_X1 U9900 ( .B1(n8123), .B2(n8241), .A(n8426), .ZN(n8243) );
  OAI21_X1 U9901 ( .B1(n8244), .B2(n8243), .A(n8359), .ZN(n8250) );
  AOI22_X1 U9902 ( .A1(n8422), .A2(n10016), .B1(n8420), .B2(n8246), .ZN(n8249)
         );
  INV_X1 U9903 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U9904 ( .A1(n8386), .A2(n5163), .ZN(n8245) );
  OAI21_X1 U9905 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8246), .A(n8245), .ZN(n8247) );
  AOI21_X1 U9906 ( .B1(n8421), .B2(n10018), .A(n8247), .ZN(n8248) );
  NAND3_X1 U9907 ( .A1(n8250), .A2(n8249), .A3(n8248), .ZN(P2_U3220) );
  OR2_X1 U9908 ( .A1(n8543), .A2(n8251), .ZN(n8252) );
  XNOR2_X1 U9909 ( .A(n8252), .B(n7176), .ZN(n8256) );
  INV_X1 U9910 ( .A(n8256), .ZN(n8257) );
  NOR3_X1 U9911 ( .A1(n4943), .A2(n8257), .A3(n8386), .ZN(n8253) );
  AOI21_X1 U9912 ( .B1(n4943), .B2(n8257), .A(n8253), .ZN(n8264) );
  NOR3_X1 U9913 ( .A1(n4943), .A2(n8256), .A3(n8386), .ZN(n8260) );
  NOR2_X1 U9914 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  OAI21_X1 U9915 ( .B1(n4943), .B2(n8425), .A(n8426), .ZN(n8261) );
  OAI211_X1 U9916 ( .C1(n8264), .C2(n8263), .A(n8262), .B(n8261), .ZN(n8268)
         );
  AOI22_X1 U9917 ( .A1(n8557), .A2(n8420), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8267) );
  INV_X1 U9918 ( .A(n8265), .ZN(n8433) );
  AOI22_X1 U9919 ( .A1(n8433), .A2(n8421), .B1(n8422), .B2(n8434), .ZN(n8266)
         );
  NAND3_X1 U9920 ( .A1(n8268), .A2(n8267), .A3(n8266), .ZN(P2_U3222) );
  AOI22_X1 U9921 ( .A1(n8422), .A2(n8451), .B1(n8421), .B2(n10016), .ZN(n8277)
         );
  AOI22_X1 U9922 ( .A1(n8386), .A2(n5123), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8269), .ZN(n8276) );
  INV_X1 U9923 ( .A(n8270), .ZN(n8274) );
  AND2_X1 U9924 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  OAI21_X1 U9925 ( .B1(n8274), .B2(n8273), .A(n8398), .ZN(n8275) );
  NAND3_X1 U9926 ( .A1(n8277), .A2(n8276), .A3(n8275), .ZN(P2_U3224) );
  XNOR2_X1 U9927 ( .A(n8279), .B(n8278), .ZN(n8287) );
  INV_X1 U9928 ( .A(n8648), .ZN(n8281) );
  OAI22_X1 U9929 ( .A1(n8412), .A2(n8281), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8280), .ZN(n8285) );
  OAI22_X1 U9930 ( .A1(n8283), .A2(n8383), .B1(n8392), .B2(n8282), .ZN(n8284)
         );
  AOI211_X1 U9931 ( .C1(n8817), .C2(n8386), .A(n8285), .B(n8284), .ZN(n8286)
         );
  OAI21_X1 U9932 ( .B1(n8287), .B2(n8426), .A(n8286), .ZN(P2_U3225) );
  XNOR2_X1 U9933 ( .A(n8289), .B(n8288), .ZN(n8290) );
  XNOR2_X1 U9934 ( .A(n8291), .B(n8290), .ZN(n8296) );
  AOI22_X1 U9935 ( .A1(n8435), .A2(n10017), .B1(n10015), .B2(n8613), .ZN(n8583) );
  NOR2_X1 U9936 ( .A1(n8583), .A2(n8292), .ZN(n8294) );
  OAI22_X1 U9937 ( .A1(n8586), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4609), .ZN(n8293) );
  AOI211_X1 U9938 ( .C1(n8799), .C2(n8386), .A(n8294), .B(n8293), .ZN(n8295)
         );
  OAI21_X1 U9939 ( .B1(n8296), .B2(n8426), .A(n8295), .ZN(P2_U3227) );
  NAND2_X1 U9940 ( .A1(n8300), .A2(n8298), .ZN(n8418) );
  INV_X1 U9941 ( .A(n8418), .ZN(n8299) );
  NOR2_X1 U9942 ( .A1(n8402), .A2(n8731), .ZN(n8431) );
  AOI21_X1 U9943 ( .B1(n8299), .B2(n8398), .A(n8431), .ZN(n8314) );
  INV_X1 U9944 ( .A(n8300), .ZN(n8302) );
  NAND2_X1 U9945 ( .A1(n8302), .A2(n8301), .ZN(n8417) );
  XNOR2_X1 U9946 ( .A(n8304), .B(n8303), .ZN(n8308) );
  NAND2_X1 U9947 ( .A1(n8417), .A2(n8308), .ZN(n8313) );
  INV_X1 U9948 ( .A(n8739), .ZN(n8306) );
  AOI22_X1 U9949 ( .A1(n8422), .A2(n8439), .B1(n8421), .B2(n8438), .ZN(n8305)
         );
  NAND2_X1 U9950 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8506) );
  OAI211_X1 U9951 ( .C1(n8412), .C2(n8306), .A(n8305), .B(n8506), .ZN(n8311)
         );
  NAND2_X1 U9952 ( .A1(n8418), .A2(n8307), .ZN(n8309) );
  AOI211_X1 U9953 ( .C1(n8309), .C2(n8417), .A(n8308), .B(n8426), .ZN(n8310)
         );
  AOI211_X1 U9954 ( .C1(n8842), .C2(n8386), .A(n8311), .B(n8310), .ZN(n8312)
         );
  OAI21_X1 U9955 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(P2_U3228) );
  AOI21_X1 U9956 ( .B1(n8316), .B2(n8315), .A(n8426), .ZN(n8317) );
  NAND2_X1 U9957 ( .A1(n8317), .A2(n8397), .ZN(n8324) );
  INV_X1 U9958 ( .A(n8318), .ZN(n8319) );
  AOI22_X1 U9959 ( .A1(n8415), .A2(n8319), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8323) );
  AOI22_X1 U9960 ( .A1(n8386), .A2(n8321), .B1(n8420), .B2(n8320), .ZN(n8322)
         );
  NAND3_X1 U9961 ( .A1(n8324), .A2(n8323), .A3(n8322), .ZN(P2_U3229) );
  NAND2_X1 U9962 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  NAND2_X1 U9963 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  OAI211_X1 U9964 ( .C1(n8330), .C2(n8329), .A(n8080), .B(n8398), .ZN(n8336)
         );
  OAI22_X1 U9965 ( .A1(n8412), .A2(n8715), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4613), .ZN(n8334) );
  OAI22_X1 U9966 ( .A1(n8332), .A2(n8383), .B1(n8392), .B2(n8331), .ZN(n8333)
         );
  AOI211_X1 U9967 ( .C1(n8838), .C2(n8386), .A(n8334), .B(n8333), .ZN(n8335)
         );
  NAND2_X1 U9968 ( .A1(n8336), .A2(n8335), .ZN(P2_U3230) );
  INV_X1 U9969 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U9970 ( .A1(n8339), .A2(n8338), .ZN(n8341) );
  XNOR2_X1 U9971 ( .A(n8341), .B(n8340), .ZN(n8342) );
  NAND3_X1 U9972 ( .A1(n8342), .A2(n8378), .A3(n8613), .ZN(n8351) );
  INV_X1 U9973 ( .A(n8342), .ZN(n8344) );
  NAND3_X1 U9974 ( .A1(n8344), .A2(n8398), .A3(n8343), .ZN(n8350) );
  INV_X1 U9975 ( .A(n8602), .ZN(n8346) );
  OAI22_X1 U9976 ( .A1(n8346), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8345), .ZN(n8348) );
  OAI22_X1 U9977 ( .A1(n8592), .A2(n8392), .B1(n8639), .B2(n8383), .ZN(n8347)
         );
  AOI211_X1 U9978 ( .C1(n8801), .C2(n8386), .A(n8348), .B(n8347), .ZN(n8349)
         );
  NAND3_X1 U9979 ( .A1(n8351), .A2(n8350), .A3(n8349), .ZN(P2_U3231) );
  INV_X1 U9980 ( .A(n8360), .ZN(n8353) );
  NAND4_X1 U9981 ( .A1(n8378), .A2(n8353), .A3(n8450), .A4(n8352), .ZN(n8365)
         );
  INV_X1 U9982 ( .A(n8354), .ZN(n8355) );
  AOI22_X1 U9983 ( .A1(n8415), .A2(n8355), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8364) );
  AOI22_X1 U9984 ( .A1(n8386), .A2(n8357), .B1(n8420), .B2(n8356), .ZN(n8363)
         );
  OAI21_X1 U9985 ( .B1(n8360), .B2(n8359), .A(n8358), .ZN(n8361) );
  NAND2_X1 U9986 ( .A1(n8361), .A2(n8398), .ZN(n8362) );
  NAND4_X1 U9987 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(
        P2_U3232) );
  XNOR2_X1 U9988 ( .A(n8367), .B(n8366), .ZN(n8373) );
  OAI22_X1 U9989 ( .A1(n8412), .A2(n8369), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8368), .ZN(n8371) );
  OAI22_X1 U9990 ( .A1(n8695), .A2(n8383), .B1(n8392), .B2(n8638), .ZN(n8370)
         );
  AOI211_X1 U9991 ( .C1(n8822), .C2(n8386), .A(n8371), .B(n8370), .ZN(n8372)
         );
  OAI21_X1 U9992 ( .B1(n8373), .B2(n8426), .A(n8372), .ZN(P2_U3235) );
  NAND2_X1 U9993 ( .A1(n8375), .A2(n8374), .ZN(n8377) );
  XNOR2_X1 U9994 ( .A(n8377), .B(n8376), .ZN(n8379) );
  NAND3_X1 U9995 ( .A1(n8379), .A2(n8378), .A3(n8654), .ZN(n8389) );
  INV_X1 U9996 ( .A(n8379), .ZN(n8381) );
  NAND3_X1 U9997 ( .A1(n8381), .A2(n8398), .A3(n8380), .ZN(n8388) );
  OAI22_X1 U9998 ( .A1(n8412), .A2(n8631), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8382), .ZN(n8385) );
  OAI22_X1 U9999 ( .A1(n8638), .A2(n8383), .B1(n8392), .B2(n8639), .ZN(n8384)
         );
  AOI211_X1 U10000 ( .C1(n8812), .C2(n8386), .A(n8385), .B(n8384), .ZN(n8387)
         );
  NAND3_X1 U10001 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(P2_U3237) );
  INV_X1 U10002 ( .A(n8390), .ZN(n8394) );
  OAI22_X1 U10003 ( .A1(n8392), .A2(n8391), .B1(n10074), .B2(n8425), .ZN(n8393) );
  AOI211_X1 U10004 ( .C1(n8395), .C2(n8420), .A(n8394), .B(n8393), .ZN(n8406)
         );
  OAI21_X1 U10005 ( .B1(n8400), .B2(n8397), .A(n8396), .ZN(n8399) );
  NAND2_X1 U10006 ( .A1(n8399), .A2(n8398), .ZN(n8405) );
  NOR3_X1 U10007 ( .A1(n8402), .A2(n8401), .A3(n8400), .ZN(n8403) );
  OAI21_X1 U10008 ( .B1(n8403), .B2(n8422), .A(n8448), .ZN(n8404) );
  NAND3_X1 U10009 ( .A1(n8406), .A2(n8405), .A3(n8404), .ZN(P2_U3241) );
  OAI22_X1 U10010 ( .A1(n8410), .A2(n10000), .B1(n8592), .B2(n9998), .ZN(n8570) );
  INV_X1 U10011 ( .A(n8574), .ZN(n8413) );
  OAI22_X1 U10012 ( .A1(n8413), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8411), .ZN(n8414) );
  AOI21_X1 U10013 ( .B1(n8570), .B2(n8415), .A(n8414), .ZN(n8416) );
  NAND2_X1 U10014 ( .A1(n8418), .A2(n8417), .ZN(n8430) );
  INV_X1 U10015 ( .A(n8754), .ZN(n8419) );
  AOI22_X1 U10016 ( .A1(n8420), .A2(n8419), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8424) );
  AOI22_X1 U10017 ( .A1(n8422), .A2(n8749), .B1(n8421), .B2(n8750), .ZN(n8423)
         );
  OAI211_X1 U10018 ( .C1(n8757), .C2(n8425), .A(n8424), .B(n8423), .ZN(n8429)
         );
  NOR3_X1 U10019 ( .A1(n8430), .A2(n8427), .A3(n8426), .ZN(n8428) );
  AOI211_X1 U10020 ( .C1(n8431), .C2(n8430), .A(n8429), .B(n8428), .ZN(n8432)
         );
  INV_X1 U10021 ( .A(n8432), .ZN(P2_U3243) );
  MUX2_X1 U10022 ( .A(n8535), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8449), .Z(
        P2_U3582) );
  MUX2_X1 U10023 ( .A(n8433), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8449), .Z(
        P2_U3581) );
  MUX2_X1 U10024 ( .A(n8537), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8449), .Z(
        P2_U3580) );
  MUX2_X1 U10025 ( .A(n8434), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8449), .Z(
        P2_U3579) );
  MUX2_X1 U10026 ( .A(n8435), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8449), .Z(
        P2_U3578) );
  MUX2_X1 U10027 ( .A(n8436), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8449), .Z(
        P2_U3577) );
  MUX2_X1 U10028 ( .A(n8613), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8449), .Z(
        P2_U3576) );
  MUX2_X1 U10029 ( .A(n8437), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8449), .Z(
        P2_U3575) );
  MUX2_X1 U10030 ( .A(n8654), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8449), .Z(
        P2_U3574) );
  MUX2_X1 U10031 ( .A(n8668), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8449), .Z(
        P2_U3573) );
  MUX2_X1 U10032 ( .A(n8686), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8449), .Z(
        P2_U3572) );
  INV_X1 U10033 ( .A(n8695), .ZN(n8667) );
  MUX2_X1 U10034 ( .A(n8667), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8449), .Z(
        P2_U3571) );
  MUX2_X1 U10035 ( .A(n8708), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8449), .Z(
        P2_U3570) );
  MUX2_X1 U10036 ( .A(n8438), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8449), .Z(
        P2_U3569) );
  MUX2_X1 U10037 ( .A(n8750), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8449), .Z(
        P2_U3568) );
  MUX2_X1 U10038 ( .A(n8439), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8449), .Z(
        P2_U3567) );
  MUX2_X1 U10039 ( .A(n8749), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8449), .Z(
        P2_U3566) );
  MUX2_X1 U10040 ( .A(n8440), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8449), .Z(
        P2_U3565) );
  MUX2_X1 U10041 ( .A(n8441), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8449), .Z(
        P2_U3564) );
  MUX2_X1 U10042 ( .A(n8442), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8449), .Z(
        P2_U3563) );
  MUX2_X1 U10043 ( .A(n8443), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8449), .Z(
        P2_U3562) );
  MUX2_X1 U10044 ( .A(n8444), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8449), .Z(
        P2_U3561) );
  MUX2_X1 U10045 ( .A(n8445), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8449), .Z(
        P2_U3560) );
  MUX2_X1 U10046 ( .A(n8446), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8449), .Z(
        P2_U3559) );
  MUX2_X1 U10047 ( .A(n8447), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8449), .Z(
        P2_U3558) );
  MUX2_X1 U10048 ( .A(n8448), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8449), .Z(
        P2_U3557) );
  MUX2_X1 U10049 ( .A(n10018), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8449), .Z(
        P2_U3556) );
  MUX2_X1 U10050 ( .A(n8450), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8449), .Z(
        P2_U3555) );
  MUX2_X1 U10051 ( .A(n10016), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8449), .Z(
        P2_U3554) );
  MUX2_X1 U10052 ( .A(n5682), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8449), .Z(
        P2_U3553) );
  MUX2_X1 U10053 ( .A(n8451), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8449), .Z(
        P2_U3552) );
  NAND2_X1 U10054 ( .A1(n8510), .A2(n8452), .ZN(n8462) );
  OAI211_X1 U10055 ( .C1(n8455), .C2(n8454), .A(n9979), .B(n8453), .ZN(n8461)
         );
  AOI22_X1 U10056 ( .A1(n9981), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8460) );
  OAI211_X1 U10057 ( .C1(n8458), .C2(n8457), .A(n9978), .B(n8456), .ZN(n8459)
         );
  NAND4_X1 U10058 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(
        P2_U3246) );
  INV_X1 U10059 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10477) );
  OAI21_X1 U10060 ( .B1(n8522), .B2(n10477), .A(n8463), .ZN(n8464) );
  AOI21_X1 U10061 ( .B1(n8510), .B2(n8465), .A(n8464), .ZN(n8474) );
  OAI211_X1 U10062 ( .C1(n8468), .C2(n8467), .A(n9978), .B(n8466), .ZN(n8473)
         );
  OAI211_X1 U10063 ( .C1(n8471), .C2(n8470), .A(n9979), .B(n8469), .ZN(n8472)
         );
  NAND3_X1 U10064 ( .A1(n8474), .A2(n8473), .A3(n8472), .ZN(P2_U3253) );
  OAI211_X1 U10065 ( .C1(n8477), .C2(n8476), .A(n8475), .B(n9979), .ZN(n8488)
         );
  INV_X1 U10066 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8480) );
  INV_X1 U10067 ( .A(n8478), .ZN(n8479) );
  OAI21_X1 U10068 ( .B1(n8522), .B2(n8480), .A(n8479), .ZN(n8481) );
  AOI21_X1 U10069 ( .B1(n8510), .B2(n8482), .A(n8481), .ZN(n8487) );
  OAI211_X1 U10070 ( .C1(n8485), .C2(n8484), .A(n9978), .B(n8483), .ZN(n8486)
         );
  NAND3_X1 U10071 ( .A1(n8488), .A2(n8487), .A3(n8486), .ZN(P2_U3254) );
  OAI211_X1 U10072 ( .C1(n8491), .C2(n8490), .A(n8489), .B(n9979), .ZN(n8501)
         );
  INV_X1 U10073 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8493) );
  OAI21_X1 U10074 ( .B1(n8522), .B2(n8493), .A(n8492), .ZN(n8494) );
  AOI21_X1 U10075 ( .B1(n8510), .B2(n8495), .A(n8494), .ZN(n8500) );
  OAI211_X1 U10076 ( .C1(n8498), .C2(n8497), .A(n8496), .B(n9978), .ZN(n8499)
         );
  NAND3_X1 U10077 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(P2_U3255) );
  OAI21_X1 U10078 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(n8505) );
  NAND2_X1 U10079 ( .A1(n8505), .A2(n9978), .ZN(n8517) );
  INV_X1 U10080 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8507) );
  OAI21_X1 U10081 ( .B1(n8522), .B2(n8507), .A(n8506), .ZN(n8508) );
  AOI21_X1 U10082 ( .B1(n8510), .B2(n8509), .A(n8508), .ZN(n8516) );
  AOI21_X1 U10083 ( .B1(n8513), .B2(n8512), .A(n8511), .ZN(n8514) );
  NAND2_X1 U10084 ( .A1(n9979), .A2(n8514), .ZN(n8515) );
  NAND3_X1 U10085 ( .A1(n8517), .A2(n8516), .A3(n8515), .ZN(P2_U3261) );
  OAI21_X1 U10086 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8532) );
  INV_X1 U10087 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10473) );
  OAI21_X1 U10088 ( .B1(n8522), .B2(n10473), .A(n8521), .ZN(n8523) );
  INV_X1 U10089 ( .A(n8523), .ZN(n8529) );
  OAI21_X1 U10090 ( .B1(n8526), .B2(n8525), .A(n8524), .ZN(n8527) );
  NAND2_X1 U10091 ( .A1(n9978), .A2(n8527), .ZN(n8528) );
  OAI211_X1 U10092 ( .C1(n9983), .C2(n8530), .A(n8529), .B(n8528), .ZN(n8531)
         );
  AOI21_X1 U10093 ( .B1(n8532), .B2(n9979), .A(n8531), .ZN(n8533) );
  INV_X1 U10094 ( .A(n8533), .ZN(P2_U3263) );
  XNOR2_X1 U10095 ( .A(n8534), .B(n8776), .ZN(n8540) );
  AOI22_X1 U10096 ( .A1(n8537), .A2(n10015), .B1(n8536), .B2(n8535), .ZN(n8538) );
  AOI21_X2 U10097 ( .B1(n8540), .B2(n10020), .A(n8539), .ZN(n8785) );
  AND2_X1 U10098 ( .A1(n4943), .A2(n8543), .ZN(n8775) );
  INV_X1 U10099 ( .A(n8775), .ZN(n8544) );
  NAND2_X1 U10100 ( .A1(n8783), .A2(n8544), .ZN(n8545) );
  XNOR2_X1 U10101 ( .A(n8545), .B(n8776), .ZN(n8546) );
  NAND2_X1 U10102 ( .A1(n8546), .A2(n10034), .ZN(n8555) );
  INV_X1 U10103 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8547) );
  OAI22_X1 U10104 ( .A1(n8548), .A2(n10026), .B1(n8547), .B2(n10027), .ZN(
        n8553) );
  NOR2_X1 U10105 ( .A1(n8779), .A2(n8551), .ZN(n8552) );
  AOI211_X1 U10106 ( .C1(n8756), .C2(n8777), .A(n8553), .B(n8552), .ZN(n8554)
         );
  OAI211_X1 U10107 ( .C1(n8785), .C2(n10036), .A(n8555), .B(n8554), .ZN(
        P2_U3267) );
  NAND2_X1 U10108 ( .A1(n8556), .A2(n10034), .ZN(n8562) );
  AOI22_X1 U10109 ( .A1(n8557), .A2(n10002), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n8766), .ZN(n8558) );
  OAI21_X1 U10110 ( .B1(n4943), .B2(n10031), .A(n8558), .ZN(n8559) );
  AOI21_X1 U10111 ( .B1(n8560), .B2(n10029), .A(n8559), .ZN(n8561) );
  OAI211_X1 U10112 ( .C1(n8563), .C2(n8766), .A(n8562), .B(n8561), .ZN(
        P2_U3268) );
  XNOR2_X1 U10113 ( .A(n8564), .B(n8568), .ZN(n8796) );
  NOR2_X1 U10114 ( .A1(n8565), .A2(n10031), .ZN(n8578) );
  AND2_X1 U10115 ( .A1(n8581), .A2(n8566), .ZN(n8569) );
  OAI21_X1 U10116 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8571) );
  INV_X1 U10117 ( .A(n8572), .ZN(n8573) );
  AOI211_X1 U10118 ( .C1(n8793), .C2(n8573), .A(n10113), .B(n5722), .ZN(n8792)
         );
  AOI22_X1 U10119 ( .A1(n8792), .A2(n8575), .B1(n10002), .B2(n8574), .ZN(n8576) );
  AOI21_X1 U10120 ( .B1(n8795), .B2(n8576), .A(n8766), .ZN(n8577) );
  OAI21_X1 U10121 ( .B1(n8796), .B2(n8763), .A(n8579), .ZN(P2_U3270) );
  XNOR2_X1 U10122 ( .A(n8580), .B(n4433), .ZN(n8800) );
  AOI22_X1 U10123 ( .A1(n8799), .A2(n8756), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8766), .ZN(n8590) );
  OAI211_X1 U10124 ( .C1(n4433), .C2(n8582), .A(n8581), .B(n10020), .ZN(n8584)
         );
  XNOR2_X1 U10125 ( .A(n8799), .B(n8601), .ZN(n8585) );
  NOR2_X1 U10126 ( .A1(n8585), .A2(n10113), .ZN(n8798) );
  INV_X1 U10127 ( .A(n8798), .ZN(n8587) );
  OAI22_X1 U10128 ( .A1(n8587), .A2(n5619), .B1(n10026), .B2(n8586), .ZN(n8588) );
  OAI21_X1 U10129 ( .B1(n8797), .B2(n8588), .A(n10027), .ZN(n8589) );
  OAI211_X1 U10130 ( .C1(n8800), .C2(n8763), .A(n8590), .B(n8589), .ZN(
        P2_U3271) );
  INV_X1 U10131 ( .A(n8599), .ZN(n8591) );
  AOI21_X1 U10132 ( .B1(n4429), .B2(n8591), .A(n9995), .ZN(n8595) );
  OAI22_X1 U10133 ( .A1(n8592), .A2(n10000), .B1(n8639), .B2(n9998), .ZN(n8593) );
  AOI21_X1 U10134 ( .B1(n8595), .B2(n8594), .A(n8593), .ZN(n8804) );
  INV_X1 U10135 ( .A(n8596), .ZN(n8597) );
  AOI21_X1 U10136 ( .B1(n8599), .B2(n8598), .A(n8597), .ZN(n8805) );
  INV_X1 U10137 ( .A(n8805), .ZN(n8607) );
  INV_X1 U10138 ( .A(n8801), .ZN(n8605) );
  NAND2_X1 U10139 ( .A1(n8801), .A2(n8618), .ZN(n8600) );
  AND2_X1 U10140 ( .A1(n8601), .A2(n8600), .ZN(n8802) );
  NAND2_X1 U10141 ( .A1(n8802), .A2(n10029), .ZN(n8604) );
  AOI22_X1 U10142 ( .A1(n10036), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8602), 
        .B2(n10002), .ZN(n8603) );
  OAI211_X1 U10143 ( .C1(n8605), .C2(n10031), .A(n8604), .B(n8603), .ZN(n8606)
         );
  AOI21_X1 U10144 ( .B1(n8607), .B2(n10034), .A(n8606), .ZN(n8608) );
  OAI21_X1 U10145 ( .B1(n10036), .B2(n8804), .A(n8608), .ZN(P2_U3272) );
  INV_X1 U10146 ( .A(n8609), .ZN(n8612) );
  OAI21_X1 U10147 ( .B1(n8612), .B2(n5975), .A(n8611), .ZN(n8614) );
  AOI222_X1 U10148 ( .A1(n10020), .A2(n8614), .B1(n8613), .B2(n10017), .C1(
        n8654), .C2(n10015), .ZN(n8810) );
  OR2_X1 U10149 ( .A1(n8616), .A2(n8615), .ZN(n8806) );
  NAND3_X1 U10150 ( .A1(n8806), .A2(n8617), .A3(n10034), .ZN(n8626) );
  INV_X1 U10151 ( .A(n8618), .ZN(n8619) );
  AOI21_X1 U10152 ( .B1(n8807), .B2(n8628), .A(n8619), .ZN(n8808) );
  NOR2_X1 U10153 ( .A1(n8620), .A2(n10031), .ZN(n8624) );
  INV_X1 U10154 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8622) );
  OAI22_X1 U10155 ( .A1(n10027), .A2(n8622), .B1(n8621), .B2(n10026), .ZN(
        n8623) );
  AOI211_X1 U10156 ( .C1(n8808), .C2(n10029), .A(n8624), .B(n8623), .ZN(n8625)
         );
  OAI211_X1 U10157 ( .C1(n10036), .C2(n8810), .A(n8626), .B(n8625), .ZN(
        P2_U3273) );
  XOR2_X1 U10158 ( .A(n8627), .B(n8637), .Z(n8816) );
  INV_X1 U10159 ( .A(n8647), .ZN(n8630) );
  INV_X1 U10160 ( .A(n8628), .ZN(n8629) );
  AOI21_X1 U10161 ( .B1(n8812), .B2(n8630), .A(n8629), .ZN(n8813) );
  INV_X1 U10162 ( .A(n8631), .ZN(n8632) );
  AOI22_X1 U10163 ( .A1(n10036), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8632), 
        .B2(n10002), .ZN(n8633) );
  OAI21_X1 U10164 ( .B1(n8634), .B2(n10031), .A(n8633), .ZN(n8644) );
  AOI21_X1 U10165 ( .B1(n8636), .B2(n8637), .A(n9995), .ZN(n8642) );
  OAI22_X1 U10166 ( .A1(n8639), .A2(n10000), .B1(n8638), .B2(n9998), .ZN(n8640) );
  AOI21_X1 U10167 ( .B1(n8642), .B2(n8641), .A(n8640), .ZN(n8815) );
  NOR2_X1 U10168 ( .A1(n8815), .A2(n8766), .ZN(n8643) );
  AOI211_X1 U10169 ( .C1(n8813), .C2(n10029), .A(n8644), .B(n8643), .ZN(n8645)
         );
  OAI21_X1 U10170 ( .B1(n8816), .B2(n8763), .A(n8645), .ZN(P2_U3274) );
  XNOR2_X1 U10171 ( .A(n8646), .B(n8653), .ZN(n8821) );
  AOI21_X1 U10172 ( .B1(n8817), .B2(n8661), .A(n8647), .ZN(n8818) );
  AOI22_X1 U10173 ( .A1(n10036), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8648), 
        .B2(n10002), .ZN(n8649) );
  OAI21_X1 U10174 ( .B1(n8650), .B2(n10031), .A(n8649), .ZN(n8657) );
  XNOR2_X1 U10175 ( .A(n8652), .B(n8653), .ZN(n8655) );
  AOI222_X1 U10176 ( .A1(n10020), .A2(n8655), .B1(n8654), .B2(n10017), .C1(
        n8686), .C2(n10015), .ZN(n8820) );
  NOR2_X1 U10177 ( .A1(n8820), .A2(n8766), .ZN(n8656) );
  AOI211_X1 U10178 ( .C1(n8818), .C2(n10029), .A(n8657), .B(n8656), .ZN(n8658)
         );
  OAI21_X1 U10179 ( .B1(n8821), .B2(n8763), .A(n8658), .ZN(P2_U3275) );
  XNOR2_X1 U10180 ( .A(n8659), .B(n8665), .ZN(n8826) );
  AOI21_X1 U10181 ( .B1(n8822), .B2(n8674), .A(n5721), .ZN(n8823) );
  INV_X1 U10182 ( .A(n8822), .ZN(n8664) );
  AOI22_X1 U10183 ( .A1(n10036), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8662), 
        .B2(n10002), .ZN(n8663) );
  OAI21_X1 U10184 ( .B1(n8664), .B2(n10031), .A(n8663), .ZN(n8671) );
  XOR2_X1 U10185 ( .A(n8666), .B(n8665), .Z(n8669) );
  AOI222_X1 U10186 ( .A1(n10020), .A2(n8669), .B1(n8668), .B2(n10017), .C1(
        n8667), .C2(n10015), .ZN(n8825) );
  NOR2_X1 U10187 ( .A1(n8825), .A2(n8766), .ZN(n8670) );
  AOI211_X1 U10188 ( .C1(n8823), .C2(n10029), .A(n8671), .B(n8670), .ZN(n8672)
         );
  OAI21_X1 U10189 ( .B1(n8763), .B2(n8826), .A(n8672), .ZN(P2_U3276) );
  XNOR2_X1 U10190 ( .A(n8673), .B(n8684), .ZN(n8831) );
  INV_X1 U10191 ( .A(n8696), .ZN(n8676) );
  INV_X1 U10192 ( .A(n8674), .ZN(n8675) );
  AOI211_X1 U10193 ( .C1(n8828), .C2(n8676), .A(n10113), .B(n8675), .ZN(n8827)
         );
  INV_X1 U10194 ( .A(n8677), .ZN(n8678) );
  AOI22_X1 U10195 ( .A1(n10036), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8678), 
        .B2(n10002), .ZN(n8679) );
  OAI21_X1 U10196 ( .B1(n8680), .B2(n10031), .A(n8679), .ZN(n8689) );
  AND2_X1 U10197 ( .A1(n8682), .A2(n8681), .ZN(n8685) );
  OAI21_X1 U10198 ( .B1(n8685), .B2(n8684), .A(n8683), .ZN(n8687) );
  AOI222_X1 U10199 ( .A1(n10020), .A2(n8687), .B1(n8686), .B2(n10017), .C1(
        n8708), .C2(n10015), .ZN(n8830) );
  NOR2_X1 U10200 ( .A1(n8830), .A2(n10036), .ZN(n8688) );
  AOI211_X1 U10201 ( .C1(n8827), .C2(n8720), .A(n8689), .B(n8688), .ZN(n8690)
         );
  OAI21_X1 U10202 ( .B1(n8763), .B2(n8831), .A(n8690), .ZN(P2_U3277) );
  XNOR2_X1 U10203 ( .A(n8691), .B(n8692), .ZN(n8836) );
  XNOR2_X1 U10204 ( .A(n8693), .B(n8692), .ZN(n8694) );
  OAI222_X1 U10205 ( .A1(n10000), .A2(n8695), .B1(n9998), .B2(n8732), .C1(
        n9995), .C2(n8694), .ZN(n8832) );
  AOI211_X1 U10206 ( .C1(n8834), .C2(n4507), .A(n10113), .B(n8696), .ZN(n8833)
         );
  NAND2_X1 U10207 ( .A1(n8833), .A2(n8720), .ZN(n8699) );
  AOI22_X1 U10208 ( .A1(n8766), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8697), .B2(
        n10002), .ZN(n8698) );
  OAI211_X1 U10209 ( .C1(n8700), .C2(n10031), .A(n8699), .B(n8698), .ZN(n8701)
         );
  AOI21_X1 U10210 ( .B1(n8832), .B2(n10027), .A(n8701), .ZN(n8702) );
  OAI21_X1 U10211 ( .B1(n8836), .B2(n8763), .A(n8702), .ZN(P2_U3278) );
  NAND2_X1 U10212 ( .A1(n8704), .A2(n8705), .ZN(n8707) );
  XNOR2_X1 U10213 ( .A(n8707), .B(n8706), .ZN(n8709) );
  AOI222_X1 U10214 ( .A1(n10020), .A2(n8709), .B1(n8708), .B2(n10017), .C1(
        n8750), .C2(n10015), .ZN(n8840) );
  OAI21_X1 U10215 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8713) );
  INV_X1 U10216 ( .A(n8713), .ZN(n8841) );
  NAND2_X1 U10217 ( .A1(n10036), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8714) );
  OAI21_X1 U10218 ( .B1(n10026), .B2(n8715), .A(n8714), .ZN(n8716) );
  AOI21_X1 U10219 ( .B1(n8838), .B2(n8756), .A(n8716), .ZN(n8722) );
  NAND2_X1 U10220 ( .A1(n8738), .A2(n8838), .ZN(n8717) );
  NAND2_X1 U10221 ( .A1(n8717), .A2(n10097), .ZN(n8718) );
  NOR2_X1 U10222 ( .A1(n8719), .A2(n8718), .ZN(n8837) );
  NAND2_X1 U10223 ( .A1(n8837), .A2(n8720), .ZN(n8721) );
  OAI211_X1 U10224 ( .C1(n8841), .C2(n8763), .A(n8722), .B(n8721), .ZN(n8723)
         );
  INV_X1 U10225 ( .A(n8723), .ZN(n8724) );
  OAI21_X1 U10226 ( .B1(n10036), .B2(n8840), .A(n8724), .ZN(P2_U3279) );
  NOR2_X1 U10227 ( .A1(n8726), .A2(n8729), .ZN(n8727) );
  NAND2_X1 U10228 ( .A1(n8728), .A2(n8729), .ZN(n8730) );
  NAND2_X1 U10229 ( .A1(n8704), .A2(n8730), .ZN(n8734) );
  OAI22_X1 U10230 ( .A1(n8732), .A2(n10000), .B1(n8731), .B2(n9998), .ZN(n8733) );
  AOI21_X1 U10231 ( .B1(n8734), .B2(n10020), .A(n8733), .ZN(n8735) );
  OAI21_X1 U10232 ( .B1(n8845), .B2(n8736), .A(n8735), .ZN(n8847) );
  NAND2_X1 U10233 ( .A1(n8847), .A2(n10027), .ZN(n8744) );
  NAND2_X1 U10234 ( .A1(n8758), .A2(n8757), .ZN(n8760) );
  NAND2_X1 U10235 ( .A1(n8760), .A2(n8842), .ZN(n8737) );
  AND2_X1 U10236 ( .A1(n8738), .A2(n8737), .ZN(n8843) );
  AOI22_X1 U10237 ( .A1(n8766), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8739), .B2(
        n10002), .ZN(n8740) );
  OAI21_X1 U10238 ( .B1(n8741), .B2(n10031), .A(n8740), .ZN(n8742) );
  AOI21_X1 U10239 ( .B1(n8843), .B2(n10029), .A(n8742), .ZN(n8743) );
  OAI211_X1 U10240 ( .C1(n8845), .C2(n10006), .A(n8744), .B(n8743), .ZN(
        P2_U3280) );
  NAND2_X1 U10241 ( .A1(n8746), .A2(n8745), .ZN(n8748) );
  XNOR2_X1 U10242 ( .A(n8748), .B(n8747), .ZN(n8751) );
  AOI222_X1 U10243 ( .A1(n10020), .A2(n8751), .B1(n8750), .B2(n10017), .C1(
        n8749), .C2(n10015), .ZN(n8850) );
  XNOR2_X1 U10244 ( .A(n8752), .B(n4718), .ZN(n8851) );
  NAND2_X1 U10245 ( .A1(n10036), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8753) );
  OAI21_X1 U10246 ( .B1(n10026), .B2(n8754), .A(n8753), .ZN(n8755) );
  AOI21_X1 U10247 ( .B1(n5704), .B2(n8756), .A(n8755), .ZN(n8762) );
  OR2_X1 U10248 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  AND2_X1 U10249 ( .A1(n8760), .A2(n8759), .ZN(n8848) );
  NAND2_X1 U10250 ( .A1(n8848), .A2(n10029), .ZN(n8761) );
  OAI211_X1 U10251 ( .C1(n8851), .C2(n8763), .A(n8762), .B(n8761), .ZN(n8764)
         );
  INV_X1 U10252 ( .A(n8764), .ZN(n8765) );
  OAI21_X1 U10253 ( .B1(n8850), .B2(n8766), .A(n8765), .ZN(P2_U3281) );
  NAND2_X1 U10254 ( .A1(n5818), .A2(n10096), .ZN(n8768) );
  NAND2_X1 U10255 ( .A1(n8769), .A2(n5057), .ZN(n8869) );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8869), .S(n10142), .Z(
        P2_U3551) );
  NAND2_X1 U10257 ( .A1(n8770), .A2(n10097), .ZN(n8772) );
  OAI211_X1 U10258 ( .C1(n8773), .C2(n10111), .A(n8772), .B(n8771), .ZN(n8870)
         );
  MUX2_X1 U10259 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8870), .S(n10142), .Z(
        P2_U3550) );
  NAND2_X1 U10260 ( .A1(n8776), .A2(n10117), .ZN(n8774) );
  NOR3_X1 U10261 ( .A1(n8776), .A2(n10085), .A3(n8775), .ZN(n8782) );
  NAND3_X1 U10262 ( .A1(n8776), .A2(n8775), .A3(n10117), .ZN(n8780) );
  NAND2_X1 U10263 ( .A1(n8777), .A2(n10096), .ZN(n8778) );
  NAND3_X1 U10264 ( .A1(n8786), .A2(n8785), .A3(n8784), .ZN(n8871) );
  MUX2_X1 U10265 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8871), .S(n10142), .Z(
        P2_U3549) );
  OAI211_X1 U10266 ( .C1(n8791), .C2(n10085), .A(n8790), .B(n8789), .ZN(n8872)
         );
  MUX2_X1 U10267 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8872), .S(n10142), .Z(
        P2_U3547) );
  AOI21_X1 U10268 ( .B1(n10096), .B2(n8793), .A(n8792), .ZN(n8794) );
  OAI211_X1 U10269 ( .C1(n8796), .C2(n10085), .A(n8795), .B(n8794), .ZN(n8873)
         );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8873), .S(n10142), .Z(
        P2_U3546) );
  AOI22_X1 U10271 ( .A1(n8802), .A2(n10097), .B1(n10096), .B2(n8801), .ZN(
        n8803) );
  OAI211_X1 U10272 ( .C1(n8805), .C2(n10085), .A(n8804), .B(n8803), .ZN(n8875)
         );
  MUX2_X1 U10273 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8875), .S(n10142), .Z(
        P2_U3544) );
  NAND3_X1 U10274 ( .A1(n8806), .A2(n8617), .A3(n10117), .ZN(n8811) );
  AOI22_X1 U10275 ( .A1(n8808), .A2(n10097), .B1(n10096), .B2(n8807), .ZN(
        n8809) );
  NAND3_X1 U10276 ( .A1(n8811), .A2(n8810), .A3(n8809), .ZN(n8876) );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8876), .S(n10142), .Z(
        P2_U3543) );
  AOI22_X1 U10278 ( .A1(n8813), .A2(n10097), .B1(n10096), .B2(n8812), .ZN(
        n8814) );
  OAI211_X1 U10279 ( .C1(n8816), .C2(n10085), .A(n8815), .B(n8814), .ZN(n8877)
         );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8877), .S(n10142), .Z(
        P2_U3542) );
  AOI22_X1 U10281 ( .A1(n8818), .A2(n10097), .B1(n10096), .B2(n8817), .ZN(
        n8819) );
  OAI211_X1 U10282 ( .C1(n8821), .C2(n10085), .A(n8820), .B(n8819), .ZN(n8878)
         );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8878), .S(n10142), .Z(
        P2_U3541) );
  AOI22_X1 U10284 ( .A1(n8823), .A2(n10097), .B1(n10096), .B2(n8822), .ZN(
        n8824) );
  OAI211_X1 U10285 ( .C1(n8826), .C2(n10085), .A(n8825), .B(n8824), .ZN(n8879)
         );
  MUX2_X1 U10286 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8879), .S(n10142), .Z(
        P2_U3540) );
  AOI21_X1 U10287 ( .B1(n10096), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI211_X1 U10288 ( .C1(n8831), .C2(n10085), .A(n8830), .B(n8829), .ZN(n8880)
         );
  MUX2_X1 U10289 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8880), .S(n10142), .Z(
        P2_U3539) );
  AOI211_X1 U10290 ( .C1(n10096), .C2(n8834), .A(n8833), .B(n8832), .ZN(n8835)
         );
  OAI21_X1 U10291 ( .B1(n10085), .B2(n8836), .A(n8835), .ZN(n8881) );
  MUX2_X1 U10292 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8881), .S(n10142), .Z(
        P2_U3538) );
  AOI21_X1 U10293 ( .B1(n10096), .B2(n8838), .A(n8837), .ZN(n8839) );
  OAI211_X1 U10294 ( .C1(n8841), .C2(n10085), .A(n8840), .B(n8839), .ZN(n8882)
         );
  MUX2_X1 U10295 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8882), .S(n10142), .Z(
        P2_U3537) );
  AOI22_X1 U10296 ( .A1(n8843), .A2(n10097), .B1(n10096), .B2(n8842), .ZN(
        n8844) );
  OAI21_X1 U10297 ( .B1(n8845), .B2(n10102), .A(n8844), .ZN(n8846) );
  OR2_X1 U10298 ( .A1(n8847), .A2(n8846), .ZN(n8883) );
  MUX2_X1 U10299 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8883), .S(n10142), .Z(
        P2_U3536) );
  AOI22_X1 U10300 ( .A1(n8848), .A2(n10097), .B1(n10096), .B2(n5704), .ZN(
        n8849) );
  OAI211_X1 U10301 ( .C1(n10085), .C2(n8851), .A(n8850), .B(n8849), .ZN(n8884)
         );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8884), .S(n10142), .Z(
        P2_U3535) );
  INV_X1 U10303 ( .A(n8852), .ZN(n8857) );
  AOI21_X1 U10304 ( .B1(n10096), .B2(n8854), .A(n8853), .ZN(n8855) );
  OAI211_X1 U10305 ( .C1(n10085), .C2(n8857), .A(n8856), .B(n8855), .ZN(n8885)
         );
  MUX2_X1 U10306 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8885), .S(n10142), .Z(
        P2_U3534) );
  AOI22_X1 U10307 ( .A1(n8859), .A2(n10097), .B1(n10096), .B2(n8858), .ZN(
        n8860) );
  OAI211_X1 U10308 ( .C1(n10102), .C2(n8862), .A(n8861), .B(n8860), .ZN(n8886)
         );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8886), .S(n10142), .Z(
        P2_U3533) );
  AND2_X1 U10310 ( .A1(n8863), .A2(n10117), .ZN(n8867) );
  OAI22_X1 U10311 ( .A1(n8865), .A2(n10113), .B1(n8864), .B2(n10111), .ZN(
        n8866) );
  MUX2_X1 U10312 ( .A(n8887), .B(P2_REG1_REG_12__SCAN_IN), .S(n10139), .Z(
        P2_U3532) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8869), .S(n10121), .Z(
        P2_U3519) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8870), .S(n10121), .Z(
        P2_U3518) );
  MUX2_X1 U10315 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8871), .S(n10121), .Z(
        P2_U3517) );
  MUX2_X1 U10316 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8872), .S(n10121), .Z(
        P2_U3515) );
  MUX2_X1 U10317 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8873), .S(n10121), .Z(
        P2_U3514) );
  MUX2_X1 U10318 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8875), .S(n10121), .Z(
        P2_U3512) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8876), .S(n10121), .Z(
        P2_U3511) );
  MUX2_X1 U10320 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8877), .S(n10121), .Z(
        P2_U3510) );
  MUX2_X1 U10321 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8878), .S(n10121), .Z(
        P2_U3509) );
  MUX2_X1 U10322 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8879), .S(n10121), .Z(
        P2_U3508) );
  MUX2_X1 U10323 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8880), .S(n10121), .Z(
        P2_U3507) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8881), .S(n10121), .Z(
        P2_U3505) );
  MUX2_X1 U10325 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8882), .S(n10121), .Z(
        P2_U3502) );
  MUX2_X1 U10326 ( .A(n8883), .B(P2_REG0_REG_16__SCAN_IN), .S(n10119), .Z(
        P2_U3499) );
  MUX2_X1 U10327 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8884), .S(n10121), .Z(
        P2_U3496) );
  MUX2_X1 U10328 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8885), .S(n10121), .Z(
        P2_U3493) );
  MUX2_X1 U10329 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8886), .S(n10121), .Z(
        P2_U3490) );
  MUX2_X1 U10330 ( .A(n8887), .B(P2_REG0_REG_12__SCAN_IN), .S(n10119), .Z(
        P2_U3487) );
  INV_X1 U10331 ( .A(n9049), .ZN(n9830) );
  INV_X1 U10332 ( .A(n8888), .ZN(n8891) );
  NOR4_X1 U10333 ( .A1(n8891), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8890), .A4(
        P2_U3152), .ZN(n8892) );
  AOI21_X1 U10334 ( .B1(n8903), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8892), .ZN(
        n8893) );
  OAI21_X1 U10335 ( .B1(n9830), .B2(n8906), .A(n8893), .ZN(P2_U3327) );
  AOI22_X1 U10336 ( .A1(n8894), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8903), .ZN(n8895) );
  OAI21_X1 U10337 ( .B1(n8896), .B2(n8906), .A(n8895), .ZN(P2_U3328) );
  INV_X1 U10338 ( .A(n9063), .ZN(n9831) );
  AOI22_X1 U10339 ( .A1(n8897), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8903), .ZN(n8898) );
  OAI21_X1 U10340 ( .B1(n9831), .B2(n8906), .A(n8898), .ZN(P2_U3329) );
  INV_X1 U10341 ( .A(n8899), .ZN(n9834) );
  AOI22_X1 U10342 ( .A1(n8900), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8903), .ZN(n8901) );
  OAI21_X1 U10343 ( .B1(n9834), .B2(n8906), .A(n8901), .ZN(P2_U3331) );
  INV_X1 U10344 ( .A(n8902), .ZN(n9839) );
  AOI22_X1 U10345 ( .A1(n8904), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8903), .ZN(n8905) );
  OAI21_X1 U10346 ( .B1(n9839), .B2(n8906), .A(n8905), .ZN(P2_U3332) );
  MUX2_X1 U10347 ( .A(n8907), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10348 ( .A(n8908), .ZN(n8911) );
  INV_X1 U10349 ( .A(n8909), .ZN(n8910) );
  OAI21_X1 U10350 ( .B1(n8913), .B2(n8912), .A(n8986), .ZN(n8918) );
  AOI22_X1 U10351 ( .A1(n8914), .A2(n9039), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8915) );
  OAI21_X1 U10352 ( .B1(n8964), .B2(n9042), .A(n8915), .ZN(n8916) );
  AOI21_X1 U10353 ( .B1(n9467), .B2(n9040), .A(n8916), .ZN(n8917) );
  OAI211_X1 U10354 ( .C1(n8919), .C2(n8996), .A(n8918), .B(n8917), .ZN(
        P1_U3212) );
  INV_X1 U10355 ( .A(n8920), .ZN(n8925) );
  AOI21_X1 U10356 ( .B1(n8922), .B2(n8924), .A(n8921), .ZN(n8923) );
  AOI21_X1 U10357 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8930) );
  OAI22_X1 U10358 ( .A1(n8926), .A2(n9042), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10261), .ZN(n8928) );
  OAI22_X1 U10359 ( .A1(n8963), .A2(n9011), .B1(n9013), .B2(n9529), .ZN(n8927)
         );
  AOI211_X1 U10360 ( .C1(n9725), .C2(n9045), .A(n8928), .B(n8927), .ZN(n8929)
         );
  OAI21_X1 U10361 ( .B1(n8930), .B2(n9047), .A(n8929), .ZN(P1_U3214) );
  INV_X1 U10362 ( .A(n8940), .ZN(n8939) );
  XNOR2_X1 U10363 ( .A(n8939), .B(n8942), .ZN(n8932) );
  XNOR2_X1 U10364 ( .A(n8931), .B(n8932), .ZN(n8938) );
  NAND2_X1 U10365 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9446) );
  OAI21_X1 U10366 ( .B1(n9042), .B2(n8933), .A(n9446), .ZN(n8936) );
  OAI22_X1 U10367 ( .A1(n9011), .A2(n8934), .B1(n9013), .B2(n9589), .ZN(n8935)
         );
  AOI211_X1 U10368 ( .C1(n9745), .C2(n9045), .A(n8936), .B(n8935), .ZN(n8937)
         );
  OAI21_X1 U10369 ( .B1(n8938), .B2(n9047), .A(n8937), .ZN(P1_U3217) );
  NOR2_X1 U10370 ( .A1(n8931), .A2(n8939), .ZN(n8943) );
  INV_X1 U10371 ( .A(n8931), .ZN(n8941) );
  OAI22_X1 U10372 ( .A1(n8943), .A2(n8942), .B1(n8941), .B2(n8940), .ZN(n8999)
         );
  NAND2_X1 U10373 ( .A1(n8944), .A2(n8945), .ZN(n9000) );
  NOR2_X1 U10374 ( .A1(n8999), .A2(n9000), .ZN(n8998) );
  INV_X1 U10375 ( .A(n8945), .ZN(n8947) );
  NOR3_X1 U10376 ( .A1(n8998), .A2(n8947), .A3(n8946), .ZN(n8950) );
  INV_X1 U10377 ( .A(n8948), .ZN(n8949) );
  OAI21_X1 U10378 ( .B1(n8950), .B2(n8949), .A(n8986), .ZN(n8955) );
  AOI22_X1 U10379 ( .A1(n9564), .A2(n9040), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8954) );
  AOI22_X1 U10380 ( .A1(n8951), .A2(n9596), .B1(n9558), .B2(n9039), .ZN(n8953)
         );
  NAND2_X1 U10381 ( .A1(n9736), .A2(n9045), .ZN(n8952) );
  NAND4_X1 U10382 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(
        P1_U3221) );
  INV_X1 U10383 ( .A(n8956), .ZN(n8958) );
  INV_X1 U10384 ( .A(n8960), .ZN(n8961) );
  OAI21_X1 U10385 ( .B1(n8962), .B2(n8961), .A(n8986), .ZN(n8968) );
  OAI22_X1 U10386 ( .A1(n8963), .A2(n9042), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10432), .ZN(n8966) );
  NOR2_X1 U10387 ( .A1(n8964), .A2(n9011), .ZN(n8965) );
  AOI211_X1 U10388 ( .C1(n9501), .C2(n9039), .A(n8966), .B(n8965), .ZN(n8967)
         );
  NOR2_X1 U10389 ( .A1(n7914), .A2(n8969), .ZN(n8970) );
  NAND2_X1 U10390 ( .A1(n7914), .A2(n8969), .ZN(n8972) );
  OAI211_X1 U10391 ( .C1(n8970), .C2(n8973), .A(n8971), .B(n8972), .ZN(n9034)
         );
  AOI211_X1 U10392 ( .C1(n8973), .C2(n8972), .A(n8971), .B(n8970), .ZN(n9036)
         );
  AOI21_X1 U10393 ( .B1(n9037), .B2(n9034), .A(n9036), .ZN(n8974) );
  AND2_X1 U10394 ( .A1(n8974), .A2(n8975), .ZN(n8984) );
  AOI21_X1 U10395 ( .B1(n8975), .B2(n8981), .A(n8974), .ZN(n8976) );
  AOI21_X1 U10396 ( .B1(n8984), .B2(n8981), .A(n8976), .ZN(n8980) );
  NAND2_X1 U10397 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9398) );
  OAI21_X1 U10398 ( .B1(n9011), .B2(n9632), .A(n9398), .ZN(n8978) );
  OAI22_X1 U10399 ( .A1(n9013), .A2(n9638), .B1(n9042), .B2(n9630), .ZN(n8977)
         );
  AOI211_X1 U10400 ( .C1(n9764), .C2(n9045), .A(n8978), .B(n8977), .ZN(n8979)
         );
  OAI21_X1 U10401 ( .B1(n8980), .B2(n9047), .A(n8979), .ZN(P1_U3224) );
  INV_X1 U10402 ( .A(n8981), .ZN(n8983) );
  NOR3_X1 U10403 ( .A1(n8984), .A2(n8983), .A3(n8982), .ZN(n8988) );
  INV_X1 U10404 ( .A(n8985), .ZN(n8987) );
  OAI21_X1 U10405 ( .B1(n8988), .B2(n8987), .A(n8986), .ZN(n8995) );
  NOR2_X1 U10406 ( .A1(n8989), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9408) );
  INV_X1 U10407 ( .A(n8990), .ZN(n8992) );
  OAI22_X1 U10408 ( .A1(n9013), .A2(n8992), .B1(n9042), .B2(n8991), .ZN(n8993)
         );
  AOI211_X1 U10409 ( .C1(n9040), .C2(n9595), .A(n9408), .B(n8993), .ZN(n8994)
         );
  OAI211_X1 U10410 ( .C1(n8997), .C2(n8996), .A(n8995), .B(n8994), .ZN(
        P1_U3226) );
  AOI21_X1 U10411 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9005) );
  OAI22_X1 U10412 ( .A1(n9042), .A2(n9001), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10321), .ZN(n9003) );
  OAI22_X1 U10413 ( .A1(n9011), .A2(n9349), .B1(n9013), .B2(n9571), .ZN(n9002)
         );
  AOI211_X1 U10414 ( .C1(n9740), .C2(n9045), .A(n9003), .B(n9002), .ZN(n9004)
         );
  OAI21_X1 U10415 ( .B1(n9005), .B2(n9047), .A(n9004), .ZN(P1_U3231) );
  NAND2_X1 U10416 ( .A1(n9006), .A2(n9007), .ZN(n9009) );
  XNOR2_X1 U10417 ( .A(n9009), .B(n9008), .ZN(n9017) );
  OAI22_X1 U10418 ( .A1(n9517), .A2(n9011), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9010), .ZN(n9015) );
  INV_X1 U10419 ( .A(n9543), .ZN(n9012) );
  OAI22_X1 U10420 ( .A1(n9349), .A2(n9042), .B1(n9013), .B2(n9012), .ZN(n9014)
         );
  AOI211_X1 U10421 ( .C1(n9731), .C2(n9045), .A(n9015), .B(n9014), .ZN(n9016)
         );
  OAI21_X1 U10422 ( .B1(n9017), .B2(n9047), .A(n9016), .ZN(P1_U3233) );
  NAND2_X1 U10423 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  XOR2_X1 U10424 ( .A(n9021), .B(n9020), .Z(n9026) );
  INV_X1 U10425 ( .A(n9613), .ZN(n9022) );
  AOI22_X1 U10426 ( .A1(n9040), .A2(n9608), .B1(n9039), .B2(n9022), .ZN(n9023)
         );
  NAND2_X1 U10427 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9429) );
  OAI211_X1 U10428 ( .C1(n9632), .C2(n9042), .A(n9023), .B(n9429), .ZN(n9024)
         );
  AOI21_X1 U10429 ( .B1(n9616), .B2(n9045), .A(n9024), .ZN(n9025) );
  OAI21_X1 U10430 ( .B1(n9026), .B2(n9047), .A(n9025), .ZN(P1_U3236) );
  NAND2_X1 U10431 ( .A1(n9489), .A2(n9040), .ZN(n9029) );
  INV_X1 U10432 ( .A(n9027), .ZN(n9481) );
  AOI22_X1 U10433 ( .A1(n9481), .A2(n9039), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9028) );
  OAI211_X1 U10434 ( .C1(n9518), .C2(n9042), .A(n9029), .B(n9028), .ZN(n9033)
         );
  INV_X1 U10435 ( .A(n9034), .ZN(n9035) );
  NOR2_X1 U10436 ( .A1(n9036), .A2(n9035), .ZN(n9038) );
  XNOR2_X1 U10437 ( .A(n9038), .B(n9037), .ZN(n9048) );
  AOI22_X1 U10438 ( .A1(n9040), .A2(n9661), .B1(n9039), .B2(n9670), .ZN(n9041)
         );
  NAND2_X1 U10439 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9366) );
  OAI211_X1 U10440 ( .C1(n9043), .C2(n9042), .A(n9041), .B(n9366), .ZN(n9044)
         );
  AOI21_X1 U10441 ( .B1(n9672), .B2(n9045), .A(n9044), .ZN(n9046) );
  OAI21_X1 U10442 ( .B1(n9048), .B2(n9047), .A(n9046), .ZN(P1_U3239) );
  NAND2_X1 U10443 ( .A1(n9049), .A2(n4377), .ZN(n9052) );
  OR2_X1 U10444 ( .A1(n9055), .A2(n9050), .ZN(n9051) );
  NAND2_X1 U10445 ( .A1(n9449), .A2(n9053), .ZN(n9169) );
  NAND2_X1 U10446 ( .A1(n9054), .A2(n4377), .ZN(n9057) );
  OR2_X1 U10447 ( .A1(n9055), .A2(n10272), .ZN(n9056) );
  INV_X1 U10448 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U10449 ( .A1(n9059), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U10450 ( .A1(n4391), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9060) );
  OAI211_X1 U10451 ( .C1(n4383), .C2(n9455), .A(n9061), .B(n9060), .ZN(n9465)
         );
  INV_X1 U10452 ( .A(n9465), .ZN(n9207) );
  NOR2_X1 U10453 ( .A1(n9683), .A2(n9207), .ZN(n9167) );
  NAND2_X1 U10454 ( .A1(n9167), .A2(n9449), .ZN(n9062) );
  AND2_X1 U10455 ( .A1(n9062), .A2(n9169), .ZN(n9163) );
  NAND2_X1 U10456 ( .A1(n9063), .A2(n4377), .ZN(n9066) );
  NAND2_X1 U10457 ( .A1(n9064), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U10458 ( .A1(n9692), .A2(n9067), .ZN(n9219) );
  INV_X1 U10459 ( .A(n9249), .ZN(n9068) );
  OR2_X1 U10460 ( .A1(n9069), .A2(n9068), .ZN(n9072) );
  AND2_X1 U10461 ( .A1(n9143), .A2(n9072), .ZN(n9273) );
  NAND2_X1 U10462 ( .A1(n9249), .A2(n9070), .ZN(n9514) );
  NAND2_X1 U10463 ( .A1(n9247), .A2(n9512), .ZN(n9534) );
  OR2_X1 U10464 ( .A1(n9514), .A2(n9534), .ZN(n9173) );
  MUX2_X1 U10465 ( .A(n9273), .B(n9073), .S(n9157), .Z(n9142) );
  MUX2_X1 U10466 ( .A(n9215), .B(n9074), .S(n9157), .Z(n9075) );
  INV_X1 U10467 ( .A(n9076), .ZN(n9243) );
  MUX2_X1 U10468 ( .A(n9222), .B(n9243), .S(n9157), .Z(n9120) );
  MUX2_X1 U10469 ( .A(n9235), .B(n9221), .S(n9157), .Z(n9119) );
  NAND2_X1 U10470 ( .A1(n4385), .A2(n9184), .ZN(n9077) );
  NAND3_X1 U10471 ( .A1(n9077), .A2(n9086), .A3(n9301), .ZN(n9080) );
  AND2_X1 U10472 ( .A1(n9090), .A2(n9157), .ZN(n9079) );
  NAND4_X1 U10473 ( .A1(n9080), .A2(n9089), .A3(n9079), .A4(n9262), .ZN(n9083)
         );
  AOI21_X1 U10474 ( .B1(n9092), .B2(n9087), .A(n9164), .ZN(n9081) );
  NAND2_X1 U10475 ( .A1(n9089), .A2(n9081), .ZN(n9082) );
  OAI211_X1 U10476 ( .C1(n9164), .C2(n9093), .A(n9083), .B(n9082), .ZN(n9084)
         );
  INV_X1 U10477 ( .A(n9084), .ZN(n9098) );
  AND2_X1 U10478 ( .A1(n9262), .A2(n9260), .ZN(n9298) );
  OAI21_X1 U10479 ( .B1(n4385), .B2(n9085), .A(n9298), .ZN(n9088) );
  AND2_X1 U10480 ( .A1(n9087), .A2(n9086), .ZN(n9252) );
  NAND2_X1 U10481 ( .A1(n9088), .A2(n9252), .ZN(n9091) );
  NAND2_X1 U10482 ( .A1(n9093), .A2(n9092), .ZN(n9095) );
  NAND2_X1 U10483 ( .A1(n9095), .A2(n9094), .ZN(n9253) );
  NAND3_X1 U10484 ( .A1(n9096), .A2(n9164), .A3(n9253), .ZN(n9097) );
  NAND4_X1 U10485 ( .A1(n9099), .A2(n9098), .A3(n9192), .A4(n9097), .ZN(n9109)
         );
  NAND2_X1 U10486 ( .A1(n9105), .A2(n9100), .ZN(n9251) );
  NAND2_X1 U10487 ( .A1(n9251), .A2(n9101), .ZN(n9102) );
  NAND3_X1 U10488 ( .A1(n9109), .A2(n9111), .A3(n9102), .ZN(n9103) );
  NAND3_X1 U10489 ( .A1(n9103), .A2(n9231), .A3(n9106), .ZN(n9104) );
  AND2_X1 U10490 ( .A1(n9104), .A2(n9112), .ZN(n9115) );
  INV_X1 U10491 ( .A(n9105), .ZN(n9107) );
  OAI21_X1 U10492 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9230) );
  INV_X1 U10493 ( .A(n9230), .ZN(n9110) );
  NAND2_X1 U10494 ( .A1(n9110), .A2(n9109), .ZN(n9113) );
  AND2_X1 U10495 ( .A1(n9112), .A2(n9111), .ZN(n9256) );
  AOI21_X1 U10496 ( .B1(n9113), .B2(n9256), .A(n4670), .ZN(n9114) );
  MUX2_X1 U10497 ( .A(n9117), .B(n8035), .S(n9164), .Z(n9118) );
  NAND3_X1 U10498 ( .A1(n9124), .A2(n9125), .A3(n9121), .ZN(n9122) );
  NAND3_X1 U10499 ( .A1(n9122), .A2(n9129), .A3(n9223), .ZN(n9128) );
  AND2_X1 U10500 ( .A1(n9223), .A2(n9123), .ZN(n9238) );
  NAND2_X1 U10501 ( .A1(n9124), .A2(n9238), .ZN(n9126) );
  AND2_X1 U10502 ( .A1(n9135), .A2(n9125), .ZN(n9240) );
  NAND2_X1 U10503 ( .A1(n9126), .A2(n9240), .ZN(n9127) );
  NAND2_X1 U10504 ( .A1(n9133), .A2(n9130), .ZN(n9239) );
  NAND2_X1 U10505 ( .A1(n9130), .A2(n4952), .ZN(n9131) );
  AND2_X1 U10506 ( .A1(n9131), .A2(n9134), .ZN(n9132) );
  NAND2_X1 U10507 ( .A1(n9132), .A2(n9137), .ZN(n9225) );
  NAND2_X1 U10508 ( .A1(n9225), .A2(n9133), .ZN(n9244) );
  OAI211_X1 U10509 ( .C1(n9136), .C2(n9239), .A(n9512), .B(n9244), .ZN(n9140)
         );
  AOI21_X1 U10510 ( .B1(n9136), .B2(n9135), .A(n4951), .ZN(n9138) );
  OAI21_X1 U10511 ( .B1(n9138), .B2(n9239), .A(n9137), .ZN(n9139) );
  INV_X1 U10512 ( .A(n9143), .ZN(n9144) );
  MUX2_X1 U10513 ( .A(n9144), .B(n9071), .S(n9164), .Z(n9149) );
  INV_X1 U10514 ( .A(n9149), .ZN(n9146) );
  MUX2_X1 U10515 ( .A(n9710), .B(n9506), .S(n9157), .Z(n9145) );
  AND2_X1 U10516 ( .A1(n9146), .A2(n9145), .ZN(n9151) );
  INV_X1 U10517 ( .A(n9171), .ZN(n9148) );
  MUX2_X1 U10518 ( .A(n9506), .B(n9710), .S(n9157), .Z(n9147) );
  AOI21_X1 U10519 ( .B1(n9149), .B2(n9148), .A(n9147), .ZN(n9150) );
  OR2_X1 U10520 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NAND2_X1 U10521 ( .A1(n9153), .A2(n9152), .ZN(n9154) );
  NAND2_X1 U10522 ( .A1(n9154), .A2(n8027), .ZN(n9156) );
  MUX2_X1 U10523 ( .A(n9274), .B(n9217), .S(n9157), .Z(n9155) );
  NAND3_X1 U10524 ( .A1(n9156), .A2(n4992), .A3(n9155), .ZN(n9159) );
  MUX2_X1 U10525 ( .A(n9461), .B(n9460), .S(n9157), .Z(n9158) );
  NAND3_X1 U10526 ( .A1(n9464), .A2(n9159), .A3(n9158), .ZN(n9161) );
  MUX2_X1 U10527 ( .A(n9219), .B(n9214), .S(n9164), .Z(n9160) );
  NAND2_X1 U10528 ( .A1(n9452), .A2(n9465), .ZN(n9162) );
  NAND2_X1 U10529 ( .A1(n9683), .A2(n9162), .ZN(n9276) );
  INV_X1 U10530 ( .A(n9163), .ZN(n9280) );
  AOI21_X1 U10531 ( .B1(n9280), .B2(n9164), .A(n9208), .ZN(n9165) );
  INV_X1 U10532 ( .A(n9167), .ZN(n9168) );
  AND2_X1 U10533 ( .A1(n9169), .A2(n9168), .ZN(n9320) );
  INV_X1 U10534 ( .A(n9170), .ZN(n9172) );
  INV_X1 U10535 ( .A(n9504), .ZN(n9496) );
  INV_X1 U10536 ( .A(n9173), .ZN(n9203) );
  INV_X1 U10537 ( .A(n9175), .ZN(n9198) );
  INV_X1 U10538 ( .A(n9652), .ZN(n9650) );
  INV_X1 U10539 ( .A(n9176), .ZN(n9191) );
  NAND4_X1 U10540 ( .A1(n9180), .A2(n9179), .A3(n9178), .A4(n9177), .ZN(n9183)
         );
  NOR3_X1 U10541 ( .A1(n9183), .A2(n9182), .A3(n9181), .ZN(n9187) );
  NAND4_X1 U10542 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n9184), .ZN(n9189)
         );
  NOR2_X1 U10543 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  NAND3_X1 U10544 ( .A1(n9192), .A2(n9191), .A3(n9190), .ZN(n9193) );
  NOR2_X1 U10545 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  NAND4_X1 U10546 ( .A1(n9650), .A2(n4394), .A3(n9196), .A4(n9195), .ZN(n9197)
         );
  NOR3_X1 U10547 ( .A1(n9198), .A2(n9116), .A3(n9197), .ZN(n9199) );
  NAND4_X1 U10548 ( .A1(n9577), .A2(n8036), .A3(n4974), .A4(n9199), .ZN(n9200)
         );
  NOR2_X1 U10549 ( .A1(n9555), .A2(n9200), .ZN(n9201) );
  AND2_X1 U10550 ( .A1(n9548), .A2(n9201), .ZN(n9202) );
  NAND4_X1 U10551 ( .A1(n9487), .A2(n9496), .A3(n9203), .A4(n9202), .ZN(n9204)
         );
  OR3_X1 U10552 ( .A1(n9205), .A2(n9204), .A3(n9316), .ZN(n9206) );
  NOR2_X1 U10553 ( .A1(n9691), .A2(n9206), .ZN(n9209) );
  NAND2_X1 U10554 ( .A1(n9683), .A2(n9207), .ZN(n9318) );
  NAND4_X1 U10555 ( .A1(n9320), .A2(n9209), .A3(n9318), .A4(n9342), .ZN(n9211)
         );
  AND2_X1 U10556 ( .A1(n9211), .A2(n9210), .ZN(n9282) );
  NOR2_X1 U10557 ( .A1(n9281), .A2(n9212), .ZN(n9324) );
  OAI211_X1 U10558 ( .C1(n9213), .C2(n9282), .A(n9340), .B(n9324), .ZN(n9347)
         );
  NAND2_X1 U10559 ( .A1(n9214), .A2(n9460), .ZN(n9317) );
  NAND2_X1 U10560 ( .A1(n9274), .A2(n4963), .ZN(n9216) );
  AND3_X1 U10561 ( .A1(n9461), .A2(n9217), .A3(n9216), .ZN(n9218) );
  OR2_X1 U10562 ( .A1(n9317), .A2(n9218), .ZN(n9220) );
  NAND2_X1 U10563 ( .A1(n9220), .A2(n9219), .ZN(n9322) );
  NAND3_X1 U10564 ( .A1(n9223), .A2(n9222), .A3(n9221), .ZN(n9224) );
  NOR2_X1 U10565 ( .A1(n9225), .A2(n9224), .ZN(n9250) );
  INV_X1 U10566 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U10567 ( .A1(n9227), .A2(n9253), .ZN(n9228) );
  NOR2_X1 U10568 ( .A1(n9251), .A2(n9228), .ZN(n9229) );
  NOR2_X1 U10569 ( .A1(n9230), .A2(n9229), .ZN(n9233) );
  INV_X1 U10570 ( .A(n9256), .ZN(n9232) );
  OAI211_X1 U10571 ( .C1(n9233), .C2(n9232), .A(n9117), .B(n9231), .ZN(n9234)
         );
  NAND2_X1 U10572 ( .A1(n9234), .A2(n8035), .ZN(n9236) );
  NAND2_X1 U10573 ( .A1(n9236), .A2(n9235), .ZN(n9237) );
  NAND2_X1 U10574 ( .A1(n9250), .A2(n9237), .ZN(n9248) );
  INV_X1 U10575 ( .A(n9238), .ZN(n9242) );
  INV_X1 U10576 ( .A(n9239), .ZN(n9241) );
  OAI211_X1 U10577 ( .C1(n9243), .C2(n9242), .A(n9241), .B(n9240), .ZN(n9245)
         );
  NAND2_X1 U10578 ( .A1(n9245), .A2(n9244), .ZN(n9246) );
  NAND4_X1 U10579 ( .A1(n9249), .A2(n9248), .A3(n9247), .A4(n9246), .ZN(n9311)
         );
  INV_X1 U10580 ( .A(n9250), .ZN(n9258) );
  INV_X1 U10581 ( .A(n9251), .ZN(n9255) );
  AND2_X1 U10582 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  NAND4_X1 U10583 ( .A1(n8035), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n9257)
         );
  NOR2_X1 U10584 ( .A1(n9258), .A2(n9257), .ZN(n9285) );
  AND3_X1 U10585 ( .A1(n9260), .A2(n9265), .A3(n9259), .ZN(n9263) );
  NAND2_X1 U10586 ( .A1(n9301), .A2(n9261), .ZN(n9303) );
  AND3_X1 U10587 ( .A1(n9263), .A2(n9262), .A3(n9303), .ZN(n9297) );
  INV_X1 U10588 ( .A(n9264), .ZN(n9267) );
  NAND3_X1 U10589 ( .A1(n9267), .A2(n9266), .A3(n9265), .ZN(n9268) );
  NAND3_X1 U10590 ( .A1(n9268), .A2(n9301), .A3(n9300), .ZN(n9269) );
  AOI22_X1 U10591 ( .A1(n9297), .A2(n9270), .B1(n9269), .B2(n9298), .ZN(n9271)
         );
  AND2_X1 U10592 ( .A1(n9285), .A2(n9271), .ZN(n9272) );
  NOR2_X1 U10593 ( .A1(n9311), .A2(n9272), .ZN(n9275) );
  INV_X1 U10594 ( .A(n9273), .ZN(n9313) );
  OAI211_X1 U10595 ( .C1(n9275), .C2(n9313), .A(n9274), .B(n9312), .ZN(n9277)
         );
  OAI21_X1 U10596 ( .B1(n9317), .B2(n9277), .A(n9276), .ZN(n9278) );
  NOR2_X1 U10597 ( .A1(n9322), .A2(n9278), .ZN(n9279) );
  OAI211_X1 U10598 ( .C1(n9280), .C2(n9279), .A(n6618), .B(n9342), .ZN(n9284)
         );
  AND2_X1 U10599 ( .A1(n9281), .A2(n9339), .ZN(n9333) );
  INV_X1 U10600 ( .A(n9282), .ZN(n9283) );
  NAND4_X1 U10601 ( .A1(n9284), .A2(n9340), .A3(n9333), .A4(n9283), .ZN(n9338)
         );
  INV_X1 U10602 ( .A(n9285), .ZN(n9309) );
  INV_X1 U10603 ( .A(n9286), .ZN(n9288) );
  NAND3_X1 U10604 ( .A1(n9288), .A2(n9287), .A3(n6618), .ZN(n9290) );
  NAND2_X1 U10605 ( .A1(n9290), .A2(n9289), .ZN(n9291) );
  OR2_X1 U10606 ( .A1(n9292), .A2(n9291), .ZN(n9296) );
  INV_X1 U10607 ( .A(n9293), .ZN(n9294) );
  AOI21_X1 U10608 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(n9307) );
  INV_X1 U10609 ( .A(n9297), .ZN(n9306) );
  INV_X1 U10610 ( .A(n9298), .ZN(n9305) );
  NAND3_X1 U10611 ( .A1(n9301), .A2(n9300), .A3(n9299), .ZN(n9302) );
  NAND2_X1 U10612 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  OAI22_X1 U10613 ( .A1(n9307), .A2(n9306), .B1(n9305), .B2(n9304), .ZN(n9308)
         );
  NOR2_X1 U10614 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  NOR2_X1 U10615 ( .A1(n9311), .A2(n9310), .ZN(n9314) );
  OAI21_X1 U10616 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9315) );
  OR3_X1 U10617 ( .A1(n9317), .A2(n9316), .A3(n9315), .ZN(n9319) );
  NAND2_X1 U10618 ( .A1(n9319), .A2(n9318), .ZN(n9321) );
  OAI21_X1 U10619 ( .B1(n9322), .B2(n9321), .A(n9320), .ZN(n9323) );
  NAND2_X1 U10620 ( .A1(n9323), .A2(n9342), .ZN(n9334) );
  NAND2_X1 U10621 ( .A1(n9324), .A2(n4378), .ZN(n9325) );
  OR2_X1 U10622 ( .A1(n9334), .A2(n9325), .ZN(n9337) );
  NAND3_X1 U10623 ( .A1(n9925), .A2(n9327), .A3(n9326), .ZN(n9330) );
  INV_X1 U10624 ( .A(P1_B_REG_SCAN_IN), .ZN(n10233) );
  AOI21_X1 U10625 ( .B1(n9328), .B2(n9339), .A(n10233), .ZN(n9329) );
  OAI21_X1 U10626 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9336) );
  NAND3_X1 U10627 ( .A1(n9334), .A2(n9333), .A3(n4378), .ZN(n9335) );
  NAND3_X1 U10628 ( .A1(n6618), .A2(n9340), .A3(n9339), .ZN(n9341) );
  NOR2_X1 U10629 ( .A1(n6084), .A2(n9341), .ZN(n9343) );
  NAND3_X1 U10630 ( .A1(n9344), .A2(n9343), .A3(n9342), .ZN(n9345) );
  NAND3_X1 U10631 ( .A1(n9347), .A2(n9346), .A3(n9345), .ZN(P1_U3240) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9465), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10634 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9467), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9489), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9506), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9488), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8024), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10639 ( .A(n9549), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9350), .Z(
        P1_U3578) );
  MUX2_X1 U10640 ( .A(n9564), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9350), .Z(
        P1_U3577) );
  INV_X1 U10641 ( .A(n9349), .ZN(n9578) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9578), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10643 ( .A(n9596), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9350), .Z(
        P1_U3575) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9608), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9595), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9607), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10647 ( .A(n9661), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9350), .Z(
        P1_U3571) );
  MUX2_X1 U10648 ( .A(n9351), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9350), .Z(
        P1_U3570) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9658), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9352), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9353), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9354), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9355), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9356), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9357), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10656 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9358), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10657 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9359), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9360), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10659 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9361), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10660 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9363), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10661 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9364), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10662 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9365), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U10663 ( .A(n9366), .ZN(n9373) );
  OAI22_X1 U10664 ( .A1(n9368), .A2(n9367), .B1(n9375), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n9914) );
  XNOR2_X1 U10665 ( .A(n9909), .B(n9369), .ZN(n9915) );
  NAND2_X1 U10666 ( .A1(n9914), .A2(n9915), .ZN(n9913) );
  OAI21_X1 U10667 ( .B1(n9909), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9913), .ZN(
        n9391) );
  XNOR2_X1 U10668 ( .A(n9392), .B(n9391), .ZN(n9371) );
  INV_X1 U10669 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9370) );
  NOR2_X1 U10670 ( .A1(n9370), .A2(n9371), .ZN(n9393) );
  AOI211_X1 U10671 ( .C1(n9371), .C2(n9370), .A(n9393), .B(n9901), .ZN(n9372)
         );
  AOI211_X1 U10672 ( .C1(n9397), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9373), .B(
        n9372), .ZN(n9384) );
  NAND2_X1 U10673 ( .A1(n9377), .A2(n9376), .ZN(n9378) );
  XNOR2_X1 U10674 ( .A(n9377), .B(n9909), .ZN(n9912) );
  NAND2_X1 U10675 ( .A1(n9912), .A2(n6392), .ZN(n9911) );
  NAND2_X1 U10676 ( .A1(n9378), .A2(n9911), .ZN(n9385) );
  XNOR2_X1 U10677 ( .A(n9392), .B(n9385), .ZN(n9380) );
  INV_X1 U10678 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9379) );
  NOR2_X1 U10679 ( .A1(n9379), .A2(n9380), .ZN(n9386) );
  AOI211_X1 U10680 ( .C1(n9380), .C2(n9379), .A(n9386), .B(n9893), .ZN(n9381)
         );
  AOI21_X1 U10681 ( .B1(n9910), .B2(n9382), .A(n9381), .ZN(n9383) );
  NAND2_X1 U10682 ( .A1(n9384), .A2(n9383), .ZN(P1_U3256) );
  NOR2_X1 U10683 ( .A1(n9392), .A2(n9385), .ZN(n9387) );
  NAND2_X1 U10684 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9413), .ZN(n9388) );
  OAI21_X1 U10685 ( .B1(n9413), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9388), .ZN(
        n9389) );
  AOI211_X1 U10686 ( .C1(n9390), .C2(n9389), .A(n9412), .B(n9893), .ZN(n9403)
         );
  NOR2_X1 U10687 ( .A1(n9392), .A2(n9391), .ZN(n9394) );
  NOR2_X1 U10688 ( .A1(n9394), .A2(n9393), .ZN(n9396) );
  XNOR2_X1 U10689 ( .A(n9413), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9395) );
  NOR2_X1 U10690 ( .A1(n9396), .A2(n9395), .ZN(n9404) );
  AOI211_X1 U10691 ( .C1(n9396), .C2(n9395), .A(n9404), .B(n9901), .ZN(n9402)
         );
  NAND2_X1 U10692 ( .A1(n9397), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9399) );
  OAI211_X1 U10693 ( .C1(n9888), .C2(n9400), .A(n9399), .B(n9398), .ZN(n9401)
         );
  OR3_X1 U10694 ( .A1(n9403), .A2(n9402), .A3(n9401), .ZN(P1_U3257) );
  INV_X1 U10695 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9411) );
  XNOR2_X1 U10696 ( .A(n9426), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9406) );
  AOI21_X1 U10697 ( .B1(n9413), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9404), .ZN(
        n9405) );
  NOR2_X1 U10698 ( .A1(n9405), .A2(n9406), .ZN(n9425) );
  AOI21_X1 U10699 ( .B1(n9406), .B2(n9405), .A(n9425), .ZN(n9407) );
  NAND2_X1 U10700 ( .A1(n9917), .A2(n9407), .ZN(n9410) );
  INV_X1 U10701 ( .A(n9408), .ZN(n9409) );
  OAI211_X1 U10702 ( .C1(n9923), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9416)
         );
  NAND2_X1 U10703 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9426), .ZN(n9418) );
  OAI21_X1 U10704 ( .B1(n9426), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9418), .ZN(
        n9414) );
  AOI211_X1 U10705 ( .C1(n4403), .C2(n9414), .A(n9419), .B(n9893), .ZN(n9415)
         );
  AOI211_X1 U10706 ( .C1(n9910), .C2(n9426), .A(n9416), .B(n9415), .ZN(n9417)
         );
  INV_X1 U10707 ( .A(n9417), .ZN(P1_U3258) );
  INV_X1 U10708 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U10709 ( .A1(n9437), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9420) );
  OAI21_X1 U10710 ( .B1(n9437), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9420), .ZN(
        n9421) );
  AOI211_X1 U10711 ( .C1(n9422), .C2(n9421), .A(n9435), .B(n9893), .ZN(n9423)
         );
  AOI21_X1 U10712 ( .B1(n9910), .B2(n9437), .A(n9423), .ZN(n9433) );
  XNOR2_X1 U10713 ( .A(n9424), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9428) );
  AOI21_X1 U10714 ( .B1(n9426), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9425), .ZN(
        n9427) );
  NAND2_X1 U10715 ( .A1(n9428), .A2(n9427), .ZN(n9436) );
  OAI21_X1 U10716 ( .B1(n9428), .B2(n9427), .A(n9436), .ZN(n9431) );
  INV_X1 U10717 ( .A(n9429), .ZN(n9430) );
  AOI21_X1 U10718 ( .B1(n9917), .B2(n9431), .A(n9430), .ZN(n9432) );
  OAI211_X1 U10719 ( .C1(n9923), .C2(n9434), .A(n9433), .B(n9432), .ZN(
        P1_U3259) );
  OAI21_X1 U10720 ( .B1(n9437), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9436), .ZN(
        n9439) );
  XNOR2_X1 U10721 ( .A(n9439), .B(n9438), .ZN(n9442) );
  OAI22_X1 U10722 ( .A1(n9441), .A2(n9893), .B1(n9442), .B2(n9901), .ZN(n9440)
         );
  AOI21_X1 U10723 ( .B1(n9442), .B2(n9917), .A(n9910), .ZN(n9443) );
  NAND2_X1 U10724 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  INV_X1 U10725 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9447) );
  OAI21_X1 U10726 ( .B1(n9923), .B2(n9447), .A(n9446), .ZN(n9448) );
  XNOR2_X1 U10727 ( .A(n9450), .B(n9449), .ZN(n9680) );
  NAND2_X1 U10728 ( .A1(n9680), .A2(n9600), .ZN(n9454) );
  NOR2_X1 U10729 ( .A1(n9835), .A2(n10233), .ZN(n9451) );
  NOR2_X1 U10730 ( .A1(n9633), .A2(n9451), .ZN(n9466) );
  NAND2_X1 U10731 ( .A1(n9466), .A2(n9452), .ZN(n9685) );
  NOR2_X1 U10732 ( .A1(n9679), .A2(n9685), .ZN(n9456) );
  AOI21_X1 U10733 ( .B1(n9679), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9456), .ZN(
        n9453) );
  OAI211_X1 U10734 ( .C1(n9682), .C2(n9635), .A(n9454), .B(n9453), .ZN(
        P1_U3261) );
  NOR2_X1 U10735 ( .A1(n7131), .A2(n9455), .ZN(n9457) );
  AOI211_X1 U10736 ( .C1(n9683), .C2(n9671), .A(n9457), .B(n9456), .ZN(n9458)
         );
  OAI21_X1 U10737 ( .B1(n9686), .B2(n9675), .A(n9458), .ZN(P1_U3262) );
  NAND2_X1 U10738 ( .A1(n9700), .A2(n9467), .ZN(n9690) );
  NAND2_X1 U10739 ( .A1(n9689), .A2(n9690), .ZN(n9459) );
  XNOR2_X1 U10740 ( .A(n9459), .B(n9691), .ZN(n9478) );
  INV_X1 U10741 ( .A(n9460), .ZN(n9462) );
  AOI22_X1 U10742 ( .A1(n9467), .A2(n9659), .B1(n9466), .B2(n9465), .ZN(n9468)
         );
  NAND2_X1 U10743 ( .A1(n9469), .A2(n9468), .ZN(n9687) );
  AOI21_X1 U10744 ( .B1(n9692), .B2(n9470), .A(n9944), .ZN(n9472) );
  NAND2_X1 U10745 ( .A1(n9472), .A2(n9471), .ZN(n9694) );
  INV_X1 U10746 ( .A(n9642), .ZN(n9618) );
  INV_X1 U10747 ( .A(n9473), .ZN(n9474) );
  AOI22_X1 U10748 ( .A1(n9474), .A2(n9669), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9679), .ZN(n9476) );
  NAND2_X1 U10749 ( .A1(n9692), .A2(n9671), .ZN(n9475) );
  OAI211_X1 U10750 ( .C1(n9694), .C2(n9618), .A(n9476), .B(n9475), .ZN(n9477)
         );
  AOI21_X1 U10751 ( .B1(n9710), .B2(n9498), .A(n9480), .ZN(n9711) );
  INV_X1 U10752 ( .A(n9710), .ZN(n9483) );
  AOI22_X1 U10753 ( .A1(n9481), .A2(n9669), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9679), .ZN(n9482) );
  OAI21_X1 U10754 ( .B1(n9483), .B2(n9635), .A(n9482), .ZN(n9494) );
  NAND2_X1 U10755 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  XOR2_X1 U10756 ( .A(n9487), .B(n9486), .Z(n9492) );
  AOI211_X1 U10757 ( .C1(n9600), .C2(n9711), .A(n9494), .B(n9493), .ZN(n9495)
         );
  OAI21_X1 U10758 ( .B1(n9714), .B2(n9645), .A(n9495), .ZN(P1_U3265) );
  XNOR2_X1 U10759 ( .A(n9497), .B(n9496), .ZN(n9719) );
  INV_X1 U10760 ( .A(n9519), .ZN(n9500) );
  INV_X1 U10761 ( .A(n9498), .ZN(n9499) );
  AOI21_X1 U10762 ( .B1(n9715), .B2(n9500), .A(n9499), .ZN(n9716) );
  AOI22_X1 U10763 ( .A1(n9501), .A2(n9669), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9679), .ZN(n9502) );
  OAI21_X1 U10764 ( .B1(n9503), .B2(n9635), .A(n9502), .ZN(n9509) );
  XNOR2_X1 U10765 ( .A(n9505), .B(n9504), .ZN(n9507) );
  AOI222_X1 U10766 ( .A1(n9656), .A2(n9507), .B1(n9506), .B2(n9660), .C1(n8024), .C2(n9659), .ZN(n9718) );
  NOR2_X1 U10767 ( .A1(n9718), .A2(n9679), .ZN(n9508) );
  AOI211_X1 U10768 ( .C1(n9716), .C2(n9600), .A(n9509), .B(n9508), .ZN(n9510)
         );
  OAI21_X1 U10769 ( .B1(n9719), .B2(n9645), .A(n9510), .ZN(P1_U3266) );
  XOR2_X1 U10770 ( .A(n9514), .B(n9511), .Z(n9724) );
  AOI22_X1 U10771 ( .A1(n9722), .A2(n9671), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9679), .ZN(n9525) );
  NAND2_X1 U10772 ( .A1(n9513), .A2(n9512), .ZN(n9515) );
  XNOR2_X1 U10773 ( .A(n9515), .B(n9514), .ZN(n9516) );
  OAI222_X1 U10774 ( .A1(n9633), .A2(n9518), .B1(n9631), .B2(n9517), .C1(n9516), .C2(n9628), .ZN(n9720) );
  AOI211_X1 U10775 ( .C1(n9722), .C2(n9527), .A(n9944), .B(n9519), .ZN(n9721)
         );
  INV_X1 U10776 ( .A(n9721), .ZN(n9522) );
  OAI22_X1 U10777 ( .A1(n9522), .A2(n9521), .B1(n9520), .B2(n9637), .ZN(n9523)
         );
  OAI21_X1 U10778 ( .B1(n9720), .B2(n9523), .A(n7131), .ZN(n9524) );
  OAI211_X1 U10779 ( .C1(n9724), .C2(n9645), .A(n9525), .B(n9524), .ZN(
        P1_U3267) );
  XNOR2_X1 U10780 ( .A(n9526), .B(n9534), .ZN(n9729) );
  INV_X1 U10781 ( .A(n9527), .ZN(n9528) );
  AOI21_X1 U10782 ( .B1(n9725), .B2(n9540), .A(n9528), .ZN(n9726) );
  INV_X1 U10783 ( .A(n9529), .ZN(n9530) );
  AOI22_X1 U10784 ( .A1(n9530), .A2(n9669), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9679), .ZN(n9531) );
  OAI21_X1 U10785 ( .B1(n9532), .B2(n9635), .A(n9531), .ZN(n9537) );
  XOR2_X1 U10786 ( .A(n9533), .B(n9534), .Z(n9535) );
  AOI211_X1 U10787 ( .C1(n9726), .C2(n9600), .A(n9537), .B(n9536), .ZN(n9538)
         );
  OAI21_X1 U10788 ( .B1(n9645), .B2(n9729), .A(n9538), .ZN(P1_U3268) );
  XOR2_X1 U10789 ( .A(n9539), .B(n9548), .Z(n9734) );
  INV_X1 U10790 ( .A(n9557), .ZN(n9542) );
  INV_X1 U10791 ( .A(n9540), .ZN(n9541) );
  AOI211_X1 U10792 ( .C1(n9731), .C2(n9542), .A(n9944), .B(n9541), .ZN(n9730)
         );
  AOI22_X1 U10793 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(n9679), .B1(n9543), .B2(
        n9669), .ZN(n9544) );
  OAI21_X1 U10794 ( .B1(n9545), .B2(n9635), .A(n9544), .ZN(n9552) );
  OAI21_X1 U10795 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9550) );
  AOI222_X1 U10796 ( .A1(n9656), .A2(n9550), .B1(n9549), .B2(n9660), .C1(n9578), .C2(n9659), .ZN(n9733) );
  NOR2_X1 U10797 ( .A1(n9733), .A2(n9679), .ZN(n9551) );
  AOI211_X1 U10798 ( .C1(n9730), .C2(n9642), .A(n9552), .B(n9551), .ZN(n9553)
         );
  OAI21_X1 U10799 ( .B1(n9734), .B2(n9645), .A(n9553), .ZN(P1_U3269) );
  OAI21_X1 U10800 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(n9739) );
  AOI211_X1 U10801 ( .C1(n9736), .C2(n5056), .A(n9944), .B(n9557), .ZN(n9735)
         );
  AOI22_X1 U10802 ( .A1(n9679), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9558), .B2(
        n9669), .ZN(n9559) );
  OAI21_X1 U10803 ( .B1(n9560), .B2(n9635), .A(n9559), .ZN(n9567) );
  OAI21_X1 U10804 ( .B1(n9563), .B2(n9562), .A(n9561), .ZN(n9565) );
  AOI222_X1 U10805 ( .A1(n9656), .A2(n9565), .B1(n9564), .B2(n9660), .C1(n9596), .C2(n9659), .ZN(n9738) );
  NOR2_X1 U10806 ( .A1(n9738), .A2(n9679), .ZN(n9566) );
  AOI211_X1 U10807 ( .C1(n9735), .C2(n9642), .A(n9567), .B(n9566), .ZN(n9568)
         );
  OAI21_X1 U10808 ( .B1(n9645), .B2(n9739), .A(n9568), .ZN(P1_U3270) );
  XOR2_X1 U10809 ( .A(n9569), .B(n9577), .Z(n9744) );
  INV_X1 U10810 ( .A(n5056), .ZN(n9570) );
  AOI21_X1 U10811 ( .B1(n9740), .B2(n9586), .A(n9570), .ZN(n9741) );
  INV_X1 U10812 ( .A(n9571), .ZN(n9572) );
  AOI22_X1 U10813 ( .A1(n9679), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9572), .B2(
        n9669), .ZN(n9573) );
  OAI21_X1 U10814 ( .B1(n9574), .B2(n9635), .A(n9573), .ZN(n9581) );
  OAI21_X1 U10815 ( .B1(n9577), .B2(n9575), .A(n9576), .ZN(n9579) );
  AOI222_X1 U10816 ( .A1(n9656), .A2(n9579), .B1(n9578), .B2(n9660), .C1(n9608), .C2(n9659), .ZN(n9743) );
  NOR2_X1 U10817 ( .A1(n9743), .A2(n9679), .ZN(n9580) );
  AOI211_X1 U10818 ( .C1(n9741), .C2(n9600), .A(n9581), .B(n9580), .ZN(n9582)
         );
  OAI21_X1 U10819 ( .B1(n9645), .B2(n9744), .A(n9582), .ZN(P1_U3271) );
  XNOR2_X1 U10820 ( .A(n9583), .B(n9584), .ZN(n9749) );
  INV_X1 U10821 ( .A(n9585), .ZN(n9588) );
  INV_X1 U10822 ( .A(n9586), .ZN(n9587) );
  AOI21_X1 U10823 ( .B1(n9745), .B2(n9588), .A(n9587), .ZN(n9746) );
  INV_X1 U10824 ( .A(n9589), .ZN(n9590) );
  AOI22_X1 U10825 ( .A1(n9679), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9590), .B2(
        n9669), .ZN(n9591) );
  OAI21_X1 U10826 ( .B1(n9592), .B2(n9635), .A(n9591), .ZN(n9599) );
  OAI21_X1 U10827 ( .B1(n4382), .B2(n8036), .A(n9593), .ZN(n9597) );
  AOI222_X1 U10828 ( .A1(n9656), .A2(n9597), .B1(n9596), .B2(n9660), .C1(n9595), .C2(n9659), .ZN(n9748) );
  NOR2_X1 U10829 ( .A1(n9748), .A2(n9679), .ZN(n9598) );
  AOI211_X1 U10830 ( .C1(n9746), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9601)
         );
  OAI21_X1 U10831 ( .B1(n9645), .B2(n9749), .A(n9601), .ZN(P1_U3272) );
  NAND2_X1 U10832 ( .A1(n4384), .A2(n9602), .ZN(n9604) );
  NAND2_X1 U10833 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  XNOR2_X1 U10834 ( .A(n9605), .B(n9174), .ZN(n9606) );
  NAND2_X1 U10835 ( .A1(n9606), .A2(n9656), .ZN(n9610) );
  AOI22_X1 U10836 ( .A1(n9608), .A2(n9660), .B1(n9659), .B2(n9607), .ZN(n9609)
         );
  NAND2_X1 U10837 ( .A1(n9610), .A2(n9609), .ZN(n9754) );
  OAI21_X1 U10838 ( .B1(n9752), .B2(n9611), .A(n9935), .ZN(n9612) );
  OR2_X1 U10839 ( .A1(n9612), .A2(n9585), .ZN(n9751) );
  INV_X1 U10840 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9614) );
  OAI22_X1 U10841 ( .A1(n7131), .A2(n9614), .B1(n9613), .B2(n9637), .ZN(n9615)
         );
  AOI21_X1 U10842 ( .B1(n9616), .B2(n9671), .A(n9615), .ZN(n9617) );
  OAI21_X1 U10843 ( .B1(n9751), .B2(n9618), .A(n9617), .ZN(n9623) );
  OR2_X1 U10844 ( .A1(n9619), .A2(n9174), .ZN(n9620) );
  NAND2_X1 U10845 ( .A1(n9621), .A2(n9620), .ZN(n9750) );
  NOR2_X1 U10846 ( .A1(n9750), .A2(n9645), .ZN(n9622) );
  AOI211_X1 U10847 ( .C1(n7131), .C2(n9754), .A(n9623), .B(n9622), .ZN(n9624)
         );
  INV_X1 U10848 ( .A(n9624), .ZN(P1_U3273) );
  XNOR2_X1 U10849 ( .A(n9116), .B(n9625), .ZN(n9766) );
  XNOR2_X1 U10850 ( .A(n9627), .B(n9626), .ZN(n9629) );
  OAI222_X1 U10851 ( .A1(n9633), .A2(n9632), .B1(n9631), .B2(n9630), .C1(n9629), .C2(n9628), .ZN(n9762) );
  NAND2_X1 U10852 ( .A1(n9762), .A2(n7131), .ZN(n9644) );
  AOI211_X1 U10853 ( .C1(n9764), .C2(n9668), .A(n9944), .B(n9634), .ZN(n9763)
         );
  INV_X1 U10854 ( .A(n9764), .ZN(n9636) );
  NOR2_X1 U10855 ( .A1(n9636), .A2(n9635), .ZN(n9641) );
  INV_X1 U10856 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9639) );
  OAI22_X1 U10857 ( .A1(n7131), .A2(n9639), .B1(n9638), .B2(n9637), .ZN(n9640)
         );
  AOI211_X1 U10858 ( .C1(n9763), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9643)
         );
  OAI211_X1 U10859 ( .C1(n9766), .C2(n9645), .A(n9644), .B(n9643), .ZN(
        P1_U3275) );
  OR2_X1 U10860 ( .A1(n9647), .A2(n9646), .ZN(n9649) );
  NAND2_X1 U10861 ( .A1(n9649), .A2(n9648), .ZN(n9651) );
  XNOR2_X1 U10862 ( .A(n9651), .B(n9650), .ZN(n9769) );
  NAND2_X1 U10863 ( .A1(n9653), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U10864 ( .A1(n9655), .A2(n9654), .ZN(n9657) );
  NAND2_X1 U10865 ( .A1(n9657), .A2(n9656), .ZN(n9663) );
  AOI22_X1 U10866 ( .A1(n9661), .A2(n9660), .B1(n9659), .B2(n9658), .ZN(n9662)
         );
  NAND2_X1 U10867 ( .A1(n9663), .A2(n9662), .ZN(n9664) );
  AOI21_X1 U10868 ( .B1(n9769), .B2(n9665), .A(n9664), .ZN(n9771) );
  OR2_X1 U10869 ( .A1(n9666), .A2(n8028), .ZN(n9667) );
  NAND2_X1 U10870 ( .A1(n9668), .A2(n9667), .ZN(n9767) );
  AOI22_X1 U10871 ( .A1(n9679), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9670), .B2(
        n9669), .ZN(n9674) );
  NAND2_X1 U10872 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  OAI211_X1 U10873 ( .C1(n9767), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  AOI21_X1 U10874 ( .B1(n9769), .B2(n9677), .A(n9676), .ZN(n9678) );
  OAI21_X1 U10875 ( .B1(n9771), .B2(n9679), .A(n9678), .ZN(P1_U3276) );
  NAND2_X1 U10876 ( .A1(n9680), .A2(n9935), .ZN(n9681) );
  OAI211_X1 U10877 ( .C1(n9682), .C2(n9965), .A(n9681), .B(n9685), .ZN(n9801)
         );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9801), .S(n9977), .Z(
        P1_U3554) );
  NAND2_X1 U10879 ( .A1(n9683), .A2(n9934), .ZN(n9684) );
  OAI211_X1 U10880 ( .C1(n9686), .C2(n9944), .A(n9685), .B(n9684), .ZN(n9802)
         );
  MUX2_X1 U10881 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9802), .S(n9977), .Z(
        P1_U3553) );
  INV_X1 U10882 ( .A(n9687), .ZN(n9699) );
  OR3_X1 U10883 ( .A1(n9689), .A2(n9691), .A3(n9962), .ZN(n9698) );
  INV_X1 U10884 ( .A(n9962), .ZN(n9958) );
  NOR2_X1 U10885 ( .A1(n5065), .A2(n5064), .ZN(n9693) );
  NAND3_X1 U10886 ( .A1(n9699), .A2(n9698), .A3(n9697), .ZN(n9803) );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9803), .S(n9977), .Z(
        P1_U3552) );
  AOI22_X1 U10888 ( .A1(n9701), .A2(n9935), .B1(n9934), .B2(n9700), .ZN(n9702)
         );
  OAI211_X1 U10889 ( .C1(n9704), .C2(n9962), .A(n9703), .B(n9702), .ZN(n9804)
         );
  MUX2_X1 U10890 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9804), .S(n9977), .Z(
        P1_U3551) );
  AOI21_X1 U10891 ( .B1(n9934), .B2(n9706), .A(n9705), .ZN(n9707) );
  OAI211_X1 U10892 ( .C1(n9709), .C2(n9962), .A(n9708), .B(n9707), .ZN(n9805)
         );
  MUX2_X1 U10893 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9805), .S(n9977), .Z(
        P1_U3550) );
  AOI22_X1 U10894 ( .A1(n9711), .A2(n9935), .B1(n9934), .B2(n9710), .ZN(n9712)
         );
  OAI211_X1 U10895 ( .C1(n9714), .C2(n9962), .A(n9713), .B(n9712), .ZN(n9806)
         );
  MUX2_X1 U10896 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9806), .S(n9977), .Z(
        P1_U3549) );
  AOI22_X1 U10897 ( .A1(n9716), .A2(n9935), .B1(n9934), .B2(n9715), .ZN(n9717)
         );
  OAI211_X1 U10898 ( .C1(n9719), .C2(n9962), .A(n9718), .B(n9717), .ZN(n9807)
         );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9807), .S(n9977), .Z(
        P1_U3548) );
  AOI22_X1 U10900 ( .A1(n9726), .A2(n9935), .B1(n9934), .B2(n9725), .ZN(n9727)
         );
  OAI211_X1 U10901 ( .C1(n9729), .C2(n9962), .A(n9728), .B(n9727), .ZN(n9809)
         );
  MUX2_X1 U10902 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9809), .S(n9977), .Z(
        P1_U3546) );
  AOI21_X1 U10903 ( .B1(n9934), .B2(n9731), .A(n9730), .ZN(n9732) );
  OAI211_X1 U10904 ( .C1(n9734), .C2(n9962), .A(n9733), .B(n9732), .ZN(n9810)
         );
  MUX2_X1 U10905 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9810), .S(n9977), .Z(
        P1_U3545) );
  AOI21_X1 U10906 ( .B1(n9934), .B2(n9736), .A(n9735), .ZN(n9737) );
  OAI211_X1 U10907 ( .C1(n9739), .C2(n9962), .A(n9738), .B(n9737), .ZN(n9811)
         );
  MUX2_X1 U10908 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9811), .S(n9977), .Z(
        P1_U3544) );
  AOI22_X1 U10909 ( .A1(n9741), .A2(n9935), .B1(n9934), .B2(n9740), .ZN(n9742)
         );
  OAI211_X1 U10910 ( .C1(n9744), .C2(n9962), .A(n9743), .B(n9742), .ZN(n9812)
         );
  MUX2_X1 U10911 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9812), .S(n9977), .Z(
        P1_U3543) );
  AOI22_X1 U10912 ( .A1(n9746), .A2(n9935), .B1(n9934), .B2(n9745), .ZN(n9747)
         );
  OAI211_X1 U10913 ( .C1(n9749), .C2(n9962), .A(n9748), .B(n9747), .ZN(n9813)
         );
  MUX2_X1 U10914 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9813), .S(n9977), .Z(
        P1_U3542) );
  OR2_X1 U10915 ( .A1(n9750), .A2(n9962), .ZN(n9756) );
  OAI21_X1 U10916 ( .B1(n9752), .B2(n9965), .A(n9751), .ZN(n9753) );
  NOR2_X1 U10917 ( .A1(n9754), .A2(n9753), .ZN(n9755) );
  NAND2_X1 U10918 ( .A1(n9756), .A2(n9755), .ZN(n9814) );
  MUX2_X1 U10919 ( .A(n9814), .B(P1_REG1_REG_18__SCAN_IN), .S(n9974), .Z(
        P1_U3541) );
  AOI211_X1 U10920 ( .C1(n9934), .C2(n9759), .A(n9758), .B(n9757), .ZN(n9760)
         );
  OAI21_X1 U10921 ( .B1(n9962), .B2(n9761), .A(n9760), .ZN(n9815) );
  MUX2_X1 U10922 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9815), .S(n9977), .Z(
        P1_U3540) );
  AOI211_X1 U10923 ( .C1(n9934), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9765)
         );
  OAI21_X1 U10924 ( .B1(n9962), .B2(n9766), .A(n9765), .ZN(n9816) );
  MUX2_X1 U10925 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9816), .S(n9977), .Z(
        P1_U3539) );
  OAI22_X1 U10926 ( .A1(n9767), .A2(n9944), .B1(n8028), .B2(n9965), .ZN(n9768)
         );
  AOI21_X1 U10927 ( .B1(n9769), .B2(n9949), .A(n9768), .ZN(n9770) );
  NAND2_X1 U10928 ( .A1(n9771), .A2(n9770), .ZN(n9817) );
  MUX2_X1 U10929 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9817), .S(n9977), .Z(
        P1_U3538) );
  AOI211_X1 U10930 ( .C1(n9934), .C2(n9774), .A(n9773), .B(n9772), .ZN(n9775)
         );
  OAI21_X1 U10931 ( .B1(n9962), .B2(n9776), .A(n9775), .ZN(n9818) );
  MUX2_X1 U10932 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9818), .S(n9977), .Z(
        P1_U3537) );
  AOI211_X1 U10933 ( .C1(n9934), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9780)
         );
  OAI21_X1 U10934 ( .B1(n9962), .B2(n9781), .A(n9780), .ZN(n9821) );
  MUX2_X1 U10935 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9821), .S(n9977), .Z(
        P1_U3535) );
  AND2_X1 U10936 ( .A1(n9782), .A2(n9949), .ZN(n9786) );
  OAI22_X1 U10937 ( .A1(n9784), .A2(n9944), .B1(n9783), .B2(n9965), .ZN(n9785)
         );
  MUX2_X1 U10938 ( .A(n9822), .B(P1_REG1_REG_11__SCAN_IN), .S(n9974), .Z(
        P1_U3534) );
  INV_X1 U10939 ( .A(n9788), .ZN(n9793) );
  AOI21_X1 U10940 ( .B1(n9934), .B2(n9790), .A(n9789), .ZN(n9791) );
  OAI211_X1 U10941 ( .C1(n9793), .C2(n9939), .A(n9792), .B(n9791), .ZN(n9823)
         );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9823), .S(n9977), .Z(
        P1_U3533) );
  INV_X1 U10943 ( .A(n9794), .ZN(n9799) );
  AOI22_X1 U10944 ( .A1(n9796), .A2(n9935), .B1(n9934), .B2(n9795), .ZN(n9797)
         );
  OAI211_X1 U10945 ( .C1(n9939), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9824)
         );
  MUX2_X1 U10946 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9824), .S(n9977), .Z(
        P1_U3532) );
  MUX2_X1 U10947 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9800), .S(n9977), .Z(
        P1_U3525) );
  MUX2_X1 U10948 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9801), .S(n10175), .Z(
        P1_U3522) );
  MUX2_X1 U10949 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9802), .S(n10175), .Z(
        P1_U3521) );
  MUX2_X1 U10950 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9803), .S(n10175), .Z(
        P1_U3520) );
  MUX2_X1 U10951 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9804), .S(n10175), .Z(
        P1_U3519) );
  MUX2_X1 U10952 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9805), .S(n10175), .Z(
        P1_U3518) );
  MUX2_X1 U10953 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9806), .S(n10175), .Z(
        P1_U3517) );
  MUX2_X1 U10954 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9807), .S(n10175), .Z(
        P1_U3516) );
  MUX2_X1 U10955 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9808), .S(n10175), .Z(
        P1_U3515) );
  MUX2_X1 U10956 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9809), .S(n10175), .Z(
        P1_U3514) );
  MUX2_X1 U10957 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9810), .S(n10175), .Z(
        P1_U3513) );
  MUX2_X1 U10958 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9811), .S(n10175), .Z(
        P1_U3512) );
  MUX2_X1 U10959 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9812), .S(n10175), .Z(
        P1_U3511) );
  MUX2_X1 U10960 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9813), .S(n10175), .Z(
        P1_U3510) );
  MUX2_X1 U10961 ( .A(n9814), .B(P1_REG0_REG_18__SCAN_IN), .S(n10173), .Z(
        P1_U3508) );
  MUX2_X1 U10962 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9815), .S(n10175), .Z(
        P1_U3505) );
  MUX2_X1 U10963 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9816), .S(n10175), .Z(
        P1_U3502) );
  MUX2_X1 U10964 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9817), .S(n10175), .Z(
        P1_U3499) );
  MUX2_X1 U10965 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9818), .S(n10175), .Z(
        P1_U3496) );
  INV_X1 U10966 ( .A(n9819), .ZN(n9820) );
  MUX2_X1 U10967 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9820), .S(n10175), .Z(
        P1_U3493) );
  MUX2_X1 U10968 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9821), .S(n10175), .Z(
        P1_U3490) );
  MUX2_X1 U10969 ( .A(n9822), .B(P1_REG0_REG_11__SCAN_IN), .S(n10173), .Z(
        P1_U3487) );
  MUX2_X1 U10970 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9823), .S(n10175), .Z(
        P1_U3484) );
  MUX2_X1 U10971 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n9824), .S(n10175), .Z(
        P1_U3481) );
  MUX2_X1 U10972 ( .A(P1_D_REG_1__SCAN_IN), .B(n9825), .S(n9925), .Z(P1_U3441)
         );
  MUX2_X1 U10973 ( .A(P1_D_REG_0__SCAN_IN), .B(n9826), .S(n9925), .Z(P1_U3440)
         );
  NOR4_X1 U10974 ( .A1(n4405), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6061), .A4(
        P1_U3084), .ZN(n9827) );
  AOI21_X1 U10975 ( .B1(n9828), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9827), .ZN(
        n9829) );
  OAI21_X1 U10976 ( .B1(n9830), .B2(n9840), .A(n9829), .ZN(P1_U3322) );
  OAI222_X1 U10977 ( .A1(n9837), .A2(n9833), .B1(P1_U3084), .B2(n9832), .C1(
        n9840), .C2(n9831), .ZN(P1_U3324) );
  OAI222_X1 U10978 ( .A1(n9837), .A2(n9836), .B1(P1_U3084), .B2(n9835), .C1(
        n9840), .C2(n9834), .ZN(P1_U3326) );
  OAI222_X1 U10979 ( .A1(n9841), .A2(P1_U3084), .B1(n9840), .B2(n9839), .C1(
        n9838), .C2(n9837), .ZN(P1_U3327) );
  MUX2_X1 U10980 ( .A(n9842), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10981 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9843) );
  AOI21_X1 U10982 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9843), .ZN(n10150) );
  NOR2_X1 U10983 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9844) );
  AOI21_X1 U10984 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9844), .ZN(n10153) );
  NOR2_X1 U10985 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9845) );
  AOI21_X1 U10986 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9845), .ZN(n10156) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9846) );
  AOI21_X1 U10988 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9846), .ZN(n10159) );
  NOR2_X1 U10989 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9847) );
  AOI21_X1 U10990 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9847), .ZN(n10162) );
  NOR2_X1 U10991 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9854) );
  XNOR2_X1 U10992 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10486) );
  NAND2_X1 U10993 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9852) );
  XOR2_X1 U10994 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10484) );
  NAND2_X1 U10995 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9850) );
  XOR2_X1 U10996 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10482) );
  AOI21_X1 U10997 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10143) );
  INV_X1 U10998 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9848) );
  NAND3_X1 U10999 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U11000 ( .A1(n10482), .A2(n10481), .ZN(n9849) );
  NAND2_X1 U11001 ( .A1(n9850), .A2(n9849), .ZN(n10483) );
  NAND2_X1 U11002 ( .A1(n10484), .A2(n10483), .ZN(n9851) );
  NAND2_X1 U11003 ( .A1(n9852), .A2(n9851), .ZN(n10485) );
  NOR2_X1 U11004 ( .A1(n10486), .A2(n10485), .ZN(n9853) );
  NOR2_X1 U11005 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9855), .ZN(n10467) );
  NAND2_X1 U11006 ( .A1(n9857), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9859) );
  XOR2_X1 U11007 ( .A(n9857), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10466) );
  NAND2_X1 U11008 ( .A1(n10466), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U11009 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9860), .ZN(n9862) );
  NAND2_X1 U11010 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10480), .ZN(n9861) );
  NAND2_X1 U11011 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9863), .ZN(n9865) );
  NAND2_X1 U11012 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10478), .ZN(n9864) );
  AND2_X1 U11013 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9866), .ZN(n9867) );
  NAND2_X1 U11014 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9868) );
  OAI21_X1 U11015 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9868), .ZN(n10170) );
  NAND2_X1 U11016 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9869) );
  OAI21_X1 U11017 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9869), .ZN(n10167) );
  NOR2_X1 U11018 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9870) );
  AOI21_X1 U11019 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9870), .ZN(n10164) );
  NAND2_X1 U11020 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  NAND2_X1 U11021 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  NAND2_X1 U11022 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  OAI21_X1 U11023 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10151), .ZN(n10149) );
  NAND2_X1 U11024 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  NOR2_X1 U11025 ( .A1(n10473), .A2(n10472), .ZN(n9871) );
  NAND2_X1 U11026 ( .A1(n10473), .A2(n10472), .ZN(n10471) );
  XNOR2_X1 U11027 ( .A(n9872), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n9873) );
  XNOR2_X1 U11028 ( .A(n9874), .B(n9873), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11029 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11030 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11031 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9876) );
  OAI22_X1 U11032 ( .A1(n9923), .A2(n9876), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9875), .ZN(n9881) );
  AOI211_X1 U11033 ( .C1(n9879), .C2(n9878), .A(n9877), .B(n9893), .ZN(n9880)
         );
  AOI211_X1 U11034 ( .C1(n9910), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9887)
         );
  OAI211_X1 U11035 ( .C1(n9885), .C2(n9884), .A(n9917), .B(n9883), .ZN(n9886)
         );
  NAND2_X1 U11036 ( .A1(n9887), .A2(n9886), .ZN(P1_U3242) );
  NAND2_X1 U11037 ( .A1(n9917), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9889) );
  OAI21_X1 U11038 ( .B1(n9889), .B2(n9902), .A(n9888), .ZN(n9898) );
  INV_X1 U11039 ( .A(n9890), .ZN(n9897) );
  MUX2_X1 U11040 ( .A(n6911), .B(P1_REG2_REG_8__SCAN_IN), .S(n9899), .Z(n9892)
         );
  NAND3_X1 U11041 ( .A1(n4809), .A2(n4487), .A3(n9892), .ZN(n9894) );
  AOI21_X1 U11042 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(n9896) );
  AOI211_X1 U11043 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9906)
         );
  AOI211_X1 U11044 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9904)
         );
  INV_X1 U11045 ( .A(n9904), .ZN(n9905) );
  OAI211_X1 U11046 ( .C1(n4523), .C2(n9923), .A(n9906), .B(n9905), .ZN(
        P1_U3249) );
  INV_X1 U11047 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9922) );
  INV_X1 U11048 ( .A(n9907), .ZN(n9908) );
  AOI21_X1 U11049 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9921) );
  OAI21_X1 U11050 ( .B1(n9912), .B2(n6392), .A(n9911), .ZN(n9919) );
  OAI21_X1 U11051 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  AOI22_X1 U11052 ( .A1(n9919), .A2(n9918), .B1(n9917), .B2(n9916), .ZN(n9920)
         );
  OAI211_X1 U11053 ( .C1(n9923), .C2(n9922), .A(n9921), .B(n9920), .ZN(
        P1_U3255) );
  AND2_X1 U11054 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9927), .ZN(P1_U3292) );
  AND2_X1 U11055 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9927), .ZN(P1_U3293) );
  AND2_X1 U11056 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9927), .ZN(P1_U3294) );
  AND2_X1 U11057 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9927), .ZN(P1_U3295) );
  AND2_X1 U11058 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9927), .ZN(P1_U3296) );
  AND2_X1 U11059 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9927), .ZN(P1_U3297) );
  AND2_X1 U11060 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9927), .ZN(P1_U3298) );
  INV_X1 U11061 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10423) );
  NOR2_X1 U11062 ( .A1(n9926), .A2(n10423), .ZN(P1_U3299) );
  AND2_X1 U11063 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9927), .ZN(P1_U3300) );
  AND2_X1 U11064 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9927), .ZN(P1_U3301) );
  AND2_X1 U11065 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9927), .ZN(P1_U3302) );
  INV_X1 U11066 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10242) );
  NOR2_X1 U11067 ( .A1(n9926), .A2(n10242), .ZN(P1_U3303) );
  INV_X1 U11068 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U11069 ( .A1(n9926), .A2(n10406), .ZN(P1_U3304) );
  INV_X1 U11070 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U11071 ( .A1(n9926), .A2(n10230), .ZN(P1_U3305) );
  AND2_X1 U11072 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9927), .ZN(P1_U3306) );
  AND2_X1 U11073 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9927), .ZN(P1_U3307) );
  INV_X1 U11074 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U11075 ( .A1(n9926), .A2(n10244), .ZN(P1_U3308) );
  AND2_X1 U11076 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9927), .ZN(P1_U3309) );
  INV_X1 U11077 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10450) );
  NOR2_X1 U11078 ( .A1(n9926), .A2(n10450), .ZN(P1_U3310) );
  AND2_X1 U11079 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9927), .ZN(P1_U3311) );
  INV_X1 U11080 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10309) );
  NOR2_X1 U11081 ( .A1(n9926), .A2(n10309), .ZN(P1_U3312) );
  AND2_X1 U11082 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9927), .ZN(P1_U3313) );
  AND2_X1 U11083 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9927), .ZN(P1_U3314) );
  AND2_X1 U11084 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9927), .ZN(P1_U3315) );
  INV_X1 U11085 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10290) );
  NOR2_X1 U11086 ( .A1(n9926), .A2(n10290), .ZN(P1_U3316) );
  AND2_X1 U11087 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9927), .ZN(P1_U3317) );
  AND2_X1 U11088 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9927), .ZN(P1_U3318) );
  AND2_X1 U11089 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9927), .ZN(P1_U3319) );
  INV_X1 U11090 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10377) );
  NOR2_X1 U11091 ( .A1(n9926), .A2(n10377), .ZN(P1_U3320) );
  AND2_X1 U11092 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9927), .ZN(P1_U3321) );
  OAI211_X1 U11093 ( .C1(n9930), .C2(n9939), .A(n9929), .B(n9928), .ZN(n9931)
         );
  NOR2_X1 U11094 ( .A1(n9932), .A2(n9931), .ZN(n9960) );
  INV_X1 U11095 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U11096 ( .A1(n10175), .A2(n9960), .B1(n10317), .B2(n10173), .ZN(
        P1_U3457) );
  AOI22_X1 U11097 ( .A1(n9936), .A2(n9935), .B1(n9934), .B2(n9933), .ZN(n9937)
         );
  OAI211_X1 U11098 ( .C1(n9940), .C2(n9939), .A(n9938), .B(n9937), .ZN(n9941)
         );
  INV_X1 U11099 ( .A(n9941), .ZN(n9961) );
  INV_X1 U11100 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U11101 ( .A1(n10175), .A2(n9961), .B1(n9942), .B2(n10173), .ZN(
        P1_U3463) );
  OAI22_X1 U11102 ( .A1(n9945), .A2(n9944), .B1(n5010), .B2(n9965), .ZN(n9947)
         );
  AOI211_X1 U11103 ( .C1(n9949), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9973)
         );
  INV_X1 U11104 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11105 ( .A1(n10175), .A2(n9973), .B1(n9950), .B2(n10173), .ZN(
        P1_U3472) );
  INV_X1 U11106 ( .A(n9951), .ZN(n9957) );
  INV_X1 U11107 ( .A(n9952), .ZN(n9953) );
  NAND3_X1 U11108 ( .A1(n9955), .A2(n9954), .A3(n9953), .ZN(n9956) );
  AOI21_X1 U11109 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9976) );
  INV_X1 U11110 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11111 ( .A1(n10175), .A2(n9976), .B1(n9959), .B2(n10173), .ZN(
        P1_U3475) );
  AOI22_X1 U11112 ( .A1(n9977), .A2(n9960), .B1(n6824), .B2(n9974), .ZN(
        P1_U3524) );
  AOI22_X1 U11113 ( .A1(n9977), .A2(n9961), .B1(n6826), .B2(n9974), .ZN(
        P1_U3526) );
  OR2_X1 U11114 ( .A1(n9963), .A2(n9962), .ZN(n9970) );
  OAI21_X1 U11115 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(n9967) );
  NOR2_X1 U11116 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  AND2_X1 U11117 ( .A1(n9970), .A2(n9969), .ZN(n10172) );
  AOI22_X1 U11118 ( .A1(n9977), .A2(n10172), .B1(n9971), .B2(n9974), .ZN(
        P1_U3528) );
  AOI22_X1 U11119 ( .A1(n9977), .A2(n9973), .B1(n9972), .B2(n9974), .ZN(
        P1_U3529) );
  AOI22_X1 U11120 ( .A1(n9977), .A2(n9976), .B1(n9975), .B2(n9974), .ZN(
        P1_U3530) );
  AOI22_X1 U11121 ( .A1(n9979), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9978), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9989) );
  AOI21_X1 U11122 ( .B1(n9981), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9980), .ZN(
        n9988) );
  NOR2_X1 U11123 ( .A1(n9982), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9986) );
  OAI21_X1 U11124 ( .B1(n9984), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9983), .ZN(
        n9985) );
  OAI21_X1 U11125 ( .B1(n9986), .B2(n9985), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9987) );
  OAI211_X1 U11126 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9989), .A(n9988), .B(
        n9987), .ZN(P2_U3245) );
  INV_X1 U11127 ( .A(n7612), .ZN(n9991) );
  OAI21_X1 U11128 ( .B1(n9991), .B2(n9990), .A(n4441), .ZN(n9992) );
  XNOR2_X1 U11129 ( .A(n9992), .B(n4399), .ZN(n10109) );
  NAND2_X1 U11130 ( .A1(n7635), .A2(n9993), .ZN(n9994) );
  XNOR2_X1 U11131 ( .A(n9994), .B(n4399), .ZN(n9996) );
  OAI222_X1 U11132 ( .A1(n10000), .A2(n9999), .B1(n9998), .B2(n9997), .C1(
        n9996), .C2(n9995), .ZN(n10107) );
  AOI21_X1 U11133 ( .B1(n10001), .B2(n10109), .A(n10107), .ZN(n10013) );
  AOI22_X1 U11134 ( .A1(n10036), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10003), 
        .B2(n10002), .ZN(n10004) );
  OAI21_X1 U11135 ( .B1(n10031), .B2(n10105), .A(n10004), .ZN(n10005) );
  INV_X1 U11136 ( .A(n10005), .ZN(n10012) );
  INV_X1 U11137 ( .A(n10006), .ZN(n10010) );
  INV_X1 U11138 ( .A(n10007), .ZN(n10008) );
  OAI21_X1 U11139 ( .B1(n10105), .B2(n4471), .A(n10008), .ZN(n10106) );
  INV_X1 U11140 ( .A(n10106), .ZN(n10009) );
  AOI22_X1 U11141 ( .A1(n10109), .A2(n10010), .B1(n10029), .B2(n10009), .ZN(
        n10011) );
  OAI211_X1 U11142 ( .C1(n10036), .C2(n10013), .A(n10012), .B(n10011), .ZN(
        P2_U3286) );
  AOI222_X1 U11143 ( .A1(n10020), .A2(n10019), .B1(n10018), .B2(n10017), .C1(
        n10016), .C2(n10015), .ZN(n10064) );
  XNOR2_X1 U11144 ( .A(n10021), .B(n10022), .ZN(n10066) );
  INV_X1 U11145 ( .A(n10023), .ZN(n10025) );
  AOI21_X1 U11146 ( .B1(n5163), .B2(n10025), .A(n10024), .ZN(n10062) );
  OAI22_X1 U11147 ( .A1(n10027), .A2(n6674), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10026), .ZN(n10028) );
  AOI21_X1 U11148 ( .B1(n10029), .B2(n10062), .A(n10028), .ZN(n10030) );
  OAI21_X1 U11149 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10033) );
  AOI21_X1 U11150 ( .B1(n10034), .B2(n10066), .A(n10033), .ZN(n10035) );
  OAI21_X1 U11151 ( .B1(n10036), .B2(n10064), .A(n10035), .ZN(P2_U3293) );
  AND2_X1 U11152 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10042), .ZN(P2_U3297) );
  AND2_X1 U11153 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10042), .ZN(P2_U3298) );
  AND2_X1 U11154 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10042), .ZN(P2_U3299) );
  AND2_X1 U11155 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10042), .ZN(P2_U3300) );
  AND2_X1 U11156 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10042), .ZN(P2_U3301) );
  AND2_X1 U11157 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10042), .ZN(P2_U3302) );
  INV_X1 U11158 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U11159 ( .A1(n10039), .A2(n10363), .ZN(P2_U3303) );
  AND2_X1 U11160 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10042), .ZN(P2_U3304) );
  AND2_X1 U11161 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10042), .ZN(P2_U3305) );
  INV_X1 U11162 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U11163 ( .A1(n10039), .A2(n10407), .ZN(P2_U3306) );
  AND2_X1 U11164 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10042), .ZN(P2_U3307) );
  AND2_X1 U11165 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10042), .ZN(P2_U3308) );
  AND2_X1 U11166 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10042), .ZN(P2_U3309) );
  INV_X1 U11167 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U11168 ( .A1(n10039), .A2(n10389), .ZN(P2_U3310) );
  INV_X1 U11169 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U11170 ( .A1(n10039), .A2(n10429), .ZN(P2_U3311) );
  INV_X1 U11171 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U11172 ( .A1(n10039), .A2(n10255), .ZN(P2_U3312) );
  AND2_X1 U11173 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10042), .ZN(P2_U3313) );
  AND2_X1 U11174 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10042), .ZN(P2_U3314) );
  AND2_X1 U11175 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10042), .ZN(P2_U3315) );
  AND2_X1 U11176 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10042), .ZN(P2_U3316) );
  AND2_X1 U11177 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10042), .ZN(P2_U3317) );
  AND2_X1 U11178 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10042), .ZN(P2_U3318) );
  INV_X1 U11179 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10303) );
  NOR2_X1 U11180 ( .A1(n10039), .A2(n10303), .ZN(P2_U3319) );
  AND2_X1 U11181 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10042), .ZN(P2_U3320) );
  AND2_X1 U11182 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10042), .ZN(P2_U3321) );
  AND2_X1 U11183 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10042), .ZN(P2_U3322) );
  AND2_X1 U11184 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10042), .ZN(P2_U3323) );
  AND2_X1 U11185 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10042), .ZN(P2_U3324) );
  AND2_X1 U11186 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10042), .ZN(P2_U3325) );
  INV_X1 U11187 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U11188 ( .A1(n10039), .A2(n10404), .ZN(P2_U3326) );
  AOI22_X1 U11189 ( .A1(n10044), .A2(n10041), .B1(n10040), .B2(n10042), .ZN(
        P2_U3437) );
  AOI22_X1 U11190 ( .A1(n10044), .A2(n10043), .B1(n10289), .B2(n10042), .ZN(
        P2_U3438) );
  NOR2_X1 U11191 ( .A1(n10046), .A2(n10045), .ZN(n10048) );
  AOI211_X1 U11192 ( .C1(n10117), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10123) );
  INV_X1 U11193 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U11194 ( .A1(n10121), .A2(n10123), .B1(n10351), .B2(n10119), .ZN(
        P2_U3451) );
  OAI21_X1 U11195 ( .B1(n10051), .B2(n10111), .A(n10050), .ZN(n10053) );
  AOI211_X1 U11196 ( .C1(n10054), .C2(n10117), .A(n10053), .B(n10052), .ZN(
        n10125) );
  INV_X1 U11197 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11198 ( .A1(n10121), .A2(n10125), .B1(n10055), .B2(n10119), .ZN(
        P2_U3454) );
  AND2_X1 U11199 ( .A1(n10056), .A2(n10117), .ZN(n10061) );
  NOR2_X1 U11200 ( .A1(n10057), .A2(n10111), .ZN(n10058) );
  NOR4_X1 U11201 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10127) );
  INV_X1 U11202 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U11203 ( .A1(n10121), .A2(n10127), .B1(n10434), .B2(n10119), .ZN(
        P2_U3457) );
  AOI22_X1 U11204 ( .A1(n10062), .A2(n10097), .B1(n10096), .B2(n5163), .ZN(
        n10063) );
  NAND2_X1 U11205 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  AOI21_X1 U11206 ( .B1(n10066), .B2(n10117), .A(n10065), .ZN(n10129) );
  INV_X1 U11207 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11208 ( .A1(n10121), .A2(n10129), .B1(n10067), .B2(n10119), .ZN(
        P2_U3460) );
  INV_X1 U11209 ( .A(n10068), .ZN(n10073) );
  OAI21_X1 U11210 ( .B1(n10070), .B2(n10111), .A(n10069), .ZN(n10071) );
  AOI211_X1 U11211 ( .C1(n10073), .C2(n10117), .A(n10072), .B(n10071), .ZN(
        n10130) );
  INV_X1 U11212 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U11213 ( .A1(n10121), .A2(n10130), .B1(n10270), .B2(n10119), .ZN(
        P2_U3463) );
  OAI22_X1 U11214 ( .A1(n10075), .A2(n10113), .B1(n10074), .B2(n10111), .ZN(
        n10077) );
  AOI211_X1 U11215 ( .C1(n10078), .C2(n10117), .A(n10077), .B(n10076), .ZN(
        n10131) );
  INV_X1 U11216 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U11217 ( .A1(n10121), .A2(n10131), .B1(n10079), .B2(n10119), .ZN(
        P2_U3469) );
  AOI21_X1 U11218 ( .B1(n10096), .B2(n10081), .A(n10080), .ZN(n10083) );
  OAI211_X1 U11219 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10086) );
  INV_X1 U11220 ( .A(n10086), .ZN(n10133) );
  INV_X1 U11221 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U11222 ( .A1(n10121), .A2(n10133), .B1(n10087), .B2(n10119), .ZN(
        P2_U3472) );
  AOI22_X1 U11223 ( .A1(n10089), .A2(n10097), .B1(n10096), .B2(n10088), .ZN(
        n10090) );
  OAI21_X1 U11224 ( .B1(n10091), .B2(n10102), .A(n10090), .ZN(n10092) );
  NOR2_X1 U11225 ( .A1(n10093), .A2(n10092), .ZN(n10135) );
  INV_X1 U11226 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11227 ( .A1(n10121), .A2(n10135), .B1(n10094), .B2(n10119), .ZN(
        P2_U3475) );
  AOI22_X1 U11228 ( .A1(n10098), .A2(n10097), .B1(n10096), .B2(n10095), .ZN(
        n10099) );
  OAI211_X1 U11229 ( .C1(n10102), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10103) );
  INV_X1 U11230 ( .A(n10103), .ZN(n10137) );
  INV_X1 U11231 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U11232 ( .A1(n10121), .A2(n10137), .B1(n10104), .B2(n10119), .ZN(
        P2_U3478) );
  OAI22_X1 U11233 ( .A1(n10106), .A2(n10113), .B1(n10105), .B2(n10111), .ZN(
        n10108) );
  AOI211_X1 U11234 ( .C1(n10117), .C2(n10109), .A(n10108), .B(n10107), .ZN(
        n10138) );
  INV_X1 U11235 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11236 ( .A1(n10121), .A2(n10138), .B1(n10110), .B2(n10119), .ZN(
        P2_U3481) );
  OAI22_X1 U11237 ( .A1(n10114), .A2(n10113), .B1(n10112), .B2(n10111), .ZN(
        n10116) );
  AOI211_X1 U11238 ( .C1(n10118), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10141) );
  INV_X1 U11239 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U11240 ( .A1(n10121), .A2(n10141), .B1(n10120), .B2(n10119), .ZN(
        P2_U3484) );
  INV_X1 U11241 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U11242 ( .A1(n10142), .A2(n10123), .B1(n10122), .B2(n10139), .ZN(
        P2_U3520) );
  INV_X1 U11243 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11244 ( .A1(n10142), .A2(n10125), .B1(n10124), .B2(n10139), .ZN(
        P2_U3521) );
  AOI22_X1 U11245 ( .A1(n10142), .A2(n10127), .B1(n10126), .B2(n10139), .ZN(
        P2_U3522) );
  AOI22_X1 U11246 ( .A1(n10142), .A2(n10129), .B1(n10128), .B2(n10139), .ZN(
        P2_U3523) );
  AOI22_X1 U11247 ( .A1(n10142), .A2(n10130), .B1(n6697), .B2(n10139), .ZN(
        P2_U3524) );
  AOI22_X1 U11248 ( .A1(n10142), .A2(n10131), .B1(n6700), .B2(n10139), .ZN(
        P2_U3526) );
  AOI22_X1 U11249 ( .A1(n10142), .A2(n10133), .B1(n10132), .B2(n10139), .ZN(
        P2_U3527) );
  AOI22_X1 U11250 ( .A1(n10142), .A2(n10135), .B1(n10134), .B2(n10139), .ZN(
        P2_U3528) );
  AOI22_X1 U11251 ( .A1(n10142), .A2(n10137), .B1(n10136), .B2(n10139), .ZN(
        P2_U3529) );
  AOI22_X1 U11252 ( .A1(n10142), .A2(n10138), .B1(n10335), .B2(n10139), .ZN(
        P2_U3530) );
  AOI22_X1 U11253 ( .A1(n10142), .A2(n10141), .B1(n10140), .B2(n10139), .ZN(
        P2_U3531) );
  INV_X1 U11254 ( .A(n10143), .ZN(n10144) );
  NAND2_X1 U11255 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  XNOR2_X1 U11256 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10146), .ZN(ADD_1071_U5)
         );
  INV_X1 U11257 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U11258 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10147), .B2(n6788), .ZN(ADD_1071_U46) );
  OAI21_X1 U11259 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(ADD_1071_U56) );
  OAI21_X1 U11260 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(ADD_1071_U57) );
  OAI21_X1 U11261 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(ADD_1071_U58) );
  OAI21_X1 U11262 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(ADD_1071_U59) );
  OAI21_X1 U11263 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(ADD_1071_U60) );
  OAI21_X1 U11264 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(ADD_1071_U61) );
  AOI21_X1 U11265 ( .B1(n10168), .B2(n10167), .A(n10166), .ZN(ADD_1071_U62) );
  AOI21_X1 U11266 ( .B1(n10171), .B2(n10170), .A(n10169), .ZN(ADD_1071_U63) );
  INV_X1 U11267 ( .A(n10172), .ZN(n10174) );
  AOI22_X1 U11268 ( .A1(n10175), .A2(n10174), .B1(P1_REG0_REG_5__SCAN_IN), 
        .B2(n10173), .ZN(n10464) );
  NAND4_X1 U11269 ( .A1(SI_27_), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P2_REG3_REG_12__SCAN_IN), .A4(n10176), .ZN(n10198) );
  NAND4_X1 U11270 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(P1_REG0_REG_14__SCAN_IN), 
        .A3(P1_REG2_REG_30__SCAN_IN), .A4(n6676), .ZN(n10197) );
  NAND4_X1 U11271 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), 
        .A3(P2_REG2_REG_24__SCAN_IN), .A4(n10256), .ZN(n10177) );
  NOR3_X1 U11272 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(n10177), .ZN(n10183) );
  NAND4_X1 U11273 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_REG3_REG_28__SCAN_IN), .A4(n10241), .ZN(n10181) );
  NAND4_X1 U11274 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .A3(n10261), .A4(n10262), .ZN(n10179) );
  NAND4_X1 U11275 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_REG0_REG_13__SCAN_IN), 
        .A3(P2_REG3_REG_7__SCAN_IN), .A4(n10233), .ZN(n10178) );
  OR4_X1 U11276 ( .A1(n10273), .A2(P2_DATAO_REG_30__SCAN_IN), .A3(n10179), 
        .A4(n10178), .ZN(n10180) );
  NOR4_X1 U11277 ( .A1(n10181), .A2(n10180), .A3(P1_DATAO_REG_28__SCAN_IN), 
        .A4(P2_IR_REG_4__SCAN_IN), .ZN(n10182) );
  INV_X1 U11278 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10258) );
  NAND4_X1 U11279 ( .A1(SI_21_), .A2(n10183), .A3(n10182), .A4(n10258), .ZN(
        n10196) );
  NAND4_X1 U11280 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), 
        .A3(P2_IR_REG_1__SCAN_IN), .A4(n10320), .ZN(n10184) );
  NOR3_X1 U11281 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), 
        .A3(n10184), .ZN(n10194) );
  NAND4_X1 U11282 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(SI_29_), .A3(n5633), 
        .A4(n10335), .ZN(n10192) );
  NAND4_X1 U11283 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(SI_19_), .A3(
        P1_REG0_REG_1__SCAN_IN), .A4(P2_REG2_REG_30__SCAN_IN), .ZN(n10191) );
  NOR4_X1 U11284 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), 
        .A3(P2_REG2_REG_23__SCAN_IN), .A4(n6433), .ZN(n10189) );
  NOR4_X1 U11285 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .A3(P2_REG2_REG_12__SCAN_IN), .A4(P2_REG0_REG_4__SCAN_IN), .ZN(n10186)
         );
  NOR4_X1 U11286 ( .A1(SI_2_), .A2(P1_REG1_REG_25__SCAN_IN), .A3(
        P2_REG2_REG_16__SCAN_IN), .A4(n10289), .ZN(n10185) );
  NAND3_X1 U11287 ( .A1(n10302), .A2(n10186), .A3(n10185), .ZN(n10187) );
  NOR4_X1 U11288 ( .A1(n10187), .A2(n10304), .A3(P1_D_REG_11__SCAN_IN), .A4(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U11289 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NOR3_X1 U11290 ( .A1(n10192), .A2(n10191), .A3(n10190), .ZN(n10193) );
  NAND4_X1 U11291 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .A3(n10194), .A4(n10193), .ZN(n10195) );
  NOR4_X1 U11292 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10225) );
  NAND4_X1 U11293 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(n10473), .A4(n10479), .ZN(n10199) );
  NOR4_X1 U11294 ( .A1(SI_14_), .A2(P2_ADDR_REG_3__SCAN_IN), .A3(
        P1_ADDR_REG_2__SCAN_IN), .A4(n10199), .ZN(n10209) );
  NAND4_X1 U11295 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(SI_6_), .A3(
        P1_REG3_REG_0__SCAN_IN), .A4(P2_REG0_REG_31__SCAN_IN), .ZN(n10203) );
  NAND4_X1 U11296 ( .A1(P1_D_REG_0__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P2_IR_REG_14__SCAN_IN), .A4(P2_REG1_REG_19__SCAN_IN), .ZN(n10202) );
  NAND4_X1 U11297 ( .A1(SI_7_), .A2(P2_DATAO_REG_7__SCAN_IN), .A3(
        P1_REG1_REG_13__SCAN_IN), .A4(n10450), .ZN(n10201) );
  NAND4_X1 U11298 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        n5543), .A4(n10404), .ZN(n10200) );
  NOR4_X1 U11299 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10208) );
  NOR4_X1 U11300 ( .A1(n10441), .A2(P1_REG3_REG_25__SCAN_IN), .A3(
        P1_IR_REG_13__SCAN_IN), .A4(n5423), .ZN(n10207) );
  AND4_X1 U11301 ( .A1(n10205), .A2(n10204), .A3(P1_DATAO_REG_1__SCAN_IN), 
        .A4(P1_REG0_REG_19__SCAN_IN), .ZN(n10206) );
  NAND4_X1 U11302 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10223) );
  NAND4_X1 U11303 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .A4(n9050), .ZN(n10222) );
  NAND4_X1 U11304 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), 
        .A3(n10430), .A4(n10210), .ZN(n10221) );
  NOR4_X1 U11305 ( .A1(SI_4_), .A2(P1_REG2_REG_11__SCAN_IN), .A3(n6507), .A4(
        n6911), .ZN(n10219) );
  NOR4_X1 U11306 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(SI_10_), .A3(
        P2_REG1_REG_14__SCAN_IN), .A4(n10211), .ZN(n10218) );
  NAND4_X1 U11307 ( .A1(P1_REG0_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(n6817), .A4(n10348), .ZN(n10216) );
  INV_X1 U11308 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10387) );
  NAND4_X1 U11309 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), 
        .A3(P2_REG1_REG_4__SCAN_IN), .A4(n10387), .ZN(n10215) );
  NAND4_X1 U11310 ( .A1(SI_3_), .A2(P1_REG1_REG_0__SCAN_IN), .A3(
        P2_REG0_REG_0__SCAN_IN), .A4(P2_REG1_REG_15__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U11311 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(n10212), .ZN(n10213) );
  INV_X1 U11312 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U11313 ( .A1(n10213), .A2(P2_REG3_REG_28__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(n10375), .ZN(n10214) );
  NOR3_X1 U11314 ( .A1(n10216), .A2(n10215), .A3(n10214), .ZN(n10217) );
  NAND3_X1 U11315 ( .A1(n10219), .A2(n10218), .A3(n10217), .ZN(n10220) );
  NOR4_X1 U11316 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10224) );
  AOI21_X1 U11317 ( .B1(n10225), .B2(n10224), .A(P2_IR_REG_24__SCAN_IN), .ZN(
        n10462) );
  AOI22_X1 U11318 ( .A1(n10479), .A2(keyinput110), .B1(n10227), .B2(keyinput46), .ZN(n10226) );
  OAI221_X1 U11319 ( .B1(n10479), .B2(keyinput110), .C1(n10227), .C2(
        keyinput46), .A(n10226), .ZN(n10239) );
  AOI22_X1 U11320 ( .A1(n10230), .A2(keyinput87), .B1(keyinput71), .B2(n10229), 
        .ZN(n10228) );
  OAI221_X1 U11321 ( .B1(n10230), .B2(keyinput87), .C1(n10229), .C2(keyinput71), .A(n10228), .ZN(n10238) );
  INV_X1 U11322 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U11323 ( .A1(n10233), .A2(keyinput2), .B1(keyinput29), .B2(n10232), 
        .ZN(n10231) );
  OAI221_X1 U11324 ( .B1(n10233), .B2(keyinput2), .C1(n10232), .C2(keyinput29), 
        .A(n10231), .ZN(n10237) );
  XNOR2_X1 U11325 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput111), .ZN(n10235)
         );
  XNOR2_X1 U11326 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput27), .ZN(n10234) );
  NAND2_X1 U11327 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  NOR4_X1 U11328 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10285) );
  AOI22_X1 U11329 ( .A1(n10242), .A2(keyinput69), .B1(keyinput99), .B2(n10241), 
        .ZN(n10240) );
  OAI221_X1 U11330 ( .B1(n10242), .B2(keyinput69), .C1(n10241), .C2(keyinput99), .A(n10240), .ZN(n10253) );
  AOI22_X1 U11331 ( .A1(n10245), .A2(keyinput116), .B1(n10244), .B2(keyinput20), .ZN(n10243) );
  OAI221_X1 U11332 ( .B1(n10245), .B2(keyinput116), .C1(n10244), .C2(
        keyinput20), .A(n10243), .ZN(n10252) );
  AOI22_X1 U11333 ( .A1(n10247), .A2(keyinput103), .B1(keyinput67), .B2(n5551), 
        .ZN(n10246) );
  OAI221_X1 U11334 ( .B1(n10247), .B2(keyinput103), .C1(n5551), .C2(keyinput67), .A(n10246), .ZN(n10251) );
  AOI22_X1 U11335 ( .A1(n10249), .A2(keyinput89), .B1(keyinput12), .B2(n5612), 
        .ZN(n10248) );
  OAI221_X1 U11336 ( .B1(n10249), .B2(keyinput89), .C1(n5612), .C2(keyinput12), 
        .A(n10248), .ZN(n10250) );
  NOR4_X1 U11337 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10284) );
  AOI22_X1 U11338 ( .A1(n10256), .A2(keyinput1), .B1(n10255), .B2(keyinput115), 
        .ZN(n10254) );
  OAI221_X1 U11339 ( .B1(n10256), .B2(keyinput1), .C1(n10255), .C2(keyinput115), .A(n10254), .ZN(n10268) );
  AOI22_X1 U11340 ( .A1(n10259), .A2(keyinput112), .B1(keyinput88), .B2(n10258), .ZN(n10257) );
  OAI221_X1 U11341 ( .B1(n10259), .B2(keyinput112), .C1(n10258), .C2(
        keyinput88), .A(n10257), .ZN(n10267) );
  AOI22_X1 U11342 ( .A1(n10262), .A2(keyinput105), .B1(n10261), .B2(keyinput14), .ZN(n10260) );
  OAI221_X1 U11343 ( .B1(n10262), .B2(keyinput105), .C1(n10261), .C2(
        keyinput14), .A(n10260), .ZN(n10266) );
  XOR2_X1 U11344 ( .A(n6037), .B(keyinput80), .Z(n10264) );
  XNOR2_X1 U11345 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput126), .ZN(n10263)
         );
  NAND2_X1 U11346 ( .A1(n10264), .A2(n10263), .ZN(n10265) );
  NOR4_X1 U11347 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10283) );
  AOI22_X1 U11348 ( .A1(n10270), .A2(keyinput93), .B1(n6681), .B2(keyinput76), 
        .ZN(n10269) );
  OAI221_X1 U11349 ( .B1(n10270), .B2(keyinput93), .C1(n6681), .C2(keyinput76), 
        .A(n10269), .ZN(n10281) );
  AOI22_X1 U11350 ( .A1(n10273), .A2(keyinput123), .B1(keyinput9), .B2(n10272), 
        .ZN(n10271) );
  OAI221_X1 U11351 ( .B1(n10273), .B2(keyinput123), .C1(n10272), .C2(keyinput9), .A(n10271), .ZN(n10280) );
  XNOR2_X1 U11352 ( .A(n10274), .B(keyinput55), .ZN(n10279) );
  XNOR2_X1 U11353 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput73), .ZN(n10277) );
  XNOR2_X1 U11354 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput13), .ZN(n10276)
         );
  XNOR2_X1 U11355 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput16), .ZN(n10275) );
  NAND3_X1 U11356 ( .A1(n10277), .A2(n10276), .A3(n10275), .ZN(n10278) );
  NOR4_X1 U11357 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND4_X1 U11358 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10460) );
  AOI22_X1 U11359 ( .A1(n6433), .A2(keyinput109), .B1(keyinput101), .B2(n10287), .ZN(n10286) );
  OAI221_X1 U11360 ( .B1(n6433), .B2(keyinput109), .C1(n10287), .C2(
        keyinput101), .A(n10286), .ZN(n10298) );
  AOI22_X1 U11361 ( .A1(n10290), .A2(keyinput63), .B1(keyinput84), .B2(n10289), 
        .ZN(n10288) );
  OAI221_X1 U11362 ( .B1(n10290), .B2(keyinput63), .C1(n10289), .C2(keyinput84), .A(n10288), .ZN(n10297) );
  XOR2_X1 U11363 ( .A(n8622), .B(keyinput102), .Z(n10295) );
  INV_X1 U11364 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10291) );
  XOR2_X1 U11365 ( .A(n10291), .B(keyinput10), .Z(n10294) );
  XNOR2_X1 U11366 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput54), .ZN(n10293) );
  XNOR2_X1 U11367 ( .A(SI_2_), .B(keyinput85), .ZN(n10292) );
  NAND4_X1 U11368 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10296) );
  NOR3_X1 U11369 ( .A1(n10298), .A2(n10297), .A3(n10296), .ZN(n10346) );
  AOI22_X1 U11370 ( .A1(n10300), .A2(keyinput70), .B1(keyinput98), .B2(n8989), 
        .ZN(n10299) );
  OAI221_X1 U11371 ( .B1(n10300), .B2(keyinput70), .C1(n8989), .C2(keyinput98), 
        .A(n10299), .ZN(n10313) );
  AOI22_X1 U11372 ( .A1(n10302), .A2(keyinput41), .B1(keyinput6), .B2(n4613), 
        .ZN(n10301) );
  OAI221_X1 U11373 ( .B1(n10302), .B2(keyinput41), .C1(n4613), .C2(keyinput6), 
        .A(n10301), .ZN(n10307) );
  XNOR2_X1 U11374 ( .A(n10303), .B(keyinput97), .ZN(n10306) );
  XNOR2_X1 U11375 ( .A(n10304), .B(keyinput121), .ZN(n10305) );
  OR3_X1 U11376 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10312) );
  AOI22_X1 U11377 ( .A1(n10310), .A2(keyinput53), .B1(n10309), .B2(keyinput48), 
        .ZN(n10308) );
  OAI221_X1 U11378 ( .B1(n10310), .B2(keyinput53), .C1(n10309), .C2(keyinput48), .A(n10308), .ZN(n10311) );
  NOR3_X1 U11379 ( .A1(n10313), .A2(n10312), .A3(n10311), .ZN(n10345) );
  AOI22_X1 U11380 ( .A1(n10315), .A2(keyinput59), .B1(keyinput37), .B2(n6788), 
        .ZN(n10314) );
  OAI221_X1 U11381 ( .B1(n10315), .B2(keyinput59), .C1(n6788), .C2(keyinput37), 
        .A(n10314), .ZN(n10328) );
  AOI22_X1 U11382 ( .A1(n10318), .A2(keyinput32), .B1(keyinput28), .B2(n10317), 
        .ZN(n10316) );
  OAI221_X1 U11383 ( .B1(n10318), .B2(keyinput32), .C1(n10317), .C2(keyinput28), .A(n10316), .ZN(n10327) );
  AOI22_X1 U11384 ( .A1(n10321), .A2(keyinput74), .B1(keyinput127), .B2(n10320), .ZN(n10319) );
  OAI221_X1 U11385 ( .B1(n10321), .B2(keyinput74), .C1(n10320), .C2(
        keyinput127), .A(n10319), .ZN(n10326) );
  INV_X1 U11386 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n10322) );
  XOR2_X1 U11387 ( .A(n10322), .B(keyinput91), .Z(n10324) );
  XNOR2_X1 U11388 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput33), .ZN(n10323)
         );
  NAND2_X1 U11389 ( .A1(n10324), .A2(n10323), .ZN(n10325) );
  NOR4_X1 U11390 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10344) );
  AOI22_X1 U11391 ( .A1(n10331), .A2(keyinput25), .B1(keyinput65), .B2(n10330), 
        .ZN(n10329) );
  OAI221_X1 U11392 ( .B1(n10331), .B2(keyinput25), .C1(n10330), .C2(keyinput65), .A(n10329), .ZN(n10342) );
  AOI22_X1 U11393 ( .A1(n6045), .A2(keyinput104), .B1(keyinput81), .B2(n10333), 
        .ZN(n10332) );
  OAI221_X1 U11394 ( .B1(n6045), .B2(keyinput104), .C1(n10333), .C2(keyinput81), .A(n10332), .ZN(n10341) );
  AOI22_X1 U11395 ( .A1(n10335), .A2(keyinput31), .B1(keyinput72), .B2(n5633), 
        .ZN(n10334) );
  OAI221_X1 U11396 ( .B1(n10335), .B2(keyinput31), .C1(n5633), .C2(keyinput72), 
        .A(n10334), .ZN(n10340) );
  AOI22_X1 U11397 ( .A1(n10338), .A2(keyinput83), .B1(n10337), .B2(keyinput75), 
        .ZN(n10336) );
  OAI221_X1 U11398 ( .B1(n10338), .B2(keyinput83), .C1(n10337), .C2(keyinput75), .A(n10336), .ZN(n10339) );
  NOR4_X1 U11399 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND4_X1 U11400 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10459) );
  AOI22_X1 U11401 ( .A1(n10348), .A2(keyinput5), .B1(n6817), .B2(keyinput35), 
        .ZN(n10347) );
  OAI221_X1 U11402 ( .B1(n10348), .B2(keyinput5), .C1(n6817), .C2(keyinput35), 
        .A(n10347), .ZN(n10358) );
  AOI22_X1 U11403 ( .A1(n6911), .A2(keyinput26), .B1(n6507), .B2(keyinput114), 
        .ZN(n10349) );
  OAI221_X1 U11404 ( .B1(n6911), .B2(keyinput26), .C1(n6507), .C2(keyinput114), 
        .A(n10349), .ZN(n10357) );
  AOI22_X1 U11405 ( .A1(n10352), .A2(keyinput95), .B1(n10351), .B2(keyinput0), 
        .ZN(n10350) );
  OAI221_X1 U11406 ( .B1(n10352), .B2(keyinput95), .C1(n10351), .C2(keyinput0), 
        .A(n10350), .ZN(n10356) );
  XOR2_X1 U11407 ( .A(n6119), .B(keyinput79), .Z(n10354) );
  XNOR2_X1 U11408 ( .A(SI_3_), .B(keyinput56), .ZN(n10353) );
  NAND2_X1 U11409 ( .A1(n10354), .A2(n10353), .ZN(n10355) );
  NOR4_X1 U11410 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10402) );
  INV_X1 U11411 ( .A(SI_4_), .ZN(n10361) );
  INV_X1 U11412 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U11413 ( .A1(n10361), .A2(keyinput21), .B1(keyinput23), .B2(n10360), 
        .ZN(n10359) );
  OAI221_X1 U11414 ( .B1(n10361), .B2(keyinput21), .C1(n10360), .C2(keyinput23), .A(n10359), .ZN(n10372) );
  AOI22_X1 U11415 ( .A1(n9050), .A2(keyinput34), .B1(n10363), .B2(keyinput61), 
        .ZN(n10362) );
  OAI221_X1 U11416 ( .B1(n9050), .B2(keyinput34), .C1(n10363), .C2(keyinput61), 
        .A(n10362), .ZN(n10371) );
  AOI22_X1 U11417 ( .A1(n10366), .A2(keyinput11), .B1(n10365), .B2(keyinput107), .ZN(n10364) );
  OAI221_X1 U11418 ( .B1(n10366), .B2(keyinput11), .C1(n10365), .C2(
        keyinput107), .A(n10364), .ZN(n10370) );
  XNOR2_X1 U11419 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput119), .ZN(n10368) );
  XNOR2_X1 U11420 ( .A(SI_12_), .B(keyinput100), .ZN(n10367) );
  NAND2_X1 U11421 ( .A1(n10368), .A2(n10367), .ZN(n10369) );
  NOR4_X1 U11422 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10401) );
  AOI22_X1 U11423 ( .A1(n10375), .A2(keyinput90), .B1(n10374), .B2(keyinput51), 
        .ZN(n10373) );
  OAI221_X1 U11424 ( .B1(n10375), .B2(keyinput90), .C1(n10374), .C2(keyinput51), .A(n10373), .ZN(n10385) );
  AOI22_X1 U11425 ( .A1(n5628), .A2(keyinput39), .B1(n10377), .B2(keyinput122), 
        .ZN(n10376) );
  OAI221_X1 U11426 ( .B1(n5628), .B2(keyinput39), .C1(n10377), .C2(keyinput122), .A(n10376), .ZN(n10384) );
  INV_X1 U11427 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U11428 ( .A1(n10380), .A2(keyinput15), .B1(keyinput124), .B2(n10379), .ZN(n10378) );
  OAI221_X1 U11429 ( .B1(n10380), .B2(keyinput15), .C1(n10379), .C2(
        keyinput124), .A(n10378), .ZN(n10383) );
  AOI22_X1 U11430 ( .A1(n6676), .A2(keyinput58), .B1(keyinput36), .B2(n9455), 
        .ZN(n10381) );
  OAI221_X1 U11431 ( .B1(n6676), .B2(keyinput58), .C1(n9455), .C2(keyinput36), 
        .A(n10381), .ZN(n10382) );
  NOR4_X1 U11432 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10400) );
  AOI22_X1 U11433 ( .A1(n10387), .A2(keyinput42), .B1(keyinput49), .B2(n6697), 
        .ZN(n10386) );
  OAI221_X1 U11434 ( .B1(n10387), .B2(keyinput42), .C1(n6697), .C2(keyinput49), 
        .A(n10386), .ZN(n10398) );
  AOI22_X1 U11435 ( .A1(n6079), .A2(keyinput77), .B1(keyinput113), .B2(n10389), 
        .ZN(n10388) );
  OAI221_X1 U11436 ( .B1(n6079), .B2(keyinput77), .C1(n10389), .C2(keyinput113), .A(n10388), .ZN(n10397) );
  INV_X1 U11437 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U11438 ( .A1(n10392), .A2(keyinput57), .B1(n10391), .B2(keyinput68), 
        .ZN(n10390) );
  OAI221_X1 U11439 ( .B1(n10392), .B2(keyinput57), .C1(n10391), .C2(keyinput68), .A(n10390), .ZN(n10396) );
  XNOR2_X1 U11440 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(keyinput60), .ZN(n10394)
         );
  XNOR2_X1 U11441 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput82), .ZN(n10393) );
  NAND2_X1 U11442 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  NOR4_X1 U11443 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10399) );
  NAND4_X1 U11444 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10458) );
  AOI22_X1 U11445 ( .A1(n10473), .A2(keyinput4), .B1(n10404), .B2(keyinput108), 
        .ZN(n10403) );
  OAI221_X1 U11446 ( .B1(n10473), .B2(keyinput4), .C1(n10404), .C2(keyinput108), .A(n10403), .ZN(n10415) );
  AOI22_X1 U11447 ( .A1(n10407), .A2(keyinput118), .B1(n10406), .B2(keyinput78), .ZN(n10405) );
  OAI221_X1 U11448 ( .B1(n10407), .B2(keyinput118), .C1(n10406), .C2(
        keyinput78), .A(n10405), .ZN(n10414) );
  INV_X1 U11449 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U11450 ( .A1(n10409), .A2(keyinput62), .B1(n5543), .B2(keyinput125), 
        .ZN(n10408) );
  OAI221_X1 U11451 ( .B1(n10409), .B2(keyinput62), .C1(n5543), .C2(keyinput125), .A(n10408), .ZN(n10413) );
  XNOR2_X1 U11452 ( .A(P1_REG1_REG_13__SCAN_IN), .B(keyinput38), .ZN(n10411)
         );
  XNOR2_X1 U11453 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput64), .ZN(n10410)
         );
  NAND2_X1 U11454 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  NOR4_X1 U11455 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10456) );
  XNOR2_X1 U11456 ( .A(n10416), .B(keyinput52), .ZN(n10417) );
  AOI21_X1 U11457 ( .B1(keyinput8), .B2(n5660), .A(n10417), .ZN(n10420) );
  XNOR2_X1 U11458 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput47), .ZN(n10419) );
  XNOR2_X1 U11459 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput24), .ZN(n10418) );
  NAND3_X1 U11460 ( .A1(n10420), .A2(n10419), .A3(n10418), .ZN(n10427) );
  AOI22_X1 U11461 ( .A1(n10423), .A2(keyinput50), .B1(keyinput17), .B2(n10422), 
        .ZN(n10421) );
  OAI221_X1 U11462 ( .B1(n10423), .B2(keyinput50), .C1(n10422), .C2(keyinput17), .A(n10421), .ZN(n10426) );
  XOR2_X1 U11463 ( .A(SI_6_), .B(keyinput94), .Z(n10425) );
  XNOR2_X1 U11464 ( .A(keyinput66), .B(n7116), .ZN(n10424) );
  NOR4_X1 U11465 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10455) );
  AOI22_X1 U11466 ( .A1(n10430), .A2(keyinput18), .B1(keyinput43), .B2(n10429), 
        .ZN(n10428) );
  OAI221_X1 U11467 ( .B1(n10430), .B2(keyinput18), .C1(n10429), .C2(keyinput43), .A(n10428), .ZN(n10440) );
  AOI22_X1 U11468 ( .A1(n10432), .A2(keyinput106), .B1(n5423), .B2(keyinput44), 
        .ZN(n10431) );
  OAI221_X1 U11469 ( .B1(n10432), .B2(keyinput106), .C1(n5423), .C2(keyinput44), .A(n10431), .ZN(n10439) );
  AOI22_X1 U11470 ( .A1(n10434), .A2(keyinput30), .B1(n7564), .B2(keyinput45), 
        .ZN(n10433) );
  OAI221_X1 U11471 ( .B1(n10434), .B2(keyinput30), .C1(n7564), .C2(keyinput45), 
        .A(n10433), .ZN(n10438) );
  XNOR2_X1 U11472 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput86), .ZN(n10436)
         );
  XNOR2_X1 U11473 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput92), .ZN(n10435) );
  NAND2_X1 U11474 ( .A1(n10436), .A2(n10435), .ZN(n10437) );
  NOR4_X1 U11475 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10454) );
  XOR2_X1 U11476 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput40), .Z(n10445) );
  XOR2_X1 U11477 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput19), .Z(n10444) );
  XNOR2_X1 U11478 ( .A(n10441), .B(keyinput117), .ZN(n10443) );
  XNOR2_X1 U11479 ( .A(keyinput96), .B(n6014), .ZN(n10442) );
  NOR4_X1 U11480 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10449) );
  XOR2_X1 U11481 ( .A(n10205), .B(keyinput3), .Z(n10448) );
  XNOR2_X1 U11482 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput120), .ZN(n10447)
         );
  XNOR2_X1 U11483 ( .A(SI_7_), .B(keyinput22), .ZN(n10446) );
  NAND4_X1 U11484 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10452) );
  XNOR2_X1 U11485 ( .A(n10450), .B(keyinput7), .ZN(n10451) );
  NOR2_X1 U11486 ( .A1(n10452), .A2(n10451), .ZN(n10453) );
  NAND4_X1 U11487 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10457) );
  NOR4_X1 U11488 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10461) );
  OAI21_X1 U11489 ( .B1(keyinput8), .B2(n10462), .A(n10461), .ZN(n10463) );
  XOR2_X1 U11490 ( .A(n10464), .B(n10463), .Z(P1_U3469) );
  XNOR2_X1 U11491 ( .A(n10466), .B(n10465), .ZN(ADD_1071_U50) );
  NOR2_X1 U11492 ( .A1(n10468), .A2(n10467), .ZN(n10470) );
  XNOR2_X1 U11493 ( .A(n10470), .B(n10469), .ZN(ADD_1071_U51) );
  OAI21_X1 U11494 ( .B1(n10473), .B2(n10472), .A(n10471), .ZN(n10474) );
  XNOR2_X1 U11495 ( .A(n10474), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11496 ( .B1(n6909), .B2(n10476), .A(n10475), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11497 ( .A(n10478), .B(n10477), .ZN(ADD_1071_U48) );
  XNOR2_X1 U11498 ( .A(n10480), .B(n10479), .ZN(ADD_1071_U49) );
  XOR2_X1 U11499 ( .A(n10482), .B(n10481), .Z(ADD_1071_U54) );
  XOR2_X1 U11500 ( .A(n10483), .B(n10484), .Z(ADD_1071_U53) );
  XNOR2_X1 U11501 ( .A(n10486), .B(n10485), .ZN(ADD_1071_U52) );
  INV_X1 U6862 ( .A(n7210), .ZN(n8447) );
  CLKBUF_X1 U4887 ( .A(n5677), .Z(n5845) );
  CLKBUF_X3 U4899 ( .A(n5193), .Z(n5791) );
  CLKBUF_X2 U4900 ( .A(n5114), .Z(n6691) );
  CLKBUF_X1 U4912 ( .A(n6393), .Z(n4383) );
  CLKBUF_X1 U4914 ( .A(n7649), .Z(n4376) );
  CLKBUF_X2 U4927 ( .A(n9332), .Z(n4378) );
endmodule

