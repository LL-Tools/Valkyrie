

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244;

  NAND2_X1 U4739 ( .A1(n5090), .A2(n5089), .ZN(n8732) );
  OR2_X1 U4740 ( .A1(n8820), .A2(n4646), .ZN(n4642) );
  NAND2_X1 U4741 ( .A1(n8813), .A2(n4838), .ZN(n8770) );
  AOI21_X1 U4742 ( .B1(n9361), .B2(n5917), .A(n5869), .ZN(n9376) );
  AND2_X1 U4743 ( .A1(n5854), .A2(n5853), .ZN(n9294) );
  NAND2_X2 U4744 ( .A1(n6322), .A2(n6321), .ZN(n9019) );
  XNOR2_X1 U4745 ( .A(n5584), .B(n5124), .ZN(n7193) );
  NAND2_X2 U4746 ( .A1(n6191), .A2(n6190), .ZN(n9066) );
  NAND2_X1 U4747 ( .A1(n8292), .A2(n8194), .ZN(n7477) );
  CLKBUF_X2 U4748 ( .A(n5207), .Z(n5746) );
  NAND2_X1 U4749 ( .A1(n4335), .A2(n4929), .ZN(n4928) );
  INV_X1 U4750 ( .A(n7522), .ZN(n7175) );
  INV_X1 U4751 ( .A(n5285), .ZN(n5640) );
  BUF_X2 U4753 ( .A(n6040), .Z(n4237) );
  INV_X1 U4754 ( .A(n6532), .ZN(n4769) );
  BUF_X2 U4755 ( .A(n5270), .Z(n4612) );
  INV_X1 U4756 ( .A(n6688), .ZN(n4236) );
  INV_X2 U4758 ( .A(n5478), .ZN(n5874) );
  INV_X1 U4759 ( .A(n6077), .ZN(n6406) );
  NAND2_X1 U4760 ( .A1(n6550), .A2(n6551), .ZN(n6688) );
  NAND2_X1 U4761 ( .A1(n7607), .A2(n7495), .ZN(n8083) );
  NAND2_X1 U4762 ( .A1(n9307), .A2(n9909), .ZN(n9918) );
  INV_X1 U4763 ( .A(n8407), .ZN(n5976) );
  NAND2_X1 U4764 ( .A1(n8463), .A2(n8219), .ZN(n9371) );
  NAND2_X1 U4765 ( .A1(n4907), .A2(n5862), .ZN(n9628) );
  INV_X1 U4766 ( .A(n9305), .ZN(n8066) );
  INV_X1 U4767 ( .A(n9307), .ZN(n9924) );
  NAND2_X1 U4768 ( .A1(n4908), .A2(n4912), .ZN(n5584) );
  AOI21_X1 U4769 ( .B1(n8732), .B2(n8352), .A(n5119), .ZN(n8715) );
  XNOR2_X1 U4770 ( .A(n4659), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U4771 ( .A1(n5692), .A2(n5691), .ZN(n9667) );
  NAND2_X1 U4772 ( .A1(n8413), .A2(n8412), .ZN(n9576) );
  XNOR2_X1 U4773 ( .A(n5354), .B(n5352), .ZN(n6723) );
  OR2_X1 U4774 ( .A1(n8986), .A2(n4454), .ZN(n4453) );
  CLKBUF_X3 U4775 ( .A(n5978), .Z(n4235) );
  NOR3_X2 U4776 ( .A1(n8145), .A2(n8167), .A3(n8433), .ZN(n8174) );
  BUF_X4 U4777 ( .A(n6010), .Z(n4234) );
  NAND2_X1 U4778 ( .A1(n5976), .A2(n5977), .ZN(n6010) );
  NAND2_X2 U4779 ( .A1(n4556), .A2(n5311), .ZN(n5354) );
  AOI21_X2 U4780 ( .B1(n4675), .B2(n4677), .A(n4674), .ZN(n4673) );
  INV_X1 U4781 ( .A(n8067), .ZN(n10209) );
  NAND2_X2 U4783 ( .A1(n5331), .A2(n5330), .ZN(n7429) );
  OR2_X2 U4784 ( .A1(n5902), .A2(n7181), .ZN(n7313) );
  NAND2_X1 U4785 ( .A1(n8141), .A2(n4282), .ZN(n4825) );
  NAND2_X1 U4786 ( .A1(n5816), .A2(n5815), .ZN(n9642) );
  NAND2_X1 U4787 ( .A1(n5844), .A2(n5843), .ZN(n9634) );
  INV_X2 U4788 ( .A(n8939), .ZN(n4777) );
  NAND2_X1 U4789 ( .A1(n5521), .A2(n5520), .ZN(n9705) );
  AND3_X1 U4790 ( .A1(n7641), .A2(n4856), .A3(n7994), .ZN(n7875) );
  NAND2_X2 U4791 ( .A1(n8275), .A2(n8083), .ZN(n7446) );
  NAND2_X1 U4792 ( .A1(n8068), .A2(n9918), .ZN(n8195) );
  NAND2_X1 U4793 ( .A1(n9305), .A2(n10209), .ZN(n8291) );
  NAND2_X1 U4794 ( .A1(n9924), .A2(n7414), .ZN(n8068) );
  XNOR2_X1 U4795 ( .A(n9892), .B(n9309), .ZN(n8192) );
  AND4_X1 U4796 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n7374)
         );
  NAND2_X1 U4797 ( .A1(n7182), .A2(n8176), .ZN(n9603) );
  CLKBUF_X1 U4798 ( .A(n8155), .Z(n4615) );
  AND2_X1 U4800 ( .A1(n5145), .A2(n5146), .ZN(n5337) );
  BUF_X2 U4801 ( .A(n6040), .Z(n4238) );
  BUF_X1 U4802 ( .A(n5285), .Z(n6779) );
  CLKBUF_X1 U4803 ( .A(n6775), .Z(n4239) );
  INV_X2 U4804 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OR2_X1 U4805 ( .A1(n6699), .A2(n4749), .ZN(n4748) );
  NOR2_X1 U4806 ( .A1(n4692), .A2(n4581), .ZN(n4635) );
  AOI21_X1 U4807 ( .B1(n4789), .B2(n4788), .A(n4786), .ZN(n8995) );
  AND2_X1 U4808 ( .A1(n4583), .A2(n4588), .ZN(n9132) );
  AOI21_X1 U4809 ( .B1(n9369), .B2(n9603), .A(n9368), .ZN(n9631) );
  NAND2_X1 U4810 ( .A1(n9407), .A2(n9414), .ZN(n9406) );
  AOI21_X1 U4811 ( .B1(n5053), .B2(n8917), .A(n4328), .ZN(n8985) );
  AOI21_X1 U4812 ( .B1(n4825), .B2(n4824), .A(n8170), .ZN(n4823) );
  AOI21_X1 U4813 ( .B1(n9402), .B2(n9603), .A(n9401), .ZN(n9644) );
  NAND2_X1 U4814 ( .A1(n8424), .A2(n8423), .ZN(n9420) );
  OAI21_X1 U4815 ( .B1(n9413), .B2(n8460), .A(n8461), .ZN(n9396) );
  XNOR2_X1 U4816 ( .A(n6346), .B(n4502), .ZN(n8496) );
  NAND2_X1 U4817 ( .A1(n4367), .A2(n4881), .ZN(n6346) );
  NAND2_X1 U4818 ( .A1(n4707), .A2(n4882), .ZN(n4367) );
  NAND2_X1 U4819 ( .A1(n4507), .A2(n5021), .ZN(n9462) );
  NAND2_X1 U4820 ( .A1(n6280), .A2(n8606), .ZN(n4707) );
  OAI21_X1 U4821 ( .B1(n8911), .B2(n5055), .A(n5054), .ZN(n8845) );
  AOI21_X1 U4822 ( .B1(n4882), .B2(n4885), .A(n4292), .ZN(n4881) );
  NAND2_X1 U4823 ( .A1(n4497), .A2(n4495), .ZN(n6280) );
  NAND2_X1 U4824 ( .A1(n9142), .A2(n4582), .ZN(n5556) );
  INV_X1 U4825 ( .A(n4380), .ZN(n4379) );
  NAND2_X1 U4826 ( .A1(n9563), .A2(n4514), .ZN(n4509) );
  XNOR2_X1 U4827 ( .A(n4832), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9344) );
  OR2_X1 U4828 ( .A1(n5058), .A2(n6633), .ZN(n5054) );
  NOR2_X1 U4829 ( .A1(n5060), .A2(n5059), .ZN(n5058) );
  AND2_X1 U4830 ( .A1(n9397), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U4831 ( .A1(n8144), .A2(n8143), .ZN(n9625) );
  NAND2_X1 U4832 ( .A1(n5532), .A2(n5531), .ZN(n9142) );
  OAI21_X1 U4833 ( .B1(n4681), .B2(n4381), .A(n8453), .ZN(n4380) );
  NAND2_X1 U4834 ( .A1(n5010), .A2(n5009), .ZN(n9421) );
  NAND2_X1 U4835 ( .A1(n6494), .A2(n6493), .ZN(n8982) );
  NAND2_X1 U4836 ( .A1(n5086), .A2(n4283), .ZN(n8903) );
  INV_X1 U4837 ( .A(n9475), .ZN(n5010) );
  AOI21_X1 U4838 ( .B1(n9517), .B2(n5026), .A(n4253), .ZN(n5025) );
  INV_X1 U4839 ( .A(n6347), .ZN(n4502) );
  OR2_X1 U4840 ( .A1(n9634), .A2(n9294), .ZN(n8463) );
  AND2_X1 U4841 ( .A1(n8942), .A2(n4843), .ZN(n8854) );
  NAND2_X1 U4842 ( .A1(n4349), .A2(n6337), .ZN(n9012) );
  INV_X1 U4843 ( .A(n9454), .ZN(n9661) );
  NAND2_X1 U4844 ( .A1(n4376), .A2(n4966), .ZN(n9578) );
  XNOR2_X1 U4845 ( .A(n6487), .B(n6486), .ZN(n8335) );
  NAND2_X1 U4846 ( .A1(n5734), .A2(n5733), .ZN(n9656) );
  NOR2_X1 U4847 ( .A1(n9034), .A2(n4845), .ZN(n4843) );
  NAND2_X1 U4848 ( .A1(n5860), .A2(n5859), .ZN(n6487) );
  NAND2_X1 U4849 ( .A1(n6353), .A2(n6352), .ZN(n9003) );
  AND2_X1 U4850 ( .A1(n5714), .A2(n5713), .ZN(n9454) );
  OR2_X1 U4851 ( .A1(n8442), .A2(n8263), .ZN(n9562) );
  XNOR2_X1 U4852 ( .A(n5858), .B(n5857), .ZN(n8054) );
  XNOR2_X1 U4853 ( .A(n5732), .B(n5759), .ZN(n7938) );
  NAND2_X1 U4854 ( .A1(n6307), .A2(n6306), .ZN(n9024) );
  OAI21_X1 U4855 ( .B1(n5727), .B2(n5726), .A(n5755), .ZN(n5732) );
  AND2_X1 U4856 ( .A1(n8430), .A2(n9610), .ZN(n9605) );
  NAND2_X1 U4857 ( .A1(n4920), .A2(n4918), .ZN(n5858) );
  NAND2_X1 U4858 ( .A1(n4360), .A2(n4280), .ZN(n7820) );
  XNOR2_X1 U4859 ( .A(n5809), .B(n5808), .ZN(n8036) );
  NOR2_X1 U4860 ( .A1(n5070), .A2(n7945), .ZN(n5069) );
  NAND2_X1 U4861 ( .A1(n5035), .A2(n5034), .ZN(n7779) );
  NAND2_X1 U4862 ( .A1(n5618), .A2(n5617), .ZN(n9681) );
  NAND2_X2 U4863 ( .A1(n6621), .A2(n6620), .ZN(n8340) );
  NAND2_X1 U4864 ( .A1(n5670), .A2(n5669), .ZN(n9672) );
  NAND2_X1 U4865 ( .A1(n7633), .A2(n7632), .ZN(n7678) );
  INV_X1 U4866 ( .A(n4245), .ZN(n5071) );
  NAND2_X1 U4867 ( .A1(n5642), .A2(n5641), .ZN(n9676) );
  NAND2_X1 U4868 ( .A1(n7638), .A2(n6595), .ZN(n7655) );
  XNOR2_X1 U4869 ( .A(n5634), .B(n5632), .ZN(n7408) );
  OAI21_X1 U4870 ( .B1(n4932), .B2(n4572), .A(n4570), .ZN(n5786) );
  NAND2_X1 U4871 ( .A1(n5568), .A2(n5567), .ZN(n9693) );
  NAND2_X1 U4872 ( .A1(n5546), .A2(n5545), .ZN(n9569) );
  NAND2_X1 U4873 ( .A1(n6242), .A2(n6241), .ZN(n9056) );
  NAND2_X1 U4874 ( .A1(n6209), .A2(n6208), .ZN(n9061) );
  NAND2_X1 U4875 ( .A1(n5499), .A2(n5498), .ZN(n9709) );
  NOR2_X1 U4876 ( .A1(n5349), .A2(n5117), .ZN(n5350) );
  OAI21_X1 U4877 ( .B1(n4878), .B2(n4874), .A(n4872), .ZN(n4501) );
  AOI21_X1 U4878 ( .B1(n7165), .B2(n7164), .A(n5256), .ZN(n7198) );
  NAND2_X1 U4879 ( .A1(n5469), .A2(n5468), .ZN(n8409) );
  NAND2_X1 U4880 ( .A1(n5438), .A2(n5437), .ZN(n7893) );
  AOI21_X1 U4881 ( .B1(n4875), .B2(n4873), .A(n4293), .ZN(n4872) );
  OR2_X1 U4882 ( .A1(n5510), .A2(n4914), .ZN(n4908) );
  NOR2_X1 U4883 ( .A1(n9089), .A2(n9083), .ZN(n4858) );
  OAI21_X1 U4884 ( .B1(n8370), .B2(n8368), .A(n8371), .ZN(n7588) );
  NAND2_X1 U4885 ( .A1(n6141), .A2(n4493), .ZN(n9077) );
  XNOR2_X1 U4886 ( .A(n4622), .B(n5411), .ZN(n6740) );
  NAND2_X2 U4887 ( .A1(n5314), .A2(n5313), .ZN(n7607) );
  NAND2_X1 U4888 ( .A1(n4905), .A2(n5412), .ZN(n4557) );
  OAI21_X1 U4889 ( .B1(n5380), .B2(n5379), .A(n5407), .ZN(n4622) );
  OR2_X2 U4890 ( .A1(n7339), .A2(n7711), .ZN(n7707) );
  NAND2_X1 U4891 ( .A1(n6792), .A2(n6793), .ZN(n6800) );
  OR2_X1 U4892 ( .A1(n7743), .A2(n9986), .ZN(n7339) );
  OR2_X1 U4893 ( .A1(n9928), .A2(n7429), .ZN(n7480) );
  INV_X1 U4894 ( .A(n7360), .ZN(n8190) );
  OR2_X1 U4895 ( .A1(n7067), .A2(n7068), .ZN(n4392) );
  NAND2_X1 U4896 ( .A1(n5289), .A2(n5288), .ZN(n8067) );
  AND2_X1 U4897 ( .A1(n4912), .A2(n4565), .ZN(n4564) );
  AND2_X1 U4898 ( .A1(n4303), .A2(n4403), .ZN(n5207) );
  NAND4_X2 U4899 ( .A1(n5280), .A2(n5279), .A3(n5278), .A4(n5277), .ZN(n9305)
         );
  AND2_X2 U4900 ( .A1(n6023), .A2(n6022), .ZN(n8391) );
  INV_X1 U4901 ( .A(n7397), .ZN(n7362) );
  INV_X1 U4902 ( .A(n7405), .ZN(n4989) );
  AND2_X1 U4903 ( .A1(n10010), .A2(n7509), .ZN(n7286) );
  NOR2_X1 U4904 ( .A1(n6907), .A2(n10000), .ZN(P2_U3966) );
  NAND4_X2 U4905 ( .A1(n5210), .A2(n5211), .A3(n5213), .A4(n5212), .ZN(n9309)
         );
  AND4_X1 U4906 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n7397)
         );
  CLKBUF_X3 U4907 ( .A(n5337), .Z(n5917) );
  OAI211_X1 U4908 ( .C1(n6779), .C2(n6836), .A(n5250), .B(n5249), .ZN(n7405)
         );
  NAND2_X1 U4909 ( .A1(n4655), .A2(n4653), .ZN(n8660) );
  NAND2_X1 U4910 ( .A1(n4337), .A2(n5283), .ZN(n5304) );
  INV_X1 U4911 ( .A(n7736), .ZN(n10010) );
  XNOR2_X1 U4912 ( .A(n5168), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U4914 ( .B1(n5309), .B2(n4906), .A(n5353), .ZN(n4343) );
  NAND2_X2 U4915 ( .A1(n5964), .A2(n4362), .ZN(n6532) );
  NAND2_X1 U4916 ( .A1(n5167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U4917 ( .A1(n5144), .A2(n9746), .ZN(n9753) );
  NAND2_X2 U4918 ( .A1(n8407), .A2(n5977), .ZN(n6025) );
  AND2_X4 U4919 ( .A1(n8407), .A2(n4235), .ZN(n6024) );
  XNOR2_X1 U4920 ( .A(n5156), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7181) );
  OR2_X1 U4921 ( .A1(n5960), .A2(n4363), .ZN(n4362) );
  OR2_X1 U4922 ( .A1(n5959), .A2(n9120), .ZN(n5960) );
  XNOR2_X1 U4923 ( .A(n4693), .B(n5171), .ZN(n6775) );
  XNOR2_X1 U4924 ( .A(n5355), .B(n4344), .ZN(n5353) );
  XNOR2_X1 U4925 ( .A(n6412), .B(n6411), .ZN(n6550) );
  OAI21_X1 U4926 ( .B1(n5961), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U4927 ( .A1(n4369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4693) );
  XNOR2_X1 U4928 ( .A(n5266), .B(SI_3_), .ZN(n5264) );
  INV_X2 U4929 ( .A(n5270), .ZN(n5180) );
  AND3_X1 U4930 ( .A1(n4494), .A2(n5956), .A3(n5955), .ZN(n4792) );
  CLKBUF_X1 U4931 ( .A(n5188), .Z(n5189) );
  NOR2_X1 U4932 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  AND4_X1 U4933 ( .A1(n5958), .A2(n4903), .A3(n6411), .A4(n5963), .ZN(n5940)
         );
  NAND3_X1 U4934 ( .A1(n9347), .A2(n4334), .A3(n4460), .ZN(n4463) );
  AND3_X1 U4935 ( .A1(n5019), .A2(n5018), .A3(n5017), .ZN(n5130) );
  AND3_X1 U4936 ( .A1(n4837), .A2(n5939), .A3(n5938), .ZN(n5941) );
  AND2_X1 U4937 ( .A1(n6018), .A2(n5945), .ZN(n5956) );
  AND4_X1 U4938 ( .A1(n5944), .A2(n6017), .A3(n5942), .A4(n5943), .ZN(n4494)
         );
  INV_X1 U4939 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6017) );
  NOR2_X2 U4940 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6018) );
  NOR2_X1 U4941 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4837) );
  NOR2_X1 U4942 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5019) );
  NOR2_X1 U4943 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5152) );
  NOR2_X1 U4944 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5018) );
  NOR2_X1 U4945 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5017) );
  NOR2_X1 U4946 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5974) );
  NOR2_X2 U4947 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4555) );
  NOR2_X1 U4948 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5939) );
  NOR2_X1 U4949 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5942) );
  INV_X1 U4950 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5171) );
  NOR2_X1 U4951 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5943) );
  NOR2_X1 U4952 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5136) );
  INV_X1 U4953 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5963) );
  NAND2_X4 U4954 ( .A1(n7626), .A2(n4368), .ZN(n6077) );
  OAI21_X1 U4955 ( .B1(n5664), .B2(n5663), .A(n5662), .ZN(n5689) );
  NAND2_X4 U4956 ( .A1(n4463), .A2(n4461), .ZN(n5270) );
  INV_X2 U4957 ( .A(n5180), .ZN(n6522) );
  INV_X1 U4958 ( .A(n5263), .ZN(n4240) );
  NAND2_X4 U4959 ( .A1(n4235), .A2(n5976), .ZN(n6009) );
  AOI21_X1 U4960 ( .B1(n5092), .B2(n5095), .A(n4290), .ZN(n5089) );
  INV_X1 U4961 ( .A(n4568), .ZN(n4567) );
  OAI21_X1 U4962 ( .B1(n4927), .B2(n4569), .A(n5116), .ZN(n4568) );
  INV_X1 U4963 ( .A(n6220), .ZN(n4892) );
  OR2_X1 U4964 ( .A1(n8729), .A2(n8740), .ZN(n6677) );
  OR2_X1 U4965 ( .A1(n5819), .A2(n5818), .ZN(n5846) );
  NAND2_X1 U4966 ( .A1(n7538), .A2(n7537), .ZN(n7723) );
  INV_X1 U4967 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U4968 ( .B1(n4347), .B2(n4345), .A(n4709), .ZN(n5664) );
  AOI21_X1 U4969 ( .B1(n5633), .B2(n4710), .A(n4291), .ZN(n4709) );
  OAI21_X1 U4970 ( .B1(n4564), .B2(n4348), .A(n4708), .ZN(n4347) );
  NOR2_X1 U4971 ( .A1(n4563), .A2(n4348), .ZN(n4345) );
  NAND2_X1 U4972 ( .A1(n6369), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6397) );
  AOI21_X1 U4973 ( .B1(n4647), .B2(n4645), .A(n4297), .ZN(n4644) );
  INV_X1 U4974 ( .A(n8819), .ZN(n4645) );
  INV_X1 U4975 ( .A(n4647), .ZN(n4646) );
  NOR2_X1 U4976 ( .A1(n8778), .A2(n4450), .ZN(n4449) );
  INV_X1 U4977 ( .A(n6651), .ZN(n4450) );
  AND2_X1 U4978 ( .A1(n6910), .A2(n5180), .ZN(n6037) );
  NAND2_X1 U4979 ( .A1(n6436), .A2(n6435), .ZN(n6534) );
  NAND2_X1 U4980 ( .A1(n9246), .A2(n9248), .ZN(n5725) );
  NAND2_X1 U4981 ( .A1(n4694), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U4982 ( .A1(n7458), .A2(n4939), .ZN(n4941) );
  AND2_X1 U4983 ( .A1(n4274), .A2(n5350), .ZN(n4939) );
  NAND2_X1 U4984 ( .A1(n4802), .A2(n4801), .ZN(n8100) );
  NOR2_X1 U4985 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  INV_X1 U4986 ( .A(n8452), .ZN(n4799) );
  NAND2_X1 U4987 ( .A1(n8112), .A2(n8113), .ZN(n8114) );
  OR2_X1 U4988 ( .A1(n8130), .A2(n8167), .ZN(n4811) );
  NAND2_X1 U4989 ( .A1(n4484), .A2(n4480), .ZN(n4479) );
  AND2_X1 U4990 ( .A1(n8796), .A2(n4268), .ZN(n4480) );
  NOR2_X1 U4991 ( .A1(n4735), .A2(n4734), .ZN(n4741) );
  NAND2_X1 U4992 ( .A1(n6674), .A2(n6673), .ZN(n4734) );
  NOR2_X1 U4993 ( .A1(n4736), .A2(n6675), .ZN(n4735) );
  NAND2_X1 U4994 ( .A1(n4825), .A2(n8142), .ZN(n8145) );
  AND2_X1 U4995 ( .A1(n4879), .A2(n4876), .ZN(n4875) );
  INV_X1 U4996 ( .A(n7525), .ZN(n4876) );
  NAND2_X1 U4997 ( .A1(n4504), .A2(n4503), .ZN(n6088) );
  INV_X1 U4998 ( .A(n6085), .ZN(n4503) );
  INV_X1 U4999 ( .A(n6086), .ZN(n4504) );
  OR2_X1 U5000 ( .A1(n8982), .A2(n4855), .ZN(n4854) );
  OR2_X1 U5001 ( .A1(n9003), .A2(n8644), .ZN(n5097) );
  INV_X1 U5002 ( .A(n5098), .ZN(n5096) );
  OR2_X1 U5003 ( .A1(n8998), .A2(n8476), .ZN(n6664) );
  NOR2_X1 U5004 ( .A1(n9019), .A2(n9012), .ZN(n4842) );
  OR2_X1 U5005 ( .A1(n9029), .A2(n8513), .ZN(n6641) );
  NOR2_X1 U5006 ( .A1(n5071), .A2(n6607), .ZN(n5070) );
  INV_X1 U5007 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5947) );
  INV_X1 U5008 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5946) );
  INV_X1 U5009 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5957) );
  OR2_X1 U5010 ( .A1(n5507), .A2(n9236), .ZN(n4960) );
  INV_X1 U5011 ( .A(n8464), .ZN(n4674) );
  OAI21_X1 U5012 ( .B1(n5038), .B2(n4680), .A(n4295), .ZN(n5037) );
  AND2_X1 U5013 ( .A1(n5027), .A2(n4247), .ZN(n5023) );
  NAND2_X1 U5014 ( .A1(n4513), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U5015 ( .A1(n5004), .A2(n9199), .ZN(n4512) );
  AND2_X1 U5016 ( .A1(n5045), .A2(n4273), .ZN(n4514) );
  OR2_X1 U5017 ( .A1(n9681), .A2(n8063), .ZN(n8187) );
  NOR2_X1 U5018 ( .A1(n7848), .A2(n8409), .ZN(n8430) );
  OR2_X1 U5019 ( .A1(n9715), .A2(n7777), .ZN(n8252) );
  NAND2_X1 U5020 ( .A1(n7429), .A2(n9926), .ZN(n8194) );
  OR2_X1 U5021 ( .A1(n6497), .A2(n6496), .ZN(n6516) );
  AOI21_X1 U5022 ( .B1(n4922), .B2(n4924), .A(n4919), .ZN(n4918) );
  NAND2_X1 U5023 ( .A1(n5786), .A2(n4922), .ZN(n4920) );
  INV_X1 U5024 ( .A(n5838), .ZN(n4919) );
  INV_X1 U5025 ( .A(n5899), .ZN(n5163) );
  INV_X1 U5026 ( .A(SI_20_), .ZN(n5665) );
  NOR2_X1 U5027 ( .A1(n5611), .A2(n4713), .ZN(n4712) );
  INV_X1 U5028 ( .A(n5585), .ZN(n4713) );
  NAND2_X1 U5029 ( .A1(n4563), .A2(n4564), .ZN(n4346) );
  INV_X1 U5030 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U5031 ( .B1(n4916), .B2(n4914), .A(n5557), .ZN(n4913) );
  AOI21_X1 U5032 ( .B1(n4889), .B2(n4892), .A(n4888), .ZN(n4887) );
  INV_X1 U5033 ( .A(n6248), .ZN(n4888) );
  OR2_X1 U5034 ( .A1(n4886), .A2(n4890), .ZN(n4500) );
  NOR2_X1 U5035 ( .A1(n7915), .A2(n7914), .ZN(n8666) );
  XNOR2_X1 U5036 ( .A(n4269), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n4415) );
  OR2_X1 U5037 ( .A1(n6397), .A2(n6396), .ZN(n6459) );
  NAND2_X1 U5038 ( .A1(n4352), .A2(n8717), .ZN(n8716) );
  OAI21_X1 U5039 ( .B1(n5074), .B2(n8776), .A(n5076), .ZN(n4353) );
  AOI21_X1 U5040 ( .B1(n8751), .B2(n8738), .A(n8737), .ZN(n4790) );
  NAND2_X1 U5041 ( .A1(n8740), .A2(n8914), .ZN(n4787) );
  OR2_X1 U5042 ( .A1(n9003), .A2(n8779), .ZN(n8750) );
  AND2_X1 U5043 ( .A1(n4644), .A2(n8778), .ZN(n4643) );
  NAND2_X1 U5044 ( .A1(n8820), .A2(n8819), .ZN(n4648) );
  AOI21_X1 U5045 ( .B1(n8845), .B2(n4782), .A(n4780), .ZN(n8797) );
  NOR2_X1 U5046 ( .A1(n5107), .A2(n4783), .ZN(n4782) );
  INV_X1 U5047 ( .A(n6645), .ZN(n4783) );
  NAND2_X1 U5048 ( .A1(n8797), .A2(n8796), .ZN(n8795) );
  AND2_X1 U5049 ( .A1(n5107), .A2(n5109), .ZN(n5106) );
  NOR2_X1 U5050 ( .A1(n4263), .A2(n5111), .ZN(n5110) );
  INV_X1 U5051 ( .A(n8347), .ZN(n5111) );
  INV_X1 U5052 ( .A(n8932), .ZN(n8912) );
  INV_X1 U5053 ( .A(n8917), .ZN(n8930) );
  AOI21_X1 U5054 ( .B1(n6455), .B2(n4278), .A(n4850), .ZN(n4849) );
  NAND2_X1 U5055 ( .A1(n6695), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5950) );
  NOR2_X1 U5056 ( .A1(n5974), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5057 ( .A1(n8716), .A2(n6673), .ZN(n8361) );
  NAND2_X1 U5058 ( .A1(n8740), .A2(n8912), .ZN(n8365) );
  OR2_X1 U5059 ( .A1(n10009), .A2(n6696), .ZN(n10020) );
  INV_X1 U5060 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5938) );
  INV_X1 U5061 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6413) );
  NOR2_X1 U5062 ( .A1(n5455), .A2(n4599), .ZN(n4598) );
  INV_X1 U5063 ( .A(n9444), .ZN(n9192) );
  NAND2_X1 U5064 ( .A1(n5556), .A2(n4955), .ZN(n4953) );
  OR2_X1 U5065 ( .A1(n5555), .A2(n9280), .ZN(n4955) );
  NAND2_X1 U5066 ( .A1(n5764), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U5067 ( .A1(n5400), .A2(n5399), .ZN(n4624) );
  AND2_X1 U5068 ( .A1(n5707), .A2(n5721), .ZN(n4961) );
  AOI21_X1 U5069 ( .B1(n4603), .B2(n5687), .A(n4602), .ZN(n4601) );
  INV_X1 U5070 ( .A(n5298), .ZN(n5299) );
  INV_X1 U5071 ( .A(n4615), .ZN(n5914) );
  INV_X1 U5072 ( .A(n5917), .ZN(n5848) );
  INV_X1 U5073 ( .A(n4626), .ZN(n8148) );
  NAND2_X1 U5074 ( .A1(n6834), .A2(n6835), .ZN(n6833) );
  NAND2_X1 U5075 ( .A1(n6768), .A2(n6767), .ZN(n6841) );
  OAI21_X1 U5076 ( .B1(n6836), .B2(P1_REG2_REG_3__SCAN_IN), .A(n4638), .ZN(
        n6767) );
  NAND2_X1 U5077 ( .A1(n6836), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4638) );
  OR2_X1 U5078 ( .A1(n9848), .A2(n4833), .ZN(n4832) );
  AND2_X1 U5079 ( .A1(n9854), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4833) );
  XNOR2_X1 U5080 ( .A(n4397), .B(n9341), .ZN(n9343) );
  NAND2_X1 U5081 ( .A1(n4399), .A2(n4398), .ZN(n4397) );
  NAND2_X1 U5082 ( .A1(n9340), .A2(n9339), .ZN(n4398) );
  OAI21_X1 U5083 ( .B1(n9420), .B2(n4519), .A(n4516), .ZN(n9360) );
  NAND2_X1 U5084 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  OR2_X1 U5085 ( .A1(n5037), .A2(n4265), .ZN(n4519) );
  INV_X1 U5086 ( .A(n5037), .ZN(n4517) );
  INV_X1 U5087 ( .A(n4515), .ZN(n9407) );
  NAND2_X1 U5088 ( .A1(n4378), .A2(n4377), .ZN(n8455) );
  AOI21_X1 U5089 ( .B1(n4379), .B2(n4381), .A(n9461), .ZN(n4377) );
  NAND2_X1 U5090 ( .A1(n4683), .A2(n4379), .ZN(n4378) );
  NAND2_X1 U5091 ( .A1(n7723), .A2(n7722), .ZN(n5035) );
  NAND2_X1 U5092 ( .A1(n7421), .A2(n7420), .ZN(n4613) );
  NAND2_X1 U5093 ( .A1(n8331), .A2(n9468), .ZN(n7176) );
  NAND2_X1 U5094 ( .A1(n5285), .A2(n4612), .ZN(n5263) );
  AND2_X1 U5095 ( .A1(n5920), .A2(n6874), .ZN(n9540) );
  OR2_X1 U5096 ( .A1(n8177), .A2(n6874), .ZN(n9927) );
  AND3_X1 U5097 ( .A1(n6895), .A2(n6894), .A3(n6893), .ZN(n7191) );
  CLKBUF_X1 U5098 ( .A(n5196), .Z(n5898) );
  XNOR2_X1 U5099 ( .A(n5900), .B(n5160), .ZN(n7934) );
  NAND2_X1 U5100 ( .A1(n7931), .A2(n6433), .ZN(n6907) );
  NAND2_X1 U5101 ( .A1(n4707), .A2(n6291), .ZN(n8505) );
  NAND2_X1 U5102 ( .A1(n4899), .A2(n4322), .ZN(n4898) );
  INV_X1 U5103 ( .A(n6447), .ZN(n4894) );
  AND2_X1 U5104 ( .A1(n9003), .A2(n8638), .ZN(n4365) );
  OAI21_X1 U5105 ( .B1(n8758), .B2(n4234), .A(n6377), .ZN(n8733) );
  NAND2_X1 U5106 ( .A1(n5910), .A2(n9566), .ZN(n9288) );
  INV_X1 U5107 ( .A(n8328), .ZN(n8325) );
  INV_X1 U5108 ( .A(n8063), .ZN(n9523) );
  NOR2_X1 U5109 ( .A1(n8069), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5110 ( .A1(n4746), .A2(n4745), .ZN(n6572) );
  OR2_X1 U5111 ( .A1(n6559), .A2(n4236), .ZN(n4745) );
  NAND2_X1 U5112 ( .A1(n6557), .A2(n4236), .ZN(n4746) );
  NAND2_X1 U5113 ( .A1(n8086), .A2(n8252), .ZN(n4805) );
  NAND2_X1 U5114 ( .A1(n8081), .A2(n8167), .ZN(n4801) );
  OAI21_X1 U5115 ( .B1(n4804), .B2(n4803), .A(n8163), .ZN(n4802) );
  NAND2_X1 U5116 ( .A1(n8435), .A2(n8088), .ZN(n4803) );
  AOI21_X1 U5117 ( .B1(n8080), .B2(n4806), .A(n4805), .ZN(n4804) );
  NOR2_X1 U5118 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U5119 ( .A1(n4492), .A2(n4489), .ZN(n6603) );
  NAND2_X1 U5120 ( .A1(n6556), .A2(n6688), .ZN(n4492) );
  AND2_X1 U5121 ( .A1(n6590), .A2(n4490), .ZN(n4489) );
  INV_X1 U5122 ( .A(n8268), .ZN(n4797) );
  AOI21_X1 U5123 ( .B1(n8268), .B2(n4249), .A(n8167), .ZN(n4796) );
  AOI21_X1 U5124 ( .B1(n4798), .B2(n4251), .A(n8163), .ZN(n4794) );
  AND2_X1 U5125 ( .A1(n6627), .A2(n8926), .ZN(n4474) );
  INV_X1 U5126 ( .A(n8136), .ZN(n4549) );
  NAND2_X1 U5127 ( .A1(n4810), .A2(n8167), .ZN(n4809) );
  NAND2_X1 U5128 ( .A1(n4486), .A2(n4485), .ZN(n4484) );
  NAND2_X1 U5129 ( .A1(n6646), .A2(n6688), .ZN(n4485) );
  NAND2_X1 U5130 ( .A1(n4487), .A2(n4236), .ZN(n4486) );
  INV_X1 U5131 ( .A(n6291), .ZN(n4884) );
  NOR2_X1 U5132 ( .A1(n4435), .A2(n5080), .ZN(n4434) );
  NOR2_X1 U5133 ( .A1(n7872), .A2(n7686), .ZN(n4436) );
  NOR2_X1 U5134 ( .A1(n6661), .A2(n6662), .ZN(n4733) );
  INV_X1 U5135 ( .A(n9363), .ZN(n8465) );
  NAND2_X1 U5136 ( .A1(n7362), .A2(n7175), .ZN(n8241) );
  INV_X1 U5137 ( .A(n5753), .ZN(n4572) );
  AND2_X1 U5138 ( .A1(n5708), .A2(n5690), .ZN(n4931) );
  AOI21_X1 U5139 ( .B1(n4912), .B2(n4914), .A(n4910), .ZN(n4909) );
  INV_X1 U5140 ( .A(n5124), .ZN(n4910) );
  INV_X1 U5141 ( .A(n5490), .ZN(n4569) );
  NAND2_X1 U5142 ( .A1(n4341), .A2(n4340), .ZN(n4339) );
  INV_X1 U5143 ( .A(n4343), .ZN(n4340) );
  OAI21_X1 U5144 ( .B1(n5180), .B2(P2_DATAO_REG_5__SCAN_IN), .A(n4336), .ZN(
        n5305) );
  NAND2_X1 U5145 ( .A1(n5180), .A2(n6718), .ZN(n4336) );
  INV_X1 U5146 ( .A(n6382), .ZN(n4721) );
  AND2_X1 U5147 ( .A1(n6331), .A2(n8660), .ZN(n6014) );
  INV_X1 U5148 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U5149 ( .A1(n5984), .A2(n6532), .ZN(n6440) );
  INV_X1 U5150 ( .A(n4235), .ZN(n5977) );
  NAND2_X1 U5151 ( .A1(n8736), .A2(n6656), .ZN(n5074) );
  NOR2_X1 U5152 ( .A1(n4841), .A2(n9007), .ZN(n4840) );
  INV_X1 U5153 ( .A(n4842), .ZN(n4841) );
  INV_X1 U5154 ( .A(n6641), .ZN(n4781) );
  NAND2_X1 U5155 ( .A1(n9050), .A2(n8647), .ZN(n5088) );
  NAND2_X1 U5156 ( .A1(n8926), .A2(n5088), .ZN(n5085) );
  NOR2_X1 U5157 ( .A1(n4778), .A2(n6588), .ZN(n4447) );
  NAND2_X1 U5158 ( .A1(n9061), .A2(n8933), .ZN(n6620) );
  NOR2_X1 U5159 ( .A1(n4857), .A2(n9077), .ZN(n4856) );
  INV_X1 U5160 ( .A(n4858), .ZN(n4857) );
  INV_X1 U5161 ( .A(n10009), .ZN(n6437) );
  AND2_X1 U5162 ( .A1(n5956), .A2(n5949), .ZN(n4729) );
  INV_X1 U5163 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6168) );
  INV_X1 U5164 ( .A(n6052), .ZN(n4427) );
  NAND2_X1 U5165 ( .A1(n5507), .A2(n9236), .ZN(n4959) );
  NOR2_X1 U5166 ( .A1(n5715), .A2(n10136), .ZN(n4694) );
  NAND2_X1 U5167 ( .A1(n8328), .A2(n5903), .ZN(n4403) );
  AOI21_X1 U5168 ( .B1(n5661), .B2(n4937), .A(n9224), .ZN(n4936) );
  INV_X1 U5169 ( .A(n5655), .ZN(n4937) );
  NAND2_X1 U5170 ( .A1(n9206), .A2(n4934), .ZN(n4933) );
  INV_X1 U5171 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U5172 ( .B1(n4936), .B2(n5687), .A(n9176), .ZN(n4604) );
  NAND2_X1 U5173 ( .A1(n4543), .A2(n4822), .ZN(n4697) );
  NOR2_X1 U5174 ( .A1(n8172), .A2(n8306), .ZN(n4822) );
  OAI21_X1 U5175 ( .B1(n8145), .B2(n4544), .A(n4823), .ZN(n4543) );
  INV_X1 U5176 ( .A(n8171), .ZN(n4544) );
  INV_X1 U5177 ( .A(n9753), .ZN(n5146) );
  OR2_X1 U5178 ( .A1(n5864), .A2(n5863), .ZN(n5911) );
  INV_X1 U5179 ( .A(n8462), .ZN(n4678) );
  INV_X1 U5180 ( .A(n8422), .ZN(n5032) );
  NAND2_X1 U5181 ( .A1(n9439), .A2(n5013), .ZN(n5012) );
  INV_X1 U5182 ( .A(n5014), .ZN(n5013) );
  NOR2_X1 U5183 ( .A1(n5643), .A2(n4704), .ZN(n4703) );
  NOR2_X1 U5184 ( .A1(n4511), .A2(n5024), .ZN(n4510) );
  NAND2_X1 U5185 ( .A1(n5025), .A2(n4247), .ZN(n5024) );
  INV_X1 U5186 ( .A(n8417), .ZN(n5028) );
  INV_X1 U5187 ( .A(n5620), .ZN(n5619) );
  NAND2_X1 U5188 ( .A1(n5008), .A2(n5007), .ZN(n5006) );
  NOR2_X1 U5189 ( .A1(n9705), .A2(n9569), .ZN(n5008) );
  AND2_X1 U5190 ( .A1(n9599), .A2(n4970), .ZN(n4969) );
  OR2_X1 U5191 ( .A1(n4972), .A2(n4971), .ZN(n4970) );
  INV_X1 U5192 ( .A(n8435), .ZN(n4971) );
  NAND2_X1 U5193 ( .A1(n4383), .A2(n4382), .ZN(n4385) );
  NAND2_X1 U5194 ( .A1(n4964), .A2(n4687), .ZN(n7436) );
  AND2_X1 U5195 ( .A1(n8247), .A2(n4965), .ZN(n4964) );
  NAND2_X1 U5196 ( .A1(n4815), .A2(n9918), .ZN(n4965) );
  AND2_X1 U5197 ( .A1(n9909), .A2(n7175), .ZN(n4987) );
  INV_X1 U5198 ( .A(SI_12_), .ZN(n10082) );
  NAND2_X1 U5199 ( .A1(n9308), .A2(n4989), .ZN(n8245) );
  NAND2_X1 U5200 ( .A1(n8241), .A2(n8240), .ZN(n7360) );
  NOR2_X1 U5201 ( .A1(n9625), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U5202 ( .A1(n4998), .A2(n9385), .ZN(n5000) );
  OR2_X1 U5203 ( .A1(n9488), .A2(n9672), .ZN(n9475) );
  AND2_X1 U5204 ( .A1(n5838), .A2(n5814), .ZN(n5836) );
  AND2_X1 U5205 ( .A1(n5690), .A2(n5668), .ZN(n5688) );
  INV_X1 U5206 ( .A(SI_16_), .ZN(n5560) );
  NAND2_X1 U5207 ( .A1(n4915), .A2(n5536), .ZN(n4914) );
  INV_X1 U5208 ( .A(n5558), .ZN(n4915) );
  NOR2_X1 U5209 ( .A1(n5537), .A2(n4917), .ZN(n4916) );
  INV_X1 U5210 ( .A(n5509), .ZN(n4917) );
  AND2_X1 U5211 ( .A1(n5489), .A2(n5459), .ZN(n4927) );
  INV_X1 U5212 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5466) );
  NOR2_X1 U5213 ( .A1(n5460), .A2(n4930), .ZN(n4929) );
  INV_X1 U5214 ( .A(n5434), .ZN(n4930) );
  NOR2_X1 U5215 ( .A1(n5435), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U5216 ( .A1(n4557), .A2(n5115), .ZN(n4335) );
  NOR2_X2 U5217 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5172) );
  INV_X1 U5218 ( .A(n7580), .ZN(n4873) );
  INV_X1 U5219 ( .A(n4875), .ZN(n4874) );
  INV_X1 U5220 ( .A(n8830), .ZN(n8513) );
  OR2_X1 U5221 ( .A1(n8555), .A2(n8559), .ZN(n4728) );
  INV_X1 U5222 ( .A(n8660), .ZN(n8599) );
  AND2_X1 U5223 ( .A1(n4887), .A2(n4499), .ZN(n4498) );
  INV_X1 U5224 ( .A(n8542), .ZN(n4499) );
  INV_X1 U5225 ( .A(n6263), .ZN(n4496) );
  OR2_X1 U5226 ( .A1(n6216), .A2(n4892), .ZN(n4891) );
  AND4_X1 U5227 ( .A1(n8737), .A2(n6546), .A3(n4241), .A4(n8717), .ZN(n4242)
         );
  AND2_X1 U5228 ( .A1(n6683), .A2(n6684), .ZN(n4742) );
  INV_X1 U5229 ( .A(n6685), .ZN(n4744) );
  NOR2_X1 U5230 ( .A1(n6440), .A2(n10009), .ZN(n6535) );
  INV_X1 U5231 ( .A(n6024), .ZN(n6327) );
  NAND2_X1 U5232 ( .A1(n4457), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5990) );
  INV_X1 U5233 ( .A(n6025), .ZN(n4457) );
  OAI22_X1 U5234 ( .A1(n4234), .A2(n7756), .B1(n6025), .B2(n6011), .ZN(n4654)
         );
  INV_X1 U5235 ( .A(n6986), .ZN(n4757) );
  NAND2_X1 U5236 ( .A1(n7136), .A2(n4425), .ZN(n4760) );
  NOR2_X1 U5237 ( .A1(n7082), .A2(n4762), .ZN(n4425) );
  NAND2_X1 U5238 ( .A1(n4423), .A2(n4422), .ZN(n4768) );
  INV_X1 U5239 ( .A(n7150), .ZN(n4422) );
  INV_X1 U5240 ( .A(n7149), .ZN(n4423) );
  NOR2_X1 U5241 ( .A1(n8666), .A2(n4330), .ZN(n8670) );
  OR2_X1 U5242 ( .A1(n8670), .A2(n8669), .ZN(n4764) );
  AND2_X1 U5243 ( .A1(n4419), .A2(n8681), .ZN(n8697) );
  INV_X1 U5244 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4334) );
  NOR2_X1 U5245 ( .A1(n8978), .A2(n4854), .ZN(n4853) );
  NAND2_X1 U5246 ( .A1(n8741), .A2(n8729), .ZN(n8723) );
  OAI21_X1 U5247 ( .B1(n5074), .B2(n8776), .A(n5076), .ZN(n4354) );
  AND2_X1 U5248 ( .A1(n6664), .A2(n8738), .ZN(n8752) );
  NOR2_X1 U5249 ( .A1(n9007), .A2(n5099), .ZN(n5098) );
  NOR2_X1 U5250 ( .A1(n8796), .A2(n4649), .ZN(n4647) );
  NAND2_X1 U5251 ( .A1(n8518), .A2(n8809), .ZN(n5101) );
  NAND2_X1 U5252 ( .A1(n5104), .A2(n5103), .ZN(n5102) );
  INV_X1 U5253 ( .A(n5105), .ZN(n5103) );
  INV_X1 U5254 ( .A(n8645), .ZN(n8810) );
  NAND2_X1 U5255 ( .A1(n5056), .A2(n5061), .ZN(n5055) );
  INV_X1 U5256 ( .A(n6480), .ZN(n5056) );
  NAND2_X1 U5257 ( .A1(n8845), .A2(n8844), .ZN(n8843) );
  OR2_X1 U5258 ( .A1(n5112), .A2(n4263), .ZN(n5109) );
  AND2_X1 U5259 ( .A1(n8348), .A2(n4272), .ZN(n5112) );
  AND2_X1 U5260 ( .A1(n8879), .A2(n6628), .ZN(n5062) );
  NAND2_X1 U5261 ( .A1(n8901), .A2(n4651), .ZN(n8888) );
  NAND2_X1 U5262 ( .A1(n8906), .A2(n8612), .ZN(n4651) );
  NAND2_X1 U5263 ( .A1(n8903), .A2(n8902), .ZN(n8901) );
  OR2_X1 U5264 ( .A1(n9056), .A2(n8913), .ZN(n8345) );
  INV_X1 U5265 ( .A(n8345), .ZN(n5087) );
  NAND2_X1 U5266 ( .A1(n8940), .A2(n8939), .ZN(n8938) );
  NAND2_X1 U5267 ( .A1(n4446), .A2(n4448), .ZN(n4443) );
  OAI211_X1 U5268 ( .C1(n7670), .C2(n4442), .A(n4441), .B(n4440), .ZN(n4446)
         );
  NAND2_X1 U5269 ( .A1(n4777), .A2(n6606), .ZN(n4442) );
  OR2_X1 U5270 ( .A1(n5069), .A2(n8939), .ZN(n4441) );
  NAND2_X1 U5271 ( .A1(n6474), .A2(n4777), .ZN(n4445) );
  AND2_X1 U5272 ( .A1(n5064), .A2(n4776), .ZN(n8931) );
  NAND2_X1 U5273 ( .A1(n4326), .A2(n7809), .ZN(n4776) );
  AND2_X1 U5274 ( .A1(n4444), .A2(n6621), .ZN(n5064) );
  AOI21_X1 U5275 ( .B1(n5069), .B2(n5071), .A(n5068), .ZN(n5067) );
  INV_X1 U5276 ( .A(n6616), .ZN(n5068) );
  NAND2_X1 U5277 ( .A1(n7865), .A2(n5069), .ZN(n5066) );
  AND2_X1 U5278 ( .A1(n5066), .A2(n4448), .ZN(n8009) );
  NAND2_X1 U5279 ( .A1(n7678), .A2(n7677), .ZN(n5082) );
  NAND2_X1 U5280 ( .A1(n7809), .A2(n6606), .ZN(n7865) );
  NAND2_X1 U5281 ( .A1(n7670), .A2(n6588), .ZN(n7809) );
  NAND2_X1 U5282 ( .A1(n7655), .A2(n7682), .ZN(n6473) );
  INV_X1 U5283 ( .A(n6093), .ZN(n5967) );
  NAND2_X1 U5284 ( .A1(n5073), .A2(n5072), .ZN(n7337) );
  AND2_X1 U5285 ( .A1(n6472), .A2(n6583), .ZN(n5072) );
  NAND2_X1 U5286 ( .A1(n7700), .A2(n7701), .ZN(n5073) );
  AND2_X1 U5287 ( .A1(n6579), .A2(n6583), .ZN(n7701) );
  AOI21_X1 U5288 ( .B1(n7237), .B2(n7238), .A(n4775), .ZN(n7747) );
  INV_X1 U5289 ( .A(n8659), .ZN(n8374) );
  OR2_X1 U5290 ( .A1(n7227), .A2(n6927), .ZN(n8932) );
  NAND2_X1 U5291 ( .A1(n9124), .A2(n6249), .ZN(n6494) );
  NAND2_X1 U5292 ( .A1(n7408), .A2(n6037), .ZN(n6266) );
  AND2_X1 U5293 ( .A1(n6437), .A2(n5984), .ZN(n9091) );
  INV_X2 U5294 ( .A(n10020), .ZN(n9090) );
  AND2_X1 U5295 ( .A1(n6419), .A2(n8049), .ZN(n9999) );
  INV_X1 U5296 ( .A(n6408), .ZN(n4730) );
  NOR2_X1 U5297 ( .A1(n6221), .A2(n4361), .ZN(n5959) );
  INV_X1 U5298 ( .A(n4901), .ZN(n4361) );
  NAND2_X1 U5299 ( .A1(n5957), .A2(n4903), .ZN(n4902) );
  NAND2_X1 U5300 ( .A1(n4792), .A2(n5957), .ZN(n6250) );
  AND2_X1 U5301 ( .A1(n6237), .A2(n6207), .ZN(n7693) );
  XNOR2_X1 U5302 ( .A(n4424), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U5303 ( .A1(n6103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U5304 ( .A1(n7607), .A2(n4633), .B1(n9303), .B2(n5252), .ZN(n5323)
         );
  NOR2_X1 U5305 ( .A1(n4947), .A2(n5803), .ZN(n4590) );
  INV_X1 U5306 ( .A(n4694), .ZN(n5735) );
  INV_X1 U5307 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5643) );
  INV_X1 U5308 ( .A(n9134), .ZN(n4587) );
  OR2_X1 U5309 ( .A1(n4945), .A2(n4589), .ZN(n4588) );
  INV_X1 U5310 ( .A(n9269), .ZN(n4589) );
  INV_X1 U5311 ( .A(n4946), .ZN(n4945) );
  OAI21_X1 U5312 ( .B1(n5802), .B2(n4947), .A(n9268), .ZN(n4946) );
  NAND2_X1 U5313 ( .A1(n4396), .A2(n4603), .ZN(n9174) );
  NAND2_X1 U5314 ( .A1(n9206), .A2(n4395), .ZN(n4396) );
  AND2_X1 U5315 ( .A1(n4934), .A2(n5686), .ZN(n4395) );
  AND2_X1 U5316 ( .A1(n5555), .A2(n9280), .ZN(n4954) );
  NAND2_X1 U5317 ( .A1(n5316), .A2(n4248), .ZN(n5388) );
  NAND2_X1 U5318 ( .A1(n4933), .A2(n4936), .ZN(n9227) );
  AND2_X1 U5319 ( .A1(n4597), .A2(n4310), .ZN(n4596) );
  NAND2_X1 U5320 ( .A1(n7793), .A2(n4598), .ZN(n4597) );
  OR2_X1 U5321 ( .A1(n5422), .A2(n5421), .ZN(n5441) );
  NAND2_X1 U5322 ( .A1(n9141), .A2(n9144), .ZN(n4582) );
  INV_X1 U5323 ( .A(n4608), .ZN(n4607) );
  OAI21_X1 U5324 ( .B1(n5155), .B2(n4609), .A(n5186), .ZN(n4608) );
  AOI21_X1 U5325 ( .B1(n9410), .B2(n5917), .A(n5795), .ZN(n8425) );
  AND2_X1 U5326 ( .A1(n5700), .A2(n5699), .ZN(n8116) );
  AND2_X1 U5327 ( .A1(n5626), .A2(n5625), .ZN(n8063) );
  NAND2_X1 U5328 ( .A1(n5917), .A2(n7196), .ZN(n5051) );
  INV_X1 U5329 ( .A(n6885), .ZN(n4406) );
  INV_X1 U5330 ( .A(n6884), .ZN(n4405) );
  NOR2_X1 U5331 ( .A1(n4836), .A2(n4575), .ZN(n4574) );
  AND2_X1 U5332 ( .A1(n6849), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4836) );
  INV_X1 U5333 ( .A(n6811), .ZN(n4575) );
  OR2_X1 U5334 ( .A1(n7348), .A2(n7349), .ZN(n4562) );
  INV_X1 U5335 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U5336 ( .A1(n4374), .A2(n4373), .ZN(n9364) );
  INV_X1 U5337 ( .A(n4677), .ZN(n4373) );
  NAND2_X1 U5338 ( .A1(n9396), .A2(n4679), .ZN(n4374) );
  NAND2_X1 U5339 ( .A1(n9398), .A2(n9540), .ZN(n9366) );
  AOI21_X1 U5340 ( .B1(n9396), .B2(n9397), .A(n8462), .ZN(n9373) );
  NOR2_X1 U5341 ( .A1(n8427), .A2(n5040), .ZN(n5039) );
  NAND2_X1 U5342 ( .A1(n4298), .A2(n5041), .ZN(n5038) );
  AND2_X1 U5343 ( .A1(n5820), .A2(n5846), .ZN(n9393) );
  AND2_X1 U5344 ( .A1(n9409), .A2(n9395), .ZN(n9391) );
  NOR2_X1 U5345 ( .A1(n4979), .A2(n8456), .ZN(n4977) );
  NAND2_X1 U5346 ( .A1(n9449), .A2(n8421), .ZN(n5033) );
  INV_X1 U5347 ( .A(n8454), .ZN(n4979) );
  OR2_X1 U5348 ( .A1(n5693), .A2(n9178), .ZN(n5715) );
  INV_X1 U5349 ( .A(n4682), .ZN(n4681) );
  AND2_X1 U5350 ( .A1(n9494), .A2(n8445), .ZN(n4684) );
  NAND2_X1 U5351 ( .A1(n4375), .A2(n4982), .ZN(n9502) );
  AOI21_X1 U5352 ( .B1(n4983), .B2(n9577), .A(n8263), .ZN(n4982) );
  NAND2_X1 U5353 ( .A1(n9578), .A2(n4983), .ZN(n4375) );
  NAND2_X1 U5354 ( .A1(n4509), .A2(n4508), .ZN(n9518) );
  INV_X1 U5355 ( .A(n4511), .ZN(n4508) );
  NAND2_X1 U5356 ( .A1(n9550), .A2(n5048), .ZN(n5047) );
  INV_X1 U5357 ( .A(n8415), .ZN(n5048) );
  AOI21_X1 U5358 ( .B1(n9550), .B2(n5046), .A(n4281), .ZN(n5045) );
  INV_X1 U5359 ( .A(n8416), .ZN(n5046) );
  INV_X1 U5360 ( .A(n9297), .ZN(n9579) );
  NAND2_X1 U5361 ( .A1(n8440), .A2(n8439), .ZN(n9582) );
  INV_X1 U5362 ( .A(n9578), .ZN(n8440) );
  AND2_X1 U5363 ( .A1(n8188), .A2(n8438), .ZN(n9599) );
  OR2_X1 U5364 ( .A1(n7840), .A2(n8205), .ZN(n8411) );
  AND2_X1 U5365 ( .A1(n7451), .A2(n4992), .ZN(n4991) );
  NAND2_X1 U5366 ( .A1(n7543), .A2(n8086), .ZN(n4661) );
  OR2_X1 U5367 ( .A1(n7539), .A2(n4975), .ZN(n4662) );
  AND2_X1 U5368 ( .A1(n7725), .A2(n7724), .ZN(n5034) );
  AND2_X1 U5369 ( .A1(n8252), .A2(n8088), .ZN(n8200) );
  NAND2_X1 U5370 ( .A1(n4976), .A2(n7539), .ZN(n7717) );
  INV_X1 U5371 ( .A(n7543), .ZN(n4976) );
  OAI21_X1 U5372 ( .B1(n7419), .B2(n7471), .A(n7418), .ZN(n7444) );
  AND2_X1 U5373 ( .A1(n5002), .A2(n5001), .ZN(n9624) );
  OAI22_X1 U5374 ( .A1(n9380), .A2(n4996), .B1(n9949), .B2(n9625), .ZN(n5002)
         );
  NAND2_X1 U5375 ( .A1(n4998), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U5376 ( .A1(n5791), .A2(n5790), .ZN(n9646) );
  AND2_X1 U5377 ( .A1(n5904), .A2(n8325), .ZN(n9893) );
  AND2_X1 U5378 ( .A1(n5140), .A2(n4617), .ZN(n5044) );
  XNOR2_X1 U5379 ( .A(n6501), .B(n6500), .ZN(n8404) );
  XNOR2_X1 U5380 ( .A(n4962), .B(n5170), .ZN(n5919) );
  NAND2_X1 U5381 ( .A1(n4963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4962) );
  AOI21_X1 U5382 ( .B1(n5163), .B2(n4634), .A(n4294), .ZN(n5167) );
  AND2_X1 U5383 ( .A1(n5123), .A2(n5160), .ZN(n4634) );
  NAND2_X1 U5384 ( .A1(n5754), .A2(n5750), .ZN(n5727) );
  NOR2_X1 U5385 ( .A1(n5189), .A2(n4258), .ZN(n5153) );
  XNOR2_X1 U5386 ( .A(n4557), .B(n5115), .ZN(n6736) );
  NAND2_X1 U5387 ( .A1(n4541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5174) );
  INV_X1 U5388 ( .A(n5172), .ZN(n4541) );
  NAND2_X1 U5389 ( .A1(n5174), .A2(n5173), .ZN(n5238) );
  OR2_X1 U5390 ( .A1(n10035), .A2(n9762), .ZN(n4531) );
  NAND2_X1 U5391 ( .A1(n9775), .A2(n9776), .ZN(n9777) );
  NAND2_X1 U5392 ( .A1(n6384), .A2(n6383), .ZN(n8992) );
  NAND2_X1 U5393 ( .A1(n8054), .A2(n6249), .ZN(n6384) );
  INV_X1 U5394 ( .A(n8649), .ZN(n8483) );
  NAND2_X1 U5395 ( .A1(n7938), .A2(n6249), .ZN(n4349) );
  NAND2_X1 U5396 ( .A1(n4898), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U5397 ( .A1(n6446), .A2(n6445), .ZN(n4896) );
  INV_X1 U5398 ( .A(n6448), .ZN(n4897) );
  NAND2_X1 U5399 ( .A1(n8505), .A2(n6319), .ZN(n8509) );
  INV_X1 U5400 ( .A(n8658), .ZN(n7590) );
  NAND2_X1 U5401 ( .A1(n6187), .A2(n8025), .ZN(n8039) );
  OR2_X1 U5402 ( .A1(n8549), .A2(n8932), .ZN(n8584) );
  AND2_X1 U5403 ( .A1(n6454), .A2(n6442), .ZN(n8631) );
  NAND2_X1 U5404 ( .A1(n6451), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8624) );
  INV_X1 U5405 ( .A(n8631), .ZN(n8627) );
  INV_X1 U5406 ( .A(n8617), .ZN(n8638) );
  NAND2_X1 U5407 ( .A1(n6550), .A2(n7806), .ZN(n10009) );
  XNOR2_X1 U5408 ( .A(n7010), .B(n7621), .ZN(n6988) );
  NAND2_X1 U5409 ( .A1(n7137), .A2(n7138), .ZN(n7136) );
  INV_X1 U5410 ( .A(n4760), .ZN(n7080) );
  NAND2_X1 U5411 ( .A1(n4421), .A2(n4420), .ZN(n4766) );
  INV_X1 U5412 ( .A(n7266), .ZN(n4420) );
  INV_X1 U5413 ( .A(n7265), .ZN(n4421) );
  AND2_X1 U5414 ( .A1(n4768), .A2(n4767), .ZN(n7265) );
  NAND2_X1 U5415 ( .A1(n7263), .A2(n7264), .ZN(n4767) );
  INV_X1 U5416 ( .A(n4771), .ZN(n4770) );
  OAI21_X1 U5417 ( .B1(n8699), .B2(n9978), .A(n9977), .ZN(n4771) );
  AND2_X1 U5418 ( .A1(n6398), .A2(n6459), .ZN(n8726) );
  NAND2_X1 U5419 ( .A1(n4327), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5420 ( .A1(n8739), .A2(n8930), .ZN(n4788) );
  INV_X1 U5421 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5422 ( .A1(n8036), .A2(n6249), .ZN(n6353) );
  INV_X1 U5423 ( .A(n10028), .ZN(n4658) );
  INV_X1 U5424 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4456) );
  XNOR2_X1 U5425 ( .A(n8361), .B(n8360), .ZN(n5053) );
  XNOR2_X1 U5426 ( .A(n8353), .B(n4439), .ZN(n8986) );
  OR2_X1 U5427 ( .A1(n4455), .A2(n4658), .ZN(n4454) );
  AND4_X1 U5428 ( .A1(n4429), .A2(n5956), .A3(n5941), .A4(n5955), .ZN(n4428)
         );
  NAND2_X1 U5429 ( .A1(n4623), .A2(n4625), .ZN(n4407) );
  NAND2_X1 U5430 ( .A1(n4949), .A2(n5802), .ZN(n9189) );
  INV_X1 U5431 ( .A(n9288), .ZN(n9235) );
  NAND2_X1 U5432 ( .A1(n5927), .A2(n6869), .ZN(n9271) );
  OR2_X1 U5433 ( .A1(n5921), .A2(n9927), .ZN(n9275) );
  INV_X1 U5434 ( .A(n9294), .ZN(n9398) );
  NAND2_X1 U5435 ( .A1(n4699), .A2(n5772), .ZN(n9444) );
  OR2_X1 U5436 ( .A1(n9423), .A2(n5848), .ZN(n4699) );
  NAND2_X1 U5437 ( .A1(n5742), .A2(n5741), .ZN(n9456) );
  OR2_X1 U5438 ( .A1(n9436), .A2(n5848), .ZN(n5742) );
  INV_X1 U5439 ( .A(n9179), .ZN(n9465) );
  INV_X1 U5440 ( .A(n8116), .ZN(n9481) );
  NAND2_X1 U5441 ( .A1(n5678), .A2(n5677), .ZN(n9496) );
  NAND2_X1 U5442 ( .A1(n7073), .A2(n7071), .ZN(n6772) );
  AOI21_X1 U5443 ( .B1(n9343), .B2(n9841), .A(n9853), .ZN(n9342) );
  XNOR2_X1 U5444 ( .A(n8429), .B(n8466), .ZN(n9627) );
  NAND2_X1 U5445 ( .A1(n4984), .A2(n8468), .ZN(n4692) );
  NAND2_X1 U5446 ( .A1(n4985), .A2(n9603), .ZN(n4984) );
  NAND2_X1 U5447 ( .A1(n9516), .A2(n8417), .ZN(n9487) );
  OR2_X1 U5448 ( .A1(n7178), .A2(n7177), .ZN(n9897) );
  OR2_X1 U5449 ( .A1(n5909), .A2(n9949), .ZN(n9566) );
  CLKBUF_X1 U5450 ( .A(n5141), .Z(n9746) );
  INV_X1 U5451 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U5452 ( .A1(n4619), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4636) );
  XNOR2_X1 U5453 ( .A(n9777), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U5454 ( .A1(n10235), .A2(n10236), .ZN(n10234) );
  NAND2_X1 U5455 ( .A1(n10040), .A2(n10041), .ZN(n10039) );
  NAND2_X1 U5456 ( .A1(n10039), .A2(n4521), .ZN(n10231) );
  NAND2_X1 U5457 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  INV_X1 U5458 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5459 ( .A1(n10231), .A2(n10232), .ZN(n10230) );
  NAND2_X1 U5460 ( .A1(n8193), .A2(n8167), .ZN(n8076) );
  INV_X1 U5461 ( .A(n8076), .ZN(n4820) );
  INV_X1 U5462 ( .A(n8089), .ZN(n4808) );
  INV_X1 U5463 ( .A(n8084), .ZN(n4807) );
  OAI22_X1 U5464 ( .A1(n6573), .A2(n6572), .B1(n4236), .B2(n6571), .ZN(n6580)
         );
  NAND2_X1 U5465 ( .A1(n4491), .A2(n4236), .ZN(n4490) );
  NAND2_X1 U5466 ( .A1(n6600), .A2(n6588), .ZN(n4491) );
  NAND2_X1 U5467 ( .A1(n4473), .A2(n8339), .ZN(n4470) );
  OAI21_X1 U5468 ( .B1(n6589), .B2(n6603), .A(n4488), .ZN(n6592) );
  AND2_X1 U5469 ( .A1(n7864), .A2(n6588), .ZN(n4488) );
  NAND2_X1 U5470 ( .A1(n4244), .A2(n6615), .ZN(n4472) );
  NAND2_X1 U5471 ( .A1(n4793), .A2(n4542), .ZN(n8121) );
  INV_X1 U5472 ( .A(n4798), .ZN(n4795) );
  NAND2_X1 U5473 ( .A1(n4751), .A2(n4750), .ZN(n6638) );
  NOR2_X1 U5474 ( .A1(n6630), .A2(n6479), .ZN(n4750) );
  AND2_X1 U5475 ( .A1(n8127), .A2(n9427), .ZN(n4813) );
  INV_X1 U5476 ( .A(n8062), .ZN(n8130) );
  NOR2_X1 U5477 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  INV_X1 U5478 ( .A(n8138), .ZN(n4547) );
  NOR2_X1 U5479 ( .A1(n4549), .A2(n4809), .ZN(n4548) );
  NAND2_X1 U5480 ( .A1(n4484), .A2(n6649), .ZN(n4483) );
  INV_X1 U5481 ( .A(n6661), .ZN(n4736) );
  NAND2_X1 U5482 ( .A1(n9309), .A2(n4974), .ZN(n8238) );
  AND2_X1 U5483 ( .A1(n9444), .A2(n4698), .ZN(n8271) );
  NAND2_X1 U5484 ( .A1(n6319), .A2(n4884), .ZN(n4883) );
  INV_X1 U5485 ( .A(n6319), .ZN(n4885) );
  NAND2_X1 U5486 ( .A1(n4481), .A2(n4478), .ZN(n6655) );
  NAND2_X1 U5487 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U5488 ( .A1(n4479), .A2(n6688), .ZN(n4478) );
  NOR2_X1 U5489 ( .A1(n6648), .A2(n6688), .ZN(n4482) );
  INV_X1 U5490 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U5491 ( .A1(n8168), .A2(n8169), .ZN(n4824) );
  INV_X1 U5492 ( .A(n9892), .ZN(n4974) );
  INV_X1 U5493 ( .A(n4923), .ZN(n4922) );
  OAI21_X1 U5494 ( .B1(n4925), .B2(n4924), .A(n5836), .ZN(n4923) );
  INV_X1 U5495 ( .A(n5807), .ZN(n4924) );
  AND2_X1 U5496 ( .A1(n4712), .A2(n5633), .ZN(n4708) );
  INV_X1 U5497 ( .A(n5610), .ZN(n4710) );
  NAND2_X1 U5498 ( .A1(n4567), .A2(n4569), .ZN(n4565) );
  NAND2_X1 U5499 ( .A1(n4864), .A2(n4863), .ZN(n4862) );
  NOR2_X1 U5500 ( .A1(n6295), .A2(n6294), .ZN(n4359) );
  XNOR2_X1 U5501 ( .A(n9024), .B(n6077), .ZN(n6332) );
  AND2_X1 U5502 ( .A1(n8656), .A2(n6331), .ZN(n6085) );
  NOR2_X1 U5503 ( .A1(n5060), .A2(n4431), .ZN(n4430) );
  NOR2_X1 U5504 ( .A1(n7945), .A2(n8939), .ZN(n4432) );
  AND2_X1 U5505 ( .A1(n4434), .A2(n8346), .ZN(n4433) );
  AOI21_X1 U5506 ( .B1(n4741), .B2(n4279), .A(n4739), .ZN(n4738) );
  INV_X1 U5507 ( .A(n6679), .ZN(n4739) );
  INV_X1 U5508 ( .A(n4741), .ZN(n4740) );
  AND2_X1 U5509 ( .A1(n5093), .A2(n8350), .ZN(n5092) );
  NAND2_X1 U5510 ( .A1(n5094), .A2(n8734), .ZN(n5093) );
  OR2_X1 U5511 ( .A1(n5114), .A2(n8349), .ZN(n5105) );
  INV_X1 U5512 ( .A(n5106), .ZN(n5104) );
  NOR2_X1 U5513 ( .A1(n6480), .A2(n4256), .ZN(n5059) );
  NOR2_X1 U5514 ( .A1(n4848), .A2(n9045), .ZN(n4847) );
  INV_X1 U5515 ( .A(n8921), .ZN(n4848) );
  NOR2_X1 U5516 ( .A1(n6231), .A2(n5970), .ZN(n6225) );
  OR2_X1 U5517 ( .A1(n5065), .A2(n5069), .ZN(n4444) );
  AND2_X1 U5518 ( .A1(n7295), .A2(n6560), .ZN(n6559) );
  NAND2_X1 U5519 ( .A1(n7590), .A2(n7746), .ZN(n6567) );
  INV_X1 U5520 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4851) );
  AND2_X1 U5521 ( .A1(n4840), .A2(n4839), .ZN(n4838) );
  INV_X1 U5522 ( .A(n9003), .ZN(n4839) );
  AOI21_X1 U5523 ( .B1(n9999), .B2(n10005), .A(n10006), .ZN(n7617) );
  OR2_X1 U5524 ( .A1(n10003), .A2(n6430), .ZN(n7225) );
  AND2_X1 U5525 ( .A1(n9999), .A2(n10002), .ZN(n6430) );
  NOR2_X1 U5526 ( .A1(n4902), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4901) );
  INV_X1 U5527 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6205) );
  OR2_X1 U5528 ( .A1(n6103), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6118) );
  OR2_X1 U5529 ( .A1(n6089), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6103) );
  INV_X1 U5530 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4426) );
  INV_X1 U5531 ( .A(n5806), .ZN(n4947) );
  NOR2_X1 U5532 ( .A1(n4938), .A2(n4935), .ZN(n4934) );
  INV_X1 U5533 ( .A(n5606), .ZN(n4935) );
  INV_X1 U5534 ( .A(n5661), .ZN(n4938) );
  INV_X1 U5535 ( .A(n5872), .ZN(n5798) );
  AND3_X1 U5536 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5315) );
  INV_X1 U5537 ( .A(n5707), .ZN(n4602) );
  NOR2_X1 U5538 ( .A1(n5547), .A2(n5523), .ZN(n4700) );
  INV_X1 U5539 ( .A(n5524), .ZN(n5522) );
  INV_X1 U5540 ( .A(n5902), .ZN(n8313) );
  NOR2_X1 U5541 ( .A1(n7978), .A2(n4829), .ZN(n9317) );
  AND2_X1 U5542 ( .A1(n7979), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4829) );
  AND2_X1 U5543 ( .A1(n9828), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5544 ( .A1(n4288), .A2(n4246), .ZN(n4518) );
  NAND2_X1 U5545 ( .A1(n9454), .A2(n5015), .ZN(n5014) );
  NOR2_X1 U5546 ( .A1(n8436), .A2(n4973), .ZN(n4972) );
  INV_X1 U5547 ( .A(n8092), .ZN(n4973) );
  NOR2_X1 U5548 ( .A1(n4994), .A2(n9715), .ZN(n4993) );
  INV_X1 U5549 ( .A(n4995), .ZN(n4994) );
  NOR2_X1 U5550 ( .A1(n9720), .A2(n7536), .ZN(n4995) );
  NOR2_X1 U5551 ( .A1(n7469), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5552 ( .A1(n8193), .A2(n8291), .ZN(n7471) );
  AND2_X1 U5553 ( .A1(n4990), .A2(n4989), .ZN(n4988) );
  INV_X1 U5554 ( .A(n7173), .ZN(n4990) );
  NOR2_X1 U5555 ( .A1(n6757), .A2(n8236), .ZN(n7316) );
  AND2_X1 U5556 ( .A1(n4988), .A2(n4987), .ZN(n9929) );
  NAND2_X1 U5557 ( .A1(n8236), .A2(n4974), .ZN(n7173) );
  NOR2_X1 U5558 ( .A1(n5189), .A2(n5157), .ZN(n5158) );
  INV_X1 U5559 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5170) );
  AND2_X1 U5560 ( .A1(n5859), .A2(n5841), .ZN(n5857) );
  NOR2_X1 U5561 ( .A1(n5808), .A2(n4926), .ZN(n4925) );
  INV_X1 U5562 ( .A(n5785), .ZN(n4926) );
  INV_X1 U5563 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5164) );
  AND2_X1 U5564 ( .A1(n4300), .A2(n4571), .ZN(n4570) );
  OR2_X1 U5565 ( .A1(n4931), .A2(n4572), .ZN(n4571) );
  OR2_X1 U5566 ( .A1(n5417), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U5567 ( .A1(n5304), .A2(n5303), .ZN(n5308) );
  XNOR2_X1 U5568 ( .A(n5305), .B(SI_5_), .ZN(n5303) );
  OAI21_X1 U5569 ( .B1(n5270), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5248), .ZN(
        n5266) );
  INV_X1 U5570 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4460) );
  INV_X1 U5571 ( .A(n6070), .ZN(n4880) );
  NOR2_X1 U5572 ( .A1(n8618), .A2(n4723), .ZN(n4722) );
  INV_X1 U5573 ( .A(n8733), .ZN(n8476) );
  NAND2_X1 U5574 ( .A1(n8482), .A2(n6216), .ZN(n8489) );
  NOR2_X1 U5575 ( .A1(n4726), .A2(n4721), .ZN(n4717) );
  INV_X1 U5576 ( .A(n4720), .ZN(n4719) );
  OAI21_X1 U5577 ( .B1(n4722), .B2(n4721), .A(n8472), .ZN(n4720) );
  NAND2_X1 U5578 ( .A1(n4359), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6323) );
  NOR2_X1 U5579 ( .A1(n4714), .A2(n8506), .ZN(n6319) );
  NAND2_X1 U5580 ( .A1(n4715), .A2(n8504), .ZN(n4714) );
  INV_X1 U5581 ( .A(n8569), .ZN(n4715) );
  XNOR2_X1 U5582 ( .A(n6332), .B(n4285), .ZN(n8506) );
  AND2_X1 U5583 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5968) );
  INV_X1 U5584 ( .A(n6177), .ZN(n5969) );
  NAND2_X1 U5585 ( .A1(n8489), .A2(n6220), .ZN(n8530) );
  OR2_X1 U5586 ( .A1(n4262), .A2(n8498), .ZN(n6357) );
  XNOR2_X1 U5587 ( .A(n6077), .B(n8391), .ZN(n6032) );
  NAND2_X1 U5588 ( .A1(n4501), .A2(n7571), .ZN(n4360) );
  NAND2_X1 U5589 ( .A1(n5971), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6295) );
  INV_X1 U5590 ( .A(n6283), .ZN(n5971) );
  INV_X1 U5591 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n6294) );
  INV_X1 U5592 ( .A(n4359), .ZN(n6309) );
  INV_X1 U5593 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8582) );
  NOR2_X1 U5594 ( .A1(n7856), .A2(n4870), .ZN(n4869) );
  INV_X1 U5595 ( .A(n6137), .ZN(n4870) );
  INV_X1 U5596 ( .A(n4864), .ZN(n8591) );
  INV_X1 U5597 ( .A(n6014), .ZN(n8593) );
  INV_X1 U5598 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U5599 ( .A1(n4358), .A2(n4357), .ZN(n6283) );
  NOR2_X1 U5600 ( .A1(n8547), .A2(n6267), .ZN(n4357) );
  INV_X1 U5601 ( .A(n6268), .ZN(n4358) );
  OR2_X1 U5602 ( .A1(n6171), .A2(n6170), .ZN(n6188) );
  INV_X1 U5603 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7159) );
  AND2_X1 U5604 ( .A1(n4766), .A2(n4765), .ZN(n7910) );
  NAND2_X1 U5605 ( .A1(n7691), .A2(n8016), .ZN(n4765) );
  NAND2_X1 U5606 ( .A1(n4764), .A2(n4763), .ZN(n4419) );
  NAND2_X1 U5607 ( .A1(n8678), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4763) );
  INV_X1 U5608 ( .A(n4854), .ZN(n4852) );
  INV_X1 U5609 ( .A(n5075), .ZN(n8739) );
  OAI21_X1 U5610 ( .B1(n8776), .B2(n5074), .A(n5076), .ZN(n5075) );
  NAND2_X1 U5611 ( .A1(n8813), .A2(n4840), .ZN(n8784) );
  NAND2_X1 U5612 ( .A1(n8813), .A2(n8355), .ZN(n8814) );
  NAND2_X1 U5613 ( .A1(n8843), .A2(n6641), .ZN(n8825) );
  NAND2_X1 U5614 ( .A1(n8942), .A2(n4847), .ZN(n8894) );
  NAND2_X1 U5615 ( .A1(n8940), .A2(n4267), .ZN(n5086) );
  NAND2_X1 U5616 ( .A1(n5087), .A2(n5088), .ZN(n5084) );
  INV_X1 U5617 ( .A(n8346), .ZN(n8902) );
  NAND2_X1 U5618 ( .A1(n6225), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6268) );
  AND2_X1 U5619 ( .A1(n8941), .A2(n8949), .ZN(n8942) );
  NAND2_X1 U5620 ( .A1(n8942), .A2(n8921), .ZN(n8918) );
  OR2_X1 U5621 ( .A1(n6192), .A2(n7159), .ZN(n6231) );
  NOR2_X2 U5622 ( .A1(n8018), .A2(n9061), .ZN(n8941) );
  NAND2_X1 U5623 ( .A1(n4652), .A2(n7945), .ZN(n8013) );
  INV_X1 U5624 ( .A(n8651), .ZN(n8030) );
  NAND2_X1 U5625 ( .A1(n4355), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6177) );
  INV_X1 U5626 ( .A(n6142), .ZN(n4355) );
  AND2_X1 U5627 ( .A1(n7869), .A2(n6604), .ZN(n5063) );
  NAND2_X1 U5628 ( .A1(n4356), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6142) );
  INV_X1 U5629 ( .A(n6125), .ZN(n4356) );
  NAND2_X1 U5630 ( .A1(n7641), .A2(n4858), .ZN(n7672) );
  OR2_X1 U5631 ( .A1(n6107), .A2(n7573), .ZN(n6125) );
  NAND2_X1 U5632 ( .A1(n7641), .A2(n7645), .ZN(n7661) );
  NAND2_X1 U5633 ( .A1(n7337), .A2(n6593), .ZN(n7636) );
  NAND2_X1 U5634 ( .A1(n7337), .A2(n4277), .ZN(n7638) );
  NAND2_X1 U5635 ( .A1(n6057), .A2(n4286), .ZN(n6093) );
  AND2_X1 U5636 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6057) );
  NAND2_X1 U5637 ( .A1(n6057), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6079) );
  INV_X1 U5638 ( .A(n6542), .ZN(n7748) );
  NAND2_X1 U5639 ( .A1(n6567), .A2(n7295), .ZN(n6542) );
  INV_X1 U5640 ( .A(n7253), .ZN(n6470) );
  NAND2_X1 U5641 ( .A1(n9091), .A2(n4769), .ZN(n7219) );
  NAND2_X1 U5642 ( .A1(n7510), .A2(n7736), .ZN(n7732) );
  INV_X1 U5643 ( .A(n7225), .ZN(n7303) );
  AND2_X1 U5644 ( .A1(n7224), .A2(n7504), .ZN(n7304) );
  INV_X1 U5645 ( .A(n9091), .ZN(n10022) );
  AND2_X1 U5646 ( .A1(n7304), .A2(n7225), .ZN(n7618) );
  XNOR2_X1 U5647 ( .A(n6457), .B(n6456), .ZN(n6927) );
  INV_X1 U5648 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U5649 ( .A(n6410), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U5650 ( .A1(n6409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6410) );
  OR2_X1 U5651 ( .A1(n6221), .A2(n6408), .ZN(n6409) );
  NAND2_X1 U5652 ( .A1(n6018), .A2(n6017), .ZN(n6038) );
  NOR2_X1 U5653 ( .A1(n5531), .A2(n4957), .ZN(n4956) );
  INV_X1 U5654 ( .A(n4959), .ZN(n4957) );
  OR2_X1 U5655 ( .A1(n5500), .A2(n7565), .ZN(n5524) );
  INV_X1 U5656 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U5657 ( .A1(n5619), .A2(n4703), .ZN(n5671) );
  NAND2_X1 U5658 ( .A1(n5316), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U5659 ( .A1(n4953), .A2(n4951), .ZN(n5583) );
  NOR2_X1 U5660 ( .A1(n4954), .A2(n4952), .ZN(n4951) );
  INV_X1 U5661 ( .A(n9196), .ZN(n4952) );
  NAND3_X1 U5662 ( .A1(n5200), .A2(n5202), .A3(n5201), .ZN(n6876) );
  NAND2_X1 U5663 ( .A1(n5252), .A2(n7387), .ZN(n5205) );
  NAND2_X1 U5664 ( .A1(n5207), .A2(n6757), .ZN(n4402) );
  INV_X1 U5665 ( .A(n4598), .ZN(n4595) );
  INV_X1 U5666 ( .A(n4303), .ZN(n5185) );
  AND2_X1 U5667 ( .A1(n5227), .A2(n5228), .ZN(n6862) );
  INV_X1 U5668 ( .A(n6863), .ZN(n4400) );
  NAND2_X1 U5669 ( .A1(n5522), .A2(n4700), .ZN(n5569) );
  NAND2_X1 U5670 ( .A1(n5522), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5548) );
  INV_X1 U5671 ( .A(n5746), .ZN(n5876) );
  NAND2_X1 U5672 ( .A1(n4697), .A2(n4821), .ZN(n4696) );
  AND2_X1 U5673 ( .A1(n8174), .A2(n8312), .ZN(n4695) );
  INV_X1 U5674 ( .A(n8173), .ZN(n4821) );
  AND2_X1 U5675 ( .A1(n9468), .A2(n8287), .ZN(n8328) );
  NAND2_X1 U5676 ( .A1(n6833), .A2(n6790), .ZN(n6884) );
  NAND2_X1 U5677 ( .A1(n4561), .A2(n6841), .ZN(n7073) );
  AND2_X1 U5678 ( .A1(n6769), .A2(n6880), .ZN(n4561) );
  AND2_X1 U5679 ( .A1(n4392), .A2(n4391), .ZN(n6792) );
  NAND2_X1 U5680 ( .A1(n7077), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4391) );
  NOR2_X1 U5681 ( .A1(n6801), .A2(n4404), .ZN(n6822) );
  AND2_X1 U5682 ( .A1(n6849), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4404) );
  AND2_X1 U5683 ( .A1(n6822), .A2(n6821), .ZN(n6819) );
  OAI21_X1 U5684 ( .B1(n6819), .B2(n6804), .A(n6803), .ZN(n7026) );
  NAND2_X1 U5685 ( .A1(n4560), .A2(n4324), .ZN(n4828) );
  INV_X1 U5686 ( .A(n7017), .ZN(n4560) );
  AOI21_X1 U5687 ( .B1(n7026), .B2(n7025), .A(n7024), .ZN(n7114) );
  NOR2_X1 U5688 ( .A1(n7101), .A2(n4826), .ZN(n7103) );
  AND2_X1 U5689 ( .A1(n7102), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U5690 ( .A1(n7103), .A2(n7104), .ZN(n7346) );
  NAND2_X1 U5691 ( .A1(n4562), .A2(n4325), .ZN(n4831) );
  OR2_X1 U5692 ( .A1(n7981), .A2(n7982), .ZN(n9315) );
  NAND2_X1 U5693 ( .A1(n9310), .A2(n4393), .ZN(n9331) );
  NAND2_X1 U5694 ( .A1(n9316), .A2(n4394), .ZN(n4393) );
  INV_X1 U5695 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n4394) );
  NOR2_X1 U5696 ( .A1(n9324), .A2(n4628), .ZN(n9825) );
  AND2_X1 U5697 ( .A1(n9325), .A2(n9333), .ZN(n4628) );
  NOR2_X1 U5698 ( .A1(n9825), .A2(n9824), .ZN(n9823) );
  INV_X1 U5699 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5564) );
  INV_X1 U5700 ( .A(n9835), .ZN(n4579) );
  OR2_X1 U5701 ( .A1(n9823), .A2(n4637), .ZN(n4580) );
  OR2_X1 U5702 ( .A1(n9856), .A2(n9857), .ZN(n4399) );
  OAI22_X1 U5703 ( .A1(n9823), .A2(n4578), .B1(n4579), .B2(n4834), .ZN(n9849)
         );
  OR2_X1 U5704 ( .A1(n4834), .A2(n4637), .ZN(n4578) );
  AND2_X1 U5705 ( .A1(n9839), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4834) );
  NOR2_X1 U5706 ( .A1(n9849), .A2(n9850), .ZN(n9848) );
  AND2_X1 U5707 ( .A1(n6781), .A2(n8055), .ZN(n9330) );
  NAND2_X1 U5708 ( .A1(n8154), .A2(n8153), .ZN(n9354) );
  INV_X1 U5709 ( .A(n5001), .ZN(n9355) );
  NAND2_X1 U5710 ( .A1(n4676), .A2(n4986), .ZN(n4671) );
  NOR2_X1 U5711 ( .A1(n4676), .A2(n4986), .ZN(n4668) );
  AND2_X1 U5712 ( .A1(n5911), .A2(n5865), .ZN(n9361) );
  NAND2_X1 U5713 ( .A1(n9398), .A2(n9542), .ZN(n9400) );
  NAND2_X1 U5714 ( .A1(n4663), .A2(n4664), .ZN(n9413) );
  AOI21_X1 U5715 ( .B1(n9427), .B2(n4665), .A(n8061), .ZN(n4664) );
  INV_X1 U5716 ( .A(n8458), .ZN(n4665) );
  NOR2_X1 U5717 ( .A1(n5012), .A2(n9652), .ZN(n5009) );
  NOR2_X1 U5718 ( .A1(n4289), .A2(n5032), .ZN(n5031) );
  AND2_X1 U5719 ( .A1(n5735), .A2(n5716), .ZN(n9452) );
  NOR2_X1 U5720 ( .A1(n9475), .A2(n9667), .ZN(n9467) );
  NOR2_X1 U5721 ( .A1(n9475), .A2(n5014), .ZN(n9450) );
  INV_X1 U5722 ( .A(n9480), .ZN(n4381) );
  INV_X1 U5723 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9178) );
  AND2_X1 U5724 ( .A1(n4703), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n4702) );
  AOI21_X1 U5725 ( .B1(n5023), .B2(n5025), .A(n5022), .ZN(n5021) );
  NOR2_X1 U5726 ( .A1(n9478), .A2(n9169), .ZN(n5022) );
  OR2_X1 U5727 ( .A1(n5593), .A2(n9209), .ZN(n5620) );
  NAND2_X1 U5728 ( .A1(n5619), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U5729 ( .A1(n5006), .A2(n9687), .ZN(n5003) );
  NAND2_X1 U5730 ( .A1(n9605), .A2(n5005), .ZN(n9545) );
  INV_X1 U5731 ( .A(n5006), .ZN(n5005) );
  NAND2_X1 U5732 ( .A1(n9605), .A2(n5008), .ZN(n9565) );
  NAND2_X1 U5733 ( .A1(n9582), .A2(n8441), .ZN(n9556) );
  AOI21_X1 U5734 ( .B1(n4969), .B2(n4971), .A(n4967), .ZN(n4966) );
  NAND2_X1 U5735 ( .A1(n7843), .A2(n4969), .ZN(n4376) );
  INV_X1 U5736 ( .A(n8438), .ZN(n4967) );
  AND2_X1 U5737 ( .A1(n9605), .A2(n9584), .ZN(n9586) );
  NAND2_X1 U5738 ( .A1(n4968), .A2(n8435), .ZN(n9596) );
  NAND2_X1 U5739 ( .A1(n7843), .A2(n4972), .ZN(n4968) );
  NAND2_X1 U5740 ( .A1(n7843), .A2(n8092), .ZN(n8437) );
  AND4_X1 U5741 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n9597)
         );
  AND2_X1 U5742 ( .A1(n8092), .A2(n8094), .ZN(n8204) );
  NAND2_X1 U5743 ( .A1(n4993), .A2(n7451), .ZN(n7781) );
  AND2_X1 U5744 ( .A1(n7451), .A2(n9948), .ZN(n7547) );
  NAND2_X1 U5745 ( .A1(n7451), .A2(n4995), .ZN(n7720) );
  NAND2_X1 U5746 ( .A1(n7541), .A2(n8084), .ZN(n7543) );
  OAI211_X1 U5747 ( .C1(n7436), .C2(n4386), .A(n4384), .B(n8085), .ZN(n7541)
         );
  NAND2_X1 U5748 ( .A1(n4385), .A2(n8083), .ZN(n4384) );
  NAND2_X1 U5749 ( .A1(n7422), .A2(n7424), .ZN(n7538) );
  NAND2_X1 U5750 ( .A1(n6723), .A2(n5327), .ZN(n5314) );
  NAND2_X1 U5751 ( .A1(n7475), .A2(n7417), .ZN(n7443) );
  INV_X1 U5752 ( .A(n4385), .ZN(n4387) );
  AND4_X1 U5753 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n9926)
         );
  NAND2_X1 U5754 ( .A1(n7396), .A2(n4814), .ZN(n9919) );
  NAND2_X1 U5755 ( .A1(n4988), .A2(n7175), .ZN(n7402) );
  NAND2_X1 U5756 ( .A1(n4990), .A2(n7175), .ZN(n7401) );
  NAND2_X1 U5757 ( .A1(n7317), .A2(n7314), .ZN(n7410) );
  NAND2_X1 U5758 ( .A1(n7312), .A2(n7311), .ZN(n7448) );
  NAND2_X1 U5759 ( .A1(n8335), .A2(n5327), .ZN(n4907) );
  INV_X1 U5760 ( .A(n7429), .ZN(n9933) );
  INV_X1 U5761 ( .A(n9719), .ZN(n9952) );
  AOI21_X1 U5762 ( .B1(n6707), .B2(n4240), .A(n5050), .ZN(n5049) );
  INV_X1 U5763 ( .A(n9893), .ZN(n9947) );
  XNOR2_X1 U5764 ( .A(n6526), .B(n6525), .ZN(n9119) );
  INV_X1 U5765 ( .A(n5781), .ZN(n4904) );
  XNOR2_X1 U5766 ( .A(n4706), .B(n5708), .ZN(n7805) );
  AND3_X1 U5767 ( .A1(n4552), .A2(n4554), .A3(n4550), .ZN(n4620) );
  AND2_X1 U5768 ( .A1(n4555), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5769 ( .A1(n4711), .A2(n5610), .ZN(n5634) );
  NAND2_X1 U5770 ( .A1(n5586), .A2(n5585), .ZN(n5612) );
  NAND2_X1 U5771 ( .A1(n4911), .A2(n5536), .ZN(n5559) );
  NAND2_X1 U5772 ( .A1(n5510), .A2(n4916), .ZN(n4911) );
  OR2_X1 U5773 ( .A1(n5514), .A2(n5513), .ZN(n5516) );
  NOR2_X1 U5774 ( .A1(n5516), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U5775 ( .A1(n5510), .A2(n5509), .ZN(n5538) );
  NAND2_X1 U5776 ( .A1(n4566), .A2(n5490), .ZN(n5508) );
  NAND2_X1 U5777 ( .A1(n4928), .A2(n5459), .ZN(n5487) );
  AND2_X1 U5778 ( .A1(n10076), .A2(n5151), .ZN(n4554) );
  INV_X1 U5779 ( .A(n4555), .ZN(n5137) );
  XNOR2_X1 U5780 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n4534) );
  AND2_X1 U5781 ( .A1(n10037), .A2(n9763), .ZN(n4529) );
  AND2_X1 U5782 ( .A1(n4528), .A2(n4525), .ZN(n9769) );
  NAND2_X1 U5783 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  INV_X1 U5784 ( .A(n10227), .ZN(n4528) );
  INV_X1 U5785 ( .A(n10228), .ZN(n4527) );
  NAND2_X1 U5786 ( .A1(n4539), .A2(n9773), .ZN(n9774) );
  NAND2_X1 U5787 ( .A1(n10238), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5788 ( .A1(n4879), .A2(n4877), .ZN(n7526) );
  NAND2_X1 U5789 ( .A1(n4878), .A2(n7580), .ZN(n4877) );
  NAND2_X1 U5790 ( .A1(n4718), .A2(n6382), .ZN(n8473) );
  NAND2_X1 U5791 ( .A1(n4724), .A2(n4722), .ZN(n4718) );
  NAND2_X1 U5792 ( .A1(n7820), .A2(n6137), .ZN(n7857) );
  NAND2_X1 U5793 ( .A1(n6736), .A2(n6249), .ZN(n4493) );
  AND2_X1 U5794 ( .A1(n6056), .A2(n6055), .ZN(n7591) );
  NAND2_X1 U5795 ( .A1(n4500), .A2(n4887), .ZN(n8543) );
  NAND2_X1 U5796 ( .A1(n4360), .A2(n6117), .ZN(n7823) );
  INV_X1 U5797 ( .A(n8608), .ZN(n8629) );
  NAND2_X1 U5798 ( .A1(n7941), .A2(n6249), .ZN(n6322) );
  AOI21_X1 U5799 ( .B1(n4498), .B2(n4890), .A(n4496), .ZN(n4495) );
  NAND2_X1 U5800 ( .A1(n4886), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U5801 ( .A1(n7580), .A2(n7579), .ZN(n7578) );
  NAND2_X1 U5802 ( .A1(n7587), .A2(n6070), .ZN(n7579) );
  NAND2_X1 U5803 ( .A1(n4724), .A2(n8526), .ZN(n8619) );
  INV_X1 U5804 ( .A(n8583), .ZN(n8636) );
  NAND2_X1 U5805 ( .A1(n6694), .A2(n6751), .ZN(n4749) );
  XNOR2_X1 U5806 ( .A(n4438), .B(n6532), .ZN(n6549) );
  INV_X1 U5807 ( .A(n6528), .ZN(n8703) );
  NAND2_X1 U5808 ( .A1(n6405), .A2(n6404), .ZN(n8740) );
  NAND4_X1 U5809 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n8658)
         );
  NAND2_X1 U5810 ( .A1(n6027), .A2(n4276), .ZN(n8659) );
  AND2_X1 U5811 ( .A1(n6012), .A2(n6013), .ZN(n4655) );
  INV_X1 U5812 ( .A(n4654), .ZN(n4653) );
  INV_X2 U5813 ( .A(P2_U3966), .ZN(n8661) );
  NAND4_X1 U5814 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n6469)
         );
  NAND2_X1 U5815 ( .A1(n6999), .A2(n6986), .ZN(n6987) );
  NAND2_X1 U5816 ( .A1(n6987), .A2(n6988), .ZN(n7011) );
  INV_X1 U5817 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7573) );
  AND2_X1 U5818 ( .A1(n4754), .A2(n7013), .ZN(n4753) );
  OR2_X1 U5819 ( .A1(n4261), .A2(n6988), .ZN(n4754) );
  INV_X1 U5820 ( .A(n6988), .ZN(n4758) );
  NAND2_X1 U5821 ( .A1(n7086), .A2(n7813), .ZN(n4759) );
  INV_X1 U5822 ( .A(n4768), .ZN(n7262) );
  OR2_X1 U5823 ( .A1(n6912), .A2(n8362), .ZN(n9978) );
  INV_X1 U5824 ( .A(n4764), .ZN(n8677) );
  NAND2_X1 U5825 ( .A1(n6929), .A2(n6927), .ZN(n9977) );
  NAND2_X1 U5826 ( .A1(n4418), .A2(n4416), .ZN(n8679) );
  INV_X1 U5827 ( .A(n8697), .ZN(n4418) );
  NAND2_X1 U5828 ( .A1(n4417), .A2(n8693), .ZN(n4416) );
  INV_X1 U5829 ( .A(n4419), .ZN(n4417) );
  INV_X1 U5830 ( .A(n8702), .ZN(n9975) );
  NAND2_X1 U5831 ( .A1(n8404), .A2(n6249), .ZN(n6503) );
  NAND2_X1 U5832 ( .A1(n8335), .A2(n6249), .ZN(n6395) );
  NAND2_X1 U5833 ( .A1(n4354), .A2(n6485), .ZN(n8718) );
  INV_X1 U5834 ( .A(n8992), .ZN(n8745) );
  NAND2_X1 U5835 ( .A1(n6397), .A2(n6372), .ZN(n8758) );
  NAND2_X1 U5836 ( .A1(n8048), .A2(n6249), .ZN(n6368) );
  NAND2_X1 U5837 ( .A1(n5091), .A2(n5094), .ZN(n8749) );
  NAND2_X1 U5838 ( .A1(n8789), .A2(n8765), .ZN(n5091) );
  NOR2_X1 U5839 ( .A1(n8789), .A2(n5098), .ZN(n8762) );
  NAND2_X1 U5840 ( .A1(n4642), .A2(n4644), .ZN(n8790) );
  NAND2_X1 U5841 ( .A1(n8795), .A2(n6651), .ZN(n8777) );
  AND2_X1 U5842 ( .A1(n4648), .A2(n4650), .ZN(n8804) );
  NAND2_X1 U5843 ( .A1(n4648), .A2(n4647), .ZN(n9014) );
  INV_X1 U5844 ( .A(n5100), .ZN(n8824) );
  AOI21_X1 U5845 ( .B1(n5108), .B2(n5106), .A(n5114), .ZN(n5100) );
  AND2_X1 U5846 ( .A1(n8849), .A2(n8848), .ZN(n9032) );
  NAND2_X1 U5847 ( .A1(n6293), .A2(n6292), .ZN(n9029) );
  NAND2_X1 U5848 ( .A1(n7788), .A2(n6037), .ZN(n6293) );
  NAND2_X1 U5849 ( .A1(n5108), .A2(n5109), .ZN(n8842) );
  AND2_X1 U5850 ( .A1(n5113), .A2(n4272), .ZN(n8862) );
  NAND2_X1 U5851 ( .A1(n8888), .A2(n8347), .ZN(n5113) );
  INV_X1 U5852 ( .A(n5057), .ZN(n8865) );
  AOI21_X1 U5853 ( .B1(n8911), .B2(n4256), .A(n6480), .ZN(n5057) );
  NAND2_X1 U5854 ( .A1(n7534), .A2(n6249), .ZN(n6282) );
  NAND2_X1 U5855 ( .A1(n8938), .A2(n8345), .ZN(n8925) );
  NOR2_X1 U5856 ( .A1(n8926), .A2(n5087), .ZN(n5083) );
  NAND2_X1 U5857 ( .A1(n4443), .A2(n4445), .ZN(n8929) );
  NAND2_X1 U5858 ( .A1(n5066), .A2(n5067), .ZN(n8010) );
  NAND2_X1 U5859 ( .A1(n9996), .A2(n9985), .ZN(n8948) );
  AOI21_X1 U5860 ( .B1(n7865), .B2(n6607), .A(n5071), .ZN(n7946) );
  NAND2_X1 U5861 ( .A1(n5081), .A2(n7873), .ZN(n7954) );
  NAND2_X1 U5862 ( .A1(n5073), .A2(n6583), .ZN(n7334) );
  INV_X1 U5863 ( .A(n8890), .ZN(n8965) );
  AND2_X1 U5864 ( .A1(n8969), .A2(n9091), .ZN(n8944) );
  AND2_X1 U5865 ( .A1(n8985), .A2(n8984), .ZN(n4351) );
  NAND2_X1 U5866 ( .A1(n8995), .A2(n4784), .ZN(n9100) );
  INV_X1 U5867 ( .A(n4785), .ZN(n4784) );
  AND2_X1 U5868 ( .A1(n6534), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10007) );
  INV_X1 U5869 ( .A(n10001), .ZN(n10004) );
  INV_X1 U5870 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U5871 ( .A1(n9121), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4505) );
  AOI21_X1 U5872 ( .B1(n4792), .B2(n4791), .A(n9120), .ZN(n4659) );
  XNOR2_X1 U5873 ( .A(n6418), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8049) );
  AND2_X1 U5874 ( .A1(n5956), .A2(n5948), .ZN(n4731) );
  INV_X1 U5875 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8038) );
  INV_X1 U5876 ( .A(n6432), .ZN(n8037) );
  XNOR2_X1 U5877 ( .A(n6415), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7931) );
  INV_X1 U5878 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10107) );
  INV_X1 U5879 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7942) );
  INV_X1 U5880 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U5881 ( .A(n5963), .B(n5962), .ZN(n7806) );
  INV_X1 U5882 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5883 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5966) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7535) );
  INV_X1 U5885 ( .A(n4902), .ZN(n4900) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7207) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10108) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10064) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6830) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10105) );
  INV_X1 U5891 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6746) );
  INV_X1 U5892 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U5893 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4774) );
  NOR2_X1 U5894 ( .A1(n5898), .A2(n6703), .ZN(n6763) );
  AND4_X1 U5895 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n7611)
         );
  NAND2_X1 U5896 ( .A1(n4586), .A2(n4584), .ZN(n5934) );
  NAND2_X1 U5897 ( .A1(n4585), .A2(n4587), .ZN(n4584) );
  INV_X1 U5898 ( .A(n4588), .ZN(n4585) );
  AND4_X1 U5899 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n7495)
         );
  NAND2_X1 U5900 ( .A1(n4944), .A2(n5350), .ZN(n7492) );
  OR2_X1 U5901 ( .A1(n7459), .A2(n5351), .ZN(n4944) );
  NAND2_X1 U5902 ( .A1(n9227), .A2(n5686), .ZN(n9175) );
  INV_X1 U5903 ( .A(n9282), .ZN(n9272) );
  NAND2_X1 U5904 ( .A1(n7795), .A2(n4598), .ZN(n4593) );
  INV_X1 U5905 ( .A(n4954), .ZN(n4950) );
  AND3_X1 U5906 ( .A1(n5573), .A2(n5572), .A3(n5571), .ZN(n9558) );
  NAND2_X1 U5907 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  AND2_X1 U5908 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  AND4_X1 U5909 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n7777)
         );
  NAND2_X1 U5910 ( .A1(n7765), .A2(n7766), .ZN(n7764) );
  NAND2_X1 U5911 ( .A1(n4941), .A2(n4942), .ZN(n7765) );
  INV_X1 U5912 ( .A(n9275), .ZN(n9284) );
  INV_X1 U5913 ( .A(n9296), .ZN(n9598) );
  OAI211_X1 U5914 ( .C1(n4596), .C2(n4594), .A(n4591), .B(n7960), .ZN(n9239)
         );
  NAND2_X1 U5915 ( .A1(n4592), .A2(n7795), .ZN(n4591) );
  NOR2_X1 U5916 ( .A1(n4595), .A2(n4594), .ZN(n4592) );
  INV_X1 U5917 ( .A(n7959), .ZN(n4594) );
  OAI21_X1 U5918 ( .B1(n7795), .B2(n7793), .A(n7792), .ZN(n7885) );
  NAND2_X1 U5919 ( .A1(n5332), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U5920 ( .A1(n7094), .A2(n7095), .ZN(n7093) );
  CLKBUF_X1 U5921 ( .A(n7458), .Z(n7459) );
  OR2_X1 U5922 ( .A1(n9382), .A2(n5848), .ZN(n5854) );
  XNOR2_X1 U5923 ( .A(n5556), .B(n5555), .ZN(n9281) );
  NAND2_X1 U5924 ( .A1(n4606), .A2(n4605), .ZN(n5187) );
  AOI21_X1 U5925 ( .B1(n4607), .B2(n4609), .A(n4609), .ZN(n4605) );
  NAND2_X1 U5926 ( .A1(n5826), .A2(n5825), .ZN(n9415) );
  INV_X1 U5927 ( .A(n9558), .ZN(n9522) );
  INV_X1 U5928 ( .A(n7495), .ZN(n9303) );
  INV_X1 U5929 ( .A(n9926), .ZN(n9304) );
  NAND4_X2 U5930 ( .A1(n5051), .A2(n5258), .A3(n5259), .A4(n5052), .ZN(n9307)
         );
  NAND2_X1 U5931 ( .A1(n5332), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5052) );
  INV_X1 U5932 ( .A(n4392), .ZN(n7066) );
  NAND2_X1 U5933 ( .A1(n4577), .A2(n4576), .ZN(n6812) );
  INV_X1 U5934 ( .A(n6777), .ZN(n4576) );
  INV_X1 U5935 ( .A(n6778), .ZN(n4577) );
  NAND2_X1 U5936 ( .A1(n6812), .A2(n6811), .ZN(n6858) );
  NAND2_X1 U5937 ( .A1(n6800), .A2(n4388), .ZN(n6851) );
  NAND2_X1 U5938 ( .A1(n4390), .A2(n4389), .ZN(n4388) );
  INV_X1 U5939 ( .A(n6810), .ZN(n4390) );
  NAND2_X1 U5940 ( .A1(n6854), .A2(n6813), .ZN(n4835) );
  NAND2_X1 U5941 ( .A1(n6777), .A2(n4574), .ZN(n4573) );
  AND2_X1 U5942 ( .A1(n4828), .A2(n4827), .ZN(n7101) );
  INV_X1 U5943 ( .A(n7019), .ZN(n4827) );
  INV_X1 U5944 ( .A(n4828), .ZN(n7020) );
  INV_X1 U5945 ( .A(n4562), .ZN(n7555) );
  AND2_X1 U5946 ( .A1(n4831), .A2(n4830), .ZN(n7978) );
  INV_X1 U5947 ( .A(n7557), .ZN(n4830) );
  INV_X1 U5948 ( .A(n4831), .ZN(n7558) );
  NAND2_X1 U5949 ( .A1(n7975), .A2(n7976), .ZN(n9310) );
  NAND2_X1 U5950 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  XNOR2_X1 U5951 ( .A(n9331), .B(n9333), .ZN(n9334) );
  INV_X1 U5952 ( .A(n4399), .ZN(n9855) );
  INV_X1 U5953 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5613) );
  INV_X1 U5954 ( .A(n8175), .ZN(n9619) );
  INV_X1 U5955 ( .A(n9354), .ZN(n9623) );
  AOI21_X1 U5956 ( .B1(n9624), .B2(n9485), .A(n8469), .ZN(n4690) );
  NAND2_X1 U5957 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  NAND2_X1 U5958 ( .A1(n9365), .A2(n9542), .ZN(n9367) );
  INV_X1 U5959 ( .A(n9634), .ZN(n9385) );
  NAND2_X1 U5960 ( .A1(n5036), .A2(n5038), .ZN(n9372) );
  NAND2_X1 U5961 ( .A1(n9407), .A2(n5039), .ZN(n5036) );
  NAND2_X1 U5962 ( .A1(n4666), .A2(n8458), .ZN(n9426) );
  NAND2_X1 U5963 ( .A1(n9441), .A2(n8457), .ZN(n4666) );
  NAND2_X1 U5964 ( .A1(n5033), .A2(n8422), .ZN(n9433) );
  NOR2_X1 U5965 ( .A1(n4978), .A2(n4979), .ZN(n4981) );
  INV_X1 U5966 ( .A(n8455), .ZN(n4978) );
  NAND2_X1 U5967 ( .A1(n4683), .A2(n4681), .ZN(n9479) );
  NAND2_X1 U5968 ( .A1(n5020), .A2(n5025), .ZN(n9474) );
  NAND2_X1 U5969 ( .A1(n9518), .A2(n5026), .ZN(n5020) );
  NAND2_X1 U5970 ( .A1(n4686), .A2(n8451), .ZN(n9495) );
  NAND2_X1 U5971 ( .A1(n5030), .A2(n5029), .ZN(n9516) );
  INV_X1 U5972 ( .A(n9518), .ZN(n5030) );
  OAI21_X1 U5973 ( .B1(n9563), .B2(n5047), .A(n5045), .ZN(n9527) );
  OAI21_X1 U5974 ( .B1(n9563), .B2(n8415), .A(n8416), .ZN(n9551) );
  NAND2_X1 U5975 ( .A1(n9582), .A2(n4983), .ZN(n9537) );
  NAND2_X1 U5976 ( .A1(n8411), .A2(n8410), .ZN(n9600) );
  NAND2_X1 U5977 ( .A1(n5035), .A2(n7724), .ZN(n7727) );
  NAND2_X1 U5978 ( .A1(n7717), .A2(n8086), .ZN(n7775) );
  NAND2_X1 U5979 ( .A1(n10221), .A2(n7315), .ZN(n9609) );
  OAI211_X2 U5980 ( .C1(n6779), .C2(n6788), .A(n5184), .B(n5183), .ZN(n7522)
         );
  OR2_X1 U5981 ( .A1(n8152), .A2(n6706), .ZN(n5183) );
  INV_X1 U5982 ( .A(n9571), .ZN(n9614) );
  INV_X1 U5983 ( .A(n9566), .ZN(n10213) );
  AND2_X2 U5984 ( .A1(n7191), .A2(n7190), .ZN(n9972) );
  INV_X1 U5985 ( .A(n9626), .ZN(n4581) );
  AND2_X2 U5986 ( .A1(n7191), .A2(n7311), .ZN(n9958) );
  AND2_X1 U5987 ( .A1(n5898), .A2(n5901), .ZN(n8327) );
  INV_X1 U5988 ( .A(n5145), .ZN(n8405) );
  NAND2_X1 U5989 ( .A1(n4618), .A2(n4616), .ZN(n5144) );
  NAND2_X1 U5990 ( .A1(n4617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4616) );
  CLKBUF_X1 U5991 ( .A(n5919), .Z(n8336) );
  INV_X1 U5992 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8051) );
  INV_X1 U5993 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8471) );
  OAI211_X1 U5994 ( .C1(n5165), .C2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_25__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  INV_X1 U5995 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7971) );
  AND2_X1 U5996 ( .A1(n4612), .A2(P1_U3084), .ZN(n7933) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7944) );
  INV_X1 U5998 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10151) );
  INV_X1 U5999 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7791) );
  INV_X1 U6000 ( .A(n7181), .ZN(n8287) );
  INV_X1 U6001 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8393) );
  INV_X1 U6002 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6832) );
  INV_X1 U6003 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6748) );
  INV_X1 U6004 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6737) );
  XNOR2_X1 U6005 ( .A(n5240), .B(n5239), .ZN(n6836) );
  OAI21_X1 U6006 ( .B1(n5174), .B2(n5173), .A(n5238), .ZN(n6788) );
  XNOR2_X1 U6007 ( .A(n4627), .B(n5220), .ZN(n6783) );
  NAND2_X1 U6008 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4627) );
  NAND2_X1 U6009 ( .A1(n4531), .A2(n10037), .ZN(n10239) );
  INV_X1 U6010 ( .A(n4534), .ZN(n10240) );
  AND2_X1 U6011 ( .A1(n9768), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n10228) );
  XNOR2_X1 U6012 ( .A(n9769), .B(n4524), .ZN(n10226) );
  XNOR2_X1 U6013 ( .A(n9772), .B(n4540), .ZN(n10238) );
  INV_X1 U6014 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4540) );
  XNOR2_X1 U6015 ( .A(n9774), .B(n4538), .ZN(n10237) );
  NOR2_X1 U6016 ( .A1(n9778), .A2(n10234), .ZN(n10062) );
  NOR2_X1 U6017 ( .A1(n10057), .A2(n4331), .ZN(n10056) );
  NAND2_X1 U6018 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  NAND2_X1 U6019 ( .A1(n10054), .A2(n4535), .ZN(n10052) );
  NAND2_X1 U6020 ( .A1(n4537), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U6021 ( .A1(n10052), .A2(n10053), .ZN(n10051) );
  OAI21_X1 U6022 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10051), .ZN(n10049) );
  OAI21_X1 U6023 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10048), .ZN(n10046) );
  OAI21_X1 U6024 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10045), .ZN(n10043) );
  NAND2_X1 U6025 ( .A1(n4893), .A2(n4321), .ZN(P2_U3222) );
  OAI211_X1 U6026 ( .C1(n4898), .C2(n4897), .A(n4895), .B(n4894), .ZN(n4893)
         );
  OAI211_X1 U6027 ( .C1(n4629), .C2(n4318), .A(n4366), .B(n4364), .ZN(P2_U3227) );
  NOR2_X1 U6028 ( .A1(n8528), .A2(n4365), .ZN(n4364) );
  NAND2_X1 U6029 ( .A1(n4629), .A2(n8527), .ZN(n4366) );
  NAND2_X1 U6030 ( .A1(n7136), .A2(n4761), .ZN(n7081) );
  INV_X1 U6031 ( .A(n4766), .ZN(n7690) );
  AND2_X1 U6032 ( .A1(n4773), .A2(n8701), .ZN(n4772) );
  NAND2_X1 U6033 ( .A1(n4657), .A2(n4656), .ZN(P2_U3549) );
  OR2_X1 U6034 ( .A1(n4333), .A2(n6463), .ZN(n4656) );
  NAND2_X1 U6035 ( .A1(n4350), .A2(n4333), .ZN(n4657) );
  OAI21_X1 U6036 ( .B1(n8986), .B2(n4658), .A(n4351), .ZN(n4350) );
  OAI211_X1 U6037 ( .C1(n8985), .C2(n4455), .A(n4453), .B(n4451), .ZN(P2_U3517) );
  INV_X1 U6038 ( .A(n4452), .ZN(n4451) );
  OAI21_X1 U6039 ( .B1(n8984), .B2(n4455), .A(n4317), .ZN(n4452) );
  OAI21_X1 U6040 ( .B1(n9412), .B2(n9235), .A(n9195), .ZN(n4631) );
  AOI21_X1 U6041 ( .B1(n9190), .B2(n9189), .A(n9278), .ZN(n4632) );
  INV_X1 U6042 ( .A(n9348), .ZN(n4639) );
  NAND2_X1 U6043 ( .A1(n9345), .A2(n9468), .ZN(n4640) );
  NAND2_X1 U6044 ( .A1(n4691), .A2(n4688), .ZN(P1_U3355) );
  NAND2_X1 U6045 ( .A1(n4692), .A2(n10221), .ZN(n4691) );
  INV_X1 U6046 ( .A(n4689), .ZN(n4688) );
  OAI21_X1 U6047 ( .B1(n9627), .B2(n9595), .A(n4690), .ZN(n4689) );
  OAI21_X1 U6048 ( .B1(n9631), .B2(n10210), .A(n4370), .ZN(P1_U3263) );
  AOI21_X1 U6049 ( .B1(n9629), .B2(n9614), .A(n4371), .ZN(n4370) );
  OAI21_X1 U6050 ( .B1(n9632), .B2(n9595), .A(n4372), .ZN(n4371) );
  INV_X1 U6051 ( .A(n9370), .ZN(n4372) );
  NAND2_X1 U6052 ( .A1(n4520), .A2(n10230), .ZN(n9783) );
  OAI21_X1 U6053 ( .B1(n10231), .B2(n10232), .A(n9863), .ZN(n4520) );
  OR2_X1 U6054 ( .A1(n8992), .A2(n8351), .ZN(n6485) );
  AND4_X1 U6055 ( .A1(n8752), .A2(n4439), .A3(n8734), .A4(n8796), .ZN(n4241)
         );
  AND2_X1 U6056 ( .A1(n7686), .A2(n7872), .ZN(n4243) );
  INV_X1 U6057 ( .A(n5252), .ZN(n5478) );
  INV_X1 U6058 ( .A(n4237), .ZN(n6239) );
  OAI21_X1 U6059 ( .B1(n4678), .B2(n9371), .A(n8463), .ZN(n4677) );
  NAND2_X1 U6060 ( .A1(n8888), .A2(n5110), .ZN(n5108) );
  OR2_X1 U6061 ( .A1(n5400), .A2(n5399), .ZN(n4625) );
  AND2_X1 U6062 ( .A1(n6619), .A2(n6618), .ZN(n4244) );
  NAND2_X1 U6063 ( .A1(n8033), .A2(n8041), .ZN(n4245) );
  AND2_X1 U6064 ( .A1(n8434), .A2(n8435), .ZN(n8205) );
  NAND2_X1 U6065 ( .A1(n9652), .A2(n9444), .ZN(n4246) );
  INV_X1 U6066 ( .A(n4676), .ZN(n4675) );
  OAI21_X1 U6067 ( .B1(n4679), .B2(n4677), .A(n8465), .ZN(n4676) );
  INV_X1 U6068 ( .A(n7446), .ZN(n4382) );
  OR2_X1 U6069 ( .A1(n9672), .A2(n9496), .ZN(n4247) );
  NAND2_X1 U6070 ( .A1(n5387), .A2(n5386), .ZN(n9720) );
  AND2_X1 U6071 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n4248) );
  NAND2_X1 U6072 ( .A1(n6253), .A2(n6252), .ZN(n9045) );
  INV_X1 U6073 ( .A(n9414), .ZN(n5040) );
  NAND2_X1 U6074 ( .A1(n8452), .A2(n8447), .ZN(n4249) );
  AND4_X1 U6075 ( .A1(n7634), .A2(n6472), .A3(n7701), .A4(n6544), .ZN(n4250)
         );
  INV_X1 U6076 ( .A(n9705), .ZN(n9584) );
  INV_X1 U6077 ( .A(n5095), .ZN(n5094) );
  OAI21_X1 U6078 ( .B1(n8734), .B2(n5096), .A(n5097), .ZN(n5095) );
  NAND2_X1 U6079 ( .A1(n6282), .A2(n6281), .ZN(n9034) );
  NAND2_X1 U6080 ( .A1(n8186), .A2(n8187), .ZN(n4251) );
  NAND2_X1 U6081 ( .A1(n5952), .A2(n5951), .ZN(n9007) );
  AND2_X1 U6082 ( .A1(n8262), .A2(n8441), .ZN(n4983) );
  AND3_X1 U6083 ( .A1(n4494), .A2(n5948), .A3(n5973), .ZN(n4252) );
  NOR2_X1 U6084 ( .A1(n9676), .A2(n9508), .ZN(n4253) );
  INV_X1 U6085 ( .A(n9628), .ZN(n4998) );
  OR2_X1 U6086 ( .A1(n6481), .A2(n6640), .ZN(n4254) );
  AND2_X1 U6087 ( .A1(n6485), .A2(n6669), .ZN(n8737) );
  NAND2_X1 U6088 ( .A1(n5599), .A2(n5598), .ZN(n9543) );
  OR2_X1 U6089 ( .A1(n9061), .A2(n8933), .ZN(n6621) );
  XNOR2_X1 U6090 ( .A(n5966), .B(n5965), .ZN(n5984) );
  AND2_X1 U6091 ( .A1(n9206), .A2(n5606), .ZN(n4255) );
  AND2_X1 U6092 ( .A1(n6631), .A2(n5062), .ZN(n4256) );
  AND2_X1 U6093 ( .A1(n4760), .A2(n4759), .ZN(n4257) );
  AND2_X1 U6094 ( .A1(n6088), .A2(n6087), .ZN(n7580) );
  NAND2_X1 U6095 ( .A1(n5152), .A2(n4551), .ZN(n4258) );
  AND2_X1 U6096 ( .A1(n4244), .A2(n4470), .ZN(n4259) );
  XNOR2_X1 U6097 ( .A(n4506), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6098 ( .A1(n8405), .A2(n9753), .ZN(n5368) );
  INV_X1 U6099 ( .A(n5368), .ZN(n5332) );
  AND2_X1 U6100 ( .A1(n8813), .A2(n4842), .ZN(n4260) );
  AND2_X1 U6101 ( .A1(n7010), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4261) );
  OR2_X1 U6102 ( .A1(n6323), .A2(n8582), .ZN(n4262) );
  INV_X1 U6103 ( .A(n4890), .ZN(n4889) );
  NAND2_X1 U6104 ( .A1(n4891), .A2(n6243), .ZN(n4890) );
  AND2_X1 U6105 ( .A1(n9034), .A2(n8846), .ZN(n4263) );
  AND2_X1 U6106 ( .A1(n4953), .A2(n4950), .ZN(n4264) );
  OAI21_X1 U6107 ( .B1(n4683), .B2(n4381), .A(n4379), .ZN(n9463) );
  OR2_X1 U6108 ( .A1(n8418), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U6109 ( .A1(n9189), .A2(n5806), .ZN(n9267) );
  INV_X1 U6110 ( .A(n8844), .ZN(n5107) );
  NOR2_X1 U6111 ( .A1(n9652), .A2(n9444), .ZN(n4265) );
  AND2_X1 U6112 ( .A1(n4590), .A2(n9269), .ZN(n4266) );
  AND2_X1 U6113 ( .A1(n8939), .A2(n5088), .ZN(n4267) );
  OR2_X1 U6114 ( .A1(n9019), .A2(n8512), .ZN(n4268) );
  INV_X1 U6115 ( .A(n8453), .ZN(n4800) );
  INV_X1 U6116 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n10120) );
  NAND2_X1 U6117 ( .A1(n6266), .A2(n6265), .ZN(n9039) );
  INV_X1 U6118 ( .A(n9039), .ZN(n4846) );
  OR2_X1 U6119 ( .A1(n8698), .A2(n8697), .ZN(n4269) );
  INV_X2 U6120 ( .A(n6910), .ZN(n5994) );
  INV_X1 U6121 ( .A(n8360), .ZN(n4439) );
  NAND2_X1 U6122 ( .A1(n4500), .A2(n4498), .ZN(n8544) );
  XOR2_X1 U6123 ( .A(n5878), .B(n5877), .Z(n4270) );
  XNOR2_X1 U6125 ( .A(n9012), .B(n8645), .ZN(n8796) );
  AND2_X1 U6126 ( .A1(n8741), .A2(n4852), .ZN(n4271) );
  NAND2_X1 U6127 ( .A1(n4846), .A2(n8546), .ZN(n4272) );
  NAND2_X1 U6128 ( .A1(n9687), .A2(n9543), .ZN(n4273) );
  NAND2_X1 U6129 ( .A1(n5378), .A2(n7489), .ZN(n4274) );
  OR2_X1 U6130 ( .A1(n8391), .A2(n8659), .ZN(n4275) );
  INV_X1 U6131 ( .A(n6606), .ZN(n4778) );
  AND3_X1 U6132 ( .A1(n6029), .A2(n6026), .A3(n6028), .ZN(n4276) );
  NAND2_X1 U6133 ( .A1(n9174), .A2(n4961), .ZN(n9246) );
  INV_X1 U6134 ( .A(n8086), .ZN(n4975) );
  AND2_X1 U6135 ( .A1(n7634), .A2(n6593), .ZN(n4277) );
  AND2_X1 U6136 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4851), .ZN(n4278) );
  OR2_X1 U6137 ( .A1(n9039), .A2(n8546), .ZN(n6631) );
  INV_X1 U6138 ( .A(n8331), .ZN(n5903) );
  XNOR2_X1 U6139 ( .A(n5187), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8331) );
  OR2_X1 U6140 ( .A1(n4733), .A2(n6675), .ZN(n4279) );
  NAND2_X1 U6141 ( .A1(n6503), .A2(n6502), .ZN(n8978) );
  AND2_X1 U6142 ( .A1(n6136), .A2(n6117), .ZN(n4280) );
  AND2_X1 U6143 ( .A1(n9693), .A2(n9522), .ZN(n4281) );
  INV_X1 U6144 ( .A(n9569), .ZN(n9698) );
  INV_X1 U6145 ( .A(n5803), .ZN(n4948) );
  OR2_X1 U6146 ( .A1(n9646), .A2(n8425), .ZN(n8461) );
  INV_X1 U6147 ( .A(n8461), .ZN(n4810) );
  AND2_X1 U6148 ( .A1(n8465), .A2(n8140), .ZN(n4282) );
  INV_X1 U6149 ( .A(n6615), .ZN(n4473) );
  AND2_X1 U6150 ( .A1(n5085), .A2(n5084), .ZN(n4283) );
  OR2_X1 U6151 ( .A1(n9007), .A2(n8557), .ZN(n6656) );
  OR2_X1 U6152 ( .A1(n4738), .A2(n8360), .ZN(n4284) );
  INV_X1 U6153 ( .A(n8456), .ZN(n4980) );
  AND2_X1 U6154 ( .A1(n8847), .A2(n6331), .ZN(n4285) );
  AND2_X1 U6155 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n4286) );
  INV_X1 U6156 ( .A(n5011), .ZN(n9434) );
  NOR2_X1 U6157 ( .A1(n9475), .A2(n5012), .ZN(n5011) );
  INV_X1 U6158 ( .A(n8427), .ZN(n5041) );
  AND2_X1 U6159 ( .A1(n4883), .A2(n6334), .ZN(n4882) );
  INV_X1 U6160 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4903) );
  NOR2_X1 U6161 ( .A1(n9380), .A2(n9628), .ZN(n4287) );
  INV_X1 U6162 ( .A(n4762), .ZN(n4761) );
  NOR2_X1 U6163 ( .A1(n7133), .A2(n7673), .ZN(n4762) );
  INV_X1 U6164 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4609) );
  AND2_X1 U6165 ( .A1(n5039), .A2(n9371), .ZN(n4288) );
  INV_X1 U6166 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6807) );
  AND2_X1 U6167 ( .A1(n9656), .A2(n9456), .ZN(n4289) );
  NOR2_X1 U6168 ( .A1(n8855), .A2(n8513), .ZN(n5114) );
  INV_X1 U6169 ( .A(n4726), .ZN(n4725) );
  OR2_X1 U6170 ( .A1(n8523), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U6171 ( .A1(n8998), .A2(n8733), .ZN(n4290) );
  INV_X1 U6172 ( .A(n4845), .ZN(n4844) );
  NAND2_X1 U6173 ( .A1(n4847), .A2(n4846), .ZN(n4845) );
  AND2_X1 U6174 ( .A1(n5635), .A2(SI_18_), .ZN(n4291) );
  INV_X1 U6175 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5958) );
  AND2_X1 U6176 ( .A1(n8577), .A2(n8579), .ZN(n4292) );
  AND2_X1 U6177 ( .A1(n6102), .A2(n6101), .ZN(n4293) );
  AND2_X1 U6178 ( .A1(n5164), .A2(n4609), .ZN(n4294) );
  INV_X1 U6179 ( .A(n9517), .ZN(n5029) );
  AND2_X1 U6180 ( .A1(n8187), .A2(n8447), .ZN(n9517) );
  NAND2_X1 U6181 ( .A1(n9385), .A2(n9294), .ZN(n4295) );
  AND2_X1 U6182 ( .A1(n7490), .A2(n5377), .ZN(n4296) );
  NOR2_X1 U6183 ( .A1(n8801), .A2(n8810), .ZN(n4297) );
  OR2_X1 U6184 ( .A1(n9628), .A2(n9376), .ZN(n8464) );
  NAND2_X1 U6185 ( .A1(n8428), .A2(n8426), .ZN(n4298) );
  INV_X1 U6186 ( .A(n4623), .ZN(n7766) );
  NAND2_X1 U6187 ( .A1(n4625), .A2(n4624), .ZN(n4623) );
  AND3_X1 U6188 ( .A1(n5989), .A2(n5988), .A3(n5121), .ZN(n7244) );
  AND3_X1 U6189 ( .A1(n4494), .A2(n5940), .A3(n10120), .ZN(n4299) );
  AND2_X1 U6190 ( .A1(n5760), .A2(n5781), .ZN(n4300) );
  NOR2_X1 U6191 ( .A1(n9709), .A2(n9297), .ZN(n4301) );
  INV_X1 U6192 ( .A(n8466), .ZN(n4986) );
  AND2_X1 U6193 ( .A1(n4901), .A2(n4837), .ZN(n4302) );
  AND2_X1 U6194 ( .A1(n7313), .A2(n5196), .ZN(n4303) );
  AND2_X1 U6195 ( .A1(n6600), .A2(n6604), .ZN(n7682) );
  AND2_X1 U6196 ( .A1(n7684), .A2(n7952), .ZN(n4304) );
  INV_X1 U6197 ( .A(n9909), .ZN(n7414) );
  AND2_X1 U6198 ( .A1(n5049), .A2(n5272), .ZN(n9909) );
  INV_X1 U6199 ( .A(n9918), .ZN(n4818) );
  INV_X1 U6200 ( .A(n6633), .ZN(n5061) );
  AND2_X1 U6201 ( .A1(n6628), .A2(n8878), .ZN(n8926) );
  AND2_X1 U6202 ( .A1(n4445), .A2(n6475), .ZN(n4305) );
  AND2_X1 U6203 ( .A1(n4853), .A2(n8745), .ZN(n4306) );
  AND2_X1 U6204 ( .A1(n9427), .A2(n8457), .ZN(n4307) );
  INV_X1 U6205 ( .A(n9494), .ZN(n4685) );
  AND2_X1 U6206 ( .A1(n8186), .A2(n8452), .ZN(n9494) );
  INV_X1 U6207 ( .A(n8717), .ZN(n8714) );
  AND2_X1 U6208 ( .A1(n6677), .A2(n6673), .ZN(n8717) );
  AND2_X1 U6209 ( .A1(n4248), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n4308) );
  AND2_X1 U6210 ( .A1(n4254), .A2(n4268), .ZN(n4309) );
  OR2_X1 U6211 ( .A1(n5454), .A2(n5453), .ZN(n4310) );
  AND2_X1 U6212 ( .A1(n4266), .A2(n4587), .ZN(n4311) );
  AND2_X1 U6213 ( .A1(n4580), .A2(n4579), .ZN(n4312) );
  INV_X1 U6214 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4551) );
  INV_X1 U6215 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4617) );
  INV_X1 U6216 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9120) );
  AND2_X1 U6217 ( .A1(n5170), .A2(n5171), .ZN(n5140) );
  NAND2_X1 U6218 ( .A1(n4573), .A2(n4835), .ZN(n4313) );
  OR2_X1 U6219 ( .A1(n4632), .A2(n4631), .ZN(P1_U3223) );
  OR2_X1 U6220 ( .A1(n7306), .A2(n7305), .ZN(n4315) );
  AND2_X1 U6221 ( .A1(n6395), .A2(n6394), .ZN(n8729) );
  INV_X1 U6222 ( .A(n8729), .ZN(n4855) );
  AND2_X1 U6223 ( .A1(n5983), .A2(n5982), .ZN(n8557) );
  INV_X1 U6224 ( .A(n8557), .ZN(n5099) );
  AND2_X1 U6225 ( .A1(n8942), .A2(n4844), .ZN(n4316) );
  NAND2_X1 U6226 ( .A1(n5082), .A2(n7684), .ZN(n7874) );
  NAND2_X1 U6227 ( .A1(n5763), .A2(n5762), .ZN(n9652) );
  INV_X1 U6228 ( .A(n9652), .ZN(n4698) );
  NAND2_X1 U6229 ( .A1(n7747), .A2(n7748), .ZN(n7294) );
  OR2_X1 U6230 ( .A1(n10030), .A2(n4456), .ZN(n4317) );
  OR3_X1 U6231 ( .A1(n4723), .A2(n8523), .A3(n8627), .ZN(n4318) );
  NAND2_X1 U6232 ( .A1(n4593), .A2(n4596), .ZN(n7961) );
  INV_X1 U6233 ( .A(n7953), .ZN(n5080) );
  INV_X1 U6234 ( .A(n8526), .ZN(n4723) );
  INV_X1 U6235 ( .A(n8234), .ZN(n4815) );
  INV_X1 U6236 ( .A(n8889), .ZN(n4437) );
  NAND2_X1 U6237 ( .A1(n4792), .A2(n4900), .ZN(n4319) );
  AOI21_X1 U6238 ( .B1(n4614), .B2(n7446), .A(n4613), .ZN(n7422) );
  INV_X1 U6239 ( .A(n6550), .ZN(n6441) );
  NAND2_X1 U6240 ( .A1(n4958), .A2(n4956), .ZN(n9141) );
  NAND2_X1 U6241 ( .A1(n6473), .A2(n6604), .ZN(n7668) );
  AND2_X1 U6242 ( .A1(n5077), .A2(n5078), .ZN(n4320) );
  NOR2_X1 U6243 ( .A1(n6466), .A2(n6467), .ZN(n4321) );
  NAND2_X1 U6244 ( .A1(n7641), .A2(n4856), .ZN(n4859) );
  AOI22_X1 U6245 ( .A1(n9293), .A2(n9540), .B1(n9351), .B2(n9291), .ZN(n8468)
         );
  NAND2_X1 U6246 ( .A1(n6393), .A2(n6392), .ZN(n4322) );
  INV_X1 U6247 ( .A(n4886), .ZN(n8482) );
  AND2_X1 U6248 ( .A1(n8039), .A2(n8040), .ZN(n4886) );
  AND2_X1 U6249 ( .A1(n5083), .A2(n8938), .ZN(n4323) );
  NAND2_X1 U6250 ( .A1(n7018), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4324) );
  NAND2_X1 U6251 ( .A1(n7556), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4325) );
  INV_X1 U6252 ( .A(n5027), .ZN(n5026) );
  NOR2_X1 U6253 ( .A1(n5065), .A2(n4778), .ZN(n4326) );
  NAND2_X1 U6254 ( .A1(n8733), .A2(n8912), .ZN(n4327) );
  NAND2_X1 U6255 ( .A1(n8365), .A2(n8364), .ZN(n4328) );
  NAND2_X1 U6256 ( .A1(n5067), .A2(n6619), .ZN(n5065) );
  INV_X1 U6257 ( .A(n5065), .ZN(n4448) );
  AND2_X1 U6258 ( .A1(n4700), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n4329) );
  NAND2_X1 U6259 ( .A1(n5941), .A2(n5940), .ZN(n6408) );
  INV_X1 U6260 ( .A(n4650), .ZN(n4649) );
  NAND2_X1 U6261 ( .A1(n8355), .A2(n8512), .ZN(n4650) );
  INV_X1 U6262 ( .A(n5760), .ZN(n4611) );
  INV_X1 U6263 ( .A(n10030), .ZN(n4455) );
  INV_X1 U6264 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U6265 ( .A1(n5592), .A2(n5591), .ZN(n9687) );
  INV_X1 U6266 ( .A(n9687), .ZN(n5004) );
  AND2_X1 U6267 ( .A1(n8667), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4330) );
  INV_X1 U6268 ( .A(n7893), .ZN(n4992) );
  INV_X1 U6269 ( .A(n9693), .ZN(n5007) );
  INV_X1 U6270 ( .A(n7792), .ZN(n4599) );
  INV_X1 U6271 ( .A(n9667), .ZN(n5015) );
  OR2_X1 U6272 ( .A1(n7378), .A2(n7181), .ZN(n9949) );
  INV_X1 U6273 ( .A(n9949), .ZN(n4997) );
  NAND3_X1 U6274 ( .A1(n4252), .A2(n4730), .A3(n4729), .ZN(n6455) );
  NAND2_X1 U6275 ( .A1(n6877), .A2(n6876), .ZN(n6875) );
  INV_X1 U6276 ( .A(n8246), .ZN(n4383) );
  INV_X1 U6277 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n4704) );
  INV_X1 U6278 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n4705) );
  OR2_X1 U6279 ( .A1(n5227), .A2(n5228), .ZN(n4401) );
  AOI21_X1 U6280 ( .B1(n6988), .B2(n4757), .A(n4261), .ZN(n4756) );
  INV_X1 U6281 ( .A(n9468), .ZN(n10220) );
  AND2_X1 U6282 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4331) );
  AND2_X1 U6283 ( .A1(n6841), .A2(n6769), .ZN(n4332) );
  INV_X1 U6284 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n4526) );
  INV_X1 U6285 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n4621) );
  INV_X1 U6286 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4524) );
  INV_X1 U6287 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n4522) );
  INV_X1 U6288 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n4537) );
  INV_X1 U6289 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n4389) );
  INV_X1 U6290 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4538) );
  INV_X1 U6291 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U6292 ( .B1(n8996), .B2(n9081), .A(n8994), .ZN(n4785) );
  INV_X2 U6293 ( .A(n4315), .ZN(n4333) );
  OR2_X1 U6294 ( .A1(n8702), .A2(n4334), .ZN(n4773) );
  NAND2_X1 U6295 ( .A1(n4335), .A2(n5434), .ZN(n5461) );
  NAND2_X1 U6296 ( .A1(n5271), .A2(n4338), .ZN(n4337) );
  INV_X1 U6297 ( .A(n5281), .ZN(n4338) );
  NAND2_X1 U6298 ( .A1(n5269), .A2(n5268), .ZN(n5271) );
  NAND2_X1 U6299 ( .A1(n4339), .A2(n5405), .ZN(n4905) );
  NAND2_X1 U6300 ( .A1(n4342), .A2(n5311), .ZN(n4341) );
  INV_X1 U6301 ( .A(n4459), .ZN(n4342) );
  NAND2_X1 U6302 ( .A1(n4459), .A2(n5309), .ZN(n4556) );
  INV_X1 U6303 ( .A(n5353), .ZN(n5352) );
  INV_X1 U6304 ( .A(SI_7_), .ZN(n4344) );
  NAND2_X1 U6305 ( .A1(n4346), .A2(n4909), .ZN(n5586) );
  INV_X1 U6306 ( .A(n4909), .ZN(n4348) );
  NAND2_X1 U6307 ( .A1(n6485), .A2(n4353), .ZN(n4352) );
  INV_X1 U6308 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U6309 ( .A1(n5960), .A2(n4363), .ZN(n5964) );
  XNOR2_X1 U6310 ( .A(n6077), .B(n8962), .ZN(n4864) );
  NAND3_X1 U6311 ( .A1(n7240), .A2(n7806), .A3(n10009), .ZN(n4368) );
  NAND3_X1 U6312 ( .A1(n5138), .A2(n5139), .A3(n5328), .ZN(n4369) );
  NAND4_X1 U6313 ( .A1(n5138), .A2(n5139), .A3(n5328), .A4(n5140), .ZN(n5142)
         );
  INV_X1 U6314 ( .A(n8083), .ZN(n4386) );
  NAND2_X1 U6315 ( .A1(n7438), .A2(n8083), .ZN(n7540) );
  NAND2_X1 U6316 ( .A1(n7436), .A2(n4387), .ZN(n7438) );
  NOR2_X2 U6317 ( .A1(n6865), .A2(n6862), .ZN(n7094) );
  AND2_X1 U6318 ( .A1(n4401), .A2(n4400), .ZN(n6865) );
  AND3_X1 U6319 ( .A1(n4402), .A2(n5206), .A3(n5205), .ZN(n6877) );
  NAND2_X1 U6320 ( .A1(n4405), .A2(n4406), .ZN(n6882) );
  NAND2_X1 U6321 ( .A1(n9807), .A2(n6789), .ZN(n6834) );
  NAND2_X2 U6322 ( .A1(n4408), .A2(n4407), .ZN(n7795) );
  NAND3_X1 U6323 ( .A1(n4941), .A2(n4625), .A3(n4942), .ZN(n4408) );
  NAND2_X1 U6324 ( .A1(n4555), .A2(n5151), .ZN(n4553) );
  INV_X1 U6325 ( .A(n5154), .ZN(n5156) );
  XNOR2_X1 U6326 ( .A(n4409), .B(n5186), .ZN(n5902) );
  OAI21_X1 U6327 ( .B1(n5154), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4409) );
  NAND3_X1 U6328 ( .A1(n4413), .A2(n4772), .A3(n4410), .ZN(P2_U3264) );
  NAND2_X1 U6329 ( .A1(n4411), .A2(n4769), .ZN(n4410) );
  NAND2_X1 U6330 ( .A1(n4412), .A2(n4770), .ZN(n4411) );
  NAND2_X1 U6331 ( .A1(n4415), .A2(n9974), .ZN(n4412) );
  NAND2_X1 U6332 ( .A1(n4414), .A2(n6532), .ZN(n4413) );
  OAI22_X1 U6333 ( .A1(n4415), .A2(n9976), .B1(n9978), .B2(n8700), .ZN(n4414)
         );
  NAND3_X1 U6334 ( .A1(n6018), .A2(n6017), .A3(n4426), .ZN(n6052) );
  NAND2_X1 U6335 ( .A1(n4427), .A2(n6053), .ZN(n6071) );
  NOR2_X1 U6336 ( .A1(n6408), .A2(n5975), .ZN(n4791) );
  NAND2_X1 U6337 ( .A1(n4428), .A2(n4299), .ZN(n9121) );
  INV_X1 U6338 ( .A(n5975), .ZN(n4429) );
  INV_X1 U6339 ( .A(n4792), .ZN(n6221) );
  NAND3_X1 U6340 ( .A1(n8926), .A2(n4430), .A3(n8844), .ZN(n6545) );
  NAND4_X1 U6341 ( .A1(n4437), .A2(n4433), .A3(n4432), .A4(n6619), .ZN(n4431)
         );
  NAND3_X1 U6342 ( .A1(n7682), .A2(n4436), .A3(n4250), .ZN(n4435) );
  NAND3_X1 U6343 ( .A1(n4242), .A2(n6548), .A3(n6547), .ZN(n4438) );
  NAND2_X1 U6344 ( .A1(n4777), .A2(n4447), .ZN(n4440) );
  AND2_X2 U6345 ( .A1(n4443), .A2(n4305), .ZN(n8911) );
  AND2_X2 U6346 ( .A1(n8795), .A2(n4449), .ZN(n8776) );
  OAI21_X1 U6347 ( .B1(n7254), .B2(n7253), .A(n6574), .ZN(n7237) );
  XNOR2_X2 U6348 ( .A(n4505), .B(n4458), .ZN(n8407) );
  XNOR2_X1 U6349 ( .A(n4459), .B(n5326), .ZN(n6711) );
  NAND2_X2 U6350 ( .A1(n5308), .A2(n5307), .ZN(n4459) );
  INV_X1 U6351 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4462) );
  NAND3_X1 U6352 ( .A1(n4462), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U6353 ( .A1(n4467), .A2(n4464), .ZN(n4471) );
  AOI21_X1 U6354 ( .B1(n4259), .B2(n4466), .A(n4465), .ZN(n4464) );
  NAND2_X1 U6355 ( .A1(n4777), .A2(n6622), .ZN(n4465) );
  NAND2_X1 U6356 ( .A1(n6611), .A2(n8339), .ZN(n4466) );
  NAND2_X1 U6357 ( .A1(n4469), .A2(n4468), .ZN(n4467) );
  NOR2_X1 U6358 ( .A1(n6612), .A2(n4472), .ZN(n4468) );
  INV_X1 U6359 ( .A(n6613), .ZN(n4469) );
  NAND2_X1 U6360 ( .A1(n4471), .A2(n4474), .ZN(n4752) );
  NAND2_X1 U6361 ( .A1(n4475), .A2(n6641), .ZN(n6634) );
  NAND2_X1 U6362 ( .A1(n4476), .A2(n5061), .ZN(n4475) );
  NAND2_X1 U6363 ( .A1(n6638), .A2(n4477), .ZN(n4476) );
  AND2_X1 U6364 ( .A1(n6632), .A2(n6631), .ZN(n4477) );
  NAND3_X1 U6365 ( .A1(n6635), .A2(n4268), .A3(n6640), .ZN(n4487) );
  AND2_X1 U6366 ( .A1(n4494), .A2(n5949), .ZN(n4732) );
  OAI21_X1 U6367 ( .B1(n4878), .B2(n4874), .A(n4872), .ZN(n7572) );
  INV_X1 U6368 ( .A(n8496), .ZN(n8497) );
  AOI21_X1 U6369 ( .B1(n7580), .B2(n4880), .A(n4871), .ZN(n4879) );
  INV_X1 U6370 ( .A(n7443), .ZN(n4614) );
  NAND2_X1 U6371 ( .A1(n9309), .A2(n5252), .ZN(n5225) );
  NAND2_X1 U6372 ( .A1(n5141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4506) );
  NAND4_X1 U6373 ( .A1(n5138), .A2(n5044), .A3(n5328), .A4(n5139), .ZN(n5141)
         );
  NAND2_X1 U6374 ( .A1(n8155), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5195) );
  AND2_X2 U6375 ( .A1(n5146), .A2(n8405), .ZN(n8155) );
  NAND2_X1 U6376 ( .A1(n4510), .A2(n4509), .ZN(n4507) );
  NAND3_X1 U6377 ( .A1(n5045), .A2(n5047), .A3(n4273), .ZN(n4513) );
  NAND2_X1 U6378 ( .A1(n9462), .A2(n9461), .ZN(n8420) );
  OAI21_X2 U6379 ( .B1(n9420), .B2(n4265), .A(n4246), .ZN(n4515) );
  NAND2_X1 U6380 ( .A1(n4531), .A2(n4529), .ZN(n4530) );
  NAND3_X1 U6381 ( .A1(n4530), .A2(n10242), .A3(n4533), .ZN(n9764) );
  NAND2_X1 U6382 ( .A1(n4532), .A2(n9763), .ZN(n10241) );
  NAND2_X1 U6383 ( .A1(n10239), .A2(n10240), .ZN(n4532) );
  NAND2_X1 U6384 ( .A1(n4534), .A2(n9763), .ZN(n4533) );
  OAI21_X1 U6385 ( .B1(n8114), .B2(n4795), .A(n4794), .ZN(n4542) );
  NAND2_X1 U6386 ( .A1(n8139), .A2(n4545), .ZN(n8141) );
  OAI21_X1 U6387 ( .B1(n8135), .B2(n4549), .A(n4546), .ZN(n4545) );
  INV_X2 U6388 ( .A(n8167), .ZN(n8163) );
  NOR2_X2 U6389 ( .A1(n9468), .A2(n8331), .ZN(n8167) );
  NAND3_X1 U6390 ( .A1(n4552), .A2(n4554), .A3(n4555), .ZN(n5361) );
  INV_X1 U6391 ( .A(n5260), .ZN(n4552) );
  NOR2_X1 U6392 ( .A1(n4553), .A2(n5260), .ZN(n5159) );
  NOR2_X2 U6393 ( .A1(n5260), .A2(n5137), .ZN(n5328) );
  NAND2_X1 U6394 ( .A1(n4558), .A2(n10220), .ZN(n4641) );
  NAND2_X1 U6395 ( .A1(n4559), .A2(n9342), .ZN(n4558) );
  NAND2_X1 U6396 ( .A1(n9344), .A2(n9330), .ZN(n4559) );
  NAND2_X1 U6397 ( .A1(n4928), .A2(n4567), .ZN(n4563) );
  NAND2_X1 U6398 ( .A1(n4928), .A2(n4927), .ZN(n4566) );
  OAI21_X2 U6399 ( .B1(n4928), .B2(n4569), .A(n4567), .ZN(n5510) );
  NAND2_X1 U6400 ( .A1(n4932), .A2(n4931), .ZN(n5754) );
  AOI21_X1 U6401 ( .B1(n5754), .B2(n5753), .A(n4611), .ZN(n5782) );
  AOI21_X1 U6402 ( .B1(n6778), .B2(n4574), .A(n4313), .ZN(n6855) );
  INV_X1 U6403 ( .A(n4580), .ZN(n9836) );
  NAND3_X1 U6404 ( .A1(n5725), .A2(n9247), .A3(n4266), .ZN(n4583) );
  NAND3_X1 U6405 ( .A1(n5725), .A2(n9247), .A3(n4311), .ZN(n4586) );
  NAND3_X1 U6406 ( .A1(n5725), .A2(n9247), .A3(n4948), .ZN(n4949) );
  NAND2_X1 U6407 ( .A1(n4600), .A2(n4601), .ZN(n5724) );
  NAND2_X1 U6408 ( .A1(n4933), .A2(n4603), .ZN(n4600) );
  NAND2_X1 U6409 ( .A1(n5156), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U6410 ( .A1(n7093), .A2(n5232), .ZN(n7165) );
  NAND2_X2 U6411 ( .A1(n9205), .A2(n9207), .ZN(n9206) );
  OR3_X1 U6412 ( .A1(n5907), .A2(n5934), .A3(n5906), .ZN(n5937) );
  NAND2_X1 U6413 ( .A1(n5724), .A2(n5723), .ZN(n9247) );
  NAND2_X1 U6414 ( .A1(n9239), .A2(n4960), .ZN(n4958) );
  NAND2_X1 U6415 ( .A1(n4921), .A2(n5807), .ZN(n5837) );
  NAND4_X1 U6416 ( .A1(n4610), .A2(n4748), .A3(n6700), .A4(n4747), .ZN(
        P2_U3244) );
  NAND2_X1 U6417 ( .A1(n6538), .A2(n6537), .ZN(n4610) );
  NAND2_X1 U6418 ( .A1(n5689), .A2(n5688), .ZN(n4932) );
  INV_X1 U6419 ( .A(n6484), .ZN(n5076) );
  AOI21_X1 U6420 ( .B1(n8205), .B2(n8410), .A(n4301), .ZN(n5043) );
  OAI21_X1 U6421 ( .B1(n9627), .B2(n9719), .A(n4635), .ZN(n5016) );
  NAND2_X1 U6422 ( .A1(n5143), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4618) );
  OAI22_X2 U6423 ( .A1(n9576), .A2(n8414), .B1(n9296), .B2(n9705), .ZN(n9563)
         );
  AND2_X2 U6424 ( .A1(n5169), .A2(n5196), .ZN(n5252) );
  INV_X1 U6425 ( .A(n4620), .ZN(n5417) );
  NAND2_X1 U6426 ( .A1(n4620), .A2(n5139), .ZN(n4619) );
  NAND3_X1 U6427 ( .A1(n4630), .A2(n5883), .A3(n5880), .ZN(n5196) );
  NAND2_X1 U6428 ( .A1(n4943), .A2(n4274), .ZN(n4942) );
  XOR2_X1 U6429 ( .A(n5872), .B(n5323), .Z(n7603) );
  NAND2_X1 U6430 ( .A1(n5130), .A2(n5129), .ZN(n5188) );
  XNOR2_X1 U6431 ( .A(n5226), .B(n5872), .ZN(n5228) );
  INV_X1 U6432 ( .A(n5879), .ZN(n4630) );
  NAND2_X1 U6433 ( .A1(n5166), .A2(n5167), .ZN(n5879) );
  NAND2_X1 U6434 ( .A1(n5204), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5201) );
  OAI22_X1 U6435 ( .A1(n6855), .A2(n6818), .B1(n6823), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n6814) );
  NAND3_X1 U6436 ( .A1(n4640), .A2(n4641), .A3(n4639), .ZN(P1_U3260) );
  NAND3_X1 U6437 ( .A1(n6351), .A2(n4728), .A3(n6350), .ZN(n4629) );
  NAND2_X1 U6438 ( .A1(n4868), .A2(n6153), .ZN(n7988) );
  INV_X1 U6439 ( .A(n5880), .ZN(n5896) );
  XNOR2_X1 U6440 ( .A(n5161), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5880) );
  AOI21_X1 U6441 ( .B1(n5350), .B2(n5351), .A(n4296), .ZN(n4940) );
  NAND2_X1 U6442 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5161) );
  NAND2_X2 U6443 ( .A1(n6775), .A2(n5919), .ZN(n5285) );
  NOR2_X1 U6444 ( .A1(n4696), .A2(n4695), .ZN(n8180) );
  AND2_X1 U6445 ( .A1(n7360), .A2(n7370), .ZN(n7412) );
  INV_X1 U6446 ( .A(n7374), .ZN(n9308) );
  XNOR2_X2 U6447 ( .A(n4636), .B(n5190), .ZN(n9468) );
  INV_X1 U6448 ( .A(n5348), .ZN(n5349) );
  NOR2_X1 U6449 ( .A1(n6814), .A2(n6815), .ZN(n7017) );
  AND2_X2 U6450 ( .A1(n4643), .A2(n4642), .ZN(n8789) );
  NAND3_X1 U6451 ( .A1(n5077), .A2(n5078), .A3(n5126), .ZN(n8344) );
  INV_X1 U6452 ( .A(n4320), .ZN(n4652) );
  NAND2_X1 U6453 ( .A1(n4320), .A2(n8339), .ZN(n7955) );
  NAND2_X1 U6454 ( .A1(n4660), .A2(n8252), .ZN(n7842) );
  NAND3_X1 U6455 ( .A1(n4662), .A2(n8200), .A3(n4661), .ZN(n4660) );
  NAND2_X1 U6456 ( .A1(n9441), .A2(n4307), .ZN(n4663) );
  INV_X1 U6457 ( .A(n9371), .ZN(n4680) );
  OAI211_X1 U6458 ( .C1(n4672), .C2(n9396), .A(n4669), .B(n4667), .ZN(n4985)
         );
  NAND2_X1 U6459 ( .A1(n9396), .A2(n4668), .ZN(n4667) );
  OAI21_X1 U6460 ( .B1(n4673), .B2(n8466), .A(n4670), .ZN(n4669) );
  NAND2_X1 U6461 ( .A1(n4673), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U6462 ( .A1(n4673), .A2(n4986), .ZN(n4672) );
  NAND2_X1 U6463 ( .A1(n9502), .A2(n8445), .ZN(n4686) );
  OAI21_X1 U6464 ( .B1(n8451), .B2(n4685), .A(n8452), .ZN(n4682) );
  NAND2_X1 U6465 ( .A1(n9502), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6466 ( .A1(n7316), .A2(n8192), .ZN(n7319) );
  NAND2_X1 U6467 ( .A1(n8243), .A2(n8190), .ZN(n7369) );
  NAND2_X1 U6468 ( .A1(n7319), .A2(n7180), .ZN(n8243) );
  NAND3_X1 U6469 ( .A1(n7395), .A2(n9918), .A3(n8191), .ZN(n4687) );
  NAND2_X1 U6470 ( .A1(n7395), .A2(n8191), .ZN(n7396) );
  NAND2_X1 U6471 ( .A1(n5316), .A2(n4308), .ZN(n5422) );
  NAND2_X1 U6472 ( .A1(n5522), .A2(n4329), .ZN(n5593) );
  NAND2_X1 U6473 ( .A1(n5619), .A2(n4702), .ZN(n5693) );
  NAND3_X1 U6474 ( .A1(n4811), .A2(n8129), .A3(n4812), .ZN(n8135) );
  NAND2_X1 U6475 ( .A1(n7805), .A2(n6249), .ZN(n6307) );
  NAND2_X1 U6476 ( .A1(n4932), .A2(n5690), .ZN(n4706) );
  NAND2_X1 U6477 ( .A1(n5586), .A2(n4712), .ZN(n4711) );
  NAND3_X1 U6478 ( .A1(n6351), .A2(n6350), .A3(n4717), .ZN(n4716) );
  NAND2_X1 U6479 ( .A1(n4716), .A2(n4719), .ZN(n4899) );
  NAND3_X1 U6480 ( .A1(n6351), .A2(n6350), .A3(n4725), .ZN(n4724) );
  NAND3_X1 U6481 ( .A1(n4730), .A2(n4732), .A3(n4731), .ZN(n6417) );
  OR2_X1 U6482 ( .A1(n6663), .A2(n8360), .ZN(n4737) );
  OAI211_X1 U6483 ( .C1(n4737), .C2(n4740), .A(n4284), .B(n4744), .ZN(n4743)
         );
  NAND2_X1 U6484 ( .A1(n4743), .A2(n4742), .ZN(n6686) );
  NAND2_X1 U6485 ( .A1(n6707), .A2(n6037), .ZN(n6042) );
  NAND4_X1 U6486 ( .A1(n6699), .A2(n7240), .A3(n6751), .A4(n10009), .ZN(n4747)
         );
  NAND3_X1 U6487 ( .A1(n4752), .A2(n8346), .A3(n6629), .ZN(n4751) );
  NAND2_X1 U6488 ( .A1(n4755), .A2(n4753), .ZN(n7056) );
  NAND2_X1 U6489 ( .A1(n6999), .A2(n4756), .ZN(n4755) );
  OAI21_X1 U6490 ( .B1(n6999), .B2(n4758), .A(n4756), .ZN(n7012) );
  XNOR2_X2 U6491 ( .A(n4774), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U6492 ( .A1(n7294), .A2(n6559), .ZN(n6471) );
  INV_X1 U6493 ( .A(n4275), .ZN(n4775) );
  NAND2_X1 U6494 ( .A1(n6645), .A2(n4781), .ZN(n4779) );
  NAND2_X1 U6495 ( .A1(n4779), .A2(n4309), .ZN(n4780) );
  XNOR2_X1 U6496 ( .A(n8659), .B(n8391), .ZN(n7236) );
  NAND2_X4 U6497 ( .A1(n5285), .A2(n5180), .ZN(n8152) );
  OAI21_X1 U6498 ( .B1(n8114), .B2(n4797), .A(n4796), .ZN(n4793) );
  INV_X1 U6499 ( .A(n8121), .ZN(n8125) );
  NAND3_X1 U6500 ( .A1(n8128), .A2(n8126), .A3(n4813), .ZN(n4812) );
  NAND2_X1 U6501 ( .A1(n7396), .A2(n8234), .ZN(n7470) );
  NAND3_X1 U6502 ( .A1(n7396), .A2(n4814), .A3(n4820), .ZN(n4819) );
  NAND3_X1 U6503 ( .A1(n4819), .A2(n8075), .A3(n4816), .ZN(n8078) );
  NAND2_X1 U6504 ( .A1(n7470), .A2(n4817), .ZN(n4816) );
  NAND2_X2 U6505 ( .A1(n5950), .A2(n4849), .ZN(n6910) );
  NAND2_X1 U6506 ( .A1(n6455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6695) );
  AND2_X1 U6507 ( .A1(n8756), .A2(n8745), .ZN(n8741) );
  NAND2_X1 U6508 ( .A1(n8756), .A2(n4306), .ZN(n8707) );
  INV_X1 U6509 ( .A(n4859), .ZN(n7812) );
  INV_X1 U6510 ( .A(n7509), .ZN(n7759) );
  AND3_X2 U6511 ( .A1(n5998), .A2(n5996), .A3(n5995), .ZN(n7509) );
  INV_X1 U6512 ( .A(n8384), .ZN(n6031) );
  NAND3_X1 U6513 ( .A1(n4866), .A2(n4861), .A3(n4860), .ZN(n8384) );
  NAND3_X1 U6514 ( .A1(n6015), .A2(n8590), .A3(n8593), .ZN(n4860) );
  INV_X1 U6515 ( .A(n7501), .ZN(n6015) );
  NAND3_X1 U6516 ( .A1(n4865), .A2(n8598), .A3(n4862), .ZN(n4861) );
  INV_X1 U6517 ( .A(n8590), .ZN(n4863) );
  NAND2_X1 U6518 ( .A1(n7501), .A2(n6014), .ZN(n4865) );
  NAND2_X1 U6519 ( .A1(n4867), .A2(n8591), .ZN(n4866) );
  OAI21_X1 U6520 ( .B1(n7501), .B2(n6014), .A(n4863), .ZN(n4867) );
  NAND2_X1 U6521 ( .A1(n7820), .A2(n4869), .ZN(n4868) );
  INV_X1 U6522 ( .A(n7587), .ZN(n4878) );
  INV_X1 U6523 ( .A(n6088), .ZN(n4871) );
  NAND2_X1 U6524 ( .A1(n4792), .A2(n4302), .ZN(n5961) );
  NAND2_X1 U6525 ( .A1(n6008), .A2(n7511), .ZN(n7501) );
  INV_X2 U6526 ( .A(n6535), .ZN(n6331) );
  NOR2_X4 U6527 ( .A1(n7707), .A2(n7631), .ZN(n7641) );
  XNOR2_X1 U6528 ( .A(n5782), .B(n4904), .ZN(n7930) );
  INV_X1 U6529 ( .A(n5311), .ZN(n4906) );
  NAND2_X1 U6530 ( .A1(n5354), .A2(n5353), .ZN(n5406) );
  NAND2_X1 U6531 ( .A1(n5786), .A2(n4925), .ZN(n4921) );
  NAND2_X1 U6532 ( .A1(n5786), .A2(n5785), .ZN(n5809) );
  INV_X1 U6533 ( .A(n4940), .ZN(n4943) );
  NAND2_X1 U6534 ( .A1(n5725), .A2(n9247), .ZN(n9151) );
  NAND2_X1 U6535 ( .A1(n4958), .A2(n4959), .ZN(n5532) );
  NAND4_X1 U6536 ( .A1(n5328), .A2(n5139), .A3(n5138), .A4(n5171), .ZN(n4963)
         );
  NAND3_X2 U6537 ( .A1(n5221), .A2(n5222), .A3(n5223), .ZN(n9892) );
  XNOR2_X1 U6538 ( .A(n9892), .B(n8236), .ZN(n7324) );
  NAND2_X1 U6539 ( .A1(n8455), .A2(n4977), .ZN(n9441) );
  XNOR2_X1 U6540 ( .A(n4981), .B(n9455), .ZN(n9457) );
  NAND3_X1 U6541 ( .A1(n4988), .A2(n4987), .A3(n10209), .ZN(n9928) );
  NAND2_X1 U6542 ( .A1(n4993), .A2(n4991), .ZN(n7848) );
  NAND2_X1 U6543 ( .A1(n9391), .A2(n9385), .ZN(n9380) );
  NAND2_X1 U6544 ( .A1(n9391), .A2(n4999), .ZN(n5001) );
  AND2_X2 U6545 ( .A1(n9605), .A2(n5003), .ZN(n9529) );
  MUX2_X1 U6546 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n5016), .S(n9972), .Z(
        P1_U3552) );
  MUX2_X1 U6547 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n5016), .S(n9958), .Z(
        P1_U3520) );
  NAND2_X1 U6548 ( .A1(n5033), .A2(n5031), .ZN(n8424) );
  NAND2_X1 U6550 ( .A1(n5042), .A2(n5043), .ZN(n8413) );
  NAND2_X1 U6551 ( .A1(n7840), .A2(n8410), .ZN(n5042) );
  NOR2_X1 U6552 ( .A1(n6779), .A2(n6881), .ZN(n5050) );
  INV_X1 U6553 ( .A(n7236), .ZN(n7238) );
  INV_X1 U6554 ( .A(n8864), .ZN(n5060) );
  NAND2_X1 U6555 ( .A1(n6473), .A2(n5063), .ZN(n7670) );
  NOR2_X1 U6556 ( .A1(n8776), .A2(n6482), .ZN(n8766) );
  NAND3_X1 U6557 ( .A1(n5082), .A2(n4243), .A3(n7684), .ZN(n5081) );
  NAND3_X1 U6558 ( .A1(n5082), .A2(n4243), .A3(n4304), .ZN(n5077) );
  NAND2_X1 U6559 ( .A1(n5079), .A2(n7952), .ZN(n5078) );
  NAND2_X1 U6560 ( .A1(n5080), .A2(n7873), .ZN(n5079) );
  NAND2_X1 U6561 ( .A1(n8789), .A2(n5092), .ZN(n5090) );
  OAI211_X2 U6562 ( .C1(n5108), .C2(n5105), .A(n5102), .B(n5101), .ZN(n8820)
         );
  AOI211_X1 U6563 ( .C1(n9077), .C2(n7672), .A(n10022), .B(n7812), .ZN(n9076)
         );
  NAND2_X1 U6564 ( .A1(n5204), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5206) );
  INV_X1 U6565 ( .A(n8813), .ZN(n8837) );
  NOR2_X2 U6566 ( .A1(n9421), .A2(n9646), .ZN(n9409) );
  OR2_X2 U6567 ( .A1(n7948), .A2(n9066), .ZN(n8018) );
  NAND2_X1 U6568 ( .A1(n8245), .A2(n8234), .ZN(n7370) );
  NAND2_X1 U6569 ( .A1(n6527), .A2(n6910), .ZN(n8977) );
  AOI21_X1 U6570 ( .B1(n5159), .B2(n5153), .A(n4609), .ZN(n5154) );
  CLKBUF_X1 U6571 ( .A(n7538), .Z(n7423) );
  NAND2_X1 U6572 ( .A1(n7198), .A2(n7197), .ZN(n7209) );
  NAND2_X1 U6573 ( .A1(n8599), .A2(n7759), .ZN(n7230) );
  NAND2_X1 U6574 ( .A1(n9892), .A2(n4303), .ZN(n5224) );
  NAND2_X1 U6575 ( .A1(n4303), .A2(n7387), .ZN(n5200) );
  AND2_X1 U6576 ( .A1(n5434), .A2(n5416), .ZN(n5115) );
  AND2_X1 U6577 ( .A1(n5509), .A2(n5494), .ZN(n5116) );
  NAND2_X1 U6578 ( .A1(n8331), .A2(n8313), .ZN(n8177) );
  INV_X1 U6579 ( .A(n8177), .ZN(n5920) );
  AND3_X1 U6580 ( .A1(n7599), .A2(n7598), .A3(n7604), .ZN(n5117) );
  INV_X1 U6581 ( .A(n7333), .ZN(n6472) );
  AND3_X1 U6582 ( .A1(n8531), .A2(n8630), .A3(n8532), .ZN(n5118) );
  AND2_X1 U6583 ( .A1(n8745), .A2(n8351), .ZN(n5119) );
  OR2_X1 U6584 ( .A1(n4998), .A2(n9376), .ZN(n5120) );
  OR2_X1 U6585 ( .A1(n6910), .A2(n5987), .ZN(n5121) );
  AND4_X1 U6586 ( .A1(n5134), .A2(n5162), .A3(n5151), .A4(n5133), .ZN(n5122)
         );
  AND2_X1 U6587 ( .A1(n5164), .A2(n5162), .ZN(n5123) );
  INV_X1 U6588 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5162) );
  AND2_X1 U6589 ( .A1(n5585), .A2(n5563), .ZN(n5124) );
  AND2_X1 U6590 ( .A1(n5180), .A2(P2_U3152), .ZN(n7937) );
  INV_X1 U6591 ( .A(n10208), .ZN(n7315) );
  AND2_X2 U6592 ( .A1(n6763), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X2 U6593 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  OR2_X1 U6594 ( .A1(n9307), .A2(n7414), .ZN(n5125) );
  AND2_X1 U6595 ( .A1(n8340), .A2(n8338), .ZN(n5126) );
  NAND2_X1 U6596 ( .A1(n7448), .A2(n9566), .ZN(n10221) );
  INV_X1 U6597 ( .A(n7471), .ZN(n7472) );
  NAND2_X1 U6598 ( .A1(n8276), .A2(n8167), .ZN(n8129) );
  INV_X1 U6599 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5972) );
  INV_X1 U6600 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5973) );
  OAI21_X1 U6601 ( .B1(n6479), .B2(n6478), .A(n6637), .ZN(n6480) );
  OAI21_X1 U6602 ( .B1(n7211), .B2(n5300), .A(n7208), .ZN(n5298) );
  INV_X1 U6603 ( .A(n5723), .ZN(n5721) );
  INV_X1 U6604 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5155) );
  INV_X1 U6605 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5151) );
  OR2_X1 U6606 ( .A1(n7227), .A2(n6696), .ZN(n7221) );
  OAI21_X1 U6607 ( .B1(n8361), .B2(n6681), .A(n6680), .ZN(n6529) );
  NAND2_X1 U6608 ( .A1(n7732), .A2(n7230), .ZN(n6565) );
  INV_X1 U6609 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6411) );
  INV_X1 U6610 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10136) );
  INV_X1 U6611 ( .A(SI_25_), .ZN(n10178) );
  INV_X1 U6612 ( .A(SI_22_), .ZN(n10154) );
  INV_X1 U6613 ( .A(SI_19_), .ZN(n5636) );
  INV_X1 U6614 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5512) );
  INV_X1 U6615 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10076) );
  INV_X1 U6616 ( .A(n7822), .ZN(n6136) );
  INV_X1 U6617 ( .A(n7221), .ZN(n7222) );
  INV_X1 U6618 ( .A(n7806), .ZN(n6563) );
  INV_X1 U6619 ( .A(n9019), .ZN(n8355) );
  NAND2_X1 U6620 ( .A1(n8704), .A2(n8643), .ZN(n8364) );
  AOI21_X1 U6621 ( .B1(n6412), .B2(n6411), .A(n9120), .ZN(n6434) );
  INV_X1 U6622 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5547) );
  INV_X1 U6623 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7565) );
  INV_X1 U6624 ( .A(SI_13_), .ZN(n10138) );
  OR2_X1 U6625 ( .A1(n8177), .A2(n8328), .ZN(n6867) );
  INV_X1 U6626 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6627 ( .A1(n5270), .A2(n6709), .ZN(n5248) );
  OAI22_X1 U6628 ( .A1(n6239), .A2(n6716), .B1(n6910), .B2(n6020), .ZN(n6021)
         );
  INV_X1 U6629 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U6630 ( .A1(n8386), .A2(n6036), .ZN(n8370) );
  NOR2_X1 U6631 ( .A1(n7223), .A2(n7222), .ZN(n7504) );
  NOR2_X1 U6632 ( .A1(n6449), .A2(n7223), .ZN(n6454) );
  AOI21_X1 U6633 ( .B1(n6531), .B2(n6530), .A(n6539), .ZN(n6533) );
  INV_X1 U6634 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U6635 ( .A1(n6441), .A2(n6563), .ZN(n7227) );
  INV_X1 U6636 ( .A(n8847), .ZN(n8809) );
  AND2_X1 U6637 ( .A1(n6614), .A2(n4245), .ZN(n7953) );
  INV_X1 U6638 ( .A(n7682), .ZN(n7654) );
  INV_X1 U6639 ( .A(n7680), .ZN(n7634) );
  OR2_X1 U6640 ( .A1(n7227), .A2(n6458), .ZN(n8934) );
  NAND2_X1 U6641 ( .A1(n6907), .A2(n10007), .ZN(n7223) );
  OR2_X1 U6642 ( .A1(n8869), .A2(n4769), .ZN(n7635) );
  INV_X1 U6643 ( .A(n7746), .ZN(n10015) );
  NAND2_X1 U6644 ( .A1(n6414), .A2(n6413), .ZN(n6435) );
  NAND2_X1 U6645 ( .A1(n6435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6415) );
  OR2_X1 U6646 ( .A1(n5921), .A2(n9925), .ZN(n9282) );
  INV_X1 U6647 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9209) );
  INV_X1 U6648 ( .A(n9496), .ZN(n9169) );
  AND2_X1 U6649 ( .A1(n9505), .A2(n9504), .ZN(n9525) );
  OR2_X1 U6650 ( .A1(n10210), .A2(n7379), .ZN(n9571) );
  NAND2_X1 U6651 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  INV_X1 U6652 ( .A(n9540), .ZN(n9925) );
  NAND2_X1 U6653 ( .A1(n5897), .A2(n7144), .ZN(n7189) );
  NAND2_X1 U6654 ( .A1(n6491), .A2(n6490), .ZN(n6497) );
  OR2_X1 U6655 ( .A1(n8549), .A2(n8934), .ZN(n8583) );
  INV_X1 U6656 ( .A(n8719), .ZN(n8351) );
  INV_X1 U6657 ( .A(n9029), .ZN(n8855) );
  INV_X1 U6658 ( .A(n8549), .ZN(n8622) );
  INV_X1 U6659 ( .A(n4234), .ZN(n6465) );
  AND2_X1 U6660 ( .A1(n6929), .A2(n6928), .ZN(n9974) );
  INV_X1 U6661 ( .A(n9978), .ZN(n9973) );
  AND2_X1 U6662 ( .A1(n6641), .A2(n6639), .ZN(n8844) );
  INV_X1 U6663 ( .A(n8934), .ZN(n8914) );
  NAND2_X1 U6664 ( .A1(n7241), .A2(n7240), .ZN(n8917) );
  OR2_X1 U6665 ( .A1(n7223), .A2(n7219), .ZN(n9990) );
  NOR2_X1 U6666 ( .A1(n7619), .A2(n4769), .ZN(n8969) );
  INV_X1 U6667 ( .A(n8948), .ZN(n8963) );
  OR2_X1 U6668 ( .A1(n7617), .A2(n7220), .ZN(n7305) );
  AND2_X1 U6669 ( .A1(n7635), .A2(n9096), .ZN(n9081) );
  INV_X1 U6670 ( .A(n9081), .ZN(n10028) );
  AND2_X1 U6671 ( .A1(n4612), .A2(P2_U3152), .ZN(n9127) );
  AND3_X1 U6672 ( .A1(n8151), .A2(n8150), .A3(n8149), .ZN(n8159) );
  AOI21_X1 U6673 ( .B1(n9452), .B2(n5917), .A(n5720), .ZN(n9179) );
  INV_X1 U6674 ( .A(n9847), .ZN(n9817) );
  AND2_X1 U6675 ( .A1(n9788), .A2(n4239), .ZN(n9841) );
  AND2_X1 U6676 ( .A1(n9330), .A2(n8336), .ZN(n9853) );
  NOR2_X1 U6677 ( .A1(n9644), .A2(n10210), .ZN(n9403) );
  AND2_X1 U6678 ( .A1(n8185), .A2(n8453), .ZN(n9480) );
  INV_X1 U6679 ( .A(n9927), .ZN(n9542) );
  INV_X1 U6680 ( .A(n9609), .ZN(n9588) );
  NAND2_X1 U6681 ( .A1(n5902), .A2(n5903), .ZN(n7378) );
  AND2_X1 U6682 ( .A1(n9897), .A2(n9896), .ZN(n9719) );
  OR2_X1 U6683 ( .A1(n8163), .A2(n7181), .ZN(n9896) );
  AND2_X1 U6684 ( .A1(n6896), .A2(n7189), .ZN(n7311) );
  AND2_X1 U6685 ( .A1(n5882), .A2(n5883), .ZN(n7142) );
  AND2_X1 U6686 ( .A1(n7934), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5901) );
  NOR2_X1 U6687 ( .A1(n4612), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9748) );
  INV_X1 U6688 ( .A(n10007), .ZN(n10000) );
  INV_X1 U6689 ( .A(n9007), .ZN(n8782) );
  AND2_X1 U6690 ( .A1(n6438), .A2(n9990), .ZN(n8617) );
  INV_X1 U6691 ( .A(n9974), .ZN(n9976) );
  NAND2_X2 U6692 ( .A1(n7619), .A2(n9990), .ZN(n9996) );
  INV_X2 U6693 ( .A(n9996), .ZN(n9998) );
  NAND2_X1 U6694 ( .A1(n9996), .A2(n9995), .ZN(n8890) );
  AND2_X2 U6695 ( .A1(n7226), .A2(n7618), .ZN(n10030) );
  NOR2_X1 U6696 ( .A1(n10000), .A2(n9999), .ZN(n10001) );
  INV_X1 U6697 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10005) );
  INV_X1 U6698 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8057) );
  INV_X1 U6699 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7789) );
  INV_X1 U6700 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6760) );
  INV_X1 U6701 ( .A(n9271), .ZN(n9286) );
  OR3_X1 U6702 ( .A1(n5908), .A2(n5920), .A3(n9893), .ZN(n9278) );
  INV_X1 U6703 ( .A(n8159), .ZN(n9350) );
  INV_X1 U6704 ( .A(n8425), .ZN(n9428) );
  INV_X1 U6705 ( .A(n9841), .ZN(n9858) );
  OR2_X1 U6706 ( .A1(n6776), .A2(n8336), .ZN(n9847) );
  OR2_X1 U6707 ( .A1(P1_U3083), .A2(n6763), .ZN(n9862) );
  INV_X1 U6708 ( .A(n10221), .ZN(n10210) );
  OR2_X1 U6709 ( .A1(n10210), .A2(n7368), .ZN(n9611) );
  NAND2_X1 U6710 ( .A1(n10221), .A2(n10214), .ZN(n9595) );
  INV_X1 U6711 ( .A(n9972), .ZN(n9969) );
  OR3_X1 U6712 ( .A1(n9702), .A2(n9701), .A3(n9700), .ZN(n9741) );
  INV_X1 U6713 ( .A(n9958), .ZN(n9956) );
  NOR2_X1 U6714 ( .A1(n7143), .A2(n7142), .ZN(n9875) );
  CLKBUF_X1 U6715 ( .A(n9875), .Z(n9891) );
  INV_X1 U6716 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7936) );
  INV_X1 U6717 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7195) );
  INV_X2 U6718 ( .A(n7933), .ZN(n9752) );
  INV_X1 U6719 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U6720 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5128) );
  NOR2_X1 U6721 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5127) );
  AND2_X1 U6722 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  INV_X1 U6723 ( .A(n5188), .ZN(n5139) );
  NOR2_X1 U6724 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U6725 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5131) );
  NAND3_X1 U6726 ( .A1(n5152), .A2(n5132), .A3(n5131), .ZN(n5157) );
  INV_X1 U6727 ( .A(n5157), .ZN(n5135) );
  NOR2_X1 U6728 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5134) );
  INV_X1 U6729 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5133) );
  AND2_X2 U6730 ( .A1(n5135), .A2(n5122), .ZN(n5138) );
  NAND2_X1 U6731 ( .A1(n5172), .A2(n5136), .ZN(n5260) );
  NAND2_X1 U6732 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6733 ( .A1(n5337), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6734 ( .A1(n8155), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5149) );
  AND2_X4 U6735 ( .A1(n9753), .A2(n5145), .ZN(n5443) );
  NAND2_X1 U6736 ( .A1(n5443), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6737 ( .A1(n5332), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5147) );
  INV_X1 U6738 ( .A(n7313), .ZN(n5169) );
  NAND2_X1 U6739 ( .A1(n5159), .A2(n5158), .ZN(n5899) );
  NAND2_X1 U6740 ( .A1(n5163), .A2(n5160), .ZN(n5165) );
  INV_X1 U6741 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5173) );
  INV_X1 U6742 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6710) );
  INV_X1 U6743 ( .A(SI_1_), .ZN(n5216) );
  NAND2_X1 U6744 ( .A1(n6710), .A2(n5216), .ZN(n5175) );
  AND2_X1 U6745 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5198) );
  AOI22_X1 U6746 ( .A1(n5175), .A2(n5198), .B1(P2_DATAO_REG_1__SCAN_IN), .B2(
        SI_1_), .ZN(n5179) );
  AND3_X1 U6747 ( .A1(SI_1_), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5177) );
  NAND2_X1 U6748 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5215) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6729) );
  AOI21_X1 U6750 ( .B1(n5216), .B2(n5215), .A(n6729), .ZN(n5176) );
  OAI21_X1 U6751 ( .B1(n5177), .B2(n5176), .A(n5180), .ZN(n5178) );
  OAI21_X1 U6752 ( .B1(n5180), .B2(n5179), .A(n5178), .ZN(n5244) );
  INV_X1 U6753 ( .A(SI_2_), .ZN(n5241) );
  XNOR2_X1 U6754 ( .A(n5244), .B(n5241), .ZN(n5182) );
  MUX2_X1 U6755 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6522), .Z(n5181) );
  XNOR2_X1 U6756 ( .A(n5182), .B(n5181), .ZN(n6728) );
  OR2_X1 U6757 ( .A1(n5263), .A2(n6728), .ZN(n5184) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6706) );
  OAI22_X1 U6759 ( .A1(n7397), .A2(n5478), .B1(n7175), .B2(n5185), .ZN(n5191)
         );
  NAND2_X4 U6760 ( .A1(n7176), .A2(n7313), .ZN(n5872) );
  XNOR2_X1 U6761 ( .A(n5191), .B(n5872), .ZN(n5229) );
  AOI22_X1 U6762 ( .A1(n7362), .A2(n5746), .B1(n5252), .B2(n7522), .ZN(n5230)
         );
  XNOR2_X1 U6763 ( .A(n5229), .B(n5230), .ZN(n7095) );
  NAND2_X1 U6764 ( .A1(n5337), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6765 ( .A1(n5443), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6766 ( .A1(n5332), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5192) );
  NAND4_X2 U6767 ( .A1(n5195), .A2(n5193), .A3(n5192), .A4(n5194), .ZN(n6757)
         );
  NAND2_X1 U6768 ( .A1(n6757), .A2(n5252), .ZN(n5202) );
  INV_X1 U6769 ( .A(n5898), .ZN(n5204) );
  INV_X1 U6770 ( .A(SI_0_), .ZN(n5999) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5197) );
  OAI21_X1 U6772 ( .B1(n5180), .B2(n5999), .A(n5197), .ZN(n5199) );
  NAND2_X1 U6773 ( .A1(n5270), .A2(n5198), .ZN(n5214) );
  AND2_X1 U6774 ( .A1(n5199), .A2(n5214), .ZN(n9756) );
  MUX2_X1 U6775 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9756), .S(n5285), .Z(n7387) );
  INV_X1 U6776 ( .A(n6876), .ZN(n5203) );
  NAND2_X1 U6777 ( .A1(n5203), .A2(n5872), .ZN(n5208) );
  AND2_X1 U6778 ( .A1(n5208), .A2(n6875), .ZN(n5227) );
  NAND2_X1 U6779 ( .A1(n8155), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6780 ( .A1(n5337), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6781 ( .A1(n5443), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5211) );
  INV_X1 U6782 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6783 ( .A1(n4626), .A2(n5209), .ZN(n5210) );
  OAI21_X1 U6784 ( .B1(n6522), .B2(n5215), .A(n5214), .ZN(n5217) );
  XNOR2_X1 U6785 ( .A(n5217), .B(n5216), .ZN(n5219) );
  MUX2_X1 U6786 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6522), .Z(n5218) );
  XNOR2_X1 U6787 ( .A(n5219), .B(n5218), .ZN(n6730) );
  OR2_X1 U6788 ( .A1(n5263), .A2(n6730), .ZN(n5223) );
  OR2_X1 U6789 ( .A1(n8152), .A2(n6710), .ZN(n5222) );
  INV_X1 U6790 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6791 ( .A1(n5285), .A2(n6783), .ZN(n5221) );
  NAND2_X1 U6792 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  AOI22_X1 U6793 ( .A1(n5746), .A2(n9309), .B1(n9892), .B2(n5252), .ZN(n6863)
         );
  INV_X1 U6794 ( .A(n5229), .ZN(n5231) );
  NAND2_X1 U6795 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  INV_X1 U6796 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6797 ( .A1(n5337), .A2(n5233), .ZN(n5237) );
  NAND2_X1 U6798 ( .A1(n8155), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6799 ( .A1(n5443), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6800 ( .A1(n5238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  INV_X1 U6801 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5239) );
  INV_X1 U6802 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U6803 ( .A1(n5270), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5242) );
  OAI211_X1 U6804 ( .C1(n5270), .C2(n6727), .A(n5242), .B(n5241), .ZN(n5243)
         );
  NAND2_X1 U6805 ( .A1(n5244), .A2(n5243), .ZN(n5247) );
  NAND2_X1 U6806 ( .A1(n5270), .A2(n6706), .ZN(n5245) );
  OAI211_X1 U6807 ( .C1(n5270), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5245), .B(
        SI_2_), .ZN(n5246) );
  NAND2_X1 U6808 ( .A1(n5247), .A2(n5246), .ZN(n5265) );
  INV_X1 U6809 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6716) );
  INV_X1 U6810 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6709) );
  XNOR2_X1 U6811 ( .A(n5265), .B(n5264), .ZN(n6715) );
  OR2_X1 U6812 ( .A1(n6715), .A2(n5263), .ZN(n5250) );
  OR2_X1 U6813 ( .A1(n8152), .A2(n6709), .ZN(n5249) );
  OAI22_X1 U6814 ( .A1(n7374), .A2(n5478), .B1(n4989), .B2(n5185), .ZN(n5251)
         );
  XNOR2_X1 U6815 ( .A(n5251), .B(n5872), .ZN(n5253) );
  AOI22_X1 U6816 ( .A1(n9308), .A2(n5746), .B1(n5252), .B2(n7405), .ZN(n5254)
         );
  XNOR2_X1 U6817 ( .A(n5253), .B(n5254), .ZN(n7164) );
  INV_X1 U6818 ( .A(n5253), .ZN(n5255) );
  NAND2_X1 U6819 ( .A1(n8155), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5259) );
  INV_X1 U6820 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U6821 ( .A(n5257), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U6822 ( .A1(n5443), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6823 ( .A1(n5260), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5261) );
  MUX2_X1 U6824 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5261), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5262) );
  OR2_X1 U6825 ( .A1(n5260), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6826 ( .A1(n5262), .A2(n5286), .ZN(n6881) );
  INV_X2 U6827 ( .A(n5263), .ZN(n5327) );
  NAND2_X1 U6828 ( .A1(n5265), .A2(n5264), .ZN(n5269) );
  INV_X1 U6829 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6830 ( .A1(n5267), .A2(SI_3_), .ZN(n5268) );
  MUX2_X1 U6831 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5270), .Z(n5282) );
  XNOR2_X1 U6832 ( .A(n5282), .B(SI_4_), .ZN(n5281) );
  XNOR2_X1 U6833 ( .A(n5271), .B(n5281), .ZN(n6707) );
  INV_X1 U6834 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6708) );
  OR2_X1 U6835 ( .A1(n8152), .A2(n6708), .ZN(n5272) );
  OAI22_X1 U6836 ( .A1(n9924), .A2(n5478), .B1(n9909), .B2(n5185), .ZN(n5273)
         );
  XNOR2_X1 U6837 ( .A(n5273), .B(n5872), .ZN(n5297) );
  AOI22_X1 U6838 ( .A1(n9307), .A2(n5746), .B1(n5252), .B2(n7414), .ZN(n5295)
         );
  XNOR2_X1 U6839 ( .A(n5297), .B(n5295), .ZN(n7197) );
  NAND2_X1 U6840 ( .A1(n8155), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5280) );
  INV_X1 U6841 ( .A(n5315), .ZN(n5334) );
  INV_X1 U6842 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6843 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5274) );
  NAND2_X1 U6844 ( .A1(n5275), .A2(n5274), .ZN(n5276) );
  AND2_X1 U6845 ( .A1(n5334), .A2(n5276), .ZN(n10212) );
  NAND2_X1 U6846 ( .A1(n5917), .A2(n10212), .ZN(n5279) );
  NAND2_X1 U6847 ( .A1(n5332), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6848 ( .A1(n5443), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6849 ( .A1(n9305), .A2(n5252), .ZN(n5291) );
  NAND2_X1 U6850 ( .A1(n5282), .A2(SI_4_), .ZN(n5283) );
  INV_X1 U6851 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6718) );
  INV_X1 U6852 ( .A(n5303), .ZN(n5284) );
  XNOR2_X1 U6853 ( .A(n5304), .B(n5284), .ZN(n6704) );
  NAND2_X1 U6854 ( .A1(n6704), .A2(n5327), .ZN(n5289) );
  INV_X2 U6855 ( .A(n8152), .ZN(n5360) );
  NAND2_X1 U6856 ( .A1(n5286), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5287) );
  XNOR2_X1 U6857 ( .A(n5287), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7077) );
  AOI22_X1 U6858 ( .A1(n5360), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5640), .B2(
        n7077), .ZN(n5288) );
  NAND2_X1 U6859 ( .A1(n8067), .A2(n4633), .ZN(n5290) );
  NAND2_X1 U6860 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  XNOR2_X1 U6861 ( .A(n5292), .B(n5798), .ZN(n7211) );
  NAND2_X1 U6862 ( .A1(n5746), .A2(n9305), .ZN(n5294) );
  NAND2_X1 U6863 ( .A1(n8067), .A2(n5874), .ZN(n5293) );
  AND2_X1 U6864 ( .A1(n5294), .A2(n5293), .ZN(n5300) );
  INV_X1 U6865 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6866 ( .A1(n5297), .A2(n5296), .ZN(n7208) );
  NAND2_X1 U6867 ( .A1(n7209), .A2(n5299), .ZN(n5302) );
  INV_X1 U6868 ( .A(n5300), .ZN(n7210) );
  NAND2_X1 U6869 ( .A1(n7211), .A2(n5300), .ZN(n5301) );
  NAND2_X1 U6870 ( .A1(n5302), .A2(n5301), .ZN(n7458) );
  INV_X1 U6871 ( .A(n5305), .ZN(n5306) );
  NAND2_X1 U6872 ( .A1(n5306), .A2(SI_5_), .ZN(n5307) );
  MUX2_X1 U6873 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6522), .Z(n5310) );
  XNOR2_X1 U6874 ( .A(n5310), .B(SI_6_), .ZN(n5326) );
  INV_X1 U6875 ( .A(n5326), .ZN(n5309) );
  NAND2_X1 U6876 ( .A1(n5310), .A2(SI_6_), .ZN(n5311) );
  MUX2_X1 U6877 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6522), .Z(n5355) );
  OR2_X1 U6878 ( .A1(n5159), .A2(n4609), .ZN(n5312) );
  XNOR2_X1 U6879 ( .A(n5312), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U6880 ( .A1(n5360), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5640), .B2(
        n6849), .ZN(n5313) );
  NAND2_X1 U6881 ( .A1(n8155), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6882 ( .A1(n5315), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5336) );
  INV_X1 U6883 ( .A(n5336), .ZN(n5316) );
  INV_X1 U6884 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6885 ( .A1(n5336), .A2(n5317), .ZN(n5318) );
  AND2_X1 U6886 ( .A1(n5366), .A2(n5318), .ZN(n7614) );
  NAND2_X1 U6887 ( .A1(n5917), .A2(n7614), .ZN(n5321) );
  NAND2_X1 U6888 ( .A1(n5332), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6889 ( .A1(n5443), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6890 ( .A1(n7607), .A2(n5252), .ZN(n5325) );
  NAND2_X1 U6891 ( .A1(n9303), .A2(n5746), .ZN(n5324) );
  NAND2_X1 U6892 ( .A1(n5325), .A2(n5324), .ZN(n7604) );
  NAND2_X1 U6893 ( .A1(n6711), .A2(n5327), .ZN(n5331) );
  OR2_X1 U6894 ( .A1(n5328), .A2(n4609), .ZN(n5329) );
  XNOR2_X1 U6895 ( .A(n5329), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U6896 ( .A1(n5360), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5640), .B2(
        n6810), .ZN(n5330) );
  NAND2_X1 U6897 ( .A1(n8155), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6898 ( .A1(n5332), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6899 ( .A1(n5443), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5339) );
  INV_X1 U6900 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6901 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  AND2_X1 U6902 ( .A1(n5336), .A2(n5335), .ZN(n7481) );
  NAND2_X1 U6903 ( .A1(n5337), .A2(n7481), .ZN(n5338) );
  NAND2_X1 U6904 ( .A1(n9304), .A2(n5252), .ZN(n5342) );
  OAI21_X1 U6905 ( .B1(n9933), .B2(n5185), .A(n5342), .ZN(n5343) );
  XNOR2_X1 U6906 ( .A(n5343), .B(n5872), .ZN(n7599) );
  OR2_X1 U6907 ( .A1(n9933), .A2(n5478), .ZN(n5346) );
  NAND2_X1 U6908 ( .A1(n5746), .A2(n9304), .ZN(n5345) );
  NAND2_X1 U6909 ( .A1(n5346), .A2(n5345), .ZN(n7598) );
  OAI22_X1 U6910 ( .A1(n7603), .A2(n7604), .B1(n7599), .B2(n7598), .ZN(n5351)
         );
  INV_X1 U6911 ( .A(n7599), .ZN(n7602) );
  INV_X1 U6912 ( .A(n7598), .ZN(n7460) );
  NOR2_X1 U6913 ( .A1(n7602), .A2(n7460), .ZN(n5347) );
  OAI21_X1 U6914 ( .B1(n5347), .B2(n7604), .A(n7603), .ZN(n5348) );
  NAND2_X1 U6915 ( .A1(n5355), .A2(SI_7_), .ZN(n5402) );
  NAND2_X1 U6916 ( .A1(n5406), .A2(n5402), .ZN(n5380) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6735) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5356) );
  MUX2_X1 U6919 ( .A(n6735), .B(n5356), .S(n6522), .Z(n5358) );
  INV_X1 U6920 ( .A(SI_8_), .ZN(n5357) );
  NAND2_X1 U6921 ( .A1(n5358), .A2(n5357), .ZN(n5407) );
  INV_X1 U6922 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6923 ( .A1(n5359), .A2(SI_8_), .ZN(n5401) );
  NAND2_X1 U6924 ( .A1(n5407), .A2(n5401), .ZN(n5379) );
  XNOR2_X1 U6925 ( .A(n5380), .B(n5379), .ZN(n6732) );
  NAND2_X1 U6926 ( .A1(n6732), .A2(n5327), .ZN(n5364) );
  NAND2_X1 U6927 ( .A1(n5361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6928 ( .A(n5362), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U6929 ( .A1(n5360), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5640), .B2(
        n6823), .ZN(n5363) );
  NAND2_X1 U6930 ( .A1(n5364), .A2(n5363), .ZN(n7536) );
  NAND2_X1 U6931 ( .A1(n7536), .A2(n4633), .ZN(n5374) );
  NAND2_X1 U6932 ( .A1(n4615), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5372) );
  INV_X1 U6933 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6934 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  AND2_X1 U6935 ( .A1(n5388), .A2(n5367), .ZN(n7498) );
  NAND2_X1 U6936 ( .A1(n5917), .A2(n7498), .ZN(n5371) );
  NAND2_X1 U6937 ( .A1(n8148), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6938 ( .A1(n5443), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5369) );
  OR2_X1 U6939 ( .A1(n7611), .A2(n5478), .ZN(n5373) );
  NAND2_X1 U6940 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  XNOR2_X1 U6941 ( .A(n5375), .B(n5798), .ZN(n7490) );
  NOR2_X1 U6942 ( .A1(n7611), .A2(n5876), .ZN(n5376) );
  AOI21_X1 U6943 ( .B1(n7536), .B2(n5874), .A(n5376), .ZN(n5377) );
  INV_X1 U6944 ( .A(n7490), .ZN(n5378) );
  INV_X1 U6945 ( .A(n5377), .ZN(n7489) );
  INV_X1 U6946 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6744) );
  INV_X1 U6947 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6742) );
  MUX2_X1 U6948 ( .A(n6744), .B(n6742), .S(n4612), .Z(n5382) );
  INV_X1 U6949 ( .A(SI_9_), .ZN(n5381) );
  NAND2_X1 U6950 ( .A1(n5382), .A2(n5381), .ZN(n5408) );
  INV_X1 U6951 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6952 ( .A1(n5383), .A2(SI_9_), .ZN(n5384) );
  NAND2_X1 U6953 ( .A1(n5408), .A2(n5384), .ZN(n5404) );
  INV_X1 U6954 ( .A(n5404), .ZN(n5411) );
  NAND2_X1 U6955 ( .A1(n6740), .A2(n5327), .ZN(n5387) );
  NAND2_X1 U6956 ( .A1(n5417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U6957 ( .A(n5385), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U6958 ( .A1(n5360), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5640), .B2(
        n7018), .ZN(n5386) );
  NAND2_X1 U6959 ( .A1(n9720), .A2(n4633), .ZN(n5395) );
  NAND2_X1 U6960 ( .A1(n4615), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6961 ( .A1(n5388), .A2(n6807), .ZN(n5389) );
  AND2_X1 U6962 ( .A1(n5422), .A2(n5389), .ZN(n7771) );
  NAND2_X1 U6963 ( .A1(n5917), .A2(n7771), .ZN(n5392) );
  NAND2_X1 U6964 ( .A1(n8148), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6965 ( .A1(n5443), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5390) );
  NAND4_X1 U6966 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n9301)
         );
  NAND2_X1 U6967 ( .A1(n9301), .A2(n5874), .ZN(n5394) );
  NAND2_X1 U6968 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  XNOR2_X1 U6969 ( .A(n5396), .B(n5872), .ZN(n5400) );
  NAND2_X1 U6970 ( .A1(n9720), .A2(n5874), .ZN(n5398) );
  NAND2_X1 U6971 ( .A1(n5746), .A2(n9301), .ZN(n5397) );
  NAND2_X1 U6972 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U6973 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NOR2_X1 U6974 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  INV_X1 U6975 ( .A(n5407), .ZN(n5410) );
  INV_X1 U6976 ( .A(n5408), .ZN(n5409) );
  AOI21_X1 U6977 ( .B1(n5411), .B2(n5410), .A(n5409), .ZN(n5412) );
  MUX2_X1 U6978 ( .A(n6739), .B(n6737), .S(n4612), .Z(n5414) );
  INV_X1 U6979 ( .A(SI_10_), .ZN(n5413) );
  NAND2_X1 U6980 ( .A1(n5414), .A2(n5413), .ZN(n5434) );
  INV_X1 U6981 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6982 ( .A1(n5415), .A2(SI_10_), .ZN(n5416) );
  NAND2_X1 U6983 ( .A1(n6736), .A2(n5327), .ZN(n5420) );
  NAND2_X1 U6984 ( .A1(n5435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U6985 ( .A(n5418), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7102) );
  AOI22_X1 U6986 ( .A1(n5360), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7102), .B2(
        n5640), .ZN(n5419) );
  NAND2_X1 U6987 ( .A1(n5420), .A2(n5419), .ZN(n9715) );
  NAND2_X1 U6988 ( .A1(n9715), .A2(n4633), .ZN(n5429) );
  NAND2_X1 U6989 ( .A1(n4615), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6990 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  AND2_X1 U6991 ( .A1(n5441), .A2(n5423), .ZN(n7802) );
  NAND2_X1 U6992 ( .A1(n5917), .A2(n7802), .ZN(n5426) );
  NAND2_X1 U6993 ( .A1(n5443), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6994 ( .A1(n8148), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5424) );
  OR2_X1 U6995 ( .A1(n7777), .A2(n5478), .ZN(n5428) );
  NAND2_X1 U6996 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  XNOR2_X1 U6997 ( .A(n5430), .B(n5798), .ZN(n5433) );
  NOR2_X1 U6998 ( .A1(n7777), .A2(n5876), .ZN(n5431) );
  AOI21_X1 U6999 ( .B1(n9715), .B2(n5874), .A(n5431), .ZN(n5432) );
  NOR2_X1 U7000 ( .A1(n5433), .A2(n5432), .ZN(n7793) );
  NAND2_X1 U7001 ( .A1(n5433), .A2(n5432), .ZN(n7792) );
  MUX2_X1 U7002 ( .A(n6746), .B(n6748), .S(n4612), .Z(n5457) );
  XNOR2_X1 U7003 ( .A(n5457), .B(SI_11_), .ZN(n5456) );
  XNOR2_X1 U7004 ( .A(n5461), .B(n5456), .ZN(n6745) );
  NAND2_X1 U7005 ( .A1(n6745), .A2(n5327), .ZN(n5438) );
  OR2_X1 U7006 ( .A1(n5467), .A2(n4609), .ZN(n5436) );
  XNOR2_X1 U7007 ( .A(n5436), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7347) );
  AOI22_X1 U7008 ( .A1(n7347), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7009 ( .A1(n7893), .A2(n4633), .ZN(n5449) );
  NAND2_X1 U7010 ( .A1(n4615), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5447) );
  INV_X1 U7011 ( .A(n5441), .ZN(n5439) );
  NAND2_X1 U7012 ( .A1(n5439), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5472) );
  INV_X1 U7013 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U7014 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  AND2_X1 U7015 ( .A1(n5472), .A2(n5442), .ZN(n7889) );
  NAND2_X1 U7016 ( .A1(n5917), .A2(n7889), .ZN(n5446) );
  NAND2_X1 U7017 ( .A1(n5443), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U7018 ( .A1(n8148), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5444) );
  NAND4_X1 U7019 ( .A1(n5447), .A2(n5446), .A3(n5445), .A4(n5444), .ZN(n9299)
         );
  NAND2_X1 U7020 ( .A1(n9299), .A2(n5874), .ZN(n5448) );
  NAND2_X1 U7021 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XNOR2_X1 U7022 ( .A(n5450), .B(n5872), .ZN(n7883) );
  NAND2_X1 U7023 ( .A1(n7893), .A2(n5874), .ZN(n5452) );
  NAND2_X1 U7024 ( .A1(n5746), .A2(n9299), .ZN(n5451) );
  NAND2_X1 U7025 ( .A1(n5452), .A2(n5451), .ZN(n7882) );
  NOR2_X1 U7026 ( .A1(n7883), .A2(n7882), .ZN(n5455) );
  INV_X1 U7027 ( .A(n7883), .ZN(n5454) );
  INV_X1 U7028 ( .A(n7882), .ZN(n5453) );
  INV_X1 U7029 ( .A(n5456), .ZN(n5460) );
  INV_X1 U7030 ( .A(n5457), .ZN(n5458) );
  NAND2_X1 U7031 ( .A1(n5458), .A2(SI_11_), .ZN(n5459) );
  INV_X1 U7032 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5462) );
  MUX2_X1 U7033 ( .A(n6760), .B(n5462), .S(n4612), .Z(n5463) );
  NAND2_X1 U7034 ( .A1(n5463), .A2(n10082), .ZN(n5490) );
  INV_X1 U7035 ( .A(n5463), .ZN(n5464) );
  NAND2_X1 U7036 ( .A1(n5464), .A2(SI_12_), .ZN(n5465) );
  NAND2_X1 U7037 ( .A1(n5490), .A2(n5465), .ZN(n5488) );
  XNOR2_X1 U7038 ( .A(n5487), .B(n5488), .ZN(n6755) );
  NAND2_X1 U7039 ( .A1(n6755), .A2(n5327), .ZN(n5469) );
  NAND2_X1 U7040 ( .A1(n5467), .A2(n5466), .ZN(n5514) );
  NAND2_X1 U7041 ( .A1(n5514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U7042 ( .A(n5495), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U7043 ( .A1(n7556), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7044 ( .A1(n8409), .A2(n4633), .ZN(n5480) );
  NAND2_X1 U7045 ( .A1(n4615), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5477) );
  INV_X1 U7046 ( .A(n5472), .ZN(n5470) );
  NAND2_X1 U7047 ( .A1(n5470), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5500) );
  INV_X1 U7048 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7049 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  AND2_X1 U7050 ( .A1(n5500), .A2(n5473), .ZN(n7967) );
  NAND2_X1 U7051 ( .A1(n5917), .A2(n7967), .ZN(n5476) );
  NAND2_X1 U7052 ( .A1(n5443), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7053 ( .A1(n8148), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5474) );
  OR2_X1 U7054 ( .A1(n9597), .A2(n5478), .ZN(n5479) );
  NAND2_X1 U7055 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  XNOR2_X1 U7056 ( .A(n5481), .B(n5798), .ZN(n5483) );
  NOR2_X1 U7057 ( .A1(n9597), .A2(n5876), .ZN(n5482) );
  AOI21_X1 U7058 ( .B1(n8409), .B2(n5874), .A(n5482), .ZN(n5484) );
  NAND2_X1 U7059 ( .A1(n5483), .A2(n5484), .ZN(n7959) );
  INV_X1 U7060 ( .A(n5483), .ZN(n5486) );
  INV_X1 U7061 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U7062 ( .A1(n5486), .A2(n5485), .ZN(n7960) );
  INV_X1 U7063 ( .A(n5488), .ZN(n5489) );
  INV_X1 U7064 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U7065 ( .A(n10105), .B(n5491), .S(n4612), .Z(n5492) );
  NAND2_X1 U7066 ( .A1(n5492), .A2(n10138), .ZN(n5509) );
  INV_X1 U7067 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U7068 ( .A1(n5493), .A2(SI_13_), .ZN(n5494) );
  XNOR2_X1 U7069 ( .A(n5508), .B(n5116), .ZN(n6761) );
  NAND2_X1 U7070 ( .A1(n6761), .A2(n5327), .ZN(n5499) );
  NAND2_X1 U7071 ( .A1(n5495), .A2(n5512), .ZN(n5496) );
  NAND2_X1 U7072 ( .A1(n5496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5497) );
  XNOR2_X1 U7073 ( .A(n5497), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7979) );
  AOI22_X1 U7074 ( .A1(n7979), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5498) );
  INV_X1 U7075 ( .A(n9709), .ZN(n9610) );
  NAND2_X1 U7076 ( .A1(n4615), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7077 ( .A1(n5500), .A2(n7565), .ZN(n5501) );
  AND2_X1 U7078 ( .A1(n5524), .A2(n5501), .ZN(n9607) );
  NAND2_X1 U7079 ( .A1(n5917), .A2(n9607), .ZN(n5504) );
  NAND2_X1 U7080 ( .A1(n5443), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7081 ( .A1(n8148), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5502) );
  NAND4_X1 U7082 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n9297)
         );
  OAI22_X1 U7083 ( .A1(n9610), .A2(n5185), .B1(n9579), .B2(n5478), .ZN(n5506)
         );
  XNOR2_X1 U7084 ( .A(n5506), .B(n5872), .ZN(n5507) );
  OAI22_X1 U7085 ( .A1(n9610), .A2(n5478), .B1(n9579), .B2(n5876), .ZN(n9236)
         );
  INV_X1 U7086 ( .A(n5507), .ZN(n9237) );
  MUX2_X1 U7087 ( .A(n6830), .B(n6832), .S(n6522), .Z(n5534) );
  XNOR2_X1 U7088 ( .A(n5534), .B(SI_14_), .ZN(n5533) );
  NAND2_X1 U7089 ( .A1(n6829), .A2(n5327), .ZN(n5521) );
  INV_X1 U7090 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7091 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U7092 ( .A1(n5516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5515) );
  MUX2_X1 U7093 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5515), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5518) );
  INV_X1 U7094 ( .A(n5565), .ZN(n5517) );
  NAND2_X1 U7095 ( .A1(n5518), .A2(n5517), .ZN(n9316) );
  OAI22_X1 U7096 ( .A1(n9316), .A2(n6779), .B1(n8152), .B2(n6832), .ZN(n5519)
         );
  INV_X1 U7097 ( .A(n5519), .ZN(n5520) );
  INV_X1 U7098 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7099 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  AND2_X1 U7100 ( .A1(n5548), .A2(n5525), .ZN(n9587) );
  NAND2_X1 U7101 ( .A1(n9587), .A2(n5917), .ZN(n5529) );
  NAND2_X1 U7102 ( .A1(n8148), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7103 ( .A1(n4615), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7104 ( .A1(n5443), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5526) );
  NAND4_X1 U7105 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n9296)
         );
  OAI22_X1 U7106 ( .A1(n9584), .A2(n5185), .B1(n9598), .B2(n5478), .ZN(n5530)
         );
  XNOR2_X1 U7107 ( .A(n5530), .B(n5872), .ZN(n5531) );
  OAI22_X1 U7108 ( .A1(n9584), .A2(n5478), .B1(n9598), .B2(n5876), .ZN(n9144)
         );
  INV_X1 U7109 ( .A(n5533), .ZN(n5537) );
  INV_X1 U7110 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7111 ( .A1(n5535), .A2(SI_14_), .ZN(n5536) );
  INV_X1 U7112 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5539) );
  MUX2_X1 U7113 ( .A(n10064), .B(n5539), .S(n6522), .Z(n5541) );
  INV_X1 U7114 ( .A(SI_15_), .ZN(n5540) );
  NAND2_X1 U7115 ( .A1(n5541), .A2(n5540), .ZN(n5557) );
  INV_X1 U7116 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7117 ( .A1(n5542), .A2(SI_15_), .ZN(n5543) );
  NAND2_X1 U7118 ( .A1(n5557), .A2(n5543), .ZN(n5558) );
  XNOR2_X1 U7119 ( .A(n5559), .B(n5558), .ZN(n7091) );
  NAND2_X1 U7120 ( .A1(n7091), .A2(n5327), .ZN(n5546) );
  OR2_X1 U7121 ( .A1(n5565), .A2(n4609), .ZN(n5544) );
  XNOR2_X1 U7122 ( .A(n5544), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9333) );
  AOI22_X1 U7123 ( .A1(n9333), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7124 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  NAND2_X1 U7125 ( .A1(n5569), .A2(n5549), .ZN(n9567) );
  NAND2_X1 U7126 ( .A1(n4615), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7127 ( .A1(n8148), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5550) );
  AND2_X1 U7128 ( .A1(n5551), .A2(n5550), .ZN(n5553) );
  NAND2_X1 U7129 ( .A1(n5443), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5552) );
  OAI211_X1 U7130 ( .C1(n9567), .C2(n5848), .A(n5553), .B(n5552), .ZN(n9541)
         );
  INV_X1 U7131 ( .A(n9541), .ZN(n9580) );
  OAI22_X1 U7132 ( .A1(n9698), .A2(n5185), .B1(n9580), .B2(n5478), .ZN(n5554)
         );
  XNOR2_X1 U7133 ( .A(n5554), .B(n5872), .ZN(n5555) );
  OAI22_X1 U7134 ( .A1(n9698), .A2(n5478), .B1(n9580), .B2(n5876), .ZN(n9280)
         );
  MUX2_X1 U7135 ( .A(n10108), .B(n7195), .S(n4612), .Z(n5561) );
  NAND2_X1 U7136 ( .A1(n5561), .A2(n5560), .ZN(n5585) );
  INV_X1 U7137 ( .A(n5561), .ZN(n5562) );
  NAND2_X1 U7138 ( .A1(n5562), .A2(SI_16_), .ZN(n5563) );
  NAND2_X1 U7139 ( .A1(n7193), .A2(n5327), .ZN(n5568) );
  NAND2_X1 U7140 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U7141 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5589) );
  XNOR2_X1 U7142 ( .A(n5589), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U7143 ( .A1(n9828), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7144 ( .A1(n9693), .A2(n4633), .ZN(n5575) );
  NAND2_X1 U7145 ( .A1(n5569), .A2(n4701), .ZN(n5570) );
  NAND2_X1 U7146 ( .A1(n5593), .A2(n5570), .ZN(n9547) );
  OR2_X1 U7147 ( .A1(n9547), .A2(n5848), .ZN(n5573) );
  AOI22_X1 U7148 ( .A1(n4615), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8148), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7149 ( .A1(n5443), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7150 ( .A1(n9522), .A2(n5874), .ZN(n5574) );
  NAND2_X1 U7151 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  XNOR2_X1 U7152 ( .A(n5576), .B(n5872), .ZN(n5579) );
  NAND2_X1 U7153 ( .A1(n9693), .A2(n5874), .ZN(n5578) );
  NAND2_X1 U7154 ( .A1(n9522), .A2(n5746), .ZN(n5577) );
  NAND2_X1 U7155 ( .A1(n5578), .A2(n5577), .ZN(n5580) );
  NAND2_X1 U7156 ( .A1(n5579), .A2(n5580), .ZN(n9196) );
  INV_X1 U7157 ( .A(n5579), .ZN(n5582) );
  INV_X1 U7158 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7159 ( .A1(n5582), .A2(n5581), .ZN(n9197) );
  NAND2_X1 U7160 ( .A1(n5583), .A2(n9197), .ZN(n9205) );
  INV_X1 U7161 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5587) );
  MUX2_X1 U7162 ( .A(n7207), .B(n5587), .S(n4612), .Z(n5608) );
  XNOR2_X1 U7163 ( .A(n5608), .B(SI_17_), .ZN(n5607) );
  XNOR2_X1 U7164 ( .A(n5612), .B(n5607), .ZN(n7204) );
  NAND2_X1 U7165 ( .A1(n7204), .A2(n5327), .ZN(n5592) );
  INV_X1 U7166 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7167 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7168 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5614) );
  XNOR2_X1 U7169 ( .A(n5614), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9839) );
  AOI22_X1 U7170 ( .A1(n9839), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7171 ( .A1(n9687), .A2(n4633), .ZN(n5601) );
  NAND2_X1 U7172 ( .A1(n5593), .A2(n9209), .ZN(n5594) );
  AND2_X1 U7173 ( .A1(n5620), .A2(n5594), .ZN(n9530) );
  NAND2_X1 U7174 ( .A1(n9530), .A2(n5917), .ZN(n5599) );
  INV_X1 U7175 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U7176 ( .A1(n5443), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7177 ( .A1(n8148), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7178 ( .C1(n5914), .C2(n9337), .A(n5596), .B(n5595), .ZN(n5597)
         );
  INV_X1 U7179 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7180 ( .A1(n9543), .A2(n5874), .ZN(n5600) );
  NAND2_X1 U7181 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  XNOR2_X1 U7182 ( .A(n5602), .B(n5872), .ZN(n5603) );
  AOI22_X1 U7183 ( .A1(n9687), .A2(n5874), .B1(n5207), .B2(n9543), .ZN(n5604)
         );
  XNOR2_X1 U7184 ( .A(n5603), .B(n5604), .ZN(n9207) );
  INV_X1 U7185 ( .A(n5603), .ZN(n5605) );
  NAND2_X1 U7186 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  INV_X1 U7187 ( .A(n5607), .ZN(n5611) );
  INV_X1 U7188 ( .A(n5608), .ZN(n5609) );
  NAND2_X1 U7189 ( .A1(n5609), .A2(SI_17_), .ZN(n5610) );
  MUX2_X1 U7190 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4612), .Z(n5635) );
  XNOR2_X1 U7191 ( .A(n5635), .B(SI_18_), .ZN(n5632) );
  NAND2_X1 U7192 ( .A1(n7408), .A2(n5327), .ZN(n5618) );
  NAND2_X1 U7193 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U7194 ( .A1(n5615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5616) );
  XNOR2_X1 U7195 ( .A(n5616), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9854) );
  AOI22_X1 U7196 ( .A1(n9854), .A2(n5640), .B1(n5360), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7197 ( .A1(n9681), .A2(n5874), .ZN(n5628) );
  NAND2_X1 U7198 ( .A1(n5620), .A2(n4704), .ZN(n5621) );
  NAND2_X1 U7199 ( .A1(n5644), .A2(n5621), .ZN(n9513) );
  OR2_X1 U7200 ( .A1(n9513), .A2(n5848), .ZN(n5626) );
  INV_X1 U7201 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U7202 ( .A1(n8148), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7203 ( .A1(n5443), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5622) );
  OAI211_X1 U7204 ( .C1(n5914), .C2(n9339), .A(n5623), .B(n5622), .ZN(n5624)
         );
  INV_X1 U7205 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7206 ( .A1(n9523), .A2(n5746), .ZN(n5627) );
  NAND2_X1 U7207 ( .A1(n5628), .A2(n5627), .ZN(n9164) );
  NAND2_X1 U7208 ( .A1(n9681), .A2(n4633), .ZN(n5630) );
  NAND2_X1 U7209 ( .A1(n9523), .A2(n5874), .ZN(n5629) );
  NAND2_X1 U7210 ( .A1(n5630), .A2(n5629), .ZN(n5631) );
  XNOR2_X1 U7211 ( .A(n5631), .B(n5872), .ZN(n9165) );
  INV_X1 U7212 ( .A(n5632), .ZN(n5633) );
  MUX2_X1 U7213 ( .A(n7535), .B(n8393), .S(n4612), .Z(n5637) );
  NAND2_X1 U7214 ( .A1(n5637), .A2(n5636), .ZN(n5662) );
  INV_X1 U7215 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7216 ( .A1(n5638), .A2(SI_19_), .ZN(n5639) );
  NAND2_X1 U7217 ( .A1(n5662), .A2(n5639), .ZN(n5663) );
  XNOR2_X1 U7218 ( .A(n5664), .B(n5663), .ZN(n7534) );
  NAND2_X1 U7219 ( .A1(n7534), .A2(n5327), .ZN(n5642) );
  AOI22_X1 U7220 ( .A1(n5360), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10220), 
        .B2(n5640), .ZN(n5641) );
  NAND2_X1 U7221 ( .A1(n9676), .A2(n4633), .ZN(n5652) );
  NAND2_X1 U7222 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  AND2_X1 U7223 ( .A1(n5671), .A2(n5645), .ZN(n9491) );
  NAND2_X1 U7224 ( .A1(n9491), .A2(n5917), .ZN(n5650) );
  INV_X1 U7225 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U7226 ( .A1(n8148), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7227 ( .A1(n5443), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7228 ( .C1(n5914), .C2(n9341), .A(n5647), .B(n5646), .ZN(n5648)
         );
  INV_X1 U7229 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U7230 ( .A1(n5650), .A2(n5649), .ZN(n9508) );
  NAND2_X1 U7231 ( .A1(n9508), .A2(n5874), .ZN(n5651) );
  NAND2_X1 U7232 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  XNOR2_X1 U7233 ( .A(n5653), .B(n5798), .ZN(n5656) );
  AND2_X1 U7234 ( .A1(n9508), .A2(n5746), .ZN(n5654) );
  AOI21_X1 U7235 ( .B1(n9676), .B2(n5874), .A(n5654), .ZN(n5657) );
  NOR2_X1 U7236 ( .A1(n5656), .A2(n5657), .ZN(n9163) );
  AOI21_X1 U7237 ( .B1(n9164), .B2(n9165), .A(n9163), .ZN(n5655) );
  NOR3_X1 U7238 ( .A1(n9163), .A2(n9164), .A3(n9165), .ZN(n5660) );
  INV_X1 U7239 ( .A(n5656), .ZN(n5659) );
  INV_X1 U7240 ( .A(n5657), .ZN(n5658) );
  NOR2_X1 U7241 ( .A1(n5659), .A2(n5658), .ZN(n9225) );
  NOR2_X1 U7242 ( .A1(n5660), .A2(n9225), .ZN(n5661) );
  MUX2_X1 U7243 ( .A(n7789), .B(n7791), .S(n4612), .Z(n5666) );
  NAND2_X1 U7244 ( .A1(n5666), .A2(n5665), .ZN(n5690) );
  INV_X1 U7245 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7246 ( .A1(n5667), .A2(SI_20_), .ZN(n5668) );
  XNOR2_X1 U7247 ( .A(n5689), .B(n5688), .ZN(n7788) );
  NAND2_X1 U7248 ( .A1(n7788), .A2(n5327), .ZN(n5670) );
  OR2_X1 U7249 ( .A1(n8152), .A2(n7791), .ZN(n5669) );
  NAND2_X1 U7250 ( .A1(n9672), .A2(n4633), .ZN(n5680) );
  NAND2_X1 U7251 ( .A1(n5671), .A2(n4705), .ZN(n5672) );
  NAND2_X1 U7252 ( .A1(n5693), .A2(n5672), .ZN(n9230) );
  OR2_X1 U7253 ( .A1(n9230), .A2(n5848), .ZN(n5678) );
  INV_X1 U7254 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7255 ( .A1(n8148), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7256 ( .A1(n5443), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5673) );
  OAI211_X1 U7257 ( .C1(n5914), .C2(n5675), .A(n5674), .B(n5673), .ZN(n5676)
         );
  INV_X1 U7258 ( .A(n5676), .ZN(n5677) );
  NAND2_X1 U7259 ( .A1(n9496), .A2(n5252), .ZN(n5679) );
  NAND2_X1 U7260 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  XNOR2_X1 U7261 ( .A(n5681), .B(n5798), .ZN(n5684) );
  AND2_X1 U7262 ( .A1(n9496), .A2(n5746), .ZN(n5682) );
  AOI21_X1 U7263 ( .B1(n9672), .B2(n5874), .A(n5682), .ZN(n5683) );
  NAND2_X1 U7264 ( .A1(n5684), .A2(n5683), .ZN(n5686) );
  OAI21_X1 U7265 ( .B1(n5684), .B2(n5683), .A(n5686), .ZN(n9224) );
  INV_X1 U7266 ( .A(n9224), .ZN(n5685) );
  INV_X1 U7267 ( .A(n5686), .ZN(n5687) );
  MUX2_X1 U7268 ( .A(n7808), .B(n10151), .S(n4612), .Z(n5709) );
  XNOR2_X1 U7269 ( .A(n5709), .B(SI_21_), .ZN(n5708) );
  NAND2_X1 U7270 ( .A1(n7805), .A2(n5327), .ZN(n5692) );
  OR2_X1 U7271 ( .A1(n8152), .A2(n10151), .ZN(n5691) );
  NAND2_X1 U7272 ( .A1(n9667), .A2(n4633), .ZN(n5702) );
  NAND2_X1 U7273 ( .A1(n5693), .A2(n9178), .ZN(n5694) );
  NAND2_X1 U7274 ( .A1(n5715), .A2(n5694), .ZN(n9470) );
  OR2_X1 U7275 ( .A1(n9470), .A2(n5848), .ZN(n5700) );
  INV_X1 U7276 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7277 ( .A1(n8148), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7278 ( .A1(n5443), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5695) );
  OAI211_X1 U7279 ( .C1(n5914), .C2(n5697), .A(n5696), .B(n5695), .ZN(n5698)
         );
  INV_X1 U7280 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7281 ( .A1(n9481), .A2(n5874), .ZN(n5701) );
  NAND2_X1 U7282 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  XNOR2_X1 U7283 ( .A(n5703), .B(n5872), .ZN(n5704) );
  AOI22_X1 U7284 ( .A1(n9667), .A2(n5874), .B1(n5746), .B2(n9481), .ZN(n5705)
         );
  XNOR2_X1 U7285 ( .A(n5704), .B(n5705), .ZN(n9176) );
  INV_X1 U7286 ( .A(n5704), .ZN(n5706) );
  NAND2_X1 U7287 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  INV_X1 U7288 ( .A(n5709), .ZN(n5710) );
  NAND2_X1 U7289 ( .A1(n5710), .A2(SI_21_), .ZN(n5750) );
  MUX2_X1 U7290 ( .A(n7942), .B(n7944), .S(n4612), .Z(n5711) );
  NAND2_X1 U7291 ( .A1(n5711), .A2(n10154), .ZN(n5755) );
  INV_X1 U7292 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7293 ( .A1(n5712), .A2(SI_22_), .ZN(n5749) );
  NAND2_X1 U7294 ( .A1(n5755), .A2(n5749), .ZN(n5726) );
  XNOR2_X1 U7295 ( .A(n5727), .B(n5726), .ZN(n7941) );
  NAND2_X1 U7296 ( .A1(n7941), .A2(n5327), .ZN(n5714) );
  OR2_X1 U7297 ( .A1(n8152), .A2(n7944), .ZN(n5713) );
  NAND2_X1 U7298 ( .A1(n5715), .A2(n10136), .ZN(n5716) );
  INV_X1 U7299 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7300 ( .A1(n5443), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7301 ( .A1(n8148), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5717) );
  OAI211_X1 U7302 ( .C1(n5914), .C2(n5719), .A(n5718), .B(n5717), .ZN(n5720)
         );
  AOI22_X1 U7303 ( .A1(n9661), .A2(n5874), .B1(n5207), .B2(n9465), .ZN(n5723)
         );
  OAI22_X1 U7304 ( .A1(n9454), .A2(n5185), .B1(n9179), .B2(n5478), .ZN(n5722)
         );
  XOR2_X1 U7305 ( .A(n5872), .B(n5722), .Z(n9248) );
  MUX2_X1 U7306 ( .A(n10107), .B(n7936), .S(n4612), .Z(n5729) );
  INV_X1 U7307 ( .A(SI_23_), .ZN(n5728) );
  NAND2_X1 U7308 ( .A1(n5729), .A2(n5728), .ZN(n5756) );
  INV_X1 U7309 ( .A(n5729), .ZN(n5730) );
  NAND2_X1 U7310 ( .A1(n5730), .A2(SI_23_), .ZN(n5731) );
  NAND2_X1 U7311 ( .A1(n5756), .A2(n5731), .ZN(n5752) );
  INV_X1 U7312 ( .A(n5752), .ZN(n5759) );
  NAND2_X1 U7313 ( .A1(n7938), .A2(n4240), .ZN(n5734) );
  OR2_X1 U7314 ( .A1(n8152), .A2(n7936), .ZN(n5733) );
  NAND2_X1 U7315 ( .A1(n9656), .A2(n4633), .ZN(n5744) );
  INV_X1 U7316 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7317 ( .A1(n5735), .A2(n9157), .ZN(n5736) );
  NAND2_X1 U7318 ( .A1(n5766), .A2(n5736), .ZN(n9436) );
  INV_X1 U7319 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7320 ( .A1(n8148), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7321 ( .A1(n5443), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U7322 ( .C1(n5914), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5740)
         );
  INV_X1 U7323 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7324 ( .A1(n9456), .A2(n5874), .ZN(n5743) );
  NAND2_X1 U7325 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  XNOR2_X1 U7326 ( .A(n5745), .B(n5872), .ZN(n9152) );
  NAND2_X1 U7327 ( .A1(n9656), .A2(n5874), .ZN(n5748) );
  NAND2_X1 U7328 ( .A1(n9456), .A2(n5746), .ZN(n5747) );
  NAND2_X1 U7329 ( .A1(n5748), .A2(n5747), .ZN(n9184) );
  NAND2_X1 U7330 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  NOR2_X1 U7331 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  INV_X1 U7332 ( .A(n5755), .ZN(n5758) );
  INV_X1 U7333 ( .A(n5756), .ZN(n5757) );
  AOI21_X1 U7334 ( .B1(n5759), .B2(n5758), .A(n5757), .ZN(n5760) );
  INV_X1 U7335 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5761) );
  MUX2_X1 U7336 ( .A(n5761), .B(n7971), .S(n4612), .Z(n5783) );
  XNOR2_X1 U7337 ( .A(n5783), .B(SI_24_), .ZN(n5781) );
  NAND2_X1 U7338 ( .A1(n7930), .A2(n5327), .ZN(n5763) );
  OR2_X1 U7339 ( .A1(n8152), .A2(n7971), .ZN(n5762) );
  NAND2_X1 U7340 ( .A1(n9652), .A2(n4633), .ZN(n5774) );
  INV_X1 U7341 ( .A(n5766), .ZN(n5764) );
  INV_X1 U7342 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7343 ( .A1(n5819), .A2(n5767), .ZN(n9423) );
  INV_X1 U7344 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7345 ( .A1(n8148), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7346 ( .A1(n5443), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5768) );
  OAI211_X1 U7347 ( .C1(n5914), .C2(n5770), .A(n5769), .B(n5768), .ZN(n5771)
         );
  INV_X1 U7348 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7349 ( .A1(n9444), .A2(n5252), .ZN(n5773) );
  NAND2_X1 U7350 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  XNOR2_X1 U7351 ( .A(n5775), .B(n5798), .ZN(n5777) );
  AND2_X1 U7352 ( .A1(n9444), .A2(n5207), .ZN(n5776) );
  AOI21_X1 U7353 ( .B1(n9652), .B2(n5874), .A(n5776), .ZN(n5778) );
  NAND2_X1 U7354 ( .A1(n5777), .A2(n5778), .ZN(n9188) );
  OAI21_X1 U7355 ( .B1(n9152), .B2(n9184), .A(n9188), .ZN(n5803) );
  INV_X1 U7356 ( .A(n9152), .ZN(n9154) );
  INV_X1 U7357 ( .A(n9184), .ZN(n9155) );
  INV_X1 U7358 ( .A(n5777), .ZN(n5780) );
  INV_X1 U7359 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U7360 ( .A1(n5780), .A2(n5779), .ZN(n9186) );
  OAI21_X1 U7361 ( .B1(n9154), .B2(n9155), .A(n9186), .ZN(n5801) );
  INV_X1 U7362 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U7363 ( .A1(n5784), .A2(SI_24_), .ZN(n5785) );
  MUX2_X1 U7364 ( .A(n8038), .B(n8471), .S(n4612), .Z(n5787) );
  NAND2_X1 U7365 ( .A1(n5787), .A2(n10178), .ZN(n5807) );
  INV_X1 U7366 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7367 ( .A1(n5788), .A2(SI_25_), .ZN(n5789) );
  NAND2_X1 U7368 ( .A1(n5807), .A2(n5789), .ZN(n5808) );
  NAND2_X1 U7369 ( .A1(n8036), .A2(n5327), .ZN(n5791) );
  OR2_X1 U7370 ( .A1(n8152), .A2(n8471), .ZN(n5790) );
  NAND2_X1 U7371 ( .A1(n9646), .A2(n4633), .ZN(n5797) );
  XNOR2_X1 U7372 ( .A(n5819), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9410) );
  INV_X1 U7373 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7374 ( .A1(n8148), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7375 ( .A1(n5443), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5792) );
  OAI211_X1 U7376 ( .C1(n5914), .C2(n5794), .A(n5793), .B(n5792), .ZN(n5795)
         );
  OR2_X1 U7377 ( .A1(n8425), .A2(n5478), .ZN(n5796) );
  NAND2_X1 U7378 ( .A1(n5797), .A2(n5796), .ZN(n5799) );
  XNOR2_X1 U7379 ( .A(n5799), .B(n5798), .ZN(n5805) );
  NOR2_X1 U7380 ( .A1(n8425), .A2(n5876), .ZN(n5800) );
  AOI21_X1 U7381 ( .B1(n9646), .B2(n5252), .A(n5800), .ZN(n5804) );
  XNOR2_X1 U7382 ( .A(n5805), .B(n5804), .ZN(n9187) );
  AOI21_X1 U7383 ( .B1(n9188), .B2(n5801), .A(n9187), .ZN(n5802) );
  NAND2_X1 U7384 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  INV_X1 U7385 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5810) );
  MUX2_X1 U7386 ( .A(n5810), .B(n8051), .S(n4612), .Z(n5812) );
  INV_X1 U7387 ( .A(SI_26_), .ZN(n5811) );
  NAND2_X1 U7388 ( .A1(n5812), .A2(n5811), .ZN(n5838) );
  INV_X1 U7389 ( .A(n5812), .ZN(n5813) );
  NAND2_X1 U7390 ( .A1(n5813), .A2(SI_26_), .ZN(n5814) );
  XNOR2_X1 U7391 ( .A(n5837), .B(n5836), .ZN(n8048) );
  NAND2_X1 U7392 ( .A1(n8048), .A2(n5327), .ZN(n5816) );
  OR2_X1 U7393 ( .A1(n8152), .A2(n8051), .ZN(n5815) );
  NAND2_X1 U7394 ( .A1(n9642), .A2(n4633), .ZN(n5828) );
  INV_X1 U7395 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9191) );
  INV_X1 U7396 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5817) );
  OAI21_X1 U7397 ( .B1(n5819), .B2(n9191), .A(n5817), .ZN(n5820) );
  NAND2_X1 U7398 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .ZN(n5818) );
  NAND2_X1 U7399 ( .A1(n9393), .A2(n5917), .ZN(n5826) );
  INV_X1 U7400 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7401 ( .A1(n5443), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7402 ( .A1(n8148), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5821) );
  OAI211_X1 U7403 ( .C1(n5914), .C2(n5823), .A(n5822), .B(n5821), .ZN(n5824)
         );
  INV_X1 U7404 ( .A(n5824), .ZN(n5825) );
  NAND2_X1 U7405 ( .A1(n9415), .A2(n5874), .ZN(n5827) );
  NAND2_X1 U7406 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  XNOR2_X1 U7407 ( .A(n5829), .B(n5872), .ZN(n5832) );
  NAND2_X1 U7408 ( .A1(n9642), .A2(n5874), .ZN(n5831) );
  NAND2_X1 U7409 ( .A1(n9415), .A2(n5207), .ZN(n5830) );
  NAND2_X1 U7410 ( .A1(n5831), .A2(n5830), .ZN(n5833) );
  NAND2_X1 U7411 ( .A1(n5832), .A2(n5833), .ZN(n9268) );
  INV_X1 U7412 ( .A(n5832), .ZN(n5835) );
  INV_X1 U7413 ( .A(n5833), .ZN(n5834) );
  NAND2_X1 U7414 ( .A1(n5835), .A2(n5834), .ZN(n9269) );
  INV_X1 U7415 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5842) );
  MUX2_X1 U7416 ( .A(n8057), .B(n5842), .S(n4612), .Z(n5839) );
  INV_X1 U7417 ( .A(SI_27_), .ZN(n10190) );
  NAND2_X1 U7418 ( .A1(n5839), .A2(n10190), .ZN(n5859) );
  INV_X1 U7419 ( .A(n5839), .ZN(n5840) );
  NAND2_X1 U7420 ( .A1(n5840), .A2(SI_27_), .ZN(n5841) );
  NAND2_X1 U7421 ( .A1(n8054), .A2(n4240), .ZN(n5844) );
  OR2_X1 U7422 ( .A1(n8152), .A2(n5842), .ZN(n5843) );
  INV_X1 U7423 ( .A(n5846), .ZN(n5845) );
  NAND2_X1 U7424 ( .A1(n5845), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5864) );
  INV_X1 U7425 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U7426 ( .A1(n5846), .A2(n10075), .ZN(n5847) );
  NAND2_X1 U7427 ( .A1(n5864), .A2(n5847), .ZN(n9382) );
  INV_X1 U7428 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7429 ( .A1(n8148), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7430 ( .A1(n5443), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5849) );
  OAI211_X1 U7431 ( .C1(n5914), .C2(n5851), .A(n5850), .B(n5849), .ZN(n5852)
         );
  INV_X1 U7432 ( .A(n5852), .ZN(n5853) );
  OAI22_X1 U7433 ( .A1(n9385), .A2(n5185), .B1(n9294), .B2(n5478), .ZN(n5855)
         );
  XOR2_X1 U7434 ( .A(n5872), .B(n5855), .Z(n9134) );
  NOR2_X1 U7435 ( .A1(n9294), .A2(n5876), .ZN(n5856) );
  AOI21_X1 U7436 ( .B1(n9634), .B2(n5252), .A(n5856), .ZN(n9133) );
  AOI21_X1 U7437 ( .B1(n9132), .B2(n9134), .A(n9133), .ZN(n5907) );
  NAND2_X1 U7438 ( .A1(n5858), .A2(n5857), .ZN(n5860) );
  INV_X1 U7439 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5861) );
  INV_X1 U7440 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8337) );
  MUX2_X1 U7441 ( .A(n5861), .B(n8337), .S(n4612), .Z(n6489) );
  XNOR2_X1 U7442 ( .A(n6489), .B(SI_28_), .ZN(n6486) );
  OR2_X1 U7443 ( .A1(n8152), .A2(n8337), .ZN(n5862) );
  NAND2_X1 U7444 ( .A1(n9628), .A2(n4633), .ZN(n5871) );
  INV_X1 U7445 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7446 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  INV_X1 U7447 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7448 ( .A1(n5443), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7449 ( .A1(n8148), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5866) );
  OAI211_X1 U7450 ( .C1(n5914), .C2(n5868), .A(n5867), .B(n5866), .ZN(n5869)
         );
  OR2_X1 U7451 ( .A1(n9376), .A2(n5478), .ZN(n5870) );
  NAND2_X1 U7452 ( .A1(n5871), .A2(n5870), .ZN(n5873) );
  XNOR2_X1 U7453 ( .A(n5873), .B(n5872), .ZN(n5878) );
  NAND2_X1 U7454 ( .A1(n9628), .A2(n5874), .ZN(n5875) );
  OAI21_X1 U7455 ( .B1(n9376), .B2(n5876), .A(n5875), .ZN(n5877) );
  NAND2_X1 U7456 ( .A1(n5879), .A2(P1_B_REG_SCAN_IN), .ZN(n5881) );
  MUX2_X1 U7457 ( .A(n5881), .B(P1_B_REG_SCAN_IN), .S(n5880), .Z(n5882) );
  INV_X1 U7458 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U7459 ( .A1(n7142), .A2(n10091), .ZN(n5885) );
  INV_X1 U7460 ( .A(n5883), .ZN(n8053) );
  NAND2_X1 U7461 ( .A1(n8053), .A2(n5879), .ZN(n5884) );
  NAND2_X1 U7462 ( .A1(n5885), .A2(n5884), .ZN(n6895) );
  INV_X1 U7463 ( .A(n6895), .ZN(n6721) );
  NOR4_X1 U7464 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5889) );
  NOR4_X1 U7465 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5888) );
  NOR4_X1 U7466 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5887) );
  NOR4_X1 U7467 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5886) );
  NAND4_X1 U7468 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n5895)
         );
  NOR2_X1 U7469 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .ZN(
        n5893) );
  NOR4_X1 U7470 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5892) );
  NOR4_X1 U7471 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5891) );
  NOR4_X1 U7472 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5890) );
  NAND4_X1 U7473 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n5894)
         );
  OAI21_X1 U7474 ( .B1(n5895), .B2(n5894), .A(n7142), .ZN(n6894) );
  NAND2_X1 U7475 ( .A1(n6721), .A2(n6894), .ZN(n7310) );
  INV_X1 U7476 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U7477 ( .A1(n7142), .A2(n7146), .ZN(n5897) );
  NAND2_X1 U7478 ( .A1(n8053), .A2(n5896), .ZN(n7144) );
  NOR2_X1 U7479 ( .A1(n7310), .A2(n7189), .ZN(n5922) );
  NAND2_X1 U7480 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7481 ( .A1(n5922), .A2(n8327), .ZN(n5908) );
  INV_X1 U7482 ( .A(n7378), .ZN(n5904) );
  INV_X1 U7483 ( .A(n9278), .ZN(n5905) );
  NAND2_X1 U7484 ( .A1(n4270), .A2(n5905), .ZN(n5906) );
  NOR2_X1 U7485 ( .A1(n4270), .A2(n9278), .ZN(n5933) );
  NAND2_X1 U7486 ( .A1(n5907), .A2(n5933), .ZN(n5936) );
  INV_X1 U7487 ( .A(n5908), .ZN(n5918) );
  OR2_X1 U7488 ( .A1(n7378), .A2(n8287), .ZN(n10208) );
  NAND2_X1 U7489 ( .A1(n5918), .A2(n7315), .ZN(n5910) );
  NAND2_X1 U7490 ( .A1(n8327), .A2(n10220), .ZN(n5909) );
  INV_X1 U7491 ( .A(n5911), .ZN(n8431) );
  INV_X1 U7492 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7493 ( .A1(n8148), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7494 ( .A1(n5443), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5912) );
  OAI211_X1 U7495 ( .C1(n5915), .C2(n5914), .A(n5913), .B(n5912), .ZN(n5916)
         );
  AOI21_X1 U7496 ( .B1(n8431), .B2(n5917), .A(n5916), .ZN(n9292) );
  NAND2_X1 U7497 ( .A1(n5918), .A2(n8328), .ZN(n5921) );
  INV_X1 U7498 ( .A(n8336), .ZN(n6874) );
  NOR2_X1 U7499 ( .A1(n9292), .A2(n9275), .ZN(n5930) );
  AND3_X1 U7500 ( .A1(n5898), .A2(n6867), .A3(n7934), .ZN(n5923) );
  INV_X1 U7501 ( .A(n5922), .ZN(n5926) );
  NAND2_X1 U7502 ( .A1(n5926), .A2(n9947), .ZN(n6868) );
  NAND2_X1 U7503 ( .A1(n5923), .A2(n6868), .ZN(n5924) );
  NAND2_X1 U7504 ( .A1(n5924), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5927) );
  AND2_X1 U7505 ( .A1(n7315), .A2(n8327), .ZN(n5925) );
  NAND2_X1 U7506 ( .A1(n5926), .A2(n5925), .ZN(n6869) );
  AOI22_X1 U7507 ( .A1(n9361), .A2(n9271), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5928) );
  OAI21_X1 U7508 ( .B1(n9294), .B2(n9282), .A(n5928), .ZN(n5929) );
  AOI211_X1 U7509 ( .C1(n9628), .C2(n9288), .A(n5930), .B(n5929), .ZN(n5931)
         );
  INV_X1 U7510 ( .A(n5931), .ZN(n5932) );
  AOI21_X1 U7511 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(n5935) );
  NAND3_X1 U7512 ( .A1(n5937), .A2(n5936), .A3(n5935), .ZN(P1_U3218) );
  NOR2_X1 U7513 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5944) );
  NOR2_X1 U7514 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5945) );
  NAND2_X1 U7515 ( .A1(n6168), .A2(n6205), .ZN(n5953) );
  NOR2_X1 U7516 ( .A1(n5953), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5949) );
  NAND3_X1 U7517 ( .A1(n5947), .A2(n5946), .A3(n6119), .ZN(n5954) );
  INV_X1 U7518 ( .A(n5954), .ZN(n5948) );
  NAND2_X1 U7519 ( .A1(n7930), .A2(n6249), .ZN(n5952) );
  NAND2_X1 U7520 ( .A1(n4237), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7521 ( .A1(n6441), .A2(n4769), .ZN(n7240) );
  NAND2_X1 U7522 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7523 ( .A1(n5984), .A2(n6563), .ZN(n7626) );
  XNOR2_X1 U7524 ( .A(n9007), .B(n6406), .ZN(n8555) );
  NAND2_X1 U7525 ( .A1(n5967), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7526 ( .A1(n5969), .A2(n5968), .ZN(n6192) );
  NAND2_X1 U7527 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n5970) );
  INV_X1 U7528 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8498) );
  XNOR2_X1 U7529 ( .A(n6357), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8785) );
  NAND3_X1 U7530 ( .A1(n5974), .A2(n5973), .A3(n5972), .ZN(n5975) );
  NAND2_X1 U7531 ( .A1(n8785), .A2(n6465), .ZN(n5983) );
  INV_X1 U7532 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8788) );
  INV_X2 U7533 ( .A(n6025), .ZN(n6399) );
  NAND2_X1 U7534 ( .A1(n6399), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7535 ( .A1(n6024), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5979) );
  OAI211_X1 U7536 ( .C1(n8788), .C2(n6009), .A(n5980), .B(n5979), .ZN(n5981)
         );
  INV_X1 U7537 ( .A(n5981), .ZN(n5982) );
  NAND2_X1 U7538 ( .A1(n5099), .A2(n6331), .ZN(n8559) );
  INV_X1 U7539 ( .A(n6728), .ZN(n5985) );
  NAND2_X1 U7540 ( .A1(n6037), .A2(n5985), .ZN(n5989) );
  NAND2_X1 U7541 ( .A1(n6040), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7542 ( .A1(n6018), .A2(n9120), .ZN(n5986) );
  XNOR2_X1 U7543 ( .A(n5986), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6923) );
  INV_X1 U7544 ( .A(n6923), .ZN(n5987) );
  NAND2_X1 U7545 ( .A1(n6024), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5993) );
  INV_X1 U7546 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8966) );
  OR2_X1 U7547 ( .A1(n6010), .A2(n8966), .ZN(n5992) );
  INV_X1 U7548 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8971) );
  OR2_X1 U7549 ( .A1(n6009), .A2(n8971), .ZN(n5991) );
  INV_X1 U7550 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6914) );
  NAND4_X2 U7551 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n6468)
         );
  NAND2_X1 U7552 ( .A1(n6331), .A2(n6468), .ZN(n8590) );
  NAND2_X1 U7553 ( .A1(n4238), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7554 ( .A1(n5994), .A2(n7040), .ZN(n5995) );
  INV_X1 U7555 ( .A(n6730), .ZN(n5997) );
  NAND2_X1 U7556 ( .A1(n6037), .A2(n5997), .ZN(n5998) );
  XNOR2_X1 U7557 ( .A(n6077), .B(n7509), .ZN(n8598) );
  NOR2_X1 U7558 ( .A1(n4612), .A2(n5999), .ZN(n6001) );
  INV_X1 U7559 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7560 ( .A(n6001), .B(n6000), .ZN(n9131) );
  MUX2_X1 U7561 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9131), .S(n6910), .Z(n7736) );
  OR2_X1 U7562 ( .A1(n6077), .A2(n7736), .ZN(n6008) );
  NAND2_X1 U7563 ( .A1(n6024), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6007) );
  INV_X1 U7564 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7565 ( .A1(n4234), .A2(n6002), .ZN(n6006) );
  INV_X1 U7566 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6003) );
  OR2_X1 U7567 ( .A1(n6009), .A2(n6003), .ZN(n6005) );
  INV_X1 U7568 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6913) );
  OR2_X1 U7569 ( .A1(n6025), .A2(n6913), .ZN(n6004) );
  AND2_X1 U7570 ( .A1(n6469), .A2(n7736), .ZN(n7279) );
  NAND2_X1 U7571 ( .A1(n6331), .A2(n7279), .ZN(n7511) );
  NAND2_X1 U7572 ( .A1(n6024), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6013) );
  INV_X1 U7573 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6921) );
  OR2_X1 U7574 ( .A1(n6009), .A2(n6921), .ZN(n6012) );
  INV_X1 U7575 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7756) );
  INV_X1 U7576 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6011) );
  INV_X1 U7577 ( .A(n6715), .ZN(n6016) );
  NAND2_X1 U7578 ( .A1(n6016), .A2(n6037), .ZN(n6023) );
  NAND2_X1 U7579 ( .A1(n6038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U7580 ( .A(n6019), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6925) );
  INV_X1 U7581 ( .A(n6925), .ZN(n6020) );
  INV_X1 U7582 ( .A(n6021), .ZN(n6022) );
  NAND2_X1 U7583 ( .A1(n6024), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6029) );
  OR2_X1 U7584 ( .A1(n4234), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6028) );
  INV_X1 U7585 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8958) );
  OR2_X1 U7586 ( .A1(n6009), .A2(n8958), .ZN(n6027) );
  INV_X1 U7587 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6915) );
  OR2_X1 U7588 ( .A1(n6025), .A2(n6915), .ZN(n6026) );
  NAND2_X1 U7589 ( .A1(n6331), .A2(n8659), .ZN(n6033) );
  XNOR2_X1 U7590 ( .A(n6032), .B(n6033), .ZN(n8383) );
  INV_X1 U7591 ( .A(n8383), .ZN(n6030) );
  NAND2_X1 U7592 ( .A1(n6031), .A2(n6030), .ZN(n8386) );
  INV_X1 U7593 ( .A(n6032), .ZN(n6035) );
  INV_X1 U7594 ( .A(n6033), .ZN(n6034) );
  NAND2_X1 U7595 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7596 ( .A1(n6052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6039) );
  XNOR2_X1 U7597 ( .A(n6039), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7598 ( .A1(n4238), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n5994), .B2(
        n6953), .ZN(n6041) );
  NAND2_X1 U7599 ( .A1(n6042), .A2(n6041), .ZN(n7746) );
  XNOR2_X1 U7600 ( .A(n6077), .B(n7746), .ZN(n8373) );
  INV_X1 U7601 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7602 ( .A1(n6327), .A2(n6043), .ZN(n6048) );
  NAND2_X1 U7603 ( .A1(n6399), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7604 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8377) );
  OR2_X1 U7605 ( .A1(n4234), .A2(n8377), .ZN(n6046) );
  INV_X1 U7606 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6044) );
  OR2_X1 U7607 ( .A1(n6009), .A2(n6044), .ZN(n6045) );
  AND2_X1 U7608 ( .A1(n6331), .A2(n8658), .ZN(n6049) );
  AND2_X1 U7609 ( .A1(n8373), .A2(n6049), .ZN(n8368) );
  INV_X1 U7610 ( .A(n8373), .ZN(n6051) );
  INV_X1 U7611 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7612 ( .A1(n6051), .A2(n6050), .ZN(n8371) );
  NAND2_X1 U7613 ( .A1(n6704), .A2(n6249), .ZN(n6056) );
  INV_X1 U7614 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7615 ( .A1(n6071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6054) );
  XNOR2_X1 U7616 ( .A(n6054), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7617 ( .A1(n4237), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5994), .B2(
        n6982), .ZN(n6055) );
  XNOR2_X1 U7618 ( .A(n6077), .B(n7591), .ZN(n6065) );
  NAND2_X1 U7619 ( .A1(n6024), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6064) );
  INV_X1 U7620 ( .A(n6057), .ZN(n6059) );
  INV_X1 U7621 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7622 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7623 ( .A1(n6079), .A2(n6060), .ZN(n9989) );
  OR2_X1 U7624 ( .A1(n4234), .A2(n9989), .ZN(n6063) );
  INV_X1 U7625 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6952) );
  OR2_X1 U7626 ( .A1(n6009), .A2(n6952), .ZN(n6062) );
  INV_X1 U7627 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6944) );
  OR2_X1 U7628 ( .A1(n6025), .A2(n6944), .ZN(n6061) );
  NAND4_X1 U7629 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n8657)
         );
  NAND2_X1 U7630 ( .A1(n6331), .A2(n8657), .ZN(n6066) );
  NAND2_X1 U7631 ( .A1(n6065), .A2(n6066), .ZN(n6070) );
  INV_X1 U7632 ( .A(n6065), .ZN(n6068) );
  INV_X1 U7633 ( .A(n6066), .ZN(n6067) );
  NAND2_X1 U7634 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  AND2_X1 U7635 ( .A1(n6070), .A2(n6069), .ZN(n7589) );
  NAND2_X1 U7636 ( .A1(n7588), .A2(n7589), .ZN(n7587) );
  NAND2_X1 U7637 ( .A1(n6711), .A2(n6249), .ZN(n6076) );
  INV_X1 U7638 ( .A(n6071), .ZN(n6073) );
  INV_X1 U7639 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7640 ( .A1(n6073), .A2(n6072), .ZN(n6089) );
  NAND2_X1 U7641 ( .A1(n6089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U7642 ( .A(n6074), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U7643 ( .A1(n4238), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5994), .B2(
        n6985), .ZN(n6075) );
  NAND2_X1 U7644 ( .A1(n6076), .A2(n6075), .ZN(n7711) );
  XNOR2_X1 U7645 ( .A(n7711), .B(n6077), .ZN(n6086) );
  NAND2_X1 U7646 ( .A1(n6024), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6084) );
  INV_X1 U7647 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6974) );
  OR2_X1 U7648 ( .A1(n6025), .A2(n6974), .ZN(n6083) );
  INV_X1 U7649 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7650 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7651 ( .A1(n6093), .A2(n6080), .ZN(n7705) );
  OR2_X1 U7652 ( .A1(n4234), .A2(n7705), .ZN(n6082) );
  INV_X1 U7653 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7706) );
  OR2_X1 U7654 ( .A1(n6009), .A2(n7706), .ZN(n6081) );
  NAND4_X1 U7655 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n8656)
         );
  NAND2_X1 U7656 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  NAND2_X1 U7657 ( .A1(n6723), .A2(n6249), .ZN(n6091) );
  AOI22_X1 U7658 ( .A1(n4237), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7010), .B2(
        n5994), .ZN(n6090) );
  NAND2_X1 U7659 ( .A1(n6091), .A2(n6090), .ZN(n7631) );
  XNOR2_X1 U7660 ( .A(n7631), .B(n6406), .ZN(n6099) );
  NAND2_X1 U7661 ( .A1(n6024), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6098) );
  INV_X1 U7662 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6976) );
  OR2_X1 U7663 ( .A1(n6025), .A2(n6976), .ZN(n6097) );
  INV_X1 U7664 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7665 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NAND2_X1 U7666 ( .A1(n6107), .A2(n6094), .ZN(n7620) );
  OR2_X1 U7667 ( .A1(n4234), .A2(n7620), .ZN(n6096) );
  INV_X1 U7668 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7621) );
  OR2_X1 U7669 ( .A1(n6009), .A2(n7621), .ZN(n6095) );
  NAND4_X1 U7670 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n8655)
         );
  NAND2_X1 U7671 ( .A1(n6331), .A2(n8655), .ZN(n6100) );
  XNOR2_X1 U7672 ( .A(n6099), .B(n6100), .ZN(n7525) );
  INV_X1 U7673 ( .A(n6099), .ZN(n6102) );
  INV_X1 U7674 ( .A(n6100), .ZN(n6101) );
  NAND2_X1 U7675 ( .A1(n6732), .A2(n6249), .ZN(n6106) );
  NAND2_X1 U7676 ( .A1(n6118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6104) );
  XNOR2_X1 U7677 ( .A(n6104), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7054) );
  AOI22_X1 U7678 ( .A1(n7054), .A2(n5994), .B1(n4238), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7679 ( .A1(n6106), .A2(n6105), .ZN(n9089) );
  XNOR2_X1 U7680 ( .A(n9089), .B(n6077), .ZN(n6116) );
  NAND2_X1 U7681 ( .A1(n6024), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6113) );
  INV_X1 U7682 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7644) );
  OR2_X1 U7683 ( .A1(n6009), .A2(n7644), .ZN(n6112) );
  NAND2_X1 U7684 ( .A1(n6107), .A2(n7573), .ZN(n6108) );
  NAND2_X1 U7685 ( .A1(n6125), .A2(n6108), .ZN(n7643) );
  OR2_X1 U7686 ( .A1(n4234), .A2(n7643), .ZN(n6111) );
  INV_X1 U7687 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7688 ( .A1(n6025), .A2(n6109), .ZN(n6110) );
  NAND4_X1 U7689 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n8654)
         );
  NAND2_X1 U7690 ( .A1(n6331), .A2(n8654), .ZN(n6114) );
  XNOR2_X1 U7691 ( .A(n6116), .B(n6114), .ZN(n7571) );
  INV_X1 U7692 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7693 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7694 ( .A1(n6740), .A2(n6249), .ZN(n6123) );
  INV_X1 U7695 ( .A(n6118), .ZN(n6120) );
  NAND2_X1 U7696 ( .A1(n6120), .A2(n6119), .ZN(n6138) );
  NAND2_X1 U7697 ( .A1(n6138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7698 ( .A(n6121), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7057) );
  AOI22_X1 U7699 ( .A1(n7057), .A2(n5994), .B1(n4237), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7700 ( .A1(n6123), .A2(n6122), .ZN(n9083) );
  XNOR2_X1 U7701 ( .A(n9083), .B(n6406), .ZN(n6131) );
  NAND2_X1 U7702 ( .A1(n6024), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7703 ( .A1(n6399), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6129) );
  INV_X1 U7704 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7705 ( .A1(n6125), .A2(n6124), .ZN(n6126) );
  NAND2_X1 U7706 ( .A1(n6142), .A2(n6126), .ZN(n7824) );
  OR2_X1 U7707 ( .A1(n4234), .A2(n7824), .ZN(n6128) );
  INV_X1 U7708 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7662) );
  OR2_X1 U7709 ( .A1(n6009), .A2(n7662), .ZN(n6127) );
  NAND4_X1 U7710 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n8653)
         );
  NAND2_X1 U7711 ( .A1(n6331), .A2(n8653), .ZN(n6132) );
  NAND2_X1 U7712 ( .A1(n6131), .A2(n6132), .ZN(n6137) );
  INV_X1 U7713 ( .A(n6131), .ZN(n6134) );
  INV_X1 U7714 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7715 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  NAND2_X1 U7716 ( .A1(n6137), .A2(n6135), .ZN(n7822) );
  INV_X1 U7717 ( .A(n6138), .ZN(n6140) );
  INV_X1 U7718 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7719 ( .A1(n6140), .A2(n6139), .ZN(n6171) );
  NAND2_X1 U7720 ( .A1(n6171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6154) );
  XNOR2_X1 U7721 ( .A(n6154), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U7722 ( .A1(n7059), .A2(n5994), .B1(n4237), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7723 ( .A(n9077), .B(n6406), .ZN(n6149) );
  NAND2_X1 U7724 ( .A1(n6024), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6148) );
  INV_X1 U7725 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7673) );
  OR2_X1 U7726 ( .A1(n6009), .A2(n7673), .ZN(n6147) );
  NAND2_X1 U7727 ( .A1(n6142), .A2(n7132), .ZN(n6143) );
  NAND2_X1 U7728 ( .A1(n6177), .A2(n6143), .ZN(n7859) );
  OR2_X1 U7729 ( .A1(n4234), .A2(n7859), .ZN(n6146) );
  INV_X1 U7730 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6144) );
  OR2_X1 U7731 ( .A1(n6025), .A2(n6144), .ZN(n6145) );
  NAND4_X1 U7732 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n8652)
         );
  NAND2_X1 U7733 ( .A1(n6331), .A2(n8652), .ZN(n6150) );
  XNOR2_X1 U7734 ( .A(n6149), .B(n6150), .ZN(n7856) );
  INV_X1 U7735 ( .A(n6149), .ZN(n6152) );
  INV_X1 U7736 ( .A(n6150), .ZN(n6151) );
  NAND2_X1 U7737 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  NAND2_X1 U7738 ( .A1(n6745), .A2(n6249), .ZN(n6158) );
  NAND2_X1 U7739 ( .A1(n6154), .A2(n6168), .ZN(n6155) );
  NAND2_X1 U7740 ( .A1(n6155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7741 ( .A(n6156), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7060) );
  AOI22_X1 U7742 ( .A1(n7060), .A2(n5994), .B1(n4238), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7743 ( .A1(n6158), .A2(n6157), .ZN(n9072) );
  XNOR2_X1 U7744 ( .A(n9072), .B(n6077), .ZN(n6165) );
  INV_X1 U7745 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U7746 ( .A(n6177), .B(n6176), .ZN(n7991) );
  OR2_X1 U7747 ( .A1(n4234), .A2(n7991), .ZN(n6162) );
  NAND2_X1 U7748 ( .A1(n6024), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6161) );
  INV_X1 U7749 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7049) );
  OR2_X1 U7750 ( .A1(n6025), .A2(n7049), .ZN(n6160) );
  INV_X1 U7751 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7752 ( .A1(n6009), .A2(n7813), .ZN(n6159) );
  NAND4_X1 U7753 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n8651)
         );
  NAND2_X1 U7754 ( .A1(n6331), .A2(n8651), .ZN(n6163) );
  XNOR2_X1 U7755 ( .A(n6165), .B(n6163), .ZN(n7987) );
  NAND2_X1 U7756 ( .A1(n7988), .A2(n7987), .ZN(n6167) );
  INV_X1 U7757 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7758 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NAND2_X1 U7759 ( .A1(n6167), .A2(n6166), .ZN(n8026) );
  NAND2_X1 U7760 ( .A1(n6755), .A2(n6249), .ZN(n6174) );
  INV_X1 U7761 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7762 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7763 ( .A1(n6188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6172) );
  XNOR2_X1 U7764 ( .A(n6172), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U7765 ( .A1(n7061), .A2(n5994), .B1(n4238), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7766 ( .A1(n6174), .A2(n6173), .ZN(n8033) );
  XNOR2_X1 U7767 ( .A(n8033), .B(n6406), .ZN(n6183) );
  NAND2_X1 U7768 ( .A1(n6399), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6182) );
  INV_X1 U7769 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8004) );
  OR2_X1 U7770 ( .A1(n6327), .A2(n8004), .ZN(n6181) );
  INV_X1 U7771 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6175) );
  OAI21_X1 U7772 ( .B1(n6177), .B2(n6176), .A(n6175), .ZN(n6178) );
  NAND2_X1 U7773 ( .A1(n6178), .A2(n6192), .ZN(n8029) );
  OR2_X1 U7774 ( .A1(n4234), .A2(n8029), .ZN(n6180) );
  INV_X1 U7775 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7877) );
  OR2_X1 U7776 ( .A1(n6009), .A2(n7877), .ZN(n6179) );
  NAND4_X1 U7777 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n8650)
         );
  NAND2_X1 U7778 ( .A1(n6331), .A2(n8650), .ZN(n6184) );
  NAND2_X1 U7779 ( .A1(n6183), .A2(n6184), .ZN(n8024) );
  NAND2_X1 U7780 ( .A1(n8026), .A2(n8024), .ZN(n6187) );
  INV_X1 U7781 ( .A(n6183), .ZN(n6186) );
  INV_X1 U7782 ( .A(n6184), .ZN(n6185) );
  NAND2_X1 U7783 ( .A1(n6186), .A2(n6185), .ZN(n8025) );
  NAND2_X1 U7784 ( .A1(n6761), .A2(n6249), .ZN(n6191) );
  OAI21_X1 U7785 ( .B1(n6188), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U7786 ( .A(n6203), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7152) );
  NOR2_X1 U7787 ( .A1(n6239), .A2(n10105), .ZN(n6189) );
  AOI21_X1 U7788 ( .B1(n7152), .B2(n5994), .A(n6189), .ZN(n6190) );
  XNOR2_X1 U7789 ( .A(n9066), .B(n6077), .ZN(n6198) );
  NAND2_X1 U7790 ( .A1(n6192), .A2(n7159), .ZN(n6193) );
  NAND2_X1 U7791 ( .A1(n6231), .A2(n6193), .ZN(n7950) );
  OR2_X1 U7792 ( .A1(n7950), .A2(n4234), .ZN(n6197) );
  NAND2_X1 U7793 ( .A1(n6399), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7794 ( .A1(n6024), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6195) );
  INV_X1 U7795 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7264) );
  OR2_X1 U7796 ( .A1(n6009), .A2(n7264), .ZN(n6194) );
  NAND4_X1 U7797 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n8649)
         );
  AND2_X1 U7798 ( .A1(n6331), .A2(n8649), .ZN(n6199) );
  NAND2_X1 U7799 ( .A1(n6198), .A2(n6199), .ZN(n6215) );
  INV_X1 U7800 ( .A(n6198), .ZN(n8484) );
  INV_X1 U7801 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7802 ( .A1(n8484), .A2(n6200), .ZN(n6201) );
  AND2_X1 U7803 ( .A1(n6215), .A2(n6201), .ZN(n8040) );
  NAND2_X1 U7804 ( .A1(n6829), .A2(n6249), .ZN(n6209) );
  INV_X1 U7805 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7806 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U7807 ( .A1(n6204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7808 ( .A1(n6206), .A2(n6205), .ZN(n6237) );
  OR2_X1 U7809 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  AOI22_X1 U7810 ( .A1(n7693), .A2(n5994), .B1(n4238), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6208) );
  XNOR2_X1 U7811 ( .A(n9061), .B(n6077), .ZN(n6217) );
  XNOR2_X1 U7812 ( .A(n6231), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U7813 ( .A1(n8015), .A2(n6465), .ZN(n6214) );
  INV_X1 U7814 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U7815 ( .A1(n6024), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6211) );
  INV_X1 U7816 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7267) );
  OR2_X1 U7817 ( .A1(n6025), .A2(n7267), .ZN(n6210) );
  OAI211_X1 U7818 ( .C1(n8016), .C2(n6009), .A(n6211), .B(n6210), .ZN(n6212)
         );
  INV_X1 U7819 ( .A(n6212), .ZN(n6213) );
  NAND2_X1 U7820 ( .A1(n6214), .A2(n6213), .ZN(n8648) );
  NAND2_X1 U7821 ( .A1(n6331), .A2(n8648), .ZN(n6218) );
  XNOR2_X1 U7822 ( .A(n6217), .B(n6218), .ZN(n8493) );
  AND2_X1 U7823 ( .A1(n8493), .A2(n6215), .ZN(n6216) );
  INV_X1 U7824 ( .A(n6217), .ZN(n6219) );
  NAND2_X1 U7825 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7826 ( .A1(n7193), .A2(n6249), .ZN(n6224) );
  NAND2_X1 U7827 ( .A1(n6221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  XNOR2_X1 U7828 ( .A(n6222), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8667) );
  AOI22_X1 U7829 ( .A1(n4237), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5994), .B2(
        n8667), .ZN(n6223) );
  NAND2_X2 U7830 ( .A1(n6224), .A2(n6223), .ZN(n9050) );
  XNOR2_X1 U7831 ( .A(n9050), .B(n6077), .ZN(n8533) );
  INV_X1 U7832 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10063) );
  INV_X1 U7833 ( .A(n6225), .ZN(n6232) );
  INV_X1 U7834 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U7835 ( .A1(n6232), .A2(n8536), .ZN(n6226) );
  NAND2_X1 U7836 ( .A1(n6268), .A2(n6226), .ZN(n8922) );
  OR2_X1 U7837 ( .A1(n8922), .A2(n4234), .ZN(n6228) );
  AOI22_X1 U7838 ( .A1(n6024), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n6399), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6227) );
  OAI211_X1 U7839 ( .C1(n6009), .C2(n10063), .A(n6228), .B(n6227), .ZN(n8647)
         );
  AND2_X1 U7840 ( .A1(n8647), .A2(n6331), .ZN(n6245) );
  INV_X1 U7841 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6236) );
  INV_X1 U7842 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6230) );
  INV_X1 U7843 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6229) );
  OAI21_X1 U7844 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(n6233) );
  AND2_X1 U7845 ( .A1(n6233), .A2(n6232), .ZN(n8945) );
  NAND2_X1 U7846 ( .A1(n8945), .A2(n6465), .ZN(n6235) );
  AOI22_X1 U7847 ( .A1(n6024), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n6399), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n6234) );
  OAI211_X1 U7848 ( .C1(n6009), .C2(n6236), .A(n6235), .B(n6234), .ZN(n8913)
         );
  AND2_X1 U7849 ( .A1(n6331), .A2(n8913), .ZN(n6244) );
  NAND2_X1 U7850 ( .A1(n7091), .A2(n6249), .ZN(n6242) );
  NAND2_X1 U7851 ( .A1(n6237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  XNOR2_X1 U7852 ( .A(n6238), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7911) );
  NOR2_X1 U7853 ( .A1(n6239), .A2(n10064), .ZN(n6240) );
  AOI21_X1 U7854 ( .B1(n7911), .B2(n5994), .A(n6240), .ZN(n6241) );
  XNOR2_X1 U7855 ( .A(n9056), .B(n6077), .ZN(n8529) );
  AOI22_X1 U7856 ( .A1(n8533), .A2(n6245), .B1(n6244), .B2(n8529), .ZN(n6243)
         );
  INV_X1 U7857 ( .A(n8533), .ZN(n6247) );
  OAI21_X1 U7858 ( .B1(n8529), .B2(n6244), .A(n6245), .ZN(n6246) );
  INV_X1 U7859 ( .A(n8529), .ZN(n8531) );
  INV_X1 U7860 ( .A(n6244), .ZN(n8630) );
  INV_X1 U7861 ( .A(n6245), .ZN(n8532) );
  AOI21_X1 U7862 ( .B1(n6247), .B2(n6246), .A(n5118), .ZN(n6248) );
  NAND2_X1 U7863 ( .A1(n7204), .A2(n6249), .ZN(n6253) );
  NAND2_X1 U7864 ( .A1(n6250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6251) );
  XNOR2_X1 U7865 ( .A(n6251), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8678) );
  AOI22_X1 U7866 ( .A1(n4238), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5994), .B2(
        n8678), .ZN(n6252) );
  XNOR2_X1 U7867 ( .A(n9045), .B(n6077), .ZN(n6259) );
  XNOR2_X1 U7868 ( .A(n6268), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U7869 ( .A1(n8904), .A2(n6465), .ZN(n6258) );
  INV_X1 U7870 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8685) );
  INV_X1 U7871 ( .A(n6009), .ZN(n6460) );
  NAND2_X1 U7872 ( .A1(n6460), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7873 ( .A1(n6024), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6254) );
  OAI211_X1 U7874 ( .C1(n6025), .C2(n8685), .A(n6255), .B(n6254), .ZN(n6256)
         );
  INV_X1 U7875 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7876 ( .A1(n6258), .A2(n6257), .ZN(n8915) );
  AND2_X1 U7877 ( .A1(n8915), .A2(n6331), .ZN(n6260) );
  NAND2_X1 U7878 ( .A1(n6259), .A2(n6260), .ZN(n6263) );
  INV_X1 U7879 ( .A(n6259), .ZN(n8609) );
  INV_X1 U7880 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7881 ( .A1(n8609), .A2(n6261), .ZN(n6262) );
  NAND2_X1 U7882 ( .A1(n6263), .A2(n6262), .ZN(n8542) );
  NAND2_X1 U7883 ( .A1(n4319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7884 ( .A(n6264), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8681) );
  AOI22_X1 U7885 ( .A1(n4237), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8681), .B2(
        n5994), .ZN(n6265) );
  XNOR2_X1 U7886 ( .A(n9039), .B(n6077), .ZN(n8394) );
  OAI21_X1 U7887 ( .B1(n6268), .B2(n8547), .A(n6267), .ZN(n6269) );
  NAND2_X1 U7888 ( .A1(n6269), .A2(n6283), .ZN(n8885) );
  OR2_X1 U7889 ( .A1(n8885), .A2(n4234), .ZN(n6275) );
  INV_X1 U7890 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7891 ( .A1(n6399), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7892 ( .A1(n6024), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U7893 ( .C1(n6272), .C2(n6009), .A(n6271), .B(n6270), .ZN(n6273)
         );
  INV_X1 U7894 ( .A(n6273), .ZN(n6274) );
  NAND2_X1 U7895 ( .A1(n6275), .A2(n6274), .ZN(n8646) );
  AND2_X1 U7896 ( .A1(n8646), .A2(n6331), .ZN(n6276) );
  NAND2_X1 U7897 ( .A1(n8394), .A2(n6276), .ZN(n6290) );
  INV_X1 U7898 ( .A(n8394), .ZN(n6278) );
  INV_X1 U7899 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7900 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  AND2_X1 U7901 ( .A1(n6290), .A2(n6279), .ZN(n8606) );
  AOI22_X1 U7902 ( .A1(n4769), .A2(n5994), .B1(n4238), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7903 ( .A(n9034), .B(n6077), .ZN(n6316) );
  INV_X1 U7904 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U7905 ( .A1(n6283), .A2(n10181), .ZN(n6284) );
  NAND2_X1 U7906 ( .A1(n6295), .A2(n6284), .ZN(n8872) );
  OR2_X1 U7907 ( .A1(n8872), .A2(n4234), .ZN(n6289) );
  INV_X1 U7908 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U7909 ( .A1(n6399), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7910 ( .A1(n6024), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6285) );
  OAI211_X1 U7911 ( .C1(n8873), .C2(n6009), .A(n6286), .B(n6285), .ZN(n6287)
         );
  INV_X1 U7912 ( .A(n6287), .ZN(n6288) );
  NAND2_X1 U7913 ( .A1(n6289), .A2(n6288), .ZN(n8846) );
  NAND2_X1 U7914 ( .A1(n8846), .A2(n6331), .ZN(n6317) );
  XNOR2_X1 U7915 ( .A(n6316), .B(n6317), .ZN(n8396) );
  AND2_X1 U7916 ( .A1(n8396), .A2(n6290), .ZN(n6291) );
  NAND2_X1 U7917 ( .A1(n4237), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U7918 ( .A(n9029), .B(n6077), .ZN(n6302) );
  NAND2_X1 U7919 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  AND2_X1 U7920 ( .A1(n6309), .A2(n6296), .ZN(n8850) );
  NAND2_X1 U7921 ( .A1(n8850), .A2(n6465), .ZN(n6301) );
  INV_X1 U7922 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U7923 ( .A1(n6399), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7924 ( .A1(n6460), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6297) );
  OAI211_X1 U7925 ( .C1(n6327), .C2(n10148), .A(n6298), .B(n6297), .ZN(n6299)
         );
  INV_X1 U7926 ( .A(n6299), .ZN(n6300) );
  NAND2_X1 U7927 ( .A1(n6301), .A2(n6300), .ZN(n8830) );
  AND2_X1 U7928 ( .A1(n8830), .A2(n6331), .ZN(n6303) );
  NAND2_X1 U7929 ( .A1(n6302), .A2(n6303), .ZN(n6320) );
  INV_X1 U7930 ( .A(n6302), .ZN(n8507) );
  INV_X1 U7931 ( .A(n6303), .ZN(n6304) );
  NAND2_X1 U7932 ( .A1(n8507), .A2(n6304), .ZN(n6305) );
  NAND2_X1 U7933 ( .A1(n6320), .A2(n6305), .ZN(n8569) );
  NAND2_X1 U7934 ( .A1(n4237), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6306) );
  INV_X1 U7935 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7936 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U7937 ( .A1(n6323), .A2(n6310), .ZN(n8833) );
  OR2_X1 U7938 ( .A1(n8833), .A2(n4234), .ZN(n6315) );
  INV_X1 U7939 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8834) );
  NAND2_X1 U7940 ( .A1(n6399), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7941 ( .A1(n6024), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6311) );
  OAI211_X1 U7942 ( .C1(n8834), .C2(n6009), .A(n6312), .B(n6311), .ZN(n6313)
         );
  INV_X1 U7943 ( .A(n6313), .ZN(n6314) );
  NAND2_X1 U7944 ( .A1(n6315), .A2(n6314), .ZN(n8847) );
  INV_X1 U7945 ( .A(n6316), .ZN(n6318) );
  NAND2_X1 U7946 ( .A1(n6318), .A2(n6317), .ZN(n8504) );
  OR2_X1 U7947 ( .A1(n8506), .A2(n6320), .ZN(n8508) );
  NAND2_X1 U7948 ( .A1(n4238), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6321) );
  XNOR2_X1 U7949 ( .A(n9019), .B(n6077), .ZN(n6335) );
  NAND2_X1 U7950 ( .A1(n6323), .A2(n8582), .ZN(n6324) );
  NAND2_X1 U7951 ( .A1(n4262), .A2(n6324), .ZN(n8816) );
  OR2_X1 U7952 ( .A1(n8816), .A2(n4234), .ZN(n6330) );
  INV_X1 U7953 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10182) );
  NAND2_X1 U7954 ( .A1(n6399), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7955 ( .A1(n6460), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U7956 ( .C1(n6327), .C2(n10182), .A(n6326), .B(n6325), .ZN(n6328)
         );
  INV_X1 U7957 ( .A(n6328), .ZN(n6329) );
  NAND2_X1 U7958 ( .A1(n6330), .A2(n6329), .ZN(n8831) );
  AND2_X1 U7959 ( .A1(n8831), .A2(n6331), .ZN(n6336) );
  AND2_X1 U7960 ( .A1(n6332), .A2(n4285), .ZN(n8574) );
  AOI21_X1 U7961 ( .B1(n6335), .B2(n6336), .A(n8574), .ZN(n6333) );
  AND2_X1 U7962 ( .A1(n8508), .A2(n6333), .ZN(n6334) );
  INV_X1 U7963 ( .A(n6335), .ZN(n8577) );
  INV_X1 U7964 ( .A(n6336), .ZN(n8579) );
  NAND2_X1 U7965 ( .A1(n4238), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6337) );
  XNOR2_X1 U7966 ( .A(n9012), .B(n6077), .ZN(n6347) );
  NAND2_X1 U7967 ( .A1(n4262), .A2(n8498), .ZN(n6338) );
  AND2_X1 U7968 ( .A1(n6357), .A2(n6338), .ZN(n8799) );
  NAND2_X1 U7969 ( .A1(n8799), .A2(n6465), .ZN(n6344) );
  INV_X1 U7970 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7971 ( .A1(n6399), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7972 ( .A1(n6024), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6339) );
  OAI211_X1 U7973 ( .C1(n6341), .C2(n6009), .A(n6340), .B(n6339), .ZN(n6342)
         );
  INV_X1 U7974 ( .A(n6342), .ZN(n6343) );
  NAND2_X1 U7975 ( .A1(n6344), .A2(n6343), .ZN(n8645) );
  NAND2_X1 U7976 ( .A1(n8645), .A2(n6331), .ZN(n8495) );
  AOI21_X1 U7977 ( .B1(n8555), .B2(n8557), .A(n8495), .ZN(n6345) );
  NAND2_X1 U7978 ( .A1(n8497), .A2(n6345), .ZN(n6351) );
  INV_X1 U7979 ( .A(n6346), .ZN(n6348) );
  AND2_X1 U7980 ( .A1(n6348), .A2(n6347), .ZN(n8553) );
  NAND2_X1 U7981 ( .A1(n8555), .A2(n8559), .ZN(n6349) );
  NAND2_X1 U7982 ( .A1(n8553), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U7983 ( .A1(n4237), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U7984 ( .A(n9003), .B(n6077), .ZN(n8524) );
  INV_X1 U7985 ( .A(n6357), .ZN(n6355) );
  AND2_X1 U7986 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6354) );
  NAND2_X1 U7987 ( .A1(n6355), .A2(n6354), .ZN(n6371) );
  INV_X1 U7988 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8561) );
  INV_X1 U7989 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7990 ( .B1(n6357), .B2(n8561), .A(n6356), .ZN(n6358) );
  AND2_X1 U7991 ( .A1(n6371), .A2(n6358), .ZN(n8519) );
  NAND2_X1 U7992 ( .A1(n8519), .A2(n6465), .ZN(n6363) );
  INV_X1 U7993 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U7994 ( .A1(n6024), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7995 ( .A1(n6399), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6359) );
  OAI211_X1 U7996 ( .C1(n6009), .C2(n8764), .A(n6360), .B(n6359), .ZN(n6361)
         );
  INV_X1 U7997 ( .A(n6361), .ZN(n6362) );
  NAND2_X1 U7998 ( .A1(n6363), .A2(n6362), .ZN(n8644) );
  AND2_X1 U7999 ( .A1(n8644), .A2(n6331), .ZN(n6364) );
  AND2_X1 U8000 ( .A1(n8524), .A2(n6364), .ZN(n8523) );
  INV_X1 U8001 ( .A(n8524), .ZN(n6366) );
  INV_X1 U8002 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U8003 ( .A1(n6366), .A2(n6365), .ZN(n8526) );
  NAND2_X1 U8004 ( .A1(n4238), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6367) );
  XNOR2_X1 U8006 ( .A(n8998), .B(n6406), .ZN(n6378) );
  INV_X1 U8007 ( .A(n6371), .ZN(n6369) );
  INV_X1 U8008 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U8009 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  INV_X1 U8010 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8011 ( .A1(n6024), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8012 ( .A1(n6399), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6373) );
  OAI211_X1 U8013 ( .C1(n6375), .C2(n6009), .A(n6374), .B(n6373), .ZN(n6376)
         );
  INV_X1 U8014 ( .A(n6376), .ZN(n6377) );
  NAND2_X1 U8015 ( .A1(n8733), .A2(n6331), .ZN(n6379) );
  XNOR2_X1 U8016 ( .A(n6378), .B(n6379), .ZN(n8618) );
  INV_X1 U8017 ( .A(n6378), .ZN(n6381) );
  INV_X1 U8018 ( .A(n6379), .ZN(n6380) );
  NAND2_X1 U8019 ( .A1(n6381), .A2(n6380), .ZN(n6382) );
  NAND2_X1 U8020 ( .A1(n4238), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6383) );
  XNOR2_X1 U8021 ( .A(n8992), .B(n6077), .ZN(n6393) );
  XNOR2_X1 U8022 ( .A(n6397), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U8023 ( .A1(n8743), .A2(n6465), .ZN(n6390) );
  INV_X1 U8024 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8025 ( .A1(n6024), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8026 ( .A1(n6399), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6385) );
  OAI211_X1 U8027 ( .C1(n6387), .C2(n6009), .A(n6386), .B(n6385), .ZN(n6388)
         );
  INV_X1 U8028 ( .A(n6388), .ZN(n6389) );
  NAND2_X1 U8029 ( .A1(n6390), .A2(n6389), .ZN(n8719) );
  NAND2_X1 U8030 ( .A1(n8719), .A2(n6331), .ZN(n6391) );
  XNOR2_X1 U8031 ( .A(n6393), .B(n6391), .ZN(n8472) );
  INV_X1 U8032 ( .A(n6391), .ZN(n6392) );
  NAND2_X1 U8033 ( .A1(n4237), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6394) );
  INV_X1 U8034 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8474) );
  INV_X1 U8035 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6452) );
  OAI21_X1 U8036 ( .B1(n6397), .B2(n8474), .A(n6452), .ZN(n6398) );
  NAND2_X1 U8037 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6396) );
  NAND2_X1 U8038 ( .A1(n8726), .A2(n6465), .ZN(n6405) );
  INV_X1 U8039 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8040 ( .A1(n6399), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8041 ( .A1(n6024), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6400) );
  OAI211_X1 U8042 ( .C1(n6402), .C2(n6009), .A(n6401), .B(n6400), .ZN(n6403)
         );
  INV_X1 U8043 ( .A(n6403), .ZN(n6404) );
  NAND2_X1 U8044 ( .A1(n8740), .A2(n6331), .ZN(n6407) );
  XNOR2_X1 U8045 ( .A(n6407), .B(n6406), .ZN(n6444) );
  INV_X1 U8046 ( .A(n6434), .ZN(n6414) );
  XOR2_X1 U8047 ( .A(n7931), .B(P2_B_REG_SCAN_IN), .Z(n6416) );
  NAND2_X1 U8048 ( .A1(n8037), .A2(n6416), .ZN(n6419) );
  NAND2_X1 U8049 ( .A1(n6417), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6418) );
  NOR2_X1 U8050 ( .A1(n8049), .A2(n6432), .ZN(n10006) );
  NOR4_X1 U8051 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6423) );
  NOR4_X1 U8052 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6422) );
  NOR4_X1 U8053 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6421) );
  NOR4_X1 U8054 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6420) );
  NAND4_X1 U8055 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n6429)
         );
  NOR2_X1 U8056 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n6427) );
  NOR4_X1 U8057 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6426) );
  NOR4_X1 U8058 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6425) );
  NOR4_X1 U8059 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6424) );
  NAND4_X1 U8060 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(n6428)
         );
  OAI21_X1 U8061 ( .B1(n6429), .B2(n6428), .A(n9999), .ZN(n7224) );
  NOR2_X1 U8062 ( .A1(n7931), .A2(n8049), .ZN(n10003) );
  INV_X1 U8063 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10002) );
  AND2_X1 U8064 ( .A1(n7224), .A2(n7303), .ZN(n6431) );
  NAND2_X1 U8065 ( .A1(n7617), .A2(n6431), .ZN(n6449) );
  AND2_X1 U8066 ( .A1(n8049), .A2(n6432), .ZN(n6433) );
  NAND2_X1 U8067 ( .A1(n6434), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6436) );
  INV_X1 U8068 ( .A(n5984), .ZN(n6691) );
  AND2_X1 U8069 ( .A1(n6437), .A2(n6691), .ZN(n9985) );
  NAND2_X1 U8070 ( .A1(n6454), .A2(n9985), .ZN(n6438) );
  NAND3_X1 U8071 ( .A1(n4855), .A2(n6444), .A3(n8617), .ZN(n6439) );
  OAI21_X1 U8072 ( .B1(n4855), .B2(n6444), .A(n6439), .ZN(n6448) );
  INV_X1 U8073 ( .A(n6440), .ZN(n6696) );
  AND2_X1 U8074 ( .A1(n10020), .A2(n7227), .ZN(n6442) );
  AOI21_X1 U8075 ( .B1(n4855), .B2(n8638), .A(n8631), .ZN(n6447) );
  INV_X1 U8076 ( .A(n6444), .ZN(n6443) );
  NAND3_X1 U8077 ( .A1(n4855), .A2(n8617), .A3(n6443), .ZN(n6446) );
  NAND2_X1 U8078 ( .A1(n8729), .A2(n6444), .ZN(n6445) );
  NAND2_X1 U8079 ( .A1(n6449), .A2(n7219), .ZN(n7505) );
  AND3_X1 U8080 ( .A1(n6907), .A2(n6534), .A3(n7221), .ZN(n6450) );
  NAND2_X1 U8081 ( .A1(n7505), .A2(n6450), .ZN(n6451) );
  INV_X1 U8082 ( .A(n8726), .ZN(n6453) );
  OAI22_X1 U8083 ( .A1(n8624), .A2(n6453), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6452), .ZN(n6467) );
  NAND2_X1 U8084 ( .A1(n6454), .A2(n6696), .ZN(n8549) );
  OAI21_X1 U8085 ( .B1(n6455), .B2(P2_IR_REG_27__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6457) );
  INV_X1 U8086 ( .A(n6927), .ZN(n6458) );
  INV_X1 U8087 ( .A(n6459), .ZN(n8356) );
  INV_X1 U8088 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8089 ( .A1(n6024), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8090 ( .A1(n6460), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6461) );
  OAI211_X1 U8091 ( .C1(n6463), .C2(n6025), .A(n6462), .B(n6461), .ZN(n6464)
         );
  AOI21_X1 U8092 ( .B1(n8356), .B2(n6465), .A(n6464), .ZN(n8722) );
  OAI22_X1 U8093 ( .A1(n8351), .A2(n8584), .B1(n8583), .B2(n8722), .ZN(n6466)
         );
  OR2_X1 U8094 ( .A1(n6468), .A2(n7244), .ZN(n6574) );
  NAND2_X1 U8095 ( .A1(n6468), .A2(n7244), .ZN(n6576) );
  NAND2_X2 U8096 ( .A1(n6574), .A2(n6576), .ZN(n7253) );
  INV_X1 U8097 ( .A(n6469), .ZN(n7510) );
  NAND2_X1 U8098 ( .A1(n8660), .A2(n7509), .ZN(n7229) );
  NAND2_X1 U8099 ( .A1(n6565), .A2(n7229), .ZN(n7254) );
  NAND2_X1 U8100 ( .A1(n10015), .A2(n8658), .ZN(n7295) );
  NAND2_X1 U8101 ( .A1(n7591), .A2(n8657), .ZN(n6560) );
  OR2_X1 U8102 ( .A1(n7591), .A2(n8657), .ZN(n6570) );
  NAND2_X1 U8103 ( .A1(n6471), .A2(n6570), .ZN(n7700) );
  INV_X1 U8104 ( .A(n8656), .ZN(n7529) );
  OR2_X1 U8105 ( .A1(n7711), .A2(n7529), .ZN(n6579) );
  NAND2_X1 U8106 ( .A1(n7711), .A2(n7529), .ZN(n6583) );
  INV_X1 U8107 ( .A(n8655), .ZN(n7702) );
  OR2_X1 U8108 ( .A1(n7631), .A2(n7702), .ZN(n6593) );
  NAND2_X1 U8109 ( .A1(n7631), .A2(n7702), .ZN(n6587) );
  NAND2_X1 U8110 ( .A1(n6593), .A2(n6587), .ZN(n7333) );
  INV_X1 U8111 ( .A(n8654), .ZN(n7335) );
  OR2_X1 U8112 ( .A1(n9089), .A2(n7335), .ZN(n6599) );
  NAND2_X1 U8113 ( .A1(n9089), .A2(n7335), .ZN(n6595) );
  NAND2_X1 U8114 ( .A1(n6599), .A2(n6595), .ZN(n7680) );
  INV_X1 U8115 ( .A(n8653), .ZN(n7669) );
  OR2_X1 U8116 ( .A1(n9083), .A2(n7669), .ZN(n6600) );
  NAND2_X1 U8117 ( .A1(n9083), .A2(n7669), .ZN(n6604) );
  INV_X1 U8118 ( .A(n8652), .ZN(n7810) );
  OR2_X1 U8119 ( .A1(n9077), .A2(n7810), .ZN(n6588) );
  NAND2_X1 U8120 ( .A1(n9077), .A2(n7810), .ZN(n6590) );
  NAND2_X1 U8121 ( .A1(n6588), .A2(n6590), .ZN(n7686) );
  NAND2_X1 U8122 ( .A1(n9072), .A2(n8030), .ZN(n6606) );
  INV_X1 U8123 ( .A(n8650), .ZN(n8041) );
  OR2_X1 U8124 ( .A1(n8033), .A2(n8041), .ZN(n6614) );
  OR2_X1 U8125 ( .A1(n9072), .A2(n8030), .ZN(n7864) );
  AND2_X1 U8126 ( .A1(n6614), .A2(n7864), .ZN(n6607) );
  OR2_X1 U8127 ( .A1(n9066), .A2(n8483), .ZN(n6617) );
  NAND2_X1 U8128 ( .A1(n9066), .A2(n8483), .ZN(n6616) );
  NAND2_X1 U8129 ( .A1(n6617), .A2(n6616), .ZN(n7945) );
  INV_X1 U8130 ( .A(n8648), .ZN(n8933) );
  INV_X1 U8131 ( .A(n6621), .ZN(n6474) );
  INV_X1 U8132 ( .A(n8913), .ZN(n8537) );
  OR2_X1 U8133 ( .A1(n9056), .A2(n8537), .ZN(n6475) );
  NAND2_X1 U8134 ( .A1(n9056), .A2(n8537), .ZN(n6623) );
  NAND2_X1 U8135 ( .A1(n6475), .A2(n6623), .ZN(n8939) );
  INV_X1 U8136 ( .A(n6475), .ZN(n6624) );
  INV_X1 U8137 ( .A(n8647), .ZN(n8935) );
  OR2_X1 U8138 ( .A1(n9050), .A2(n8935), .ZN(n6628) );
  INV_X1 U8139 ( .A(n8646), .ZN(n8546) );
  INV_X1 U8140 ( .A(n8915), .ZN(n8612) );
  OR2_X1 U8141 ( .A1(n9045), .A2(n8612), .ZN(n8879) );
  INV_X1 U8142 ( .A(n6631), .ZN(n6479) );
  NAND2_X1 U8143 ( .A1(n9050), .A2(n8935), .ZN(n8878) );
  NOR2_X1 U8144 ( .A1(n8878), .A2(n8915), .ZN(n6477) );
  INV_X1 U8145 ( .A(n8878), .ZN(n6476) );
  OAI22_X1 U8146 ( .A1(n6477), .A2(n9045), .B1(n6476), .B2(n8612), .ZN(n6478)
         );
  NAND2_X1 U8147 ( .A1(n9039), .A2(n8546), .ZN(n6637) );
  INV_X1 U8148 ( .A(n8846), .ZN(n8613) );
  NOR2_X1 U8149 ( .A1(n9034), .A2(n8613), .ZN(n6636) );
  AND2_X1 U8150 ( .A1(n9034), .A2(n8613), .ZN(n6633) );
  NOR2_X1 U8151 ( .A1(n6636), .A2(n6633), .ZN(n8864) );
  NAND2_X1 U8152 ( .A1(n9029), .A2(n8513), .ZN(n6639) );
  INV_X1 U8153 ( .A(n8831), .ZN(n8512) );
  AND2_X1 U8154 ( .A1(n9019), .A2(n8512), .ZN(n6481) );
  INV_X1 U8155 ( .A(n6481), .ZN(n6647) );
  NAND2_X1 U8156 ( .A1(n9024), .A2(n8809), .ZN(n8807) );
  AND2_X1 U8157 ( .A1(n6647), .A2(n8807), .ZN(n6645) );
  OR2_X1 U8158 ( .A1(n9024), .A2(n8809), .ZN(n6640) );
  NAND2_X1 U8159 ( .A1(n9012), .A2(n8810), .ZN(n6651) );
  NAND2_X1 U8160 ( .A1(n9007), .A2(n8557), .ZN(n6650) );
  NAND2_X1 U8161 ( .A1(n6656), .A2(n6650), .ZN(n8778) );
  INV_X1 U8162 ( .A(n6656), .ZN(n6482) );
  NAND2_X1 U8163 ( .A1(n8998), .A2(n8476), .ZN(n8738) );
  INV_X1 U8164 ( .A(n8644), .ZN(n8779) );
  NAND2_X1 U8165 ( .A1(n8752), .A2(n8750), .ZN(n6483) );
  INV_X1 U8166 ( .A(n6483), .ZN(n8736) );
  NAND2_X1 U8167 ( .A1(n9003), .A2(n8779), .ZN(n6658) );
  NAND2_X1 U8168 ( .A1(n8992), .A2(n8351), .ZN(n6669) );
  OAI211_X1 U8169 ( .C1(n6483), .C2(n6658), .A(n8737), .B(n8738), .ZN(n6484)
         );
  INV_X1 U8170 ( .A(n6485), .ZN(n6670) );
  NAND2_X1 U8171 ( .A1(n8729), .A2(n8740), .ZN(n6673) );
  NAND2_X1 U8172 ( .A1(n6487), .A2(n6486), .ZN(n6491) );
  INV_X1 U8173 ( .A(SI_28_), .ZN(n6488) );
  NAND2_X1 U8174 ( .A1(n6489), .A2(n6488), .ZN(n6490) );
  INV_X1 U8175 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9126) );
  INV_X1 U8176 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9754) );
  MUX2_X1 U8177 ( .A(n9126), .B(n9754), .S(n4612), .Z(n6498) );
  XNOR2_X1 U8178 ( .A(n6498), .B(SI_29_), .ZN(n6492) );
  XNOR2_X1 U8179 ( .A(n6497), .B(n6492), .ZN(n9124) );
  NAND2_X1 U8180 ( .A1(n4238), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6493) );
  NOR2_X1 U8181 ( .A1(n8982), .A2(n8722), .ZN(n6681) );
  NAND2_X1 U8182 ( .A1(n8982), .A2(n8722), .ZN(n6680) );
  INV_X1 U8183 ( .A(SI_29_), .ZN(n6495) );
  AND2_X1 U8184 ( .A1(n6498), .A2(n6495), .ZN(n6496) );
  INV_X1 U8185 ( .A(n6498), .ZN(n6499) );
  NAND2_X1 U8186 ( .A1(n6499), .A2(SI_29_), .ZN(n6514) );
  NAND2_X1 U8187 ( .A1(n6516), .A2(n6514), .ZN(n6501) );
  MUX2_X1 U8188 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4612), .Z(n6517) );
  XNOR2_X1 U8189 ( .A(n6517), .B(SI_30_), .ZN(n6500) );
  NAND2_X1 U8190 ( .A1(n4237), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8191 ( .A1(n6024), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6508) );
  INV_X1 U8192 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6504) );
  OR2_X1 U8193 ( .A1(n6025), .A2(n6504), .ZN(n6507) );
  INV_X1 U8194 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6505) );
  OR2_X1 U8195 ( .A1(n6009), .A2(n6505), .ZN(n6506) );
  AND3_X1 U8196 ( .A1(n6508), .A2(n6507), .A3(n6506), .ZN(n6528) );
  OAI211_X1 U8197 ( .C1(n6529), .C2(n8978), .A(n6528), .B(n6563), .ZN(n6531)
         );
  NAND2_X1 U8198 ( .A1(n6024), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6512) );
  INV_X1 U8199 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6509) );
  OR2_X1 U8200 ( .A1(n6025), .A2(n6509), .ZN(n6511) );
  INV_X1 U8201 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8709) );
  OR2_X1 U8202 ( .A1(n6009), .A2(n8709), .ZN(n6510) );
  AND3_X1 U8203 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(n8363) );
  OR2_X1 U8204 ( .A1(n8978), .A2(n8363), .ZN(n6683) );
  NAND2_X1 U8205 ( .A1(n6517), .A2(SI_30_), .ZN(n6513) );
  AND2_X1 U8206 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U8207 ( .A1(n6516), .A2(n6515), .ZN(n6521) );
  INV_X1 U8208 ( .A(n6517), .ZN(n6519) );
  INV_X1 U8209 ( .A(SI_30_), .ZN(n6518) );
  NAND2_X1 U8210 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NAND2_X1 U8211 ( .A1(n6521), .A2(n6520), .ZN(n6526) );
  MUX2_X1 U8212 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4612), .Z(n6524) );
  INV_X1 U8213 ( .A(SI_31_), .ZN(n6523) );
  XNOR2_X1 U8214 ( .A(n6524), .B(n6523), .ZN(n6525) );
  MUX2_X1 U8215 ( .A(n9119), .B(P1_DATAO_REG_31__SCAN_IN), .S(n4612), .Z(n6527) );
  NAND2_X1 U8216 ( .A1(n8977), .A2(n8703), .ZN(n6689) );
  NAND2_X1 U8217 ( .A1(n8978), .A2(n8363), .ZN(n6684) );
  NAND2_X1 U8218 ( .A1(n6689), .A2(n6684), .ZN(n6552) );
  AOI21_X1 U8219 ( .B1(n6529), .B2(n6683), .A(n6552), .ZN(n6530) );
  NOR2_X1 U8220 ( .A1(n8977), .A2(n8703), .ZN(n6539) );
  XNOR2_X1 U8221 ( .A(n6533), .B(n6532), .ZN(n6538) );
  NOR2_X1 U8222 ( .A1(n5984), .A2(n7806), .ZN(n7239) );
  NOR2_X1 U8223 ( .A1(n6534), .A2(P2_U3152), .ZN(n6751) );
  OAI21_X1 U8224 ( .B1(n6535), .B2(n7239), .A(n6751), .ZN(n6536) );
  INV_X1 U8225 ( .A(n6536), .ZN(n6537) );
  INV_X1 U8226 ( .A(n6539), .ZN(n6690) );
  NAND2_X1 U8227 ( .A1(n6690), .A2(n6683), .ZN(n6553) );
  INV_X1 U8228 ( .A(n6553), .ZN(n6548) );
  INV_X1 U8229 ( .A(n6552), .ZN(n6547) );
  INV_X1 U8230 ( .A(n6681), .ZN(n6540) );
  NAND2_X1 U8231 ( .A1(n6540), .A2(n6680), .ZN(n8360) );
  INV_X1 U8232 ( .A(n8737), .ZN(n8352) );
  NAND2_X1 U8233 ( .A1(n8750), .A2(n6658), .ZN(n8765) );
  INV_X1 U8234 ( .A(n8765), .ZN(n8734) );
  NAND2_X1 U8235 ( .A1(n4268), .A2(n6647), .ZN(n8819) );
  XNOR2_X1 U8236 ( .A(n9024), .B(n8809), .ZN(n8826) );
  NAND2_X1 U8237 ( .A1(n6631), .A2(n6637), .ZN(n8889) );
  INV_X1 U8238 ( .A(n8340), .ZN(n6619) );
  INV_X1 U8239 ( .A(n7945), .ZN(n8339) );
  NAND2_X1 U8240 ( .A1(n7864), .A2(n6606), .ZN(n7872) );
  INV_X1 U8241 ( .A(n7229), .ZN(n6541) );
  NOR2_X1 U8242 ( .A1(n6565), .A2(n6541), .ZN(n7280) );
  NAND2_X1 U8243 ( .A1(n6469), .A2(n10010), .ZN(n7731) );
  NAND4_X1 U8244 ( .A1(n7280), .A2(n6470), .A3(n6691), .A4(n7731), .ZN(n6543)
         );
  NAND2_X1 U8245 ( .A1(n6570), .A2(n6560), .ZN(n7296) );
  NOR4_X1 U8246 ( .A1(n6543), .A2(n7296), .A3(n7236), .A4(n6542), .ZN(n6544)
         );
  XNOR2_X1 U8247 ( .A(n9045), .B(n8915), .ZN(n8346) );
  NOR4_X1 U8248 ( .A1(n8778), .A2(n8819), .A3(n8826), .A4(n6545), .ZN(n6546)
         );
  OAI22_X1 U8249 ( .A1(n6549), .A2(n6563), .B1(n6691), .B2(n7240), .ZN(n6694)
         );
  NOR2_X1 U8250 ( .A1(n6532), .A2(n7806), .ZN(n6551) );
  MUX2_X1 U8251 ( .A(n6553), .B(n6552), .S(n4236), .Z(n6554) );
  INV_X1 U8252 ( .A(n6554), .ZN(n6687) );
  INV_X1 U8253 ( .A(n8879), .ZN(n8880) );
  INV_X1 U8254 ( .A(n9045), .ZN(n8906) );
  OAI21_X1 U8255 ( .B1(n8906), .B2(n8915), .A(n6637), .ZN(n6555) );
  MUX2_X1 U8256 ( .A(n8880), .B(n6555), .S(n4236), .Z(n6630) );
  INV_X1 U8257 ( .A(n6604), .ZN(n6556) );
  NAND2_X1 U8258 ( .A1(n6570), .A2(n6567), .ZN(n6557) );
  NAND2_X1 U8259 ( .A1(n8391), .A2(n8659), .ZN(n6558) );
  AOI22_X1 U8260 ( .A1(n6572), .A2(n6560), .B1(n6559), .B2(n6558), .ZN(n6562)
         );
  INV_X1 U8261 ( .A(n6579), .ZN(n6561) );
  OAI21_X1 U8262 ( .B1(n6562), .B2(n6561), .A(n4236), .ZN(n6582) );
  AND2_X1 U8263 ( .A1(n7731), .A2(n6563), .ZN(n6564) );
  OAI211_X1 U8264 ( .C1(n6565), .C2(n6564), .A(n7229), .B(n6576), .ZN(n6566)
         );
  NAND3_X1 U8265 ( .A1(n6566), .A2(n6574), .A3(n6688), .ZN(n6569) );
  AOI21_X1 U8266 ( .B1(n6567), .B2(n4275), .A(n4236), .ZN(n6568) );
  AOI21_X1 U8267 ( .B1(n6569), .B2(n7238), .A(n6568), .ZN(n6573) );
  AND2_X1 U8268 ( .A1(n6583), .A2(n6570), .ZN(n6571) );
  NAND2_X1 U8269 ( .A1(n7229), .A2(n7731), .ZN(n6575) );
  NAND3_X1 U8270 ( .A1(n7230), .A2(n6575), .A3(n6574), .ZN(n6577) );
  NAND3_X1 U8271 ( .A1(n6577), .A2(n4236), .A3(n6576), .ZN(n6578) );
  NAND3_X1 U8272 ( .A1(n6580), .A2(n6579), .A3(n6578), .ZN(n6581) );
  NAND2_X1 U8273 ( .A1(n6582), .A2(n6581), .ZN(n6586) );
  NOR2_X1 U8274 ( .A1(n6583), .A2(n6688), .ZN(n6584) );
  NOR2_X1 U8275 ( .A1(n7333), .A2(n6584), .ZN(n6585) );
  NAND2_X1 U8276 ( .A1(n6586), .A2(n6585), .ZN(n6598) );
  NAND3_X1 U8277 ( .A1(n6598), .A2(n7634), .A3(n6587), .ZN(n6589) );
  NAND2_X1 U8278 ( .A1(n6606), .A2(n6590), .ZN(n6591) );
  MUX2_X1 U8279 ( .A(n6592), .B(n6591), .S(n4236), .Z(n6613) );
  INV_X1 U8280 ( .A(n6593), .ZN(n6594) );
  NOR2_X1 U8281 ( .A1(n7680), .A2(n6594), .ZN(n6597) );
  INV_X1 U8282 ( .A(n6595), .ZN(n6596) );
  AOI21_X1 U8283 ( .B1(n6598), .B2(n6597), .A(n6596), .ZN(n6602) );
  AND2_X1 U8284 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  MUX2_X1 U8285 ( .A(n6602), .B(n6601), .S(n6688), .Z(n6605) );
  AOI21_X1 U8286 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6612) );
  NAND2_X1 U8287 ( .A1(n4245), .A2(n6606), .ZN(n6609) );
  INV_X1 U8288 ( .A(n6607), .ZN(n6608) );
  MUX2_X1 U8289 ( .A(n6609), .B(n6608), .S(n4236), .Z(n6610) );
  INV_X1 U8290 ( .A(n6610), .ZN(n6611) );
  MUX2_X1 U8291 ( .A(n6614), .B(n4245), .S(n4236), .Z(n6615) );
  MUX2_X1 U8292 ( .A(n6617), .B(n6616), .S(n4236), .Z(n6618) );
  MUX2_X1 U8293 ( .A(n6621), .B(n6620), .S(n6688), .Z(n6622) );
  INV_X1 U8294 ( .A(n6623), .ZN(n6625) );
  MUX2_X1 U8295 ( .A(n6625), .B(n6624), .S(n6688), .Z(n6626) );
  INV_X1 U8296 ( .A(n6626), .ZN(n6627) );
  MUX2_X1 U8297 ( .A(n6628), .B(n8878), .S(n6688), .Z(n6629) );
  INV_X1 U8298 ( .A(n6636), .ZN(n6632) );
  NAND3_X1 U8299 ( .A1(n6634), .A2(n6639), .A3(n8807), .ZN(n6635) );
  AOI21_X1 U8300 ( .B1(n6638), .B2(n6637), .A(n6636), .ZN(n6643) );
  NAND2_X1 U8301 ( .A1(n6639), .A2(n5061), .ZN(n6642) );
  OAI211_X1 U8302 ( .C1(n6643), .C2(n6642), .A(n6641), .B(n6640), .ZN(n6644)
         );
  NAND2_X1 U8303 ( .A1(n6645), .A2(n6644), .ZN(n6646) );
  AND2_X1 U8304 ( .A1(n8796), .A2(n6647), .ZN(n6649) );
  INV_X1 U8305 ( .A(n8778), .ZN(n8791) );
  OAI21_X1 U8306 ( .B1(n8810), .B2(n9012), .A(n8791), .ZN(n6648) );
  INV_X1 U8307 ( .A(n6650), .ZN(n6654) );
  NAND2_X1 U8308 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND2_X1 U8309 ( .A1(n6652), .A2(n6688), .ZN(n6653) );
  OAI21_X1 U8310 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(n6663) );
  NOR2_X1 U8311 ( .A1(n6656), .A2(n4236), .ZN(n6657) );
  NOR2_X1 U8312 ( .A1(n8765), .A2(n6657), .ZN(n6662) );
  NAND2_X1 U8313 ( .A1(n6664), .A2(n8750), .ZN(n6660) );
  NAND2_X1 U8314 ( .A1(n8752), .A2(n6658), .ZN(n6659) );
  MUX2_X1 U8315 ( .A(n6660), .B(n6659), .S(n6688), .Z(n6661) );
  INV_X1 U8316 ( .A(n8738), .ZN(n6666) );
  INV_X1 U8317 ( .A(n6664), .ZN(n6665) );
  MUX2_X1 U8318 ( .A(n6666), .B(n6665), .S(n6688), .Z(n6667) );
  INV_X1 U8319 ( .A(n6667), .ZN(n6668) );
  NAND2_X1 U8320 ( .A1(n8737), .A2(n6668), .ZN(n6675) );
  NAND2_X1 U8321 ( .A1(n6677), .A2(n6669), .ZN(n6671) );
  MUX2_X1 U8322 ( .A(n6671), .B(n6670), .S(n4236), .Z(n6672) );
  INV_X1 U8323 ( .A(n6672), .ZN(n6674) );
  NAND2_X1 U8324 ( .A1(n8729), .A2(n6688), .ZN(n6676) );
  NAND2_X1 U8325 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  OAI21_X1 U8326 ( .B1(n4236), .B2(n8740), .A(n6678), .ZN(n6679) );
  INV_X1 U8327 ( .A(n6680), .ZN(n6682) );
  MUX2_X1 U8328 ( .A(n6682), .B(n6681), .S(n6688), .Z(n6685) );
  NAND2_X1 U8329 ( .A1(n6687), .A2(n6686), .ZN(n6693) );
  MUX2_X1 U8330 ( .A(n6690), .B(n6689), .S(n6688), .Z(n6692) );
  AOI21_X1 U8331 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6699) );
  INV_X1 U8332 ( .A(n6751), .ZN(n7939) );
  INV_X1 U8333 ( .A(n7223), .ZN(n6697) );
  XNOR2_X1 U8334 ( .A(n6695), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8362) );
  NAND4_X1 U8335 ( .A1(n6697), .A2(n8912), .A3(n8362), .A4(n6696), .ZN(n6698)
         );
  OAI211_X1 U8336 ( .C1(n6441), .C2(n7939), .A(n6698), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6700) );
  NAND2_X1 U8337 ( .A1(n8177), .A2(n5898), .ZN(n6701) );
  NAND2_X1 U8338 ( .A1(n6701), .A2(n7934), .ZN(n6781) );
  NAND2_X1 U8339 ( .A1(n6781), .A2(n6779), .ZN(n6702) );
  NAND2_X1 U8340 ( .A1(n6702), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8341 ( .A(n7934), .ZN(n6703) );
  INV_X1 U8342 ( .A(n6704), .ZN(n6717) );
  AOI22_X1 U8343 ( .A1(n7077), .A2(P1_STATE_REG_SCAN_IN), .B1(n9748), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n6705) );
  OAI21_X1 U8344 ( .B1(n6717), .B2(n9752), .A(n6705), .ZN(P1_U3348) );
  INV_X1 U8345 ( .A(n9748), .ZN(n9755) );
  OAI222_X1 U8346 ( .A1(n6788), .A2(P1_U3084), .B1(n9752), .B2(n6728), .C1(
        n6706), .C2(n9755), .ZN(P1_U3351) );
  INV_X1 U8347 ( .A(n6707), .ZN(n6719) );
  OAI222_X1 U8348 ( .A1(n9755), .A2(n6708), .B1(n9752), .B2(n6719), .C1(
        P1_U3084), .C2(n6881), .ZN(P1_U3349) );
  OAI222_X1 U8349 ( .A1(n9755), .A2(n6709), .B1(n9752), .B2(n6715), .C1(
        P1_U3084), .C2(n6836), .ZN(P1_U3350) );
  OAI222_X1 U8350 ( .A1(n6783), .A2(P1_U3084), .B1(n9752), .B2(n6730), .C1(
        n6710), .C2(n9755), .ZN(P1_U3352) );
  INV_X1 U8351 ( .A(n6711), .ZN(n6713) );
  AOI22_X1 U8352 ( .A1(n6810), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9748), .ZN(n6712) );
  OAI21_X1 U8353 ( .B1(n6713), .B2(n9752), .A(n6712), .ZN(P1_U3347) );
  INV_X2 U8354 ( .A(n9127), .ZN(n9125) );
  INV_X1 U8355 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6714) );
  INV_X1 U8356 ( .A(n6985), .ZN(n7004) );
  OAI222_X1 U8357 ( .A1(n9125), .A2(n6714), .B1(n7807), .B2(n6713), .C1(
        P2_U3152), .C2(n7004), .ZN(P2_U3352) );
  OAI222_X1 U8358 ( .A1(n9125), .A2(n6716), .B1(n7807), .B2(n6715), .C1(
        P2_U3152), .C2(n6020), .ZN(P2_U3355) );
  INV_X1 U8359 ( .A(n6982), .ZN(n6960) );
  OAI222_X1 U8360 ( .A1(n9125), .A2(n6718), .B1(n7807), .B2(n6717), .C1(
        P2_U3152), .C2(n6960), .ZN(P2_U3353) );
  INV_X1 U8361 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6720) );
  INV_X1 U8362 ( .A(n6953), .ZN(n6943) );
  OAI222_X1 U8363 ( .A1(n9125), .A2(n6720), .B1(n7807), .B2(n6719), .C1(
        P2_U3152), .C2(n6943), .ZN(P2_U3354) );
  NAND2_X1 U8364 ( .A1(n6721), .A2(n8327), .ZN(n6722) );
  OAI21_X1 U8365 ( .B1(n10091), .B2(n8327), .A(n6722), .ZN(P1_U3441) );
  INV_X1 U8366 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6724) );
  INV_X1 U8367 ( .A(n6723), .ZN(n6725) );
  INV_X1 U8368 ( .A(n6849), .ZN(n6854) );
  OAI222_X1 U8369 ( .A1(n9755), .A2(n6724), .B1(n9752), .B2(n6725), .C1(
        P1_U3084), .C2(n6854), .ZN(P1_U3346) );
  INV_X1 U8370 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6726) );
  INV_X1 U8371 ( .A(n7010), .ZN(n6991) );
  OAI222_X1 U8372 ( .A1(n9125), .A2(n6726), .B1(n7807), .B2(n6725), .C1(
        P2_U3152), .C2(n6991), .ZN(P2_U3351) );
  OAI222_X1 U8373 ( .A1(n5987), .A2(P2_U3152), .B1(n7807), .B2(n6728), .C1(
        n6727), .C2(n9125), .ZN(P2_U3356) );
  INV_X1 U8374 ( .A(n7040), .ZN(n6731) );
  INV_X2 U8375 ( .A(n7937), .ZN(n7807) );
  OAI222_X1 U8376 ( .A1(n6731), .A2(P2_U3152), .B1(n7807), .B2(n6730), .C1(
        n6729), .C2(n9125), .ZN(P2_U3357) );
  INV_X1 U8377 ( .A(n6732), .ZN(n6734) );
  AOI22_X1 U8378 ( .A1(n6823), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9748), .ZN(n6733) );
  OAI21_X1 U8379 ( .B1(n6734), .B2(n9752), .A(n6733), .ZN(P1_U3345) );
  INV_X1 U8380 ( .A(n7054), .ZN(n7016) );
  OAI222_X1 U8381 ( .A1(n9125), .A2(n6735), .B1(n7807), .B2(n6734), .C1(
        P2_U3152), .C2(n7016), .ZN(P2_U3350) );
  INV_X1 U8382 ( .A(n6736), .ZN(n6738) );
  INV_X1 U8383 ( .A(n7102), .ZN(n7022) );
  OAI222_X1 U8384 ( .A1(n9755), .A2(n6737), .B1(n9752), .B2(n6738), .C1(n7022), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8385 ( .A(n7059), .ZN(n7133) );
  OAI222_X1 U8386 ( .A1(n9125), .A2(n6739), .B1(n7807), .B2(n6738), .C1(n7133), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8387 ( .A(n6740), .ZN(n6743) );
  INV_X1 U8388 ( .A(n7018), .ZN(n6741) );
  OAI222_X1 U8389 ( .A1(n9755), .A2(n6742), .B1(n9752), .B2(n6743), .C1(n6741), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8390 ( .A(n7057), .ZN(n7122) );
  OAI222_X1 U8391 ( .A1(n9125), .A2(n6744), .B1(n7807), .B2(n6743), .C1(n7122), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8392 ( .A(n6745), .ZN(n6747) );
  INV_X1 U8393 ( .A(n7060), .ZN(n7086) );
  OAI222_X1 U8394 ( .A1(n9125), .A2(n6746), .B1(n7807), .B2(n6747), .C1(n7086), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8395 ( .A(n7347), .ZN(n7110) );
  OAI222_X1 U8396 ( .A1(n9755), .A2(n6748), .B1(n9752), .B2(n6747), .C1(n7110), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8397 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U8398 ( .A1(n8703), .A2(P2_U3966), .ZN(n6749) );
  OAI21_X1 U8399 ( .B1(P2_U3966), .B2(n6750), .A(n6749), .ZN(P2_U3583) );
  NAND2_X1 U8400 ( .A1(n6751), .A2(n5994), .ZN(n6752) );
  NAND2_X1 U8401 ( .A1(n7223), .A2(n6752), .ZN(n6754) );
  NAND2_X1 U8402 ( .A1(n7227), .A2(n6910), .ZN(n6753) );
  NAND2_X1 U8403 ( .A1(n6754), .A2(n6753), .ZN(n8702) );
  NOR2_X1 U8404 ( .A1(n9975), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8405 ( .A(n6755), .ZN(n6759) );
  AOI22_X1 U8406 ( .A1(n7556), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9748), .ZN(n6756) );
  OAI21_X1 U8407 ( .B1(n6759), .B2(n9752), .A(n6756), .ZN(P1_U3341) );
  NAND2_X1 U8408 ( .A1(P1_U4006), .A2(n6757), .ZN(n6758) );
  OAI21_X1 U8409 ( .B1(P1_U4006), .B2(n6000), .A(n6758), .ZN(P1_U3555) );
  INV_X1 U8410 ( .A(n7061), .ZN(n7148) );
  OAI222_X1 U8411 ( .A1(n9125), .A2(n6760), .B1(n7807), .B2(n6759), .C1(
        P2_U3152), .C2(n7148), .ZN(P2_U3346) );
  INV_X1 U8412 ( .A(n6761), .ZN(n6799) );
  AOI22_X1 U8413 ( .A1(n7979), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9748), .ZN(n6762) );
  OAI21_X1 U8414 ( .B1(n6799), .B2(n9752), .A(n6762), .ZN(P1_U3340) );
  INV_X1 U8415 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6764) );
  MUX2_X1 U8416 ( .A(n6764), .B(P1_REG2_REG_2__SCAN_IN), .S(n6788), .Z(n9818)
         );
  XNOR2_X1 U8417 ( .A(n6783), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9804) );
  AND2_X1 U8418 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6765) );
  NAND2_X1 U8419 ( .A1(n9804), .A2(n6765), .ZN(n9803) );
  INV_X1 U8420 ( .A(n6783), .ZN(n9793) );
  NAND2_X1 U8421 ( .A1(n9793), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8422 ( .A1(n9803), .A2(n6766), .ZN(n9819) );
  NAND2_X1 U8423 ( .A1(n9818), .A2(n9819), .ZN(n9816) );
  INV_X1 U8424 ( .A(n6788), .ZN(n9810) );
  NAND2_X1 U8425 ( .A1(n9810), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8426 ( .A1(n9816), .A2(n6838), .ZN(n6768) );
  INV_X1 U8427 ( .A(n6836), .ZN(n6842) );
  NAND2_X1 U8428 ( .A1(n6842), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6769) );
  INV_X1 U8429 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6770) );
  MUX2_X1 U8430 ( .A(n6770), .B(P1_REG2_REG_4__SCAN_IN), .S(n6881), .Z(n6880)
         );
  NAND2_X1 U8431 ( .A1(n6881), .A2(n6770), .ZN(n7071) );
  INV_X1 U8432 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6771) );
  MUX2_X1 U8433 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6771), .S(n7077), .Z(n7070)
         );
  NAND2_X1 U8434 ( .A1(n6772), .A2(n7070), .ZN(n7075) );
  OR2_X1 U8435 ( .A1(n7077), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8436 ( .A1(n7075), .A2(n6773), .ZN(n6778) );
  INV_X1 U8437 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6774) );
  MUX2_X1 U8438 ( .A(n6774), .B(P1_REG2_REG_6__SCAN_IN), .S(n6810), .Z(n6777)
         );
  NOR2_X1 U8439 ( .A1(n4239), .A2(P1_U3084), .ZN(n8055) );
  INV_X1 U8440 ( .A(n9330), .ZN(n6776) );
  AOI21_X1 U8441 ( .B1(n6778), .B2(n6777), .A(n9847), .ZN(n6795) );
  AND2_X1 U8442 ( .A1(n6779), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6780) );
  AND2_X1 U8443 ( .A1(n6781), .A2(n6780), .ZN(n9788) );
  XOR2_X1 U8444 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6810), .Z(n6793) );
  INV_X1 U8445 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6782) );
  OR2_X1 U8446 ( .A1(n6783), .A2(n6782), .ZN(n6787) );
  NAND2_X1 U8447 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  NAND2_X1 U8448 ( .A1(n6787), .A2(n6784), .ZN(n9795) );
  INV_X1 U8449 ( .A(n9795), .ZN(n6786) );
  AND2_X1 U8450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6785) );
  NAND2_X1 U8451 ( .A1(n6786), .A2(n6785), .ZN(n9797) );
  NAND2_X1 U8452 ( .A1(n9797), .A2(n6787), .ZN(n9808) );
  XNOR2_X1 U8453 ( .A(n6788), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U8454 ( .A1(n9808), .A2(n9809), .ZN(n9807) );
  NAND2_X1 U8455 ( .A1(n9810), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6789) );
  XNOR2_X1 U8456 ( .A(n6836), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8457 ( .A1(n6842), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6790) );
  INV_X1 U8458 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9962) );
  MUX2_X1 U8459 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9962), .S(n6881), .Z(n6885)
         );
  NAND2_X1 U8460 ( .A1(n6881), .A2(n9962), .ZN(n6791) );
  NAND2_X1 U8461 ( .A1(n6882), .A2(n6791), .ZN(n7067) );
  XNOR2_X1 U8462 ( .A(n7077), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n7068) );
  OAI21_X1 U8463 ( .B1(n6793), .B2(n6792), .A(n6800), .ZN(n6794) );
  AOI22_X1 U8464 ( .A1(n6795), .A2(n6812), .B1(n9841), .B2(n6794), .ZN(n6798)
         );
  NAND2_X1 U8465 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7463) );
  INV_X1 U8466 ( .A(n7463), .ZN(n6796) );
  AOI21_X1 U8467 ( .B1(n9853), .B2(n6810), .A(n6796), .ZN(n6797) );
  OAI211_X1 U8468 ( .C1(n4524), .C2(n9862), .A(n6798), .B(n6797), .ZN(P1_U3247) );
  INV_X1 U8469 ( .A(n7152), .ZN(n7263) );
  OAI222_X1 U8470 ( .A1(n9125), .A2(n10105), .B1(n7807), .B2(n6799), .C1(n7263), .C2(P2_U3152), .ZN(P2_U3345) );
  AOI21_X1 U8471 ( .B1(n6854), .B2(n9967), .A(n6851), .ZN(n6801) );
  INV_X1 U8472 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U8473 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9970), .S(n6823), .Z(n6821)
         );
  NOR2_X1 U8474 ( .A1(n6823), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6804) );
  OR2_X1 U8475 ( .A1(n7018), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8476 ( .A1(n7018), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6802) );
  AND2_X1 U8477 ( .A1(n7025), .A2(n6802), .ZN(n6803) );
  INV_X1 U8478 ( .A(n7026), .ZN(n6806) );
  NOR3_X1 U8479 ( .A1(n6819), .A2(n6804), .A3(n6803), .ZN(n6805) );
  OAI21_X1 U8480 ( .B1(n6806), .B2(n6805), .A(n9841), .ZN(n6809) );
  NOR2_X1 U8481 ( .A1(n6807), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7768) );
  AOI21_X1 U8482 ( .B1(n9853), .B2(n7018), .A(n7768), .ZN(n6808) );
  OAI211_X1 U8483 ( .C1(n10236), .C2(n9862), .A(n6809), .B(n6808), .ZN(n6817)
         );
  XNOR2_X1 U8484 ( .A(n7018), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6815) );
  INV_X1 U8485 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8486 ( .A1(n6810), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6811) );
  XNOR2_X1 U8487 ( .A(n6823), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6818) );
  AOI211_X1 U8488 ( .C1(n6815), .C2(n6814), .A(n9847), .B(n7017), .ZN(n6816)
         );
  OR2_X1 U8489 ( .A1(n6817), .A2(n6816), .ZN(P1_U3250) );
  XOR2_X1 U8490 ( .A(n6818), .B(n6855), .Z(n6828) );
  INV_X1 U8491 ( .A(n6819), .ZN(n6820) );
  OAI21_X1 U8492 ( .B1(n6822), .B2(n6821), .A(n6820), .ZN(n6826) );
  NAND2_X1 U8493 ( .A1(n9853), .A2(n6823), .ZN(n6824) );
  NAND2_X1 U8494 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7493) );
  OAI211_X1 U8495 ( .C1(n9862), .C2(n4538), .A(n6824), .B(n7493), .ZN(n6825)
         );
  AOI21_X1 U8496 ( .B1(n6826), .B2(n9841), .A(n6825), .ZN(n6827) );
  OAI21_X1 U8497 ( .B1(n9847), .B2(n6828), .A(n6827), .ZN(P1_U3249) );
  INV_X1 U8498 ( .A(n6829), .ZN(n6831) );
  INV_X1 U8499 ( .A(n7693), .ZN(n7691) );
  OAI222_X1 U8500 ( .A1(n9125), .A2(n6830), .B1(n7807), .B2(n6831), .C1(n7691), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U8501 ( .A1(n9755), .A2(n6832), .B1(n9752), .B2(n6831), .C1(n9316), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8502 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6848) );
  OAI211_X1 U8503 ( .C1(n6835), .C2(n6834), .A(n9841), .B(n6833), .ZN(n6846)
         );
  INV_X1 U8504 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U8505 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6837), .S(n6836), .Z(n6839)
         );
  NAND3_X1 U8506 ( .A1(n6839), .A2(n9816), .A3(n6838), .ZN(n6840) );
  NAND3_X1 U8507 ( .A1(n9817), .A2(n6841), .A3(n6840), .ZN(n6845) );
  NAND2_X1 U8508 ( .A1(n9853), .A2(n6842), .ZN(n6844) );
  NOR2_X1 U8509 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5233), .ZN(n7168) );
  INV_X1 U8510 ( .A(n7168), .ZN(n6843) );
  AND4_X1 U8511 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  OAI21_X1 U8512 ( .B1(n6848), .B2(n9862), .A(n6847), .ZN(P1_U3244) );
  XNOR2_X1 U8513 ( .A(n6849), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6850) );
  XNOR2_X1 U8514 ( .A(n6851), .B(n6850), .ZN(n6861) );
  INV_X1 U8515 ( .A(n9862), .ZN(n9789) );
  AND2_X1 U8516 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7608) );
  INV_X1 U8517 ( .A(n9853), .ZN(n7106) );
  NAND3_X1 U8518 ( .A1(n9330), .A2(P1_REG2_REG_7__SCAN_IN), .A3(n6858), .ZN(
        n6852) );
  AOI21_X1 U8519 ( .B1(n7106), .B2(n6852), .A(n6854), .ZN(n6853) );
  AOI211_X1 U8520 ( .C1(n9789), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7608), .B(
        n6853), .ZN(n6860) );
  NAND2_X1 U8521 ( .A1(n6854), .A2(n6813), .ZN(n6857) );
  INV_X1 U8522 ( .A(n6855), .ZN(n6856) );
  OAI211_X1 U8523 ( .C1(n6858), .C2(n6857), .A(n6856), .B(n9817), .ZN(n6859)
         );
  OAI211_X1 U8524 ( .C1(n6861), .C2(n9858), .A(n6860), .B(n6859), .ZN(P1_U3248) );
  INV_X1 U8525 ( .A(n6862), .ZN(n6864) );
  AOI21_X1 U8526 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6866) );
  AOI21_X1 U8527 ( .B1(n7094), .B2(n4401), .A(n6866), .ZN(n6873) );
  NAND2_X1 U8528 ( .A1(n6867), .A2(n8327), .ZN(n7188) );
  INV_X1 U8529 ( .A(n7188), .ZN(n6896) );
  AND3_X1 U8530 ( .A1(n6869), .A2(n6868), .A3(n6896), .ZN(n7096) );
  INV_X1 U8531 ( .A(n7096), .ZN(n6870) );
  AOI22_X1 U8532 ( .A1(n6870), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9288), .B2(
        n9892), .ZN(n6872) );
  AOI22_X1 U8533 ( .A1(n9284), .A2(n7362), .B1(n9272), .B2(n6757), .ZN(n6871)
         );
  OAI211_X1 U8534 ( .C1(n6873), .C2(n9278), .A(n6872), .B(n6871), .ZN(P1_U3220) );
  INV_X1 U8535 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6892) );
  INV_X1 U8536 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9785) );
  OAI21_X1 U8537 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n4239), .A(n6874), .ZN(
        n9784) );
  INV_X1 U8538 ( .A(P1_U4006), .ZN(n9295) );
  NAND2_X1 U8539 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9802) );
  OAI21_X1 U8540 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6904) );
  MUX2_X1 U8541 ( .A(n9802), .B(n6904), .S(n4239), .Z(n6878) );
  NOR2_X1 U8542 ( .A1(n6878), .A2(n8336), .ZN(n6879) );
  AOI211_X1 U8543 ( .C1(n9785), .C2(n9784), .A(n9295), .B(n6879), .ZN(n9815)
         );
  INV_X1 U8544 ( .A(n9815), .ZN(n6891) );
  OAI21_X1 U8545 ( .B1(n4332), .B2(n6880), .A(n7073), .ZN(n6889) );
  NOR2_X1 U8546 ( .A1(n7106), .A2(n6881), .ZN(n6888) );
  INV_X1 U8547 ( .A(n6882), .ZN(n6883) );
  AOI21_X1 U8548 ( .B1(n6885), .B2(n6884), .A(n6883), .ZN(n6886) );
  NAND2_X1 U8549 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U8550 ( .B1(n9858), .B2(n6886), .A(n7199), .ZN(n6887) );
  AOI211_X1 U8551 ( .C1(n9817), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6890)
         );
  OAI211_X1 U8552 ( .C1(n6892), .C2(n9862), .A(n6891), .B(n6890), .ZN(P1_U3245) );
  OR2_X1 U8553 ( .A1(n9949), .A2(n9468), .ZN(n6893) );
  INV_X1 U8554 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6903) );
  INV_X1 U8555 ( .A(n7387), .ZN(n8236) );
  AND2_X1 U8556 ( .A1(n6757), .A2(n7387), .ZN(n7314) );
  INV_X1 U8557 ( .A(n7314), .ZN(n6899) );
  INV_X1 U8558 ( .A(n6757), .ZN(n6897) );
  NAND2_X1 U8559 ( .A1(n6897), .A2(n8236), .ZN(n6898) );
  NAND2_X1 U8560 ( .A1(n6899), .A2(n6898), .ZN(n8189) );
  OR2_X1 U8561 ( .A1(n8177), .A2(n8325), .ZN(n6900) );
  NAND2_X1 U8562 ( .A1(n6900), .A2(n7378), .ZN(n7178) );
  INV_X1 U8563 ( .A(n9309), .ZN(n7179) );
  OAI22_X1 U8564 ( .A1(n8189), .A2(n7178), .B1(n7179), .B2(n9927), .ZN(n7386)
         );
  INV_X1 U8565 ( .A(n7386), .ZN(n6901) );
  OAI21_X1 U8566 ( .B1(n7378), .B2(n8236), .A(n6901), .ZN(n9725) );
  NAND2_X1 U8567 ( .A1(n9725), .A2(n9958), .ZN(n6902) );
  OAI21_X1 U8568 ( .B1(n9958), .B2(n6903), .A(n6902), .ZN(P1_U3454) );
  INV_X1 U8569 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9791) );
  AOI22_X1 U8570 ( .A1(n9284), .A2(n9309), .B1(n7387), .B2(n9288), .ZN(n6906)
         );
  NAND2_X1 U8571 ( .A1(n5905), .A2(n6904), .ZN(n6905) );
  OAI211_X1 U8572 ( .C1(n7096), .C2(n9791), .A(n6906), .B(n6905), .ZN(P1_U3230) );
  INV_X1 U8573 ( .A(n7227), .ZN(n6909) );
  OR2_X1 U8574 ( .A1(n6927), .A2(P2_U3152), .ZN(n9129) );
  OR2_X1 U8575 ( .A1(n6907), .A2(n9129), .ZN(n6908) );
  OAI211_X1 U8576 ( .C1(n7223), .C2(n6909), .A(n6908), .B(n7939), .ZN(n6911)
         );
  NAND2_X1 U8577 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8578 ( .A1(n6912), .A2(n8661), .ZN(n6929) );
  INV_X1 U8579 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U8580 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10175), .ZN(n6920) );
  MUX2_X1 U8581 ( .A(n6011), .B(P2_REG1_REG_1__SCAN_IN), .S(n7040), .Z(n7037)
         );
  INV_X1 U8582 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7034) );
  NOR3_X1 U8583 ( .A1(n7037), .A2(n6913), .A3(n7034), .ZN(n7035) );
  AOI21_X1 U8584 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n7040), .A(n7035), .ZN(
        n6935) );
  MUX2_X1 U8585 ( .A(n6914), .B(P2_REG1_REG_2__SCAN_IN), .S(n6923), .Z(n6934)
         );
  NOR2_X1 U8586 ( .A1(n6935), .A2(n6934), .ZN(n6964) );
  NOR2_X1 U8587 ( .A1(n5987), .A2(n6914), .ZN(n6963) );
  MUX2_X1 U8588 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6915), .S(n6925), .Z(n6962)
         );
  OAI21_X1 U8589 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6961) );
  NAND2_X1 U8590 ( .A1(n6925), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6917) );
  INV_X1 U8591 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10032) );
  MUX2_X1 U8592 ( .A(n10032), .B(P2_REG1_REG_4__SCAN_IN), .S(n6953), .Z(n6916)
         );
  AOI21_X1 U8593 ( .B1(n6961), .B2(n6917), .A(n6916), .ZN(n6947) );
  AND3_X1 U8594 ( .A1(n6961), .A2(n6917), .A3(n6916), .ZN(n6918) );
  NOR3_X1 U8595 ( .A1(n9978), .A2(n6947), .A3(n6918), .ZN(n6919) );
  AOI211_X1 U8596 ( .C1(n9975), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6920), .B(
        n6919), .ZN(n6933) );
  MUX2_X1 U8597 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6044), .S(n6953), .Z(n6931)
         );
  XNOR2_X1 U8598 ( .A(n6923), .B(n8971), .ZN(n6940) );
  XNOR2_X1 U8599 ( .A(n7040), .B(n6921), .ZN(n7043) );
  AND2_X1 U8600 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7042) );
  NAND2_X1 U8601 ( .A1(n7043), .A2(n7042), .ZN(n7041) );
  NAND2_X1 U8602 ( .A1(n7040), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U8603 ( .A1(n7041), .A2(n6922), .ZN(n6939) );
  NAND2_X1 U8604 ( .A1(n6940), .A2(n6939), .ZN(n6938) );
  NAND2_X1 U8605 ( .A1(n6923), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U8606 ( .A1(n6938), .A2(n6924), .ZN(n6970) );
  XNOR2_X1 U8607 ( .A(n6925), .B(n8958), .ZN(n6971) );
  NAND2_X1 U8608 ( .A1(n6970), .A2(n6971), .ZN(n6969) );
  NAND2_X1 U8609 ( .A1(n6925), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U8610 ( .A1(n6969), .A2(n6926), .ZN(n6930) );
  INV_X1 U8611 ( .A(n8362), .ZN(n8059) );
  NOR2_X1 U8612 ( .A1(n8059), .A2(n6927), .ZN(n6928) );
  NAND2_X1 U8613 ( .A1(n6930), .A2(n6931), .ZN(n6955) );
  OAI211_X1 U8614 ( .C1(n6931), .C2(n6930), .A(n9974), .B(n6955), .ZN(n6932)
         );
  OAI211_X1 U8615 ( .C1(n9977), .C2(n6943), .A(n6933), .B(n6932), .ZN(P2_U3249) );
  NOR2_X1 U8616 ( .A1(n8966), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6937) );
  AOI211_X1 U8617 ( .C1(n6935), .C2(n6934), .A(n6964), .B(n9978), .ZN(n6936)
         );
  AOI211_X1 U8618 ( .C1(n9975), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n6937), .B(
        n6936), .ZN(n6942) );
  OAI211_X1 U8619 ( .C1(n6940), .C2(n6939), .A(n9974), .B(n6938), .ZN(n6941)
         );
  OAI211_X1 U8620 ( .C1(n9977), .C2(n5987), .A(n6942), .B(n6941), .ZN(P2_U3247) );
  NAND2_X1 U8621 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7592) );
  INV_X1 U8622 ( .A(n7592), .ZN(n6951) );
  NOR2_X1 U8623 ( .A1(n6943), .A2(n10032), .ZN(n6946) );
  MUX2_X1 U8624 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6944), .S(n6982), .Z(n6945)
         );
  OAI21_X1 U8625 ( .B1(n6947), .B2(n6946), .A(n6945), .ZN(n6994) );
  INV_X1 U8626 ( .A(n6994), .ZN(n6949) );
  NOR3_X1 U8627 ( .A1(n6947), .A2(n6946), .A3(n6945), .ZN(n6948) );
  NOR3_X1 U8628 ( .A1(n9978), .A2(n6949), .A3(n6948), .ZN(n6950) );
  AOI211_X1 U8629 ( .C1(n9975), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6951), .B(
        n6950), .ZN(n6959) );
  XNOR2_X1 U8630 ( .A(n6982), .B(n6952), .ZN(n6957) );
  NAND2_X1 U8631 ( .A1(n6953), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8632 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  NAND2_X1 U8633 ( .A1(n6956), .A2(n6957), .ZN(n6984) );
  OAI211_X1 U8634 ( .C1(n6957), .C2(n6956), .A(n9974), .B(n6984), .ZN(n6958)
         );
  OAI211_X1 U8635 ( .C1(n9977), .C2(n6960), .A(n6959), .B(n6958), .ZN(P2_U3250) );
  INV_X1 U8636 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8954) );
  NOR2_X1 U8637 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8954), .ZN(n6968) );
  INV_X1 U8638 ( .A(n6961), .ZN(n6966) );
  NOR3_X1 U8639 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n6965) );
  NOR3_X1 U8640 ( .A1(n9978), .A2(n6966), .A3(n6965), .ZN(n6967) );
  AOI211_X1 U8641 ( .C1(n9975), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6968), .B(
        n6967), .ZN(n6973) );
  OAI211_X1 U8642 ( .C1(n6971), .C2(n6970), .A(n9974), .B(n6969), .ZN(n6972)
         );
  OAI211_X1 U8643 ( .C1(n9977), .C2(n6020), .A(n6973), .B(n6972), .ZN(P2_U3248) );
  NOR2_X1 U8644 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6092), .ZN(n7527) );
  NAND2_X1 U8645 ( .A1(n6982), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6993) );
  MUX2_X1 U8646 ( .A(n6974), .B(P2_REG1_REG_6__SCAN_IN), .S(n6985), .Z(n6992)
         );
  AOI21_X1 U8647 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n6996) );
  NOR2_X1 U8648 ( .A1(n7004), .A2(n6974), .ZN(n6978) );
  NAND2_X1 U8649 ( .A1(n7010), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U8650 ( .A1(n6991), .A2(n6976), .ZN(n6975) );
  OAI211_X1 U8651 ( .C1(n6996), .C2(n6978), .A(n7005), .B(n6975), .ZN(n7006)
         );
  INV_X1 U8652 ( .A(n7006), .ZN(n6980) );
  MUX2_X1 U8653 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6976), .S(n7010), .Z(n6977)
         );
  NOR3_X1 U8654 ( .A1(n6996), .A2(n6978), .A3(n6977), .ZN(n6979) );
  NOR3_X1 U8655 ( .A1(n6980), .A2(n6979), .A3(n9978), .ZN(n6981) );
  AOI211_X1 U8656 ( .C1(n9975), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7527), .B(
        n6981), .ZN(n6990) );
  NAND2_X1 U8657 ( .A1(n6982), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U8658 ( .A1(n6984), .A2(n6983), .ZN(n7000) );
  XNOR2_X1 U8659 ( .A(n6985), .B(n7706), .ZN(n7001) );
  NAND2_X1 U8660 ( .A1(n7000), .A2(n7001), .ZN(n6999) );
  NAND2_X1 U8661 ( .A1(n6985), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6986) );
  OAI211_X1 U8662 ( .C1(n6988), .C2(n6987), .A(n9974), .B(n7011), .ZN(n6989)
         );
  OAI211_X1 U8663 ( .C1(n9977), .C2(n6991), .A(n6990), .B(n6989), .ZN(P2_U3252) );
  NAND2_X1 U8664 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7581) );
  INV_X1 U8665 ( .A(n7581), .ZN(n6998) );
  AND3_X1 U8666 ( .A1(n6994), .A2(n6993), .A3(n6992), .ZN(n6995) );
  NOR3_X1 U8667 ( .A1(n9978), .A2(n6996), .A3(n6995), .ZN(n6997) );
  AOI211_X1 U8668 ( .C1(n9975), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6998), .B(
        n6997), .ZN(n7003) );
  OAI211_X1 U8669 ( .C1(n7001), .C2(n7000), .A(n9974), .B(n6999), .ZN(n7002)
         );
  OAI211_X1 U8670 ( .C1(n9977), .C2(n7004), .A(n7003), .B(n7002), .ZN(P2_U3251) );
  NOR2_X1 U8671 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7573), .ZN(n7009) );
  NAND2_X1 U8672 ( .A1(n7006), .A2(n7005), .ZN(n7047) );
  XOR2_X1 U8673 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7054), .Z(n7046) );
  XNOR2_X1 U8674 ( .A(n7047), .B(n7046), .ZN(n7007) );
  NOR2_X1 U8675 ( .A1(n7007), .A2(n9978), .ZN(n7008) );
  AOI211_X1 U8676 ( .C1(n9975), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7009), .B(
        n7008), .ZN(n7015) );
  XNOR2_X1 U8677 ( .A(n7054), .B(n7644), .ZN(n7013) );
  OAI211_X1 U8678 ( .C1(n7013), .C2(n7012), .A(n9974), .B(n7056), .ZN(n7014)
         );
  OAI211_X1 U8679 ( .C1(n9977), .C2(n7016), .A(n7015), .B(n7014), .ZN(P2_U3253) );
  XNOR2_X1 U8680 ( .A(n7102), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7019) );
  AOI211_X1 U8681 ( .C1(n7020), .C2(n7019), .A(n9847), .B(n7101), .ZN(n7033)
         );
  INV_X1 U8682 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8683 ( .A1(n7022), .A2(n7021), .ZN(n7108) );
  NAND2_X1 U8684 ( .A1(n7102), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U8685 ( .A1(n7108), .A2(n7023), .ZN(n7024) );
  INV_X1 U8686 ( .A(n7114), .ZN(n7028) );
  NAND3_X1 U8687 ( .A1(n7026), .A2(n7025), .A3(n7024), .ZN(n7027) );
  AOI21_X1 U8688 ( .B1(n7028), .B2(n7027), .A(n9858), .ZN(n7032) );
  INV_X1 U8689 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8690 ( .A1(n9853), .A2(n7102), .ZN(n7029) );
  NAND2_X1 U8691 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7797) );
  OAI211_X1 U8692 ( .C1(n9862), .C2(n7030), .A(n7029), .B(n7797), .ZN(n7031)
         );
  OR3_X1 U8693 ( .A1(n7033), .A2(n7032), .A3(n7031), .ZN(P1_U3251) );
  INV_X1 U8694 ( .A(n9977), .ZN(n7053) );
  INV_X1 U8695 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9762) );
  OAI22_X1 U8696 ( .A1(n8702), .A2(n9762), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7756), .ZN(n7039) );
  OR2_X1 U8697 ( .A1(n7034), .A2(n6913), .ZN(n7036) );
  AOI211_X1 U8698 ( .C1(n7037), .C2(n7036), .A(n7035), .B(n9978), .ZN(n7038)
         );
  AOI211_X1 U8699 ( .C1(n7053), .C2(n7040), .A(n7039), .B(n7038), .ZN(n7045)
         );
  OAI211_X1 U8700 ( .C1(n7043), .C2(n7042), .A(n9974), .B(n7041), .ZN(n7044)
         );
  NAND2_X1 U8701 ( .A1(n7045), .A2(n7044), .ZN(P2_U3246) );
  INV_X1 U8702 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U8703 ( .A1(n7148), .A2(n8007), .ZN(n7151) );
  OAI21_X1 U8704 ( .B1(n8007), .B2(n7148), .A(n7151), .ZN(n7051) );
  AOI22_X1 U8705 ( .A1(n7047), .A2(n7046), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7054), .ZN(n7121) );
  XNOR2_X1 U8706 ( .A(n7057), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7120) );
  INV_X1 U8707 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7048) );
  OAI22_X1 U8708 ( .A1(n7121), .A2(n7120), .B1(n7122), .B2(n7048), .ZN(n7131)
         );
  XOR2_X1 U8709 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7059), .Z(n7130) );
  AOI22_X1 U8710 ( .A1(n7131), .A2(n7130), .B1(n7059), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7083) );
  XNOR2_X1 U8711 ( .A(n7060), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7084) );
  OAI22_X1 U8712 ( .A1(n7083), .A2(n7084), .B1(n7086), .B2(n7049), .ZN(n7050)
         );
  NOR2_X1 U8713 ( .A1(n7050), .A2(n7051), .ZN(n7156) );
  AOI21_X1 U8714 ( .B1(n7051), .B2(n7050), .A(n7156), .ZN(n7065) );
  NAND2_X1 U8715 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8028) );
  OAI21_X1 U8716 ( .B1(n8702), .B2(n4537), .A(n8028), .ZN(n7052) );
  AOI21_X1 U8717 ( .B1(n7053), .B2(n7061), .A(n7052), .ZN(n7064) );
  NAND2_X1 U8718 ( .A1(n7054), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8719 ( .A1(n7056), .A2(n7055), .ZN(n7125) );
  XNOR2_X1 U8720 ( .A(n7057), .B(n7662), .ZN(n7126) );
  NAND2_X1 U8721 ( .A1(n7125), .A2(n7126), .ZN(n7124) );
  NAND2_X1 U8722 ( .A1(n7057), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8723 ( .A1(n7124), .A2(n7058), .ZN(n7137) );
  XNOR2_X1 U8724 ( .A(n7059), .B(n7673), .ZN(n7138) );
  XNOR2_X1 U8725 ( .A(n7060), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n7082) );
  XNOR2_X1 U8726 ( .A(n7061), .B(n7877), .ZN(n7062) );
  NAND2_X1 U8727 ( .A1(n4257), .A2(n7062), .ZN(n7147) );
  OAI211_X1 U8728 ( .C1(n4257), .C2(n7062), .A(n7147), .B(n9974), .ZN(n7063)
         );
  OAI211_X1 U8729 ( .C1(n7065), .C2(n9978), .A(n7064), .B(n7063), .ZN(P2_U3257) );
  AOI211_X1 U8730 ( .C1(n7068), .C2(n7067), .A(n7066), .B(n9858), .ZN(n7069)
         );
  AND2_X1 U8731 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7215) );
  NOR2_X1 U8732 ( .A1(n7069), .A2(n7215), .ZN(n7079) );
  INV_X1 U8733 ( .A(n7070), .ZN(n7072) );
  NAND3_X1 U8734 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7074) );
  AOI21_X1 U8735 ( .B1(n7075), .B2(n7074), .A(n9847), .ZN(n7076) );
  AOI21_X1 U8736 ( .B1(n9853), .B2(n7077), .A(n7076), .ZN(n7078) );
  OAI211_X1 U8737 ( .C1(n4526), .C2(n9862), .A(n7079), .B(n7078), .ZN(P1_U3246) );
  AOI21_X1 U8738 ( .B1(n7082), .B2(n7081), .A(n7080), .ZN(n7090) );
  XOR2_X1 U8739 ( .A(n7084), .B(n7083), .Z(n7088) );
  AND2_X1 U8740 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7989) );
  AOI21_X1 U8741 ( .B1(n9975), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7989), .ZN(
        n7085) );
  OAI21_X1 U8742 ( .B1(n9977), .B2(n7086), .A(n7085), .ZN(n7087) );
  AOI21_X1 U8743 ( .B1(n7088), .B2(n9973), .A(n7087), .ZN(n7089) );
  OAI21_X1 U8744 ( .B1(n7090), .B2(n9976), .A(n7089), .ZN(P2_U3256) );
  INV_X1 U8745 ( .A(n7091), .ZN(n7171) );
  AOI22_X1 U8746 ( .A1(n9333), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9748), .ZN(n7092) );
  OAI21_X1 U8747 ( .B1(n7171), .B2(n9752), .A(n7092), .ZN(P1_U3338) );
  OAI21_X1 U8748 ( .B1(n7095), .B2(n7094), .A(n7093), .ZN(n7099) );
  INV_X1 U8749 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9822) );
  OAI22_X1 U8750 ( .A1(n9235), .A2(n7175), .B1(n9822), .B2(n7096), .ZN(n7098)
         );
  OAI22_X1 U8751 ( .A1(n7374), .A2(n9275), .B1(n9282), .B2(n7179), .ZN(n7097)
         );
  AOI211_X1 U8752 ( .C1(n7099), .C2(n5905), .A(n7098), .B(n7097), .ZN(n7100)
         );
  INV_X1 U8753 ( .A(n7100), .ZN(P1_U3235) );
  XOR2_X1 U8754 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7347), .Z(n7104) );
  OAI21_X1 U8755 ( .B1(n7104), .B2(n7103), .A(n7346), .ZN(n7105) );
  INV_X1 U8756 ( .A(n7105), .ZN(n7119) );
  NAND2_X1 U8757 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7886) );
  OAI21_X1 U8758 ( .B1(n7106), .B2(n7110), .A(n7886), .ZN(n7107) );
  AOI21_X1 U8759 ( .B1(n9789), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7107), .ZN(
        n7118) );
  INV_X1 U8760 ( .A(n7108), .ZN(n7113) );
  INV_X1 U8761 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8762 ( .A1(n7110), .A2(n7109), .ZN(n7352) );
  NAND2_X1 U8763 ( .A1(n7347), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7111) );
  AND2_X1 U8764 ( .A1(n7352), .A2(n7111), .ZN(n7112) );
  OAI21_X1 U8765 ( .B1(n7114), .B2(n7113), .A(n7112), .ZN(n7353) );
  INV_X1 U8766 ( .A(n7353), .ZN(n7116) );
  NOR3_X1 U8767 ( .A1(n7114), .A2(n7113), .A3(n7112), .ZN(n7115) );
  OAI21_X1 U8768 ( .B1(n7116), .B2(n7115), .A(n9841), .ZN(n7117) );
  OAI211_X1 U8769 ( .C1(n7119), .C2(n9847), .A(n7118), .B(n7117), .ZN(P1_U3252) );
  XNOR2_X1 U8770 ( .A(n7121), .B(n7120), .ZN(n7129) );
  AND2_X1 U8771 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7826) );
  NOR2_X1 U8772 ( .A1(n9977), .A2(n7122), .ZN(n7123) );
  AOI211_X1 U8773 ( .C1(n9975), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7826), .B(
        n7123), .ZN(n7128) );
  OAI211_X1 U8774 ( .C1(n7126), .C2(n7125), .A(n9974), .B(n7124), .ZN(n7127)
         );
  OAI211_X1 U8775 ( .C1(n7129), .C2(n9978), .A(n7128), .B(n7127), .ZN(P2_U3254) );
  XNOR2_X1 U8776 ( .A(n7131), .B(n7130), .ZN(n7141) );
  NOR2_X1 U8777 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7132), .ZN(n7135) );
  NOR2_X1 U8778 ( .A1(n9977), .A2(n7133), .ZN(n7134) );
  AOI211_X1 U8779 ( .C1(n9975), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7135), .B(
        n7134), .ZN(n7140) );
  OAI211_X1 U8780 ( .C1(n7138), .C2(n7137), .A(n9974), .B(n7136), .ZN(n7139)
         );
  OAI211_X1 U8781 ( .C1(n7141), .C2(n9978), .A(n7140), .B(n7139), .ZN(P2_U3255) );
  INV_X1 U8782 ( .A(n8327), .ZN(n7143) );
  OAI21_X1 U8783 ( .B1(n9891), .B2(P1_D_REG_0__SCAN_IN), .A(n7144), .ZN(n7145)
         );
  OAI21_X1 U8784 ( .B1(n8327), .B2(n7146), .A(n7145), .ZN(P1_U3440) );
  XNOR2_X1 U8785 ( .A(n7152), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n7150) );
  OAI21_X1 U8786 ( .B1(n7877), .B2(n7148), .A(n7147), .ZN(n7149) );
  AOI21_X1 U8787 ( .B1(n7150), .B2(n7149), .A(n7262), .ZN(n7163) );
  INV_X1 U8788 ( .A(n7151), .ZN(n7155) );
  OR2_X1 U8789 ( .A1(n7152), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7268) );
  NAND2_X1 U8790 ( .A1(n7152), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7153) );
  AND2_X1 U8791 ( .A1(n7268), .A2(n7153), .ZN(n7154) );
  OAI21_X1 U8792 ( .B1(n7156), .B2(n7155), .A(n7154), .ZN(n7269) );
  INV_X1 U8793 ( .A(n7269), .ZN(n7158) );
  NOR3_X1 U8794 ( .A1(n7156), .A2(n7155), .A3(n7154), .ZN(n7157) );
  OAI21_X1 U8795 ( .B1(n7158), .B2(n7157), .A(n9973), .ZN(n7162) );
  NOR2_X1 U8796 ( .A1(n7159), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8043) );
  NOR2_X1 U8797 ( .A1(n9977), .A2(n7263), .ZN(n7160) );
  AOI211_X1 U8798 ( .C1(n9975), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8043), .B(
        n7160), .ZN(n7161) );
  OAI211_X1 U8799 ( .C1(n7163), .C2(n9976), .A(n7162), .B(n7161), .ZN(P2_U3258) );
  XNOR2_X1 U8800 ( .A(n7165), .B(n7164), .ZN(n7166) );
  NAND2_X1 U8801 ( .A1(n7166), .A2(n5905), .ZN(n7170) );
  OAI22_X1 U8802 ( .A1(n7397), .A2(n9282), .B1(n9275), .B2(n9924), .ZN(n7167)
         );
  AOI211_X1 U8803 ( .C1(n7405), .C2(n9288), .A(n7168), .B(n7167), .ZN(n7169)
         );
  OAI211_X1 U8804 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9286), .A(n7170), .B(
        n7169), .ZN(P1_U3216) );
  INV_X1 U8805 ( .A(n7911), .ZN(n7903) );
  OAI222_X1 U8806 ( .A1(n9125), .A2(n10064), .B1(n7807), .B2(n7171), .C1(
        P2_U3152), .C2(n7903), .ZN(P2_U3343) );
  INV_X1 U8807 ( .A(n9896), .ZN(n9912) );
  NAND2_X1 U8808 ( .A1(n7397), .A2(n7522), .ZN(n8240) );
  INV_X1 U8809 ( .A(n8192), .ZN(n7317) );
  NAND2_X1 U8810 ( .A1(n9309), .A2(n9892), .ZN(n7411) );
  AND2_X1 U8811 ( .A1(n7410), .A2(n7411), .ZN(n7361) );
  INV_X1 U8812 ( .A(n7361), .ZN(n7172) );
  NOR2_X1 U8813 ( .A1(n7172), .A2(n8190), .ZN(n7393) );
  AOI21_X1 U8814 ( .B1(n8190), .B2(n7172), .A(n7393), .ZN(n7519) );
  INV_X1 U8815 ( .A(n7519), .ZN(n7187) );
  NAND2_X1 U8816 ( .A1(n7173), .A2(n7522), .ZN(n7174) );
  NAND2_X1 U8817 ( .A1(n7401), .A2(n7174), .ZN(n7518) );
  OAI22_X1 U8818 ( .A1(n7518), .A2(n9949), .B1(n9947), .B2(n7175), .ZN(n7186)
         );
  AND2_X1 U8819 ( .A1(n7176), .A2(n8325), .ZN(n7177) );
  AOI22_X1 U8820 ( .A1(n9308), .A2(n9542), .B1(n9540), .B2(n9309), .ZN(n7185)
         );
  NAND2_X1 U8821 ( .A1(n7179), .A2(n9892), .ZN(n7180) );
  XNOR2_X1 U8822 ( .A(n8243), .B(n8190), .ZN(n7183) );
  NAND2_X1 U8823 ( .A1(n8331), .A2(n10220), .ZN(n7182) );
  NAND2_X1 U8824 ( .A1(n8313), .A2(n7181), .ZN(n8176) );
  NAND2_X1 U8825 ( .A1(n7183), .A2(n9603), .ZN(n7184) );
  OAI211_X1 U8826 ( .C1(n7519), .C2(n9897), .A(n7185), .B(n7184), .ZN(n7515)
         );
  AOI211_X1 U8827 ( .C1(n9912), .C2(n7187), .A(n7186), .B(n7515), .ZN(n9902)
         );
  NOR2_X1 U8828 ( .A1(n7189), .A2(n7188), .ZN(n7190) );
  NAND2_X1 U8829 ( .A1(n9969), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U8830 ( .B1(n9902), .B2(n9969), .A(n7192), .ZN(P1_U3525) );
  INV_X1 U8831 ( .A(n7193), .ZN(n7194) );
  INV_X1 U8832 ( .A(n8667), .ZN(n8663) );
  OAI222_X1 U8833 ( .A1(n9125), .A2(n10108), .B1(n7807), .B2(n7194), .C1(n8663), .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8834 ( .A(n9828), .ZN(n9336) );
  OAI222_X1 U8835 ( .A1(n9755), .A2(n7195), .B1(n9752), .B2(n7194), .C1(n9336), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8836 ( .A(n7196), .ZN(n7381) );
  OAI211_X1 U8837 ( .C1(n7198), .C2(n7197), .A(n7209), .B(n5905), .ZN(n7203)
         );
  INV_X1 U8838 ( .A(n7199), .ZN(n7201) );
  OAI22_X1 U8839 ( .A1(n7374), .A2(n9282), .B1(n9275), .B2(n8066), .ZN(n7200)
         );
  AOI211_X1 U8840 ( .C1(n7414), .C2(n9288), .A(n7201), .B(n7200), .ZN(n7202)
         );
  OAI211_X1 U8841 ( .C1(n9286), .C2(n7381), .A(n7203), .B(n7202), .ZN(P1_U3228) );
  INV_X1 U8842 ( .A(n7204), .ZN(n7206) );
  AOI22_X1 U8843 ( .A1(n9839), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9748), .ZN(n7205) );
  OAI21_X1 U8844 ( .B1(n7206), .B2(n9752), .A(n7205), .ZN(P1_U3336) );
  INV_X1 U8845 ( .A(n8678), .ZN(n8684) );
  OAI222_X1 U8846 ( .A1(n9125), .A2(n7207), .B1(n7807), .B2(n7206), .C1(n8684), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8847 ( .A1(n7209), .A2(n7208), .ZN(n7213) );
  XNOR2_X1 U8848 ( .A(n7211), .B(n7210), .ZN(n7212) );
  XNOR2_X1 U8849 ( .A(n7213), .B(n7212), .ZN(n7218) );
  OAI22_X1 U8850 ( .A1(n9924), .A2(n9282), .B1(n9275), .B2(n9926), .ZN(n7214)
         );
  AOI211_X1 U8851 ( .C1(n8067), .C2(n9288), .A(n7215), .B(n7214), .ZN(n7217)
         );
  NAND2_X1 U8852 ( .A1(n9271), .A2(n10212), .ZN(n7216) );
  OAI211_X1 U8853 ( .C1(n7218), .C2(n9278), .A(n7217), .B(n7216), .ZN(P1_U3225) );
  INV_X1 U8854 ( .A(n7219), .ZN(n7220) );
  INV_X1 U8855 ( .A(n7305), .ZN(n7226) );
  INV_X1 U8856 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U8857 ( .A1(n6550), .A2(n7626), .ZN(n7228) );
  NAND2_X1 U8858 ( .A1(n7228), .A2(n7227), .ZN(n8869) );
  NAND3_X1 U8859 ( .A1(n6550), .A2(n4769), .A3(n5984), .ZN(n9096) );
  NAND2_X1 U8860 ( .A1(n7230), .A2(n7229), .ZN(n7281) );
  INV_X1 U8861 ( .A(n7279), .ZN(n7231) );
  NAND3_X1 U8862 ( .A1(n7281), .A2(n7253), .A3(n7231), .ZN(n7234) );
  NOR2_X1 U8863 ( .A1(n7759), .A2(n8660), .ZN(n7251) );
  INV_X1 U8864 ( .A(n7244), .ZN(n8962) );
  NOR2_X1 U8865 ( .A1(n8962), .A2(n6468), .ZN(n7232) );
  AOI21_X1 U8866 ( .B1(n7253), .B2(n7251), .A(n7232), .ZN(n7233) );
  NAND2_X1 U8867 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  NAND2_X1 U8868 ( .A1(n7235), .A2(n7236), .ZN(n7291) );
  OAI21_X1 U8869 ( .B1(n7235), .B2(n7236), .A(n7291), .ZN(n8953) );
  INV_X1 U8870 ( .A(n8953), .ZN(n7248) );
  XNOR2_X1 U8871 ( .A(n7238), .B(n7237), .ZN(n7243) );
  INV_X1 U8872 ( .A(n7239), .ZN(n7241) );
  INV_X1 U8873 ( .A(n6468), .ZN(n7242) );
  OAI22_X1 U8874 ( .A1(n7242), .A2(n8932), .B1(n8934), .B2(n7590), .ZN(n8388)
         );
  AOI21_X1 U8875 ( .B1(n7243), .B2(n8917), .A(n8388), .ZN(n8957) );
  INV_X1 U8876 ( .A(n8391), .ZN(n8952) );
  NAND2_X1 U8877 ( .A1(n7286), .A2(n7244), .ZN(n7258) );
  NOR2_X2 U8878 ( .A1(n7258), .A2(n8952), .ZN(n7742) );
  NAND2_X1 U8879 ( .A1(n7258), .A2(n8952), .ZN(n7245) );
  NAND2_X1 U8880 ( .A1(n9091), .A2(n7245), .ZN(n7246) );
  NOR2_X1 U8881 ( .A1(n7742), .A2(n7246), .ZN(n8956) );
  AOI21_X1 U8882 ( .B1(n9090), .B2(n8952), .A(n8956), .ZN(n7247) );
  OAI211_X1 U8883 ( .C1(n9081), .C2(n7248), .A(n8957), .B(n7247), .ZN(n7832)
         );
  NAND2_X1 U8884 ( .A1(n10030), .A2(n7832), .ZN(n7249) );
  OAI21_X1 U8885 ( .B1(n10030), .B2(n7250), .A(n7249), .ZN(P2_U3460) );
  INV_X1 U8886 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10121) );
  INV_X1 U8887 ( .A(n7281), .ZN(n7278) );
  NOR2_X1 U8888 ( .A1(n7278), .A2(n7279), .ZN(n7277) );
  NOR2_X1 U8889 ( .A1(n7277), .A2(n7251), .ZN(n7252) );
  XNOR2_X1 U8890 ( .A(n7252), .B(n6470), .ZN(n8964) );
  INV_X1 U8891 ( .A(n8964), .ZN(n7260) );
  XNOR2_X1 U8892 ( .A(n7254), .B(n7253), .ZN(n7255) );
  OAI22_X1 U8893 ( .A1(n8599), .A2(n8932), .B1(n8934), .B2(n8374), .ZN(n8597)
         );
  AOI21_X1 U8894 ( .B1(n7255), .B2(n8917), .A(n8597), .ZN(n8970) );
  INV_X1 U8895 ( .A(n7286), .ZN(n7256) );
  NAND2_X1 U8896 ( .A1(n7256), .A2(n8962), .ZN(n7257) );
  AND3_X1 U8897 ( .A1(n9091), .A2(n7258), .A3(n7257), .ZN(n8968) );
  AOI21_X1 U8898 ( .B1(n9090), .B2(n8962), .A(n8968), .ZN(n7259) );
  OAI211_X1 U8899 ( .C1(n7260), .C2(n9081), .A(n8970), .B(n7259), .ZN(n7834)
         );
  NAND2_X1 U8900 ( .A1(n10030), .A2(n7834), .ZN(n7261) );
  OAI21_X1 U8901 ( .B1(n10030), .B2(n10121), .A(n7261), .ZN(P2_U3457) );
  MUX2_X1 U8902 ( .A(n8016), .B(P2_REG2_REG_14__SCAN_IN), .S(n7693), .Z(n7266)
         );
  AOI21_X1 U8903 ( .B1(n7266), .B2(n7265), .A(n7690), .ZN(n7276) );
  XNOR2_X1 U8904 ( .A(n7693), .B(n7267), .ZN(n7271) );
  NAND2_X1 U8905 ( .A1(n7269), .A2(n7268), .ZN(n7270) );
  NAND2_X1 U8906 ( .A1(n7270), .A2(n7271), .ZN(n7692) );
  OAI21_X1 U8907 ( .B1(n7271), .B2(n7270), .A(n7692), .ZN(n7274) );
  NAND2_X1 U8908 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U8909 ( .A1(n9975), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7272) );
  OAI211_X1 U8910 ( .C1(n9977), .C2(n7691), .A(n8486), .B(n7272), .ZN(n7273)
         );
  AOI21_X1 U8911 ( .B1(n7274), .B2(n9973), .A(n7273), .ZN(n7275) );
  OAI21_X1 U8912 ( .B1(n7276), .B2(n9976), .A(n7275), .ZN(P2_U3259) );
  INV_X1 U8913 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7289) );
  AOI21_X1 U8914 ( .B1(n7279), .B2(n7278), .A(n7277), .ZN(n7763) );
  NOR2_X1 U8915 ( .A1(n8932), .A2(n7510), .ZN(n7284) );
  INV_X1 U8916 ( .A(n7732), .ZN(n7282) );
  AOI211_X1 U8917 ( .C1(n7282), .C2(n7281), .A(n8930), .B(n7280), .ZN(n7283)
         );
  AOI211_X1 U8918 ( .C1(n8914), .C2(n6468), .A(n7284), .B(n7283), .ZN(n7757)
         );
  NOR2_X1 U8919 ( .A1(n7509), .A2(n10010), .ZN(n7285) );
  NOR2_X1 U8920 ( .A1(n7286), .A2(n7285), .ZN(n7760) );
  AOI22_X1 U8921 ( .A1(n7760), .A2(n9091), .B1(n9090), .B2(n7759), .ZN(n7287)
         );
  OAI211_X1 U8922 ( .C1(n9081), .C2(n7763), .A(n7757), .B(n7287), .ZN(n7830)
         );
  NAND2_X1 U8923 ( .A1(n7830), .A2(n10030), .ZN(n7288) );
  OAI21_X1 U8924 ( .B1(n10030), .B2(n7289), .A(n7288), .ZN(P2_U3454) );
  INV_X1 U8925 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U8926 ( .A1(n8374), .A2(n8391), .ZN(n7290) );
  NAND2_X1 U8927 ( .A1(n7291), .A2(n7290), .ZN(n7741) );
  NAND2_X1 U8928 ( .A1(n7741), .A2(n6542), .ZN(n7740) );
  NAND2_X1 U8929 ( .A1(n10015), .A2(n7590), .ZN(n7292) );
  NAND2_X1 U8930 ( .A1(n7740), .A2(n7292), .ZN(n7293) );
  NAND2_X1 U8931 ( .A1(n7293), .A2(n7296), .ZN(n7330) );
  OAI21_X1 U8932 ( .B1(n7293), .B2(n7296), .A(n7330), .ZN(n9994) );
  INV_X1 U8933 ( .A(n9994), .ZN(n7300) );
  NAND2_X1 U8934 ( .A1(n7294), .A2(n7295), .ZN(n7297) );
  XNOR2_X1 U8935 ( .A(n7297), .B(n7296), .ZN(n7298) );
  AOI222_X1 U8936 ( .A1(n8917), .A2(n7298), .B1(n8656), .B2(n8914), .C1(n8658), 
        .C2(n8912), .ZN(n9991) );
  INV_X1 U8937 ( .A(n7591), .ZN(n9986) );
  NAND2_X1 U8938 ( .A1(n7742), .A2(n10015), .ZN(n7743) );
  INV_X1 U8939 ( .A(n7339), .ZN(n7708) );
  AOI211_X1 U8940 ( .C1(n9986), .C2(n7743), .A(n10022), .B(n7708), .ZN(n9984)
         );
  AOI21_X1 U8941 ( .B1(n9090), .B2(n9986), .A(n9984), .ZN(n7299) );
  OAI211_X1 U8942 ( .C1(n9081), .C2(n7300), .A(n9991), .B(n7299), .ZN(n7307)
         );
  NAND2_X1 U8943 ( .A1(n7307), .A2(n10030), .ZN(n7301) );
  OAI21_X1 U8944 ( .B1(n10030), .B2(n7302), .A(n7301), .ZN(P2_U3466) );
  NAND2_X1 U8945 ( .A1(n7304), .A2(n7303), .ZN(n7306) );
  NAND2_X1 U8946 ( .A1(n7307), .A2(n4333), .ZN(n7308) );
  OAI21_X1 U8947 ( .B1(n4333), .B2(n6944), .A(n7308), .ZN(P2_U3525) );
  NAND2_X1 U8948 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8661), .ZN(n7309) );
  OAI21_X1 U8949 ( .B1(n8722), .B2(n8661), .A(n7309), .ZN(P2_U3581) );
  INV_X1 U8950 ( .A(n7310), .ZN(n7312) );
  OR2_X1 U8951 ( .A1(n7313), .A2(n9468), .ZN(n7368) );
  NAND2_X1 U8952 ( .A1(n9897), .A2(n7368), .ZN(n10214) );
  OAI21_X1 U8953 ( .B1(n7317), .B2(n7314), .A(n7410), .ZN(n9898) );
  INV_X2 U8954 ( .A(n10221), .ZN(n9616) );
  AOI22_X1 U8955 ( .A1(n9588), .A2(n9892), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9616), .ZN(n7328) );
  INV_X1 U8956 ( .A(n7316), .ZN(n7318) );
  NAND2_X1 U8957 ( .A1(n7318), .A2(n7317), .ZN(n7320) );
  NAND2_X1 U8958 ( .A1(n7320), .A2(n7319), .ZN(n7321) );
  NAND2_X1 U8959 ( .A1(n7321), .A2(n9603), .ZN(n7323) );
  AOI22_X1 U8960 ( .A1(n7362), .A2(n9542), .B1(n9540), .B2(n6757), .ZN(n7322)
         );
  NAND2_X1 U8961 ( .A1(n7323), .A2(n7322), .ZN(n9901) );
  NAND2_X1 U8962 ( .A1(n7324), .A2(n4997), .ZN(n9895) );
  INV_X1 U8963 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7325) );
  OAI22_X1 U8964 ( .A1(n9895), .A2(n10220), .B1(n9566), .B2(n7325), .ZN(n7326)
         );
  OAI21_X1 U8965 ( .B1(n9901), .B2(n7326), .A(n10221), .ZN(n7327) );
  OAI211_X1 U8966 ( .C1(n9595), .C2(n9898), .A(n7328), .B(n7327), .ZN(P1_U3290) );
  INV_X1 U8967 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7343) );
  INV_X1 U8968 ( .A(n8657), .ZN(n8376) );
  NAND2_X1 U8969 ( .A1(n7591), .A2(n8376), .ZN(n7329) );
  NAND2_X1 U8970 ( .A1(n7330), .A2(n7329), .ZN(n7714) );
  INV_X1 U8971 ( .A(n7701), .ZN(n7713) );
  NAND2_X1 U8972 ( .A1(n7714), .A2(n7713), .ZN(n7712) );
  OR2_X1 U8973 ( .A1(n7711), .A2(n8656), .ZN(n7331) );
  NAND2_X1 U8974 ( .A1(n7712), .A2(n7331), .ZN(n7332) );
  NAND2_X1 U8975 ( .A1(n7332), .A2(n7333), .ZN(n7633) );
  OAI21_X1 U8976 ( .B1(n7332), .B2(n7333), .A(n7633), .ZN(n7627) );
  INV_X1 U8977 ( .A(n7627), .ZN(n7341) );
  AOI21_X1 U8978 ( .B1(n7334), .B2(n7333), .A(n8930), .ZN(n7338) );
  OAI22_X1 U8979 ( .A1(n7335), .A2(n8934), .B1(n8932), .B2(n7529), .ZN(n7336)
         );
  AOI21_X1 U8980 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7630) );
  AOI21_X1 U8981 ( .B1(n7631), .B2(n7707), .A(n7641), .ZN(n7625) );
  AOI22_X1 U8982 ( .A1(n7625), .A2(n9091), .B1(n9090), .B2(n7631), .ZN(n7340)
         );
  OAI211_X1 U8983 ( .C1(n7341), .C2(n9081), .A(n7630), .B(n7340), .ZN(n7344)
         );
  NAND2_X1 U8984 ( .A1(n7344), .A2(n10030), .ZN(n7342) );
  OAI21_X1 U8985 ( .B1(n10030), .B2(n7343), .A(n7342), .ZN(P2_U3472) );
  NAND2_X1 U8986 ( .A1(n7344), .A2(n4333), .ZN(n7345) );
  OAI21_X1 U8987 ( .B1(n4333), .B2(n6976), .A(n7345), .ZN(P2_U3527) );
  XNOR2_X1 U8988 ( .A(n7556), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7349) );
  OAI21_X1 U8989 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7347), .A(n7346), .ZN(
        n7348) );
  AOI211_X1 U8990 ( .C1(n7349), .C2(n7348), .A(n9847), .B(n7555), .ZN(n7359)
         );
  OR2_X1 U8991 ( .A1(n7556), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U8992 ( .A1(n7556), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U8993 ( .A1(n7559), .A2(n7350), .ZN(n7351) );
  AOI21_X1 U8994 ( .B1(n7353), .B2(n7352), .A(n7351), .ZN(n7563) );
  INV_X1 U8995 ( .A(n7563), .ZN(n7355) );
  NAND3_X1 U8996 ( .A1(n7353), .A2(n7352), .A3(n7351), .ZN(n7354) );
  AOI21_X1 U8997 ( .B1(n7355), .B2(n7354), .A(n9858), .ZN(n7358) );
  NAND2_X1 U8998 ( .A1(n9853), .A2(n7556), .ZN(n7356) );
  NAND2_X1 U8999 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7963) );
  OAI211_X1 U9000 ( .C1(n9862), .C2(n4536), .A(n7356), .B(n7963), .ZN(n7357)
         );
  OR3_X1 U9001 ( .A1(n7359), .A2(n7358), .A3(n7357), .ZN(P1_U3253) );
  NAND2_X1 U9002 ( .A1(n7374), .A2(n7405), .ZN(n8234) );
  NAND2_X1 U9003 ( .A1(n7361), .A2(n7412), .ZN(n7366) );
  NOR2_X1 U9004 ( .A1(n7362), .A2(n7522), .ZN(n7392) );
  NAND2_X1 U9005 ( .A1(n7370), .A2(n7392), .ZN(n7364) );
  NAND2_X1 U9006 ( .A1(n7374), .A2(n4989), .ZN(n7363) );
  NAND2_X1 U9007 ( .A1(n7364), .A2(n7363), .ZN(n7413) );
  INV_X1 U9008 ( .A(n7413), .ZN(n7365) );
  NAND2_X1 U9009 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  XNOR2_X1 U9010 ( .A(n8195), .B(n7367), .ZN(n9913) );
  INV_X1 U9011 ( .A(n9913), .ZN(n7385) );
  NAND2_X1 U9012 ( .A1(n7369), .A2(n8240), .ZN(n7395) );
  INV_X1 U9013 ( .A(n7370), .ZN(n8191) );
  INV_X1 U9014 ( .A(n8195), .ZN(n7371) );
  XNOR2_X1 U9015 ( .A(n7470), .B(n7371), .ZN(n7372) );
  NAND2_X1 U9016 ( .A1(n7372), .A2(n9603), .ZN(n7377) );
  INV_X1 U9017 ( .A(n9897), .ZN(n7546) );
  NAND2_X1 U9018 ( .A1(n9305), .A2(n9542), .ZN(n7373) );
  OAI21_X1 U9019 ( .B1(n7374), .B2(n9925), .A(n7373), .ZN(n7375) );
  AOI21_X1 U9020 ( .B1(n9913), .B2(n7546), .A(n7375), .ZN(n7376) );
  AND2_X1 U9021 ( .A1(n7377), .A2(n7376), .ZN(n9915) );
  MUX2_X1 U9022 ( .A(n9915), .B(n6770), .S(n9616), .Z(n7384) );
  OR2_X1 U9023 ( .A1(n8325), .A2(n7378), .ZN(n7379) );
  AND2_X1 U9024 ( .A1(n7402), .A2(n7414), .ZN(n7380) );
  OR2_X1 U9025 ( .A1(n7380), .A2(n9929), .ZN(n9910) );
  OAI22_X1 U9026 ( .A1(n9571), .A2(n9910), .B1(n7381), .B2(n9566), .ZN(n7382)
         );
  AOI21_X1 U9027 ( .B1(n9588), .B2(n7414), .A(n7382), .ZN(n7383) );
  OAI211_X1 U9028 ( .C1(n7385), .C2(n9611), .A(n7384), .B(n7383), .ZN(P1_U3287) );
  AOI21_X1 U9029 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10213), .A(n7386), .ZN(
        n7391) );
  OAI21_X1 U9030 ( .B1(n9614), .B2(n9588), .A(n7387), .ZN(n7390) );
  INV_X1 U9031 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7388) );
  OR2_X1 U9032 ( .A1(n10221), .A2(n7388), .ZN(n7389) );
  OAI211_X1 U9033 ( .C1(n9616), .C2(n7391), .A(n7390), .B(n7389), .ZN(P1_U3291) );
  NOR2_X1 U9034 ( .A1(n7393), .A2(n7392), .ZN(n7394) );
  XNOR2_X1 U9035 ( .A(n7370), .B(n7394), .ZN(n9903) );
  OAI21_X1 U9036 ( .B1(n8191), .B2(n7395), .A(n7396), .ZN(n7400) );
  OAI22_X1 U9037 ( .A1(n7397), .A2(n9925), .B1(n9924), .B2(n9927), .ZN(n7399)
         );
  NOR2_X1 U9038 ( .A1(n9903), .A2(n9897), .ZN(n7398) );
  AOI211_X1 U9039 ( .C1(n9603), .C2(n7400), .A(n7399), .B(n7398), .ZN(n9905)
         );
  MUX2_X1 U9040 ( .A(n6837), .B(n9905), .S(n10221), .Z(n7407) );
  INV_X1 U9041 ( .A(n7401), .ZN(n7403) );
  OAI21_X1 U9042 ( .B1(n7403), .B2(n4989), .A(n7402), .ZN(n9904) );
  OAI22_X1 U9043 ( .A1(n9571), .A2(n9904), .B1(n9566), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7404) );
  AOI21_X1 U9044 ( .B1(n9588), .B2(n7405), .A(n7404), .ZN(n7406) );
  OAI211_X1 U9045 ( .C1(n9903), .C2(n9611), .A(n7407), .B(n7406), .ZN(P1_U3288) );
  INV_X1 U9046 ( .A(n7408), .ZN(n7487) );
  AOI22_X1 U9047 ( .A1(n8681), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9127), .ZN(n7409) );
  OAI21_X1 U9048 ( .B1(n7487), .B2(n7807), .A(n7409), .ZN(P2_U3340) );
  NAND4_X1 U9049 ( .A1(n7412), .A2(n8195), .A3(n7411), .A4(n7410), .ZN(n7416)
         );
  NAND2_X1 U9050 ( .A1(n7413), .A2(n8195), .ZN(n7415) );
  NAND3_X1 U9051 ( .A1(n7416), .A2(n7415), .A3(n5125), .ZN(n7475) );
  NAND2_X2 U9052 ( .A1(n9933), .A2(n9304), .ZN(n8292) );
  NAND2_X1 U9053 ( .A1(n9305), .A2(n8067), .ZN(n7476) );
  AND2_X1 U9054 ( .A1(n7477), .A2(n7476), .ZN(n7417) );
  OR2_X2 U9055 ( .A1(n7607), .A2(n7495), .ZN(n8275) );
  NAND2_X1 U9056 ( .A1(n7477), .A2(n7476), .ZN(n7419) );
  NAND2_X1 U9057 ( .A1(n8066), .A2(n8067), .ZN(n8193) );
  NAND2_X1 U9058 ( .A1(n9933), .A2(n9926), .ZN(n7418) );
  NAND2_X1 U9059 ( .A1(n7444), .A2(n7446), .ZN(n7421) );
  OR2_X1 U9060 ( .A1(n7607), .A2(n9303), .ZN(n7420) );
  OR2_X1 U9061 ( .A1(n7536), .A2(n7611), .ZN(n8085) );
  NAND2_X1 U9062 ( .A1(n7536), .A2(n7611), .ZN(n8084) );
  NAND2_X1 U9063 ( .A1(n8085), .A2(n8084), .ZN(n7424) );
  OAI21_X1 U9064 ( .B1(n7422), .B2(n7424), .A(n7423), .ZN(n9946) );
  AND3_X1 U9065 ( .A1(n8194), .A2(n8193), .A3(n8068), .ZN(n8247) );
  NAND2_X1 U9066 ( .A1(n8292), .A2(n8291), .ZN(n8196) );
  AND2_X1 U9067 ( .A1(n8194), .A2(n8196), .ZN(n8246) );
  INV_X1 U9068 ( .A(n7424), .ZN(n8198) );
  XNOR2_X1 U9069 ( .A(n7540), .B(n8198), .ZN(n7427) );
  NAND2_X1 U9070 ( .A1(n9301), .A2(n9542), .ZN(n7425) );
  OAI21_X1 U9071 ( .B1(n7495), .B2(n9925), .A(n7425), .ZN(n7426) );
  AOI21_X1 U9072 ( .B1(n7427), .B2(n9603), .A(n7426), .ZN(n9955) );
  OAI21_X1 U9073 ( .B1(n9897), .B2(n9946), .A(n9955), .ZN(n7428) );
  NAND2_X1 U9074 ( .A1(n7428), .A2(n10221), .ZN(n7435) );
  NOR2_X2 U9075 ( .A1(n7480), .A2(n7607), .ZN(n7451) );
  INV_X1 U9076 ( .A(n7536), .ZN(n9948) );
  NOR2_X1 U9077 ( .A1(n7451), .A2(n9948), .ZN(n7430) );
  OR2_X1 U9078 ( .A1(n7547), .A2(n7430), .ZN(n9950) );
  INV_X1 U9079 ( .A(n9950), .ZN(n7433) );
  AOI22_X1 U9080 ( .A1(n9616), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7498), .B2(
        n10213), .ZN(n7431) );
  OAI21_X1 U9081 ( .B1(n9948), .B2(n9609), .A(n7431), .ZN(n7432) );
  AOI21_X1 U9082 ( .B1(n7433), .B2(n9614), .A(n7432), .ZN(n7434) );
  OAI211_X1 U9083 ( .C1(n9946), .C2(n9611), .A(n7435), .B(n7434), .ZN(P1_U3283) );
  NAND2_X1 U9084 ( .A1(n7436), .A2(n4383), .ZN(n7437) );
  NAND2_X1 U9085 ( .A1(n7437), .A2(n7446), .ZN(n7439) );
  NAND2_X1 U9086 ( .A1(n7439), .A2(n7438), .ZN(n7440) );
  NAND2_X1 U9087 ( .A1(n7440), .A2(n9603), .ZN(n7442) );
  INV_X1 U9088 ( .A(n7611), .ZN(n9302) );
  AOI22_X1 U9089 ( .A1(n9302), .A2(n9542), .B1(n9540), .B2(n9304), .ZN(n7441)
         );
  NAND2_X1 U9090 ( .A1(n7442), .A2(n7441), .ZN(n9944) );
  INV_X1 U9091 ( .A(n9944), .ZN(n7457) );
  INV_X1 U9092 ( .A(n9595), .ZN(n9573) );
  INV_X1 U9093 ( .A(n7444), .ZN(n7445) );
  NAND2_X1 U9094 ( .A1(n7443), .A2(n7445), .ZN(n7447) );
  XNOR2_X1 U9095 ( .A(n7447), .B(n7446), .ZN(n9939) );
  NOR2_X1 U9096 ( .A1(n7448), .A2(n10220), .ZN(n9554) );
  INV_X1 U9097 ( .A(n9554), .ZN(n9591) );
  NAND2_X1 U9098 ( .A1(n7480), .A2(n7607), .ZN(n7449) );
  NAND2_X1 U9099 ( .A1(n7449), .A2(n4997), .ZN(n7450) );
  OR2_X1 U9100 ( .A1(n7451), .A2(n7450), .ZN(n9940) );
  INV_X1 U9101 ( .A(n7614), .ZN(n7452) );
  OAI22_X1 U9102 ( .A1(n10221), .A2(n6813), .B1(n7452), .B2(n9566), .ZN(n7453)
         );
  AOI21_X1 U9103 ( .B1(n9588), .B2(n7607), .A(n7453), .ZN(n7454) );
  OAI21_X1 U9104 ( .B1(n9591), .B2(n9940), .A(n7454), .ZN(n7455) );
  AOI21_X1 U9105 ( .B1(n9573), .B2(n9939), .A(n7455), .ZN(n7456) );
  OAI21_X1 U9106 ( .B1(n7457), .B2(n9616), .A(n7456), .ZN(P1_U3284) );
  XNOR2_X1 U9107 ( .A(n7599), .B(n7460), .ZN(n7461) );
  XNOR2_X1 U9108 ( .A(n7459), .B(n7461), .ZN(n7467) );
  AOI22_X1 U9109 ( .A1(n9272), .A2(n9305), .B1(n7429), .B2(n9288), .ZN(n7465)
         );
  NAND2_X1 U9110 ( .A1(n9271), .A2(n7481), .ZN(n7464) );
  NAND2_X1 U9111 ( .A1(n9284), .A2(n9303), .ZN(n7462) );
  NAND4_X1 U9112 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .ZN(n7466)
         );
  AOI21_X1 U9113 ( .B1(n7467), .B2(n5905), .A(n7466), .ZN(n7468) );
  INV_X1 U9114 ( .A(n7468), .ZN(P1_U3237) );
  INV_X1 U9115 ( .A(n8068), .ZN(n7469) );
  NAND3_X1 U9116 ( .A1(n9919), .A2(n7472), .A3(n9918), .ZN(n9917) );
  NAND2_X1 U9117 ( .A1(n9917), .A2(n8193), .ZN(n7473) );
  XNOR2_X1 U9118 ( .A(n7473), .B(n7477), .ZN(n7474) );
  INV_X1 U9119 ( .A(n9603), .ZN(n9923) );
  OAI222_X1 U9120 ( .A1(n9927), .A2(n7495), .B1(n9925), .B2(n8066), .C1(n7474), 
        .C2(n9923), .ZN(n9935) );
  INV_X1 U9121 ( .A(n9935), .ZN(n7486) );
  OR2_X1 U9122 ( .A1(n7475), .A2(n7472), .ZN(n10216) );
  NAND2_X1 U9123 ( .A1(n10216), .A2(n7476), .ZN(n7478) );
  INV_X1 U9124 ( .A(n7477), .ZN(n8077) );
  XNOR2_X1 U9125 ( .A(n7478), .B(n8077), .ZN(n9937) );
  NAND2_X1 U9126 ( .A1(n9928), .A2(n7429), .ZN(n7479) );
  NAND2_X1 U9127 ( .A1(n7480), .A2(n7479), .ZN(n9934) );
  NAND2_X1 U9128 ( .A1(n9588), .A2(n7429), .ZN(n7483) );
  AOI22_X1 U9129 ( .A1(n9616), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7481), .B2(
        n10213), .ZN(n7482) );
  OAI211_X1 U9130 ( .C1(n9571), .C2(n9934), .A(n7483), .B(n7482), .ZN(n7484)
         );
  AOI21_X1 U9131 ( .B1(n9937), .B2(n9573), .A(n7484), .ZN(n7485) );
  OAI21_X1 U9132 ( .B1(n7486), .B2(n9616), .A(n7485), .ZN(P1_U3285) );
  INV_X1 U9133 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7488) );
  INV_X1 U9134 ( .A(n9854), .ZN(n9340) );
  OAI222_X1 U9135 ( .A1(n9755), .A2(n7488), .B1(n9752), .B2(n7487), .C1(
        P1_U3084), .C2(n9340), .ZN(P1_U3335) );
  XNOR2_X1 U9136 ( .A(n7490), .B(n7489), .ZN(n7491) );
  XNOR2_X1 U9137 ( .A(n7492), .B(n7491), .ZN(n7500) );
  NOR2_X1 U9138 ( .A1(n9235), .A2(n9948), .ZN(n7497) );
  NAND2_X1 U9139 ( .A1(n9284), .A2(n9301), .ZN(n7494) );
  OAI211_X1 U9140 ( .C1(n7495), .C2(n9282), .A(n7494), .B(n7493), .ZN(n7496)
         );
  AOI211_X1 U9141 ( .C1(n7498), .C2(n9271), .A(n7497), .B(n7496), .ZN(n7499)
         );
  OAI21_X1 U9142 ( .B1(n7500), .B2(n9278), .A(n7499), .ZN(P1_U3219) );
  INV_X1 U9143 ( .A(n8584), .ZN(n8637) );
  AOI22_X1 U9144 ( .A1(n8637), .A2(n6469), .B1(n8636), .B2(n6468), .ZN(n7508)
         );
  XNOR2_X1 U9145 ( .A(n8598), .B(n8593), .ZN(n7502) );
  INV_X1 U9146 ( .A(n7502), .ZN(n7503) );
  NOR2_X1 U9147 ( .A1(n7502), .A2(n7501), .ZN(n8592) );
  INV_X1 U9148 ( .A(n8592), .ZN(n8600) );
  OAI21_X1 U9149 ( .B1(n6015), .B2(n7503), .A(n8600), .ZN(n7506) );
  NAND2_X1 U9150 ( .A1(n7505), .A2(n7504), .ZN(n8596) );
  AOI22_X1 U9151 ( .A1(n8631), .A2(n7506), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8596), .ZN(n7507) );
  OAI211_X1 U9152 ( .C1(n7509), .C2(n8617), .A(n7508), .B(n7507), .ZN(P2_U3224) );
  NAND2_X1 U9153 ( .A1(n8631), .A2(n6331), .ZN(n8608) );
  OAI22_X1 U9154 ( .A1(n7510), .A2(n8608), .B1(n8627), .B2(n10010), .ZN(n7512)
         );
  NAND2_X1 U9155 ( .A1(n7512), .A2(n7511), .ZN(n7514) );
  NOR2_X1 U9156 ( .A1(n8934), .A2(n8599), .ZN(n7733) );
  AOI22_X1 U9157 ( .A1(n8622), .A2(n7733), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8596), .ZN(n7513) );
  OAI211_X1 U9158 ( .C1(n8617), .C2(n10010), .A(n7514), .B(n7513), .ZN(
        P2_U3234) );
  INV_X1 U9159 ( .A(n7515), .ZN(n7524) );
  NOR2_X1 U9160 ( .A1(n9566), .A2(n9822), .ZN(n7516) );
  AOI21_X1 U9161 ( .B1(n9616), .B2(P1_REG2_REG_2__SCAN_IN), .A(n7516), .ZN(
        n7517) );
  OAI21_X1 U9162 ( .B1(n9571), .B2(n7518), .A(n7517), .ZN(n7521) );
  NOR2_X1 U9163 ( .A1(n7519), .A2(n9611), .ZN(n7520) );
  AOI211_X1 U9164 ( .C1(n9588), .C2(n7522), .A(n7521), .B(n7520), .ZN(n7523)
         );
  OAI21_X1 U9165 ( .B1(n9616), .B2(n7524), .A(n7523), .ZN(P1_U3289) );
  XNOR2_X1 U9166 ( .A(n7526), .B(n7525), .ZN(n7533) );
  INV_X1 U9167 ( .A(n7527), .ZN(n7528) );
  OAI21_X1 U9168 ( .B1(n8624), .B2(n7620), .A(n7528), .ZN(n7531) );
  INV_X1 U9169 ( .A(n7631), .ZN(n7622) );
  OAI22_X1 U9170 ( .A1(n7622), .A2(n8617), .B1(n8584), .B2(n7529), .ZN(n7530)
         );
  AOI211_X1 U9171 ( .C1(n8636), .C2(n8654), .A(n7531), .B(n7530), .ZN(n7532)
         );
  OAI21_X1 U9172 ( .B1(n7533), .B2(n8627), .A(n7532), .ZN(P2_U3215) );
  INV_X1 U9173 ( .A(n7534), .ZN(n8392) );
  OAI222_X1 U9174 ( .A1(n9125), .A2(n7535), .B1(n7807), .B2(n8392), .C1(
        P2_U3152), .C2(n6532), .ZN(P2_U3339) );
  NAND2_X1 U9175 ( .A1(n7536), .A2(n9302), .ZN(n7537) );
  INV_X1 U9176 ( .A(n9301), .ZN(n7799) );
  OR2_X1 U9177 ( .A1(n9720), .A2(n7799), .ZN(n8086) );
  NAND2_X1 U9178 ( .A1(n9720), .A2(n7799), .ZN(n8089) );
  NAND2_X1 U9179 ( .A1(n8086), .A2(n8089), .ZN(n8201) );
  INV_X1 U9180 ( .A(n8201), .ZN(n7539) );
  XNOR2_X1 U9181 ( .A(n7723), .B(n7539), .ZN(n7551) );
  OAI22_X1 U9182 ( .A1(n7611), .A2(n9925), .B1(n7777), .B2(n9927), .ZN(n7545)
         );
  INV_X1 U9183 ( .A(n7717), .ZN(n7542) );
  AOI211_X1 U9184 ( .C1(n8201), .C2(n7543), .A(n9923), .B(n7542), .ZN(n7544)
         );
  AOI211_X1 U9185 ( .C1(n7551), .C2(n7546), .A(n7545), .B(n7544), .ZN(n9723)
         );
  INV_X1 U9186 ( .A(n7547), .ZN(n7549) );
  INV_X1 U9187 ( .A(n9720), .ZN(n7774) );
  INV_X1 U9188 ( .A(n7720), .ZN(n7548) );
  AOI21_X1 U9189 ( .B1(n9720), .B2(n7549), .A(n7548), .ZN(n9721) );
  AOI22_X1 U9190 ( .A1(n9616), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7771), .B2(
        n10213), .ZN(n7550) );
  OAI21_X1 U9191 ( .B1(n7774), .B2(n9609), .A(n7550), .ZN(n7553) );
  INV_X1 U9192 ( .A(n7551), .ZN(n9724) );
  NOR2_X1 U9193 ( .A1(n9724), .A2(n9611), .ZN(n7552) );
  AOI211_X1 U9194 ( .C1(n9721), .C2(n9614), .A(n7553), .B(n7552), .ZN(n7554)
         );
  OAI21_X1 U9195 ( .B1(n9723), .B2(n9616), .A(n7554), .ZN(P1_U3282) );
  XNOR2_X1 U9196 ( .A(n7979), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7557) );
  AOI211_X1 U9197 ( .C1(n7558), .C2(n7557), .A(n9847), .B(n7978), .ZN(n7570)
         );
  INV_X1 U9198 ( .A(n7559), .ZN(n7562) );
  OR2_X1 U9199 ( .A1(n7979), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7973) );
  NAND2_X1 U9200 ( .A1(n7979), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7560) );
  AND2_X1 U9201 ( .A1(n7973), .A2(n7560), .ZN(n7561) );
  OAI21_X1 U9202 ( .B1(n7563), .B2(n7562), .A(n7561), .ZN(n7974) );
  OR3_X1 U9203 ( .A1(n7563), .A2(n7562), .A3(n7561), .ZN(n7564) );
  AOI21_X1 U9204 ( .B1(n7974), .B2(n7564), .A(n9858), .ZN(n7569) );
  INV_X1 U9205 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U9206 ( .A1(n7565), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9240) );
  AOI21_X1 U9207 ( .B1(n9853), .B2(n7979), .A(n9240), .ZN(n7566) );
  OAI21_X1 U9208 ( .B1(n7567), .B2(n9862), .A(n7566), .ZN(n7568) );
  OR3_X1 U9209 ( .A1(n7570), .A2(n7569), .A3(n7568), .ZN(P1_U3254) );
  XNOR2_X1 U9210 ( .A(n7572), .B(n7571), .ZN(n7577) );
  OAI22_X1 U9211 ( .A1(n8624), .A2(n7643), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7573), .ZN(n7575) );
  INV_X1 U9212 ( .A(n9089), .ZN(n7645) );
  OAI22_X1 U9213 ( .A1(n7645), .A2(n8617), .B1(n8584), .B2(n7702), .ZN(n7574)
         );
  AOI211_X1 U9214 ( .C1(n8636), .C2(n8653), .A(n7575), .B(n7574), .ZN(n7576)
         );
  OAI21_X1 U9215 ( .B1(n8627), .B2(n7577), .A(n7576), .ZN(P2_U3223) );
  OAI21_X1 U9216 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(n7585) );
  INV_X1 U9217 ( .A(n7711), .ZN(n10021) );
  OAI22_X1 U9218 ( .A1(n10021), .A2(n8617), .B1(n8584), .B2(n8376), .ZN(n7584)
         );
  NAND2_X1 U9219 ( .A1(n8636), .A2(n8655), .ZN(n7582) );
  OAI211_X1 U9220 ( .C1(n8624), .C2(n7705), .A(n7582), .B(n7581), .ZN(n7583)
         );
  AOI211_X1 U9221 ( .C1(n8631), .C2(n7585), .A(n7584), .B(n7583), .ZN(n7586)
         );
  INV_X1 U9222 ( .A(n7586), .ZN(P2_U3241) );
  OAI21_X1 U9223 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7596) );
  OAI22_X1 U9224 ( .A1(n7591), .A2(n8617), .B1(n8584), .B2(n7590), .ZN(n7595)
         );
  NAND2_X1 U9225 ( .A1(n8636), .A2(n8656), .ZN(n7593) );
  OAI211_X1 U9226 ( .C1(n8624), .C2(n9989), .A(n7593), .B(n7592), .ZN(n7594)
         );
  AOI211_X1 U9227 ( .C1(n8631), .C2(n7596), .A(n7595), .B(n7594), .ZN(n7597)
         );
  INV_X1 U9228 ( .A(n7597), .ZN(P2_U3229) );
  INV_X1 U9229 ( .A(n7459), .ZN(n7600) );
  OAI21_X1 U9230 ( .B1(n7600), .B2(n7599), .A(n7598), .ZN(n7601) );
  OAI21_X1 U9231 ( .B1(n7602), .B2(n7459), .A(n7601), .ZN(n7606) );
  XOR2_X1 U9232 ( .A(n7604), .B(n7603), .Z(n7605) );
  XNOR2_X1 U9233 ( .A(n7606), .B(n7605), .ZN(n7616) );
  INV_X1 U9234 ( .A(n7607), .ZN(n9941) );
  NOR2_X1 U9235 ( .A1(n9235), .A2(n9941), .ZN(n7613) );
  NAND2_X1 U9236 ( .A1(n9272), .A2(n9304), .ZN(n7610) );
  INV_X1 U9237 ( .A(n7608), .ZN(n7609) );
  OAI211_X1 U9238 ( .C1(n7611), .C2(n9275), .A(n7610), .B(n7609), .ZN(n7612)
         );
  AOI211_X1 U9239 ( .C1(n7614), .C2(n9271), .A(n7613), .B(n7612), .ZN(n7615)
         );
  OAI21_X1 U9240 ( .B1(n7616), .B2(n9278), .A(n7615), .ZN(P1_U3211) );
  NAND2_X1 U9241 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  OAI22_X1 U9242 ( .A1(n9996), .A2(n7621), .B1(n7620), .B2(n9990), .ZN(n7624)
         );
  NOR2_X1 U9243 ( .A1(n8948), .A2(n7622), .ZN(n7623) );
  AOI211_X1 U9244 ( .C1(n7625), .C2(n8944), .A(n7624), .B(n7623), .ZN(n7629)
         );
  OR2_X1 U9245 ( .A1(n7626), .A2(n6532), .ZN(n7648) );
  NAND2_X1 U9246 ( .A1(n7635), .A2(n7648), .ZN(n9995) );
  NAND2_X1 U9247 ( .A1(n8965), .A2(n7627), .ZN(n7628) );
  OAI211_X1 U9248 ( .C1(n9998), .C2(n7630), .A(n7629), .B(n7628), .ZN(P2_U3289) );
  OR2_X1 U9249 ( .A1(n7631), .A2(n8655), .ZN(n7632) );
  NOR2_X1 U9250 ( .A1(n7678), .A2(n7634), .ZN(n7652) );
  AOI21_X1 U9251 ( .B1(n7634), .B2(n7678), .A(n7652), .ZN(n9088) );
  INV_X1 U9252 ( .A(n7635), .ZN(n7659) );
  NAND2_X1 U9253 ( .A1(n7636), .A2(n7680), .ZN(n7637) );
  AOI21_X1 U9254 ( .B1(n7638), .B2(n7637), .A(n8930), .ZN(n7640) );
  OAI22_X1 U9255 ( .A1(n7669), .A2(n8934), .B1(n8932), .B2(n7702), .ZN(n7639)
         );
  AOI211_X1 U9256 ( .C1(n9088), .C2(n7659), .A(n7640), .B(n7639), .ZN(n9094)
         );
  OR2_X1 U9257 ( .A1(n7641), .A2(n7645), .ZN(n7642) );
  AND2_X1 U9258 ( .A1(n7642), .A2(n7661), .ZN(n9092) );
  OAI22_X1 U9259 ( .A1(n9996), .A2(n7644), .B1(n7643), .B2(n9990), .ZN(n7647)
         );
  NOR2_X1 U9260 ( .A1(n8948), .A2(n7645), .ZN(n7646) );
  AOI211_X1 U9261 ( .C1(n9092), .C2(n8944), .A(n7647), .B(n7646), .ZN(n7651)
         );
  INV_X1 U9262 ( .A(n7648), .ZN(n7649) );
  AND2_X1 U9263 ( .A1(n9996), .A2(n7649), .ZN(n8863) );
  NAND2_X1 U9264 ( .A1(n9088), .A2(n8863), .ZN(n7650) );
  OAI211_X1 U9265 ( .C1(n9094), .C2(n9998), .A(n7651), .B(n7650), .ZN(P2_U3288) );
  AND2_X1 U9266 ( .A1(n9089), .A2(n8654), .ZN(n7679) );
  NOR2_X1 U9267 ( .A1(n7652), .A2(n7679), .ZN(n7653) );
  XNOR2_X1 U9268 ( .A(n7653), .B(n7654), .ZN(n9082) );
  XNOR2_X1 U9269 ( .A(n7655), .B(n7654), .ZN(n7657) );
  AOI22_X1 U9270 ( .A1(n8914), .A2(n8652), .B1(n8912), .B2(n8654), .ZN(n7656)
         );
  OAI21_X1 U9271 ( .B1(n7657), .B2(n8930), .A(n7656), .ZN(n7658) );
  AOI21_X1 U9272 ( .B1(n9082), .B2(n7659), .A(n7658), .ZN(n9086) );
  INV_X1 U9273 ( .A(n7672), .ZN(n7660) );
  AOI21_X1 U9274 ( .B1(n9083), .B2(n7661), .A(n7660), .ZN(n9084) );
  OAI22_X1 U9275 ( .A1(n9996), .A2(n7662), .B1(n7824), .B2(n9990), .ZN(n7665)
         );
  INV_X1 U9276 ( .A(n9083), .ZN(n7663) );
  NOR2_X1 U9277 ( .A1(n8948), .A2(n7663), .ZN(n7664) );
  AOI211_X1 U9278 ( .C1(n9084), .C2(n8944), .A(n7665), .B(n7664), .ZN(n7667)
         );
  NAND2_X1 U9279 ( .A1(n9082), .A2(n8863), .ZN(n7666) );
  OAI211_X1 U9280 ( .C1(n9086), .C2(n9998), .A(n7667), .B(n7666), .ZN(P2_U3287) );
  AOI21_X1 U9281 ( .B1(n7668), .B2(n7686), .A(n8930), .ZN(n7671) );
  OAI22_X1 U9282 ( .A1(n8030), .A2(n8934), .B1(n8932), .B2(n7669), .ZN(n7858)
         );
  AOI21_X1 U9283 ( .B1(n7671), .B2(n7670), .A(n7858), .ZN(n9079) );
  OAI22_X1 U9284 ( .A1(n9996), .A2(n7673), .B1(n7859), .B2(n9990), .ZN(n7676)
         );
  INV_X1 U9285 ( .A(n9077), .ZN(n7674) );
  NOR2_X1 U9286 ( .A1(n8948), .A2(n7674), .ZN(n7675) );
  AOI211_X1 U9287 ( .C1(n9076), .C2(n8969), .A(n7676), .B(n7675), .ZN(n7689)
         );
  NOR2_X1 U9288 ( .A1(n7682), .A2(n7679), .ZN(n7677) );
  OR2_X1 U9289 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  OAI22_X1 U9290 ( .A1(n7682), .A2(n7681), .B1(n9083), .B2(n8653), .ZN(n7683)
         );
  INV_X1 U9291 ( .A(n7683), .ZN(n7684) );
  INV_X1 U9292 ( .A(n7874), .ZN(n7687) );
  INV_X1 U9293 ( .A(n7686), .ZN(n7869) );
  NOR2_X1 U9294 ( .A1(n7874), .A2(n7869), .ZN(n7816) );
  INV_X1 U9295 ( .A(n7816), .ZN(n7685) );
  OAI21_X1 U9296 ( .B1(n7687), .B2(n7686), .A(n7685), .ZN(n9080) );
  OR2_X1 U9297 ( .A1(n9080), .A2(n8890), .ZN(n7688) );
  OAI211_X1 U9298 ( .C1(n9079), .C2(n9998), .A(n7689), .B(n7688), .ZN(P2_U3286) );
  XNOR2_X1 U9299 ( .A(n7910), .B(n7911), .ZN(n7912) );
  XNOR2_X1 U9300 ( .A(n7912), .B(n6236), .ZN(n7699) );
  OAI21_X1 U9301 ( .B1(n7693), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7692), .ZN(
        n7902) );
  XOR2_X1 U9302 ( .A(n7911), .B(n7902), .Z(n7905) );
  XNOR2_X1 U9303 ( .A(n7905), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n7697) );
  AND2_X1 U9304 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7694) );
  AOI21_X1 U9305 ( .B1(n9975), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7694), .ZN(
        n7695) );
  OAI21_X1 U9306 ( .B1(n9977), .B2(n7903), .A(n7695), .ZN(n7696) );
  AOI21_X1 U9307 ( .B1(n7697), .B2(n9973), .A(n7696), .ZN(n7698) );
  OAI21_X1 U9308 ( .B1(n7699), .B2(n9976), .A(n7698), .ZN(P2_U3260) );
  XNOR2_X1 U9309 ( .A(n7700), .B(n7701), .ZN(n7704) );
  OAI22_X1 U9310 ( .A1(n8376), .A2(n8932), .B1(n8934), .B2(n7702), .ZN(n7703)
         );
  AOI21_X1 U9311 ( .B1(n7704), .B2(n8917), .A(n7703), .ZN(n10024) );
  OAI22_X1 U9312 ( .A1(n9996), .A2(n7706), .B1(n7705), .B2(n9990), .ZN(n7710)
         );
  INV_X1 U9313 ( .A(n8944), .ZN(n8713) );
  OAI21_X1 U9314 ( .B1(n7708), .B2(n10021), .A(n7707), .ZN(n10023) );
  NOR2_X1 U9315 ( .A1(n8713), .A2(n10023), .ZN(n7709) );
  AOI211_X1 U9316 ( .C1(n8963), .C2(n7711), .A(n7710), .B(n7709), .ZN(n7716)
         );
  OAI21_X1 U9317 ( .B1(n7714), .B2(n7713), .A(n7712), .ZN(n10027) );
  NAND2_X1 U9318 ( .A1(n8965), .A2(n10027), .ZN(n7715) );
  OAI211_X1 U9319 ( .C1(n9998), .C2(n10024), .A(n7716), .B(n7715), .ZN(
        P2_U3290) );
  NAND2_X1 U9320 ( .A1(n9715), .A2(n7777), .ZN(n8088) );
  XOR2_X1 U9321 ( .A(n7775), .B(n8200), .Z(n7718) );
  AOI222_X1 U9322 ( .A1(n9603), .A2(n7718), .B1(n9301), .B2(n9540), .C1(n9299), 
        .C2(n9542), .ZN(n9717) );
  INV_X1 U9323 ( .A(n7781), .ZN(n7719) );
  AOI211_X1 U9324 ( .C1(n9715), .C2(n7720), .A(n9949), .B(n7719), .ZN(n9714)
         );
  INV_X1 U9325 ( .A(n9715), .ZN(n7796) );
  AOI22_X1 U9326 ( .A1(n9616), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7802), .B2(
        n10213), .ZN(n7721) );
  OAI21_X1 U9327 ( .B1(n7796), .B2(n9609), .A(n7721), .ZN(n7729) );
  OR2_X1 U9328 ( .A1(n9720), .A2(n9301), .ZN(n7722) );
  NAND2_X1 U9329 ( .A1(n9720), .A2(n9301), .ZN(n7724) );
  INV_X1 U9330 ( .A(n8200), .ZN(n7725) );
  INV_X1 U9331 ( .A(n7779), .ZN(n7726) );
  AOI21_X1 U9332 ( .B1(n8200), .B2(n7727), .A(n7726), .ZN(n9718) );
  NOR2_X1 U9333 ( .A1(n9718), .A2(n9595), .ZN(n7728) );
  AOI211_X1 U9334 ( .C1(n9714), .C2(n9554), .A(n7729), .B(n7728), .ZN(n7730)
         );
  OAI21_X1 U9335 ( .B1(n9616), .B2(n9717), .A(n7730), .ZN(P1_U3281) );
  NAND2_X1 U9336 ( .A1(n7732), .A2(n7731), .ZN(n10012) );
  INV_X1 U9337 ( .A(n10012), .ZN(n7739) );
  AOI21_X1 U9338 ( .B1(n8917), .B2(n10012), .A(n7733), .ZN(n10008) );
  INV_X1 U9339 ( .A(n9990), .ZN(n8955) );
  NAND2_X1 U9340 ( .A1(n8955), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7734) );
  AOI21_X1 U9341 ( .B1(n10008), .B2(n7734), .A(n9998), .ZN(n7735) );
  AOI21_X1 U9342 ( .B1(n9998), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7735), .ZN(
        n7738) );
  OAI21_X1 U9343 ( .B1(n8944), .B2(n8963), .A(n7736), .ZN(n7737) );
  OAI211_X1 U9344 ( .C1(n7739), .C2(n8890), .A(n7738), .B(n7737), .ZN(P2_U3296) );
  OAI21_X1 U9345 ( .B1(n7741), .B2(n6542), .A(n7740), .ZN(n10019) );
  INV_X1 U9346 ( .A(n10019), .ZN(n7755) );
  INV_X1 U9347 ( .A(n7742), .ZN(n7745) );
  INV_X1 U9348 ( .A(n7743), .ZN(n7744) );
  AOI21_X1 U9349 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n10014) );
  AOI22_X1 U9350 ( .A1(n8944), .A2(n10014), .B1(n8963), .B2(n7746), .ZN(n7754)
         );
  OAI211_X1 U9351 ( .C1(n7748), .C2(n7747), .A(n7294), .B(n8917), .ZN(n7751)
         );
  OAI22_X1 U9352 ( .A1(n8374), .A2(n8932), .B1(n8934), .B2(n8376), .ZN(n7749)
         );
  INV_X1 U9353 ( .A(n7749), .ZN(n7750) );
  NAND2_X1 U9354 ( .A1(n7751), .A2(n7750), .ZN(n10018) );
  OAI22_X1 U9355 ( .A1(n9996), .A2(n6044), .B1(n8377), .B2(n9990), .ZN(n7752)
         );
  AOI21_X1 U9356 ( .B1(n9996), .B2(n10018), .A(n7752), .ZN(n7753) );
  OAI211_X1 U9357 ( .C1(n7755), .C2(n8890), .A(n7754), .B(n7753), .ZN(P2_U3292) );
  OAI22_X1 U9358 ( .A1(n9998), .A2(n7757), .B1(n7756), .B2(n9990), .ZN(n7758)
         );
  AOI21_X1 U9359 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n9998), .A(n7758), .ZN(
        n7762) );
  AOI22_X1 U9360 ( .A1(n8944), .A2(n7760), .B1(n8963), .B2(n7759), .ZN(n7761)
         );
  OAI211_X1 U9361 ( .C1(n7763), .C2(n8890), .A(n7762), .B(n7761), .ZN(P2_U3295) );
  OAI21_X1 U9362 ( .B1(n7766), .B2(n7765), .A(n7764), .ZN(n7767) );
  NAND2_X1 U9363 ( .A1(n7767), .A2(n5905), .ZN(n7773) );
  AOI21_X1 U9364 ( .B1(n9272), .B2(n9302), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9365 ( .B1(n7777), .B2(n9275), .A(n7769), .ZN(n7770) );
  AOI21_X1 U9366 ( .B1(n7771), .B2(n9271), .A(n7770), .ZN(n7772) );
  OAI211_X1 U9367 ( .C1(n7774), .C2(n9235), .A(n7773), .B(n7772), .ZN(P1_U3229) );
  INV_X1 U9368 ( .A(n9299), .ZN(n7965) );
  OR2_X1 U9369 ( .A1(n7893), .A2(n7965), .ZN(n8092) );
  NAND2_X1 U9370 ( .A1(n7893), .A2(n7965), .ZN(n8094) );
  XNOR2_X1 U9371 ( .A(n7842), .B(n8204), .ZN(n7776) );
  OAI222_X1 U9372 ( .A1(n9927), .A2(n9597), .B1(n9925), .B2(n7777), .C1(n9923), 
        .C2(n7776), .ZN(n7895) );
  INV_X1 U9373 ( .A(n7895), .ZN(n7787) );
  INV_X1 U9374 ( .A(n7777), .ZN(n9300) );
  OR2_X1 U9375 ( .A1(n9715), .A2(n9300), .ZN(n7778) );
  NAND2_X1 U9376 ( .A1(n7779), .A2(n7778), .ZN(n7837) );
  INV_X1 U9377 ( .A(n8204), .ZN(n7780) );
  XNOR2_X1 U9378 ( .A(n7837), .B(n7780), .ZN(n7897) );
  NAND2_X1 U9379 ( .A1(n7781), .A2(n7893), .ZN(n7782) );
  NAND2_X1 U9380 ( .A1(n7848), .A2(n7782), .ZN(n7894) );
  AOI22_X1 U9381 ( .A1(n9616), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7889), .B2(
        n10213), .ZN(n7784) );
  NAND2_X1 U9382 ( .A1(n9588), .A2(n7893), .ZN(n7783) );
  OAI211_X1 U9383 ( .C1(n7894), .C2(n9571), .A(n7784), .B(n7783), .ZN(n7785)
         );
  AOI21_X1 U9384 ( .B1(n7897), .B2(n9573), .A(n7785), .ZN(n7786) );
  OAI21_X1 U9385 ( .B1(n7787), .B2(n9616), .A(n7786), .ZN(P1_U3280) );
  INV_X1 U9386 ( .A(n7788), .ZN(n7790) );
  OAI222_X1 U9387 ( .A1(n9125), .A2(n7789), .B1(n7807), .B2(n7790), .C1(n5984), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U9388 ( .A1(n9755), .A2(n7791), .B1(P1_U3084), .B2(n8287), .C1(
        n9752), .C2(n7790), .ZN(P1_U3333) );
  NOR2_X1 U9389 ( .A1(n7793), .A2(n4599), .ZN(n7794) );
  XNOR2_X1 U9390 ( .A(n7795), .B(n7794), .ZN(n7804) );
  NOR2_X1 U9391 ( .A1(n9235), .A2(n7796), .ZN(n7801) );
  NAND2_X1 U9392 ( .A1(n9284), .A2(n9299), .ZN(n7798) );
  OAI211_X1 U9393 ( .C1(n7799), .C2(n9282), .A(n7798), .B(n7797), .ZN(n7800)
         );
  AOI211_X1 U9394 ( .C1(n7802), .C2(n9271), .A(n7801), .B(n7800), .ZN(n7803)
         );
  OAI21_X1 U9395 ( .B1(n7804), .B2(n9278), .A(n7803), .ZN(P1_U3215) );
  INV_X1 U9396 ( .A(n7805), .ZN(n7901) );
  OAI222_X1 U9397 ( .A1(n9125), .A2(n7808), .B1(n7807), .B2(n7901), .C1(n7806), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XNOR2_X1 U9398 ( .A(n7809), .B(n7872), .ZN(n7811) );
  OAI22_X1 U9399 ( .A1(n7810), .A2(n8932), .B1(n8934), .B2(n8041), .ZN(n7990)
         );
  AOI21_X1 U9400 ( .B1(n7811), .B2(n8917), .A(n7990), .ZN(n9074) );
  INV_X1 U9401 ( .A(n9072), .ZN(n7994) );
  AOI211_X1 U9402 ( .C1(n9072), .C2(n4859), .A(n10022), .B(n7875), .ZN(n9071)
         );
  NOR2_X1 U9403 ( .A1(n8948), .A2(n7994), .ZN(n7815) );
  OAI22_X1 U9404 ( .A1(n9996), .A2(n7813), .B1(n7991), .B2(n9990), .ZN(n7814)
         );
  AOI211_X1 U9405 ( .C1(n9071), .C2(n8969), .A(n7815), .B(n7814), .ZN(n7819)
         );
  AND2_X1 U9406 ( .A1(n9077), .A2(n8652), .ZN(n7871) );
  NOR2_X1 U9407 ( .A1(n7816), .A2(n7871), .ZN(n7817) );
  INV_X1 U9408 ( .A(n7872), .ZN(n7870) );
  XNOR2_X1 U9409 ( .A(n7817), .B(n7870), .ZN(n9075) );
  OR2_X1 U9410 ( .A1(n9075), .A2(n8890), .ZN(n7818) );
  OAI211_X1 U9411 ( .C1(n9074), .C2(n9998), .A(n7819), .B(n7818), .ZN(P2_U3285) );
  INV_X1 U9412 ( .A(n7820), .ZN(n7821) );
  AOI21_X1 U9413 ( .B1(n7823), .B2(n7822), .A(n7821), .ZN(n7829) );
  AOI22_X1 U9414 ( .A1(n8636), .A2(n8652), .B1(n8637), .B2(n8654), .ZN(n7828)
         );
  NOR2_X1 U9415 ( .A1(n8624), .A2(n7824), .ZN(n7825) );
  AOI211_X1 U9416 ( .C1(n9083), .C2(n8638), .A(n7826), .B(n7825), .ZN(n7827)
         );
  OAI211_X1 U9417 ( .C1(n7829), .C2(n8627), .A(n7828), .B(n7827), .ZN(P2_U3233) );
  NAND2_X1 U9418 ( .A1(n7830), .A2(n4333), .ZN(n7831) );
  OAI21_X1 U9419 ( .B1(n4333), .B2(n6011), .A(n7831), .ZN(P2_U3521) );
  NAND2_X1 U9420 ( .A1(n4333), .A2(n7832), .ZN(n7833) );
  OAI21_X1 U9421 ( .B1(n4333), .B2(n6915), .A(n7833), .ZN(P2_U3523) );
  NAND2_X1 U9422 ( .A1(n4333), .A2(n7834), .ZN(n7835) );
  OAI21_X1 U9423 ( .B1(n4333), .B2(n6914), .A(n7835), .ZN(P2_U3522) );
  NAND2_X1 U9424 ( .A1(n7893), .A2(n9299), .ZN(n7836) );
  NAND2_X1 U9425 ( .A1(n7837), .A2(n7836), .ZN(n7839) );
  OR2_X1 U9426 ( .A1(n7893), .A2(n9299), .ZN(n7838) );
  NAND2_X1 U9427 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  OR2_X1 U9428 ( .A1(n8409), .A2(n9597), .ZN(n8434) );
  NAND2_X1 U9429 ( .A1(n8409), .A2(n9597), .ZN(n8435) );
  NAND2_X1 U9430 ( .A1(n7840), .A2(n8205), .ZN(n7841) );
  NAND2_X1 U9431 ( .A1(n8411), .A2(n7841), .ZN(n7922) );
  NAND2_X1 U9432 ( .A1(n7842), .A2(n8094), .ZN(n7843) );
  INV_X1 U9433 ( .A(n8205), .ZN(n7844) );
  XNOR2_X1 U9434 ( .A(n8437), .B(n7844), .ZN(n7845) );
  NAND2_X1 U9435 ( .A1(n7845), .A2(n9603), .ZN(n7847) );
  AOI22_X1 U9436 ( .A1(n9542), .A2(n9297), .B1(n9299), .B2(n9540), .ZN(n7846)
         );
  OAI211_X1 U9437 ( .C1(n9897), .C2(n7922), .A(n7847), .B(n7846), .ZN(n7924)
         );
  NAND2_X1 U9438 ( .A1(n7924), .A2(n10221), .ZN(n7855) );
  INV_X1 U9439 ( .A(n8430), .ZN(n9606) );
  AOI21_X1 U9440 ( .B1(n7848), .B2(n8409), .A(n9949), .ZN(n7849) );
  NAND2_X1 U9441 ( .A1(n9606), .A2(n7849), .ZN(n7920) );
  INV_X1 U9442 ( .A(n7920), .ZN(n7853) );
  INV_X1 U9443 ( .A(n8409), .ZN(n7851) );
  AOI22_X1 U9444 ( .A1(n9616), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7967), .B2(
        n10213), .ZN(n7850) );
  OAI21_X1 U9445 ( .B1(n7851), .B2(n9609), .A(n7850), .ZN(n7852) );
  AOI21_X1 U9446 ( .B1(n7853), .B2(n9554), .A(n7852), .ZN(n7854) );
  OAI211_X1 U9447 ( .C1(n9611), .C2(n7922), .A(n7855), .B(n7854), .ZN(P1_U3279) );
  XNOR2_X1 U9448 ( .A(n7857), .B(n7856), .ZN(n7863) );
  AOI22_X1 U9449 ( .A1(n8622), .A2(n7858), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7862) );
  INV_X1 U9450 ( .A(n8624), .ZN(n8635) );
  INV_X1 U9451 ( .A(n7859), .ZN(n7860) );
  AOI22_X1 U9452 ( .A1(n8638), .A2(n9077), .B1(n8635), .B2(n7860), .ZN(n7861)
         );
  OAI211_X1 U9453 ( .C1(n7863), .C2(n8627), .A(n7862), .B(n7861), .ZN(P2_U3219) );
  NAND2_X1 U9454 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  XNOR2_X1 U9455 ( .A(n7866), .B(n5080), .ZN(n7868) );
  OAI22_X1 U9456 ( .A1(n8483), .A2(n8934), .B1(n8932), .B2(n8030), .ZN(n7867)
         );
  AOI21_X1 U9457 ( .B1(n7868), .B2(n8917), .A(n7867), .ZN(n8003) );
  AOI22_X1 U9458 ( .A1(n7872), .A2(n7871), .B1(n9072), .B2(n8651), .ZN(n7873)
         );
  XNOR2_X1 U9459 ( .A(n7954), .B(n7953), .ZN(n8001) );
  INV_X1 U9460 ( .A(n8033), .ZN(n7998) );
  NAND2_X1 U9461 ( .A1(n7875), .A2(n7998), .ZN(n7948) );
  OR2_X1 U9462 ( .A1(n7875), .A2(n7998), .ZN(n7876) );
  NAND2_X1 U9463 ( .A1(n7948), .A2(n7876), .ZN(n7999) );
  OAI22_X1 U9464 ( .A1(n9996), .A2(n7877), .B1(n8029), .B2(n9990), .ZN(n7878)
         );
  AOI21_X1 U9465 ( .B1(n8963), .B2(n8033), .A(n7878), .ZN(n7879) );
  OAI21_X1 U9466 ( .B1(n8713), .B2(n7999), .A(n7879), .ZN(n7880) );
  AOI21_X1 U9467 ( .B1(n8965), .B2(n8001), .A(n7880), .ZN(n7881) );
  OAI21_X1 U9468 ( .B1(n8003), .B2(n9998), .A(n7881), .ZN(P2_U3284) );
  XNOR2_X1 U9469 ( .A(n7883), .B(n7882), .ZN(n7884) );
  XNOR2_X1 U9470 ( .A(n7885), .B(n7884), .ZN(n7892) );
  NAND2_X1 U9471 ( .A1(n9272), .A2(n9300), .ZN(n7887) );
  OAI211_X1 U9472 ( .C1(n9597), .C2(n9275), .A(n7887), .B(n7886), .ZN(n7888)
         );
  AOI21_X1 U9473 ( .B1(n7889), .B2(n9271), .A(n7888), .ZN(n7891) );
  NAND2_X1 U9474 ( .A1(n9288), .A2(n7893), .ZN(n7890) );
  OAI211_X1 U9475 ( .C1(n7892), .C2(n9278), .A(n7891), .B(n7890), .ZN(P1_U3234) );
  OAI22_X1 U9476 ( .A1(n7894), .A2(n9949), .B1(n4992), .B2(n9947), .ZN(n7896)
         );
  AOI211_X1 U9477 ( .C1(n9952), .C2(n7897), .A(n7896), .B(n7895), .ZN(n7900)
         );
  NAND2_X1 U9478 ( .A1(n9969), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7898) );
  OAI21_X1 U9479 ( .B1(n7900), .B2(n9969), .A(n7898), .ZN(P1_U3534) );
  NAND2_X1 U9480 ( .A1(n9956), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7899) );
  OAI21_X1 U9481 ( .B1(n7900), .B2(n9956), .A(n7899), .ZN(P1_U3487) );
  OAI222_X1 U9482 ( .A1(n9755), .A2(n10151), .B1(P1_U3084), .B2(n5902), .C1(
        n9752), .C2(n7901), .ZN(P1_U3332) );
  XNOR2_X1 U9483 ( .A(n8667), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7907) );
  INV_X1 U9484 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7904) );
  OAI22_X1 U9485 ( .A1(n7905), .A2(n7904), .B1(n7903), .B2(n7902), .ZN(n7906)
         );
  NOR2_X1 U9486 ( .A1(n7906), .A2(n7907), .ZN(n8662) );
  AOI21_X1 U9487 ( .B1(n7907), .B2(n7906), .A(n8662), .ZN(n7919) );
  NOR2_X1 U9488 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8536), .ZN(n7909) );
  NOR2_X1 U9489 ( .A1(n9977), .A2(n8663), .ZN(n7908) );
  AOI211_X1 U9490 ( .C1(n9975), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7909), .B(
        n7908), .ZN(n7918) );
  OAI22_X1 U9491 ( .A1(n7912), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7911), .B2(
        n7910), .ZN(n7915) );
  NAND2_X1 U9492 ( .A1(n8667), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7913) );
  OAI21_X1 U9493 ( .B1(n8667), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7913), .ZN(
        n7914) );
  AOI211_X1 U9494 ( .C1(n7915), .C2(n7914), .A(n8666), .B(n9976), .ZN(n7916)
         );
  INV_X1 U9495 ( .A(n7916), .ZN(n7917) );
  OAI211_X1 U9496 ( .C1(n7919), .C2(n9978), .A(n7918), .B(n7917), .ZN(P2_U3261) );
  INV_X1 U9497 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U9498 ( .A1(n8409), .A2(n9893), .ZN(n7921) );
  OAI211_X1 U9499 ( .C1(n7922), .C2(n9896), .A(n7921), .B(n7920), .ZN(n7923)
         );
  NOR2_X1 U9500 ( .A1(n7924), .A2(n7923), .ZN(n7927) );
  MUX2_X1 U9501 ( .A(n7925), .B(n7927), .S(n9958), .Z(n7926) );
  INV_X1 U9502 ( .A(n7926), .ZN(P1_U3490) );
  INV_X1 U9503 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7928) );
  MUX2_X1 U9504 ( .A(n7928), .B(n7927), .S(n9972), .Z(n7929) );
  INV_X1 U9505 ( .A(n7929), .ZN(P1_U3535) );
  INV_X1 U9506 ( .A(n7930), .ZN(n7972) );
  AOI22_X1 U9507 ( .A1(n7931), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9127), .ZN(n7932) );
  OAI21_X1 U9508 ( .B1(n7972), .B2(n7807), .A(n7932), .ZN(P2_U3334) );
  NAND2_X1 U9509 ( .A1(n7938), .A2(n7933), .ZN(n7935) );
  NOR2_X1 U9510 ( .A1(n7934), .A2(P1_U3084), .ZN(n8324) );
  INV_X1 U9511 ( .A(n8324), .ZN(n8330) );
  OAI211_X1 U9512 ( .C1(n7936), .C2(n9755), .A(n7935), .B(n8330), .ZN(P1_U3330) );
  NAND2_X1 U9513 ( .A1(n7938), .A2(n7937), .ZN(n7940) );
  OAI211_X1 U9514 ( .C1(n10107), .C2(n9125), .A(n7940), .B(n7939), .ZN(
        P2_U3335) );
  INV_X1 U9515 ( .A(n7941), .ZN(n7943) );
  OAI222_X1 U9516 ( .A1(n9125), .A2(n7942), .B1(n7807), .B2(n7943), .C1(
        P2_U3152), .C2(n6550), .ZN(P2_U3336) );
  OAI222_X1 U9517 ( .A1(n9755), .A2(n7944), .B1(n9752), .B2(n7943), .C1(n5903), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  XNOR2_X1 U9518 ( .A(n7946), .B(n7945), .ZN(n7947) );
  AOI222_X1 U9519 ( .A1(n8917), .A2(n7947), .B1(n8650), .B2(n8912), .C1(n8648), 
        .C2(n8914), .ZN(n9069) );
  NAND2_X1 U9520 ( .A1(n7948), .A2(n9066), .ZN(n7949) );
  AND2_X1 U9521 ( .A1(n8018), .A2(n7949), .ZN(n9067) );
  INV_X1 U9522 ( .A(n9066), .ZN(n8047) );
  INV_X1 U9523 ( .A(n7950), .ZN(n8044) );
  AOI22_X1 U9524 ( .A1(n9998), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8044), .B2(
        n8955), .ZN(n7951) );
  OAI21_X1 U9525 ( .B1(n8047), .B2(n8948), .A(n7951), .ZN(n7957) );
  OR2_X1 U9526 ( .A1(n8033), .A2(n8650), .ZN(n7952) );
  NAND2_X1 U9527 ( .A1(n8013), .A2(n7955), .ZN(n9070) );
  NOR2_X1 U9528 ( .A1(n9070), .A2(n8890), .ZN(n7956) );
  AOI211_X1 U9529 ( .C1(n9067), .C2(n8944), .A(n7957), .B(n7956), .ZN(n7958)
         );
  OAI21_X1 U9530 ( .B1(n9069), .B2(n9998), .A(n7958), .ZN(P2_U3283) );
  NAND2_X1 U9531 ( .A1(n7960), .A2(n7959), .ZN(n7962) );
  XOR2_X1 U9532 ( .A(n7962), .B(n7961), .Z(n7970) );
  NAND2_X1 U9533 ( .A1(n9284), .A2(n9297), .ZN(n7964) );
  OAI211_X1 U9534 ( .C1(n7965), .C2(n9282), .A(n7964), .B(n7963), .ZN(n7966)
         );
  AOI21_X1 U9535 ( .B1(n7967), .B2(n9271), .A(n7966), .ZN(n7969) );
  NAND2_X1 U9536 ( .A1(n8409), .A2(n9288), .ZN(n7968) );
  OAI211_X1 U9537 ( .C1(n7970), .C2(n9278), .A(n7969), .B(n7968), .ZN(P1_U3222) );
  OAI222_X1 U9538 ( .A1(P1_U3084), .A2(n5896), .B1(n9752), .B2(n7972), .C1(
        n7971), .C2(n9755), .ZN(P1_U3329) );
  XNOR2_X1 U9539 ( .A(n9316), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7976) );
  OAI21_X1 U9540 ( .B1(n7976), .B2(n7975), .A(n9310), .ZN(n7985) );
  INV_X1 U9541 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10110) );
  INV_X1 U9542 ( .A(n9316), .ZN(n9311) );
  NAND2_X1 U9543 ( .A1(n9853), .A2(n9311), .ZN(n7977) );
  NAND2_X1 U9544 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9145) );
  OAI211_X1 U9545 ( .C1(n9862), .C2(n10110), .A(n7977), .B(n9145), .ZN(n7984)
         );
  INV_X1 U9546 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7982) );
  XNOR2_X1 U9547 ( .A(n9317), .B(n9316), .ZN(n7981) );
  INV_X1 U9548 ( .A(n9315), .ZN(n7980) );
  AOI211_X1 U9549 ( .C1(n7982), .C2(n7981), .A(n9847), .B(n7980), .ZN(n7983)
         );
  AOI211_X1 U9550 ( .C1(n9841), .C2(n7985), .A(n7984), .B(n7983), .ZN(n7986)
         );
  INV_X1 U9551 ( .A(n7986), .ZN(P1_U3255) );
  XOR2_X1 U9552 ( .A(n7988), .B(n7987), .Z(n7996) );
  AOI21_X1 U9553 ( .B1(n8622), .B2(n7990), .A(n7989), .ZN(n7993) );
  OR2_X1 U9554 ( .A1(n8624), .A2(n7991), .ZN(n7992) );
  OAI211_X1 U9555 ( .C1(n7994), .C2(n8617), .A(n7993), .B(n7992), .ZN(n7995)
         );
  AOI21_X1 U9556 ( .B1(n7996), .B2(n8631), .A(n7995), .ZN(n7997) );
  INV_X1 U9557 ( .A(n7997), .ZN(P2_U3238) );
  OAI22_X1 U9558 ( .A1(n7999), .A2(n10022), .B1(n7998), .B2(n10020), .ZN(n8000) );
  AOI21_X1 U9559 ( .B1(n8001), .B2(n10028), .A(n8000), .ZN(n8002) );
  AND2_X1 U9560 ( .A1(n8003), .A2(n8002), .ZN(n8006) );
  MUX2_X1 U9561 ( .A(n8004), .B(n8006), .S(n10030), .Z(n8005) );
  INV_X1 U9562 ( .A(n8005), .ZN(P2_U3487) );
  MUX2_X1 U9563 ( .A(n8007), .B(n8006), .S(n4333), .Z(n8008) );
  INV_X1 U9564 ( .A(n8008), .ZN(P2_U3532) );
  AOI211_X1 U9565 ( .C1(n8340), .C2(n8010), .A(n8930), .B(n8009), .ZN(n8012)
         );
  OAI22_X1 U9566 ( .A1(n8537), .A2(n8934), .B1(n8932), .B2(n8483), .ZN(n8011)
         );
  NOR2_X1 U9567 ( .A1(n8012), .A2(n8011), .ZN(n9064) );
  NAND2_X1 U9568 ( .A1(n9066), .A2(n8649), .ZN(n8338) );
  NAND2_X1 U9569 ( .A1(n8013), .A2(n8338), .ZN(n8014) );
  XNOR2_X1 U9570 ( .A(n8014), .B(n8340), .ZN(n9065) );
  INV_X1 U9571 ( .A(n8015), .ZN(n8488) );
  OAI22_X1 U9572 ( .A1(n9996), .A2(n8016), .B1(n8488), .B2(n9990), .ZN(n8017)
         );
  AOI21_X1 U9573 ( .B1(n8963), .B2(n9061), .A(n8017), .ZN(n8021) );
  AND2_X1 U9574 ( .A1(n8018), .A2(n9061), .ZN(n8019) );
  NOR2_X1 U9575 ( .A1(n8941), .A2(n8019), .ZN(n9062) );
  NAND2_X1 U9576 ( .A1(n9062), .A2(n8944), .ZN(n8020) );
  OAI211_X1 U9577 ( .C1(n9065), .C2(n8890), .A(n8021), .B(n8020), .ZN(n8022)
         );
  INV_X1 U9578 ( .A(n8022), .ZN(n8023) );
  OAI21_X1 U9579 ( .B1(n9064), .B2(n9998), .A(n8023), .ZN(P2_U3282) );
  NAND2_X1 U9580 ( .A1(n8025), .A2(n8024), .ZN(n8027) );
  XOR2_X1 U9581 ( .A(n8027), .B(n8026), .Z(n8035) );
  OAI21_X1 U9582 ( .B1(n8624), .B2(n8029), .A(n8028), .ZN(n8032) );
  OAI22_X1 U9583 ( .A1(n8483), .A2(n8583), .B1(n8584), .B2(n8030), .ZN(n8031)
         );
  AOI211_X1 U9584 ( .C1(n8033), .C2(n8638), .A(n8032), .B(n8031), .ZN(n8034)
         );
  OAI21_X1 U9585 ( .B1(n8035), .B2(n8627), .A(n8034), .ZN(P2_U3226) );
  INV_X1 U9586 ( .A(n8036), .ZN(n8470) );
  OAI222_X1 U9587 ( .A1(n9125), .A2(n8038), .B1(n7807), .B2(n8470), .C1(
        P2_U3152), .C2(n8037), .ZN(P2_U3333) );
  OAI211_X1 U9588 ( .C1(n8040), .C2(n8039), .A(n8482), .B(n8631), .ZN(n8046)
         );
  OAI22_X1 U9589 ( .A1(n8933), .A2(n8583), .B1(n8584), .B2(n8041), .ZN(n8042)
         );
  AOI211_X1 U9590 ( .C1(n8635), .C2(n8044), .A(n8043), .B(n8042), .ZN(n8045)
         );
  OAI211_X1 U9591 ( .C1(n8047), .C2(n8617), .A(n8046), .B(n8045), .ZN(P2_U3236) );
  INV_X1 U9592 ( .A(n8048), .ZN(n8052) );
  AOI22_X1 U9593 ( .A1(n8049), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9127), .ZN(n8050) );
  OAI21_X1 U9594 ( .B1(n8052), .B2(n7807), .A(n8050), .ZN(P2_U3332) );
  OAI222_X1 U9595 ( .A1(P1_U3084), .A2(n8053), .B1(n9752), .B2(n8052), .C1(
        n8051), .C2(n9755), .ZN(P1_U3327) );
  INV_X1 U9596 ( .A(n8054), .ZN(n8058) );
  AOI21_X1 U9597 ( .B1(n9748), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8055), .ZN(
        n8056) );
  OAI21_X1 U9598 ( .B1(n8058), .B2(n9752), .A(n8056), .ZN(P1_U3326) );
  OAI222_X1 U9599 ( .A1(P2_U3152), .A2(n8059), .B1(n7807), .B2(n8058), .C1(
        n8057), .C2(n9125), .ZN(P2_U3331) );
  NAND2_X1 U9600 ( .A1(n9652), .A2(n9192), .ZN(n8459) );
  INV_X1 U9601 ( .A(n8459), .ZN(n8061) );
  INV_X1 U9602 ( .A(n9456), .ZN(n9252) );
  OR2_X1 U9603 ( .A1(n9656), .A2(n9252), .ZN(n8250) );
  INV_X1 U9604 ( .A(n8271), .ZN(n8060) );
  OAI211_X1 U9605 ( .C1(n8061), .C2(n8250), .A(n8461), .B(n8060), .ZN(n8062)
         );
  INV_X1 U9606 ( .A(n9543), .ZN(n9199) );
  OR2_X1 U9607 ( .A1(n9687), .A2(n9199), .ZN(n9505) );
  NAND2_X1 U9608 ( .A1(n8187), .A2(n9505), .ZN(n8446) );
  NAND2_X1 U9609 ( .A1(n9681), .A2(n8063), .ZN(n8447) );
  NAND2_X1 U9610 ( .A1(n9687), .A2(n9199), .ZN(n9504) );
  NAND2_X1 U9611 ( .A1(n8447), .A2(n9504), .ZN(n8064) );
  MUX2_X1 U9612 ( .A(n8446), .B(n8064), .S(n8167), .Z(n8065) );
  INV_X1 U9613 ( .A(n8065), .ZN(n8113) );
  NAND2_X1 U9614 ( .A1(n8205), .A2(n8252), .ZN(n8081) );
  NAND2_X1 U9615 ( .A1(n8291), .A2(n8163), .ZN(n8069) );
  AOI21_X1 U9616 ( .B1(n8066), .B2(n8163), .A(n10209), .ZN(n8073) );
  AOI21_X1 U9617 ( .B1(n9305), .B2(n8167), .A(n8067), .ZN(n8072) );
  OR2_X1 U9618 ( .A1(n8076), .A2(n9918), .ZN(n8071) );
  OR2_X1 U9619 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  OAI211_X1 U9620 ( .C1(n8073), .C2(n8072), .A(n8071), .B(n8070), .ZN(n8074)
         );
  INV_X1 U9621 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U9622 ( .A1(n8078), .A2(n8077), .ZN(n8082) );
  NAND3_X1 U9623 ( .A1(n8082), .A2(n8083), .A3(n8194), .ZN(n8079) );
  NAND3_X1 U9624 ( .A1(n8079), .A2(n8085), .A3(n8275), .ZN(n8080) );
  NAND3_X1 U9625 ( .A1(n8082), .A2(n8275), .A3(n8292), .ZN(n8087) );
  AND2_X1 U9626 ( .A1(n8084), .A2(n8083), .ZN(n8230) );
  NAND2_X1 U9627 ( .A1(n8086), .A2(n8085), .ZN(n8254) );
  AOI21_X1 U9628 ( .B1(n8087), .B2(n8230), .A(n8254), .ZN(n8090) );
  NAND2_X1 U9629 ( .A1(n8089), .A2(n8088), .ZN(n8227) );
  OR3_X1 U9630 ( .A1(n8090), .A2(n8163), .A3(n8227), .ZN(n8091) );
  NAND2_X1 U9631 ( .A1(n8091), .A2(n8204), .ZN(n8099) );
  OR2_X1 U9632 ( .A1(n9705), .A2(n9598), .ZN(n8441) );
  OR2_X1 U9633 ( .A1(n9709), .A2(n9579), .ZN(n8188) );
  NAND2_X1 U9634 ( .A1(n8434), .A2(n8092), .ZN(n8093) );
  NAND2_X1 U9635 ( .A1(n8093), .A2(n8435), .ZN(n8255) );
  AND3_X1 U9636 ( .A1(n8441), .A2(n8188), .A3(n8255), .ZN(n8097) );
  NAND2_X1 U9637 ( .A1(n9705), .A2(n9598), .ZN(n8102) );
  NAND2_X1 U9638 ( .A1(n9709), .A2(n9579), .ZN(n8438) );
  NAND2_X1 U9639 ( .A1(n8102), .A2(n8438), .ZN(n8226) );
  NAND2_X1 U9640 ( .A1(n8435), .A2(n8094), .ZN(n8229) );
  AND2_X1 U9641 ( .A1(n8229), .A2(n8434), .ZN(n8095) );
  NOR2_X1 U9642 ( .A1(n8226), .A2(n8095), .ZN(n8096) );
  MUX2_X1 U9643 ( .A(n8097), .B(n8096), .S(n8167), .Z(n8098) );
  OAI21_X1 U9644 ( .B1(n8100), .B2(n8099), .A(n8098), .ZN(n8107) );
  AND2_X1 U9645 ( .A1(n9698), .A2(n9541), .ZN(n8442) );
  NAND2_X1 U9646 ( .A1(n9569), .A2(n9580), .ZN(n9536) );
  INV_X1 U9647 ( .A(n9536), .ZN(n8263) );
  INV_X1 U9648 ( .A(n9562), .ZN(n8106) );
  INV_X1 U9649 ( .A(n8188), .ZN(n8101) );
  NAND2_X1 U9650 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  AND2_X1 U9651 ( .A1(n8103), .A2(n8441), .ZN(n8258) );
  NAND2_X1 U9652 ( .A1(n8226), .A2(n8441), .ZN(n8104) );
  MUX2_X1 U9653 ( .A(n8258), .B(n8104), .S(n8163), .Z(n8105) );
  NAND3_X1 U9654 ( .A1(n8107), .A2(n8106), .A3(n8105), .ZN(n8109) );
  OR2_X1 U9655 ( .A1(n9693), .A2(n9558), .ZN(n8443) );
  NAND2_X1 U9656 ( .A1(n9693), .A2(n9558), .ZN(n9503) );
  NAND2_X1 U9657 ( .A1(n8443), .A2(n9503), .ZN(n9550) );
  INV_X1 U9658 ( .A(n9550), .ZN(n9501) );
  INV_X1 U9659 ( .A(n8442), .ZN(n8262) );
  MUX2_X1 U9660 ( .A(n8262), .B(n9536), .S(n8167), .Z(n8108) );
  NAND3_X1 U9661 ( .A1(n8109), .A2(n9501), .A3(n8108), .ZN(n8111) );
  MUX2_X1 U9662 ( .A(n8443), .B(n9503), .S(n8163), .Z(n8110) );
  NAND3_X1 U9663 ( .A1(n8111), .A2(n9525), .A3(n8110), .ZN(n8112) );
  INV_X1 U9664 ( .A(n9508), .ZN(n9261) );
  OR2_X1 U9665 ( .A1(n9676), .A2(n9261), .ZN(n8186) );
  NAND2_X1 U9666 ( .A1(n9672), .A2(n9169), .ZN(n8453) );
  NAND2_X1 U9667 ( .A1(n9676), .A2(n9261), .ZN(n8452) );
  OR2_X1 U9668 ( .A1(n9672), .A2(n9169), .ZN(n8185) );
  AND2_X1 U9669 ( .A1(n8185), .A2(n8186), .ZN(n8268) );
  OR2_X1 U9670 ( .A1(n9667), .A2(n8116), .ZN(n8269) );
  INV_X1 U9671 ( .A(n8269), .ZN(n8115) );
  NOR2_X1 U9672 ( .A1(n8121), .A2(n8115), .ZN(n8119) );
  AND2_X1 U9673 ( .A1(n9661), .A2(n9179), .ZN(n8456) );
  NAND2_X1 U9674 ( .A1(n8269), .A2(n4800), .ZN(n8117) );
  NAND2_X1 U9675 ( .A1(n9667), .A2(n8116), .ZN(n8454) );
  NAND2_X1 U9676 ( .A1(n8117), .A2(n8454), .ZN(n8118) );
  OR2_X1 U9677 ( .A1(n8456), .A2(n8118), .ZN(n8225) );
  OR2_X1 U9678 ( .A1(n9661), .A2(n9179), .ZN(n9440) );
  OAI211_X1 U9679 ( .C1(n8119), .C2(n8225), .A(n8163), .B(n9440), .ZN(n8128)
         );
  NAND2_X1 U9680 ( .A1(n9656), .A2(n9252), .ZN(n8458) );
  NAND2_X1 U9681 ( .A1(n8250), .A2(n8458), .ZN(n9442) );
  NOR2_X1 U9682 ( .A1(n9440), .A2(n8163), .ZN(n8120) );
  NOR2_X1 U9683 ( .A1(n9442), .A2(n8120), .ZN(n8127) );
  XNOR2_X1 U9684 ( .A(n9652), .B(n9444), .ZN(n9427) );
  NAND2_X1 U9685 ( .A1(n8269), .A2(n8185), .ZN(n8124) );
  NAND2_X1 U9686 ( .A1(n8454), .A2(n8167), .ZN(n8122) );
  NOR2_X1 U9687 ( .A1(n8456), .A2(n8122), .ZN(n8123) );
  OAI21_X1 U9688 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8126) );
  NAND2_X1 U9689 ( .A1(n9646), .A2(n8425), .ZN(n8184) );
  OAI211_X1 U9690 ( .C1(n8271), .C2(n8458), .A(n8184), .B(n8459), .ZN(n8276)
         );
  NAND2_X1 U9691 ( .A1(n9634), .A2(n9294), .ZN(n8219) );
  INV_X1 U9692 ( .A(n9415), .ZN(n9375) );
  INV_X1 U9693 ( .A(n8184), .ZN(n8460) );
  OAI21_X1 U9694 ( .B1(n9375), .B2(n8460), .A(n8463), .ZN(n8133) );
  NAND2_X1 U9695 ( .A1(n9642), .A2(n8461), .ZN(n8131) );
  NAND2_X1 U9696 ( .A1(n8219), .A2(n8131), .ZN(n8132) );
  MUX2_X1 U9697 ( .A(n8133), .B(n8132), .S(n8167), .Z(n8134) );
  OAI21_X1 U9698 ( .B1(n8135), .B2(n9371), .A(n8134), .ZN(n8139) );
  INV_X1 U9699 ( .A(n9642), .ZN(n9395) );
  MUX2_X1 U9700 ( .A(n9375), .B(n9395), .S(n8167), .Z(n8136) );
  AOI21_X1 U9701 ( .B1(n9375), .B2(n8460), .A(n9642), .ZN(n8137) );
  MUX2_X1 U9702 ( .A(n9375), .B(n8137), .S(n8163), .Z(n8138) );
  NAND2_X1 U9703 ( .A1(n9628), .A2(n9376), .ZN(n8222) );
  NAND2_X2 U9704 ( .A1(n8464), .A2(n8222), .ZN(n9363) );
  MUX2_X1 U9705 ( .A(n8463), .B(n8219), .S(n8163), .Z(n8140) );
  MUX2_X1 U9706 ( .A(n8464), .B(n8222), .S(n8167), .Z(n8142) );
  NAND2_X1 U9707 ( .A1(n9124), .A2(n4240), .ZN(n8144) );
  OR2_X1 U9708 ( .A1(n8152), .A2(n9754), .ZN(n8143) );
  INV_X1 U9709 ( .A(n9625), .ZN(n8433) );
  NAND2_X1 U9710 ( .A1(n9119), .A2(n5327), .ZN(n8147) );
  OR2_X1 U9711 ( .A1(n8152), .A2(n6750), .ZN(n8146) );
  NAND2_X1 U9712 ( .A1(n8147), .A2(n8146), .ZN(n8175) );
  NAND2_X1 U9713 ( .A1(n4615), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U9714 ( .A1(n5443), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U9715 ( .A1(n8148), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U9716 ( .A1(n8175), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U9717 ( .A1(n8404), .A2(n5327), .ZN(n8154) );
  INV_X1 U9718 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8406) );
  OR2_X1 U9719 ( .A1(n8152), .A2(n8406), .ZN(n8153) );
  INV_X1 U9720 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U9721 ( .A1(n4615), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U9722 ( .A1(n5443), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8156) );
  OAI211_X1 U9723 ( .C1(n4626), .C2(n10165), .A(n8157), .B(n8156), .ZN(n9291)
         );
  INV_X1 U9724 ( .A(n9291), .ZN(n8182) );
  OR2_X1 U9725 ( .A1(n9354), .A2(n8182), .ZN(n8158) );
  NAND2_X1 U9726 ( .A1(n8161), .A2(n8158), .ZN(n8284) );
  AND2_X1 U9727 ( .A1(n8284), .A2(n8175), .ZN(n8172) );
  INV_X1 U9728 ( .A(n8172), .ZN(n8312) );
  NAND2_X1 U9729 ( .A1(n9350), .A2(n9291), .ZN(n8160) );
  AND2_X1 U9730 ( .A1(n9354), .A2(n8160), .ZN(n8306) );
  NAND3_X1 U9731 ( .A1(n8161), .A2(n8306), .A3(n8163), .ZN(n8162) );
  OAI21_X1 U9732 ( .B1(n8312), .B2(n8163), .A(n8162), .ZN(n8173) );
  NOR2_X1 U9733 ( .A1(n9292), .A2(n8163), .ZN(n8171) );
  AND2_X1 U9734 ( .A1(n9292), .A2(n8163), .ZN(n8166) );
  INV_X1 U9735 ( .A(n8166), .ZN(n8165) );
  NOR2_X1 U9736 ( .A1(n9625), .A2(n8171), .ZN(n8164) );
  AOI21_X1 U9737 ( .B1(n9625), .B2(n8165), .A(n8164), .ZN(n8170) );
  NAND2_X1 U9738 ( .A1(n8464), .A2(n8166), .ZN(n8169) );
  NAND3_X1 U9739 ( .A1(n8433), .A2(n8167), .A3(n8222), .ZN(n8168) );
  AND2_X1 U9740 ( .A1(n9619), .A2(n9350), .ZN(n8181) );
  NOR4_X1 U9741 ( .A1(n8180), .A2(n8331), .A3(n8181), .A4(n8176), .ZN(n8322)
         );
  INV_X1 U9742 ( .A(n8181), .ZN(n8179) );
  OR2_X1 U9743 ( .A1(n9468), .A2(n8287), .ZN(n8318) );
  INV_X1 U9744 ( .A(n8318), .ZN(n8178) );
  AND4_X1 U9745 ( .A1(n8180), .A2(n8179), .A3(n5920), .A4(n8178), .ZN(n8321)
         );
  NAND2_X1 U9746 ( .A1(n9354), .A2(n8182), .ZN(n8183) );
  NAND2_X1 U9747 ( .A1(n8179), .A2(n8183), .ZN(n8283) );
  INV_X1 U9748 ( .A(n8283), .ZN(n8216) );
  INV_X1 U9749 ( .A(n8284), .ZN(n8215) );
  OR2_X1 U9750 ( .A1(n9625), .A2(n9292), .ZN(n8223) );
  NAND2_X1 U9751 ( .A1(n9625), .A2(n9292), .ZN(n8308) );
  NAND2_X1 U9752 ( .A1(n8223), .A2(n8308), .ZN(n8466) );
  NAND2_X1 U9753 ( .A1(n8461), .A2(n8184), .ZN(n9414) );
  INV_X1 U9754 ( .A(n9442), .ZN(n8211) );
  NAND2_X1 U9755 ( .A1(n4980), .A2(n9440), .ZN(n9455) );
  NAND2_X1 U9756 ( .A1(n8269), .A2(n8454), .ZN(n9461) );
  INV_X1 U9757 ( .A(n9461), .ZN(n9464) );
  XNOR2_X1 U9758 ( .A(n9705), .B(n9598), .ZN(n9577) );
  NAND4_X1 U9759 ( .A1(n8192), .A2(n8191), .A3(n8190), .A4(n8189), .ZN(n8197)
         );
  NAND2_X1 U9760 ( .A1(n8194), .A2(n8193), .ZN(n8294) );
  NOR4_X1 U9761 ( .A1(n8197), .A2(n8196), .A3(n8294), .A4(n8195), .ZN(n8199)
         );
  NAND4_X1 U9762 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n4382), .ZN(n8202)
         );
  NOR2_X1 U9763 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  NAND4_X1 U9764 ( .A1(n9599), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(n8206)
         );
  NOR3_X1 U9765 ( .A1(n9562), .A2(n9577), .A3(n8206), .ZN(n8207) );
  AND4_X1 U9766 ( .A1(n9517), .A2(n9501), .A3(n9525), .A4(n8207), .ZN(n8208)
         );
  NAND4_X1 U9767 ( .A1(n9464), .A2(n9480), .A3(n9494), .A4(n8208), .ZN(n8209)
         );
  NOR2_X1 U9768 ( .A1(n9455), .A2(n8209), .ZN(n8210) );
  AND4_X1 U9769 ( .A1(n5040), .A2(n8211), .A3(n8210), .A4(n9427), .ZN(n8212)
         );
  XNOR2_X1 U9770 ( .A(n9642), .B(n9415), .ZN(n9397) );
  NAND3_X1 U9771 ( .A1(n4680), .A2(n8212), .A3(n9397), .ZN(n8213) );
  NOR2_X1 U9772 ( .A1(n8213), .A2(n9363), .ZN(n8214) );
  NAND4_X1 U9773 ( .A1(n8216), .A2(n8215), .A3(n4986), .A4(n8214), .ZN(n8217)
         );
  NAND2_X1 U9774 ( .A1(n8217), .A2(n5902), .ZN(n8319) );
  NAND2_X1 U9775 ( .A1(n9642), .A2(n9375), .ZN(n8218) );
  NAND2_X1 U9776 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  NAND2_X1 U9777 ( .A1(n8220), .A2(n8463), .ZN(n8221) );
  NAND2_X1 U9778 ( .A1(n8222), .A2(n8221), .ZN(n8304) );
  NOR2_X1 U9779 ( .A1(n9642), .A2(n9375), .ZN(n8462) );
  NOR2_X1 U9780 ( .A1(n8462), .A2(n4810), .ZN(n8224) );
  OAI211_X1 U9781 ( .C1(n8304), .C2(n8224), .A(n8223), .B(n8464), .ZN(n8310)
         );
  INV_X1 U9782 ( .A(n8304), .ZN(n8280) );
  INV_X1 U9783 ( .A(n8225), .ZN(n8273) );
  NAND2_X1 U9784 ( .A1(n9504), .A2(n9503), .ZN(n8449) );
  INV_X1 U9785 ( .A(n8226), .ZN(n8261) );
  AND2_X1 U9786 ( .A1(n8227), .A2(n8252), .ZN(n8228) );
  NOR2_X1 U9787 ( .A1(n8229), .A2(n8228), .ZN(n8251) );
  NAND4_X1 U9788 ( .A1(n9536), .A2(n8261), .A3(n8230), .A4(n8251), .ZN(n8231)
         );
  OR2_X1 U9789 ( .A1(n8449), .A2(n8231), .ZN(n8232) );
  NOR2_X1 U9790 ( .A1(n4249), .A2(n8232), .ZN(n8233) );
  NAND2_X1 U9791 ( .A1(n8273), .A2(n8233), .ZN(n8290) );
  INV_X1 U9792 ( .A(n8247), .ZN(n8235) );
  OR3_X1 U9793 ( .A1(n8290), .A2(n4815), .A3(n8235), .ZN(n8299) );
  NAND2_X1 U9794 ( .A1(n6757), .A2(n8236), .ZN(n8237) );
  NAND3_X1 U9795 ( .A1(n8238), .A2(n8237), .A3(n8313), .ZN(n8239) );
  NAND2_X1 U9796 ( .A1(n8240), .A2(n8239), .ZN(n8242) );
  OAI21_X1 U9797 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8244) );
  INV_X1 U9798 ( .A(n8244), .ZN(n8249) );
  NAND2_X1 U9799 ( .A1(n9918), .A2(n8245), .ZN(n8288) );
  AOI21_X1 U9800 ( .B1(n8247), .B2(n8288), .A(n8246), .ZN(n8248) );
  OAI22_X1 U9801 ( .A1(n8299), .A2(n8249), .B1(n8248), .B2(n8290), .ZN(n8277)
         );
  AND2_X1 U9802 ( .A1(n8250), .A2(n9440), .ZN(n8457) );
  INV_X1 U9803 ( .A(n8251), .ZN(n8257) );
  INV_X1 U9804 ( .A(n8252), .ZN(n8253) );
  NOR2_X1 U9805 ( .A1(n8254), .A2(n8253), .ZN(n8256) );
  OAI21_X1 U9806 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(n8260) );
  INV_X1 U9807 ( .A(n8258), .ZN(n8259) );
  AOI21_X1 U9808 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8264) );
  OAI211_X1 U9809 ( .C1(n8264), .C2(n8263), .A(n8443), .B(n8262), .ZN(n8265)
         );
  INV_X1 U9810 ( .A(n8265), .ZN(n8266) );
  NOR2_X1 U9811 ( .A1(n8449), .A2(n8266), .ZN(n8267) );
  NOR2_X1 U9812 ( .A1(n8446), .A2(n8267), .ZN(n8270) );
  OAI211_X1 U9813 ( .C1(n8270), .C2(n4249), .A(n8269), .B(n8268), .ZN(n8272)
         );
  AOI21_X1 U9814 ( .B1(n8273), .B2(n8272), .A(n8271), .ZN(n8274) );
  OAI211_X1 U9815 ( .C1(n8290), .C2(n8275), .A(n8457), .B(n8274), .ZN(n8301)
         );
  INV_X1 U9816 ( .A(n8276), .ZN(n8300) );
  OAI21_X1 U9817 ( .B1(n8277), .B2(n8301), .A(n8300), .ZN(n8278) );
  NAND2_X1 U9818 ( .A1(n4680), .A2(n8278), .ZN(n8279) );
  AND2_X1 U9819 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  OAI21_X1 U9820 ( .B1(n8310), .B2(n8281), .A(n8308), .ZN(n8282) );
  OR2_X1 U9821 ( .A1(n8283), .A2(n8282), .ZN(n8286) );
  NAND2_X1 U9822 ( .A1(n8284), .A2(n8179), .ZN(n8285) );
  NAND2_X1 U9823 ( .A1(n8286), .A2(n8285), .ZN(n8323) );
  OAI21_X1 U9824 ( .B1(n8323), .B2(n9468), .A(n8287), .ZN(n8317) );
  INV_X1 U9825 ( .A(n8288), .ZN(n8289) );
  AND2_X1 U9826 ( .A1(n7395), .A2(n8289), .ZN(n8298) );
  INV_X1 U9827 ( .A(n8290), .ZN(n8296) );
  AND2_X1 U9828 ( .A1(n8291), .A2(n9918), .ZN(n8293) );
  OAI21_X1 U9829 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n8295) );
  NAND2_X1 U9830 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  OAI21_X1 U9831 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8302) );
  OAI21_X1 U9832 ( .B1(n8302), .B2(n8301), .A(n8300), .ZN(n8303) );
  AND2_X1 U9833 ( .A1(n8303), .A2(n8463), .ZN(n8305) );
  NOR2_X1 U9834 ( .A1(n8305), .A2(n8304), .ZN(n8309) );
  INV_X1 U9835 ( .A(n8306), .ZN(n8307) );
  OAI211_X1 U9836 ( .C1(n8310), .C2(n8309), .A(n8308), .B(n8307), .ZN(n8311)
         );
  NAND2_X1 U9837 ( .A1(n8312), .A2(n8311), .ZN(n8314) );
  NAND3_X1 U9838 ( .A1(n8314), .A2(n8313), .A3(n8179), .ZN(n8315) );
  NAND3_X1 U9839 ( .A1(n8319), .A2(n8315), .A3(n9468), .ZN(n8316) );
  OAI211_X1 U9840 ( .C1(n8319), .C2(n8318), .A(n8317), .B(n8316), .ZN(n8320)
         );
  NOR3_X1 U9841 ( .A1(n8322), .A2(n8321), .A3(n8320), .ZN(n8334) );
  INV_X1 U9842 ( .A(n8323), .ZN(n8326) );
  OAI21_X1 U9843 ( .B1(n8326), .B2(n8325), .A(n8324), .ZN(n8333) );
  INV_X1 U9844 ( .A(n4239), .ZN(n8467) );
  NAND4_X1 U9845 ( .A1(n8328), .A2(n9540), .A3(n8467), .A4(n8327), .ZN(n8329)
         );
  OAI211_X1 U9846 ( .C1(n8331), .C2(n8330), .A(n8329), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8332) );
  OAI21_X1 U9847 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(P1_U3240) );
  INV_X1 U9848 ( .A(n8335), .ZN(n9130) );
  OAI222_X1 U9849 ( .A1(n9755), .A2(n8337), .B1(P1_U3084), .B2(n8336), .C1(
        n9752), .C2(n9130), .ZN(P1_U3325) );
  INV_X1 U9850 ( .A(n9012), .ZN(n8801) );
  NAND3_X1 U9851 ( .A1(n8340), .A2(n8339), .A3(n8338), .ZN(n8341) );
  OAI21_X1 U9852 ( .B1(n8648), .B2(n9061), .A(n8341), .ZN(n8342) );
  INV_X1 U9853 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U9854 ( .A1(n8344), .A2(n8343), .ZN(n8940) );
  NAND2_X1 U9855 ( .A1(n9039), .A2(n8646), .ZN(n8347) );
  INV_X1 U9856 ( .A(n9034), .ZN(n8354) );
  NAND2_X1 U9857 ( .A1(n8354), .A2(n8613), .ZN(n8348) );
  INV_X1 U9858 ( .A(n9024), .ZN(n8518) );
  NOR2_X1 U9859 ( .A1(n8518), .A2(n8809), .ZN(n8349) );
  INV_X1 U9860 ( .A(n8796), .ZN(n8803) );
  INV_X1 U9861 ( .A(n8752), .ZN(n8350) );
  OAI22_X1 U9862 ( .A1(n8715), .A2(n8717), .B1(n4855), .B2(n8740), .ZN(n8353)
         );
  INV_X1 U9863 ( .A(n9056), .ZN(n8949) );
  INV_X1 U9864 ( .A(n9050), .ZN(n8921) );
  NAND2_X1 U9865 ( .A1(n8855), .A2(n8854), .ZN(n8857) );
  NOR2_X2 U9866 ( .A1(n8857), .A2(n9024), .ZN(n8813) );
  AOI21_X1 U9868 ( .B1(n8982), .B2(n8723), .A(n4271), .ZN(n8983) );
  INV_X1 U9869 ( .A(n8982), .ZN(n8358) );
  AOI22_X1 U9870 ( .A1(n9998), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8356), .B2(
        n8955), .ZN(n8357) );
  OAI21_X1 U9871 ( .B1(n8358), .B2(n8948), .A(n8357), .ZN(n8359) );
  AOI21_X1 U9872 ( .B1(n8983), .B2(n8944), .A(n8359), .ZN(n8367) );
  AOI21_X1 U9873 ( .B1(n8362), .B2(P2_B_REG_SCAN_IN), .A(n8934), .ZN(n8704) );
  INV_X1 U9874 ( .A(n8363), .ZN(n8643) );
  OR2_X1 U9875 ( .A1(n8985), .A2(n9998), .ZN(n8366) );
  OAI211_X1 U9876 ( .C1(n8986), .C2(n8890), .A(n8367), .B(n8366), .ZN(P2_U3267) );
  INV_X1 U9877 ( .A(n8368), .ZN(n8369) );
  NAND2_X1 U9878 ( .A1(n8369), .A2(n8371), .ZN(n8372) );
  MUX2_X1 U9879 ( .A(n8372), .B(n8371), .S(n8370), .Z(n8382) );
  NAND3_X1 U9880 ( .A1(n8370), .A2(n8658), .A3(n8373), .ZN(n8375) );
  OAI22_X1 U9881 ( .A1(n8375), .A2(n8608), .B1(n8584), .B2(n8374), .ZN(n8380)
         );
  OAI22_X1 U9882 ( .A1(n10015), .A2(n8617), .B1(n8583), .B2(n8376), .ZN(n8379)
         );
  OAI22_X1 U9883 ( .A1(n8624), .A2(n8377), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10175), .ZN(n8378) );
  NOR3_X1 U9884 ( .A1(n8380), .A2(n8379), .A3(n8378), .ZN(n8381) );
  OAI21_X1 U9885 ( .B1(n8382), .B2(n8627), .A(n8381), .ZN(P2_U3232) );
  NAND2_X1 U9886 ( .A1(n8384), .A2(n8383), .ZN(n8385) );
  AND2_X1 U9887 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  AOI22_X1 U9888 ( .A1(n8622), .A2(n8388), .B1(n8631), .B2(n8387), .ZN(n8390)
         );
  MUX2_X1 U9889 ( .A(n8624), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8389) );
  OAI211_X1 U9890 ( .C1(n8391), .C2(n8617), .A(n8390), .B(n8389), .ZN(P2_U3220) );
  OAI222_X1 U9891 ( .A1(n9755), .A2(n8393), .B1(n9752), .B2(n8392), .C1(n9468), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  NAND3_X1 U9892 ( .A1(n8394), .A2(n8629), .A3(n8646), .ZN(n8395) );
  OAI21_X1 U9893 ( .B1(n4707), .B2(n8627), .A(n8395), .ZN(n8398) );
  INV_X1 U9894 ( .A(n8396), .ZN(n8397) );
  NAND2_X1 U9895 ( .A1(n8398), .A2(n8397), .ZN(n8403) );
  NOR2_X1 U9896 ( .A1(n8624), .A2(n8872), .ZN(n8401) );
  AND2_X1 U9897 ( .A1(n8646), .A2(n8912), .ZN(n8399) );
  AOI21_X1 U9898 ( .B1(n8830), .B2(n8914), .A(n8399), .ZN(n8866) );
  OAI22_X1 U9899 ( .A1(n8549), .A2(n8866), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10181), .ZN(n8400) );
  AOI211_X1 U9900 ( .C1(n9034), .C2(n8638), .A(n8401), .B(n8400), .ZN(n8402)
         );
  OAI211_X1 U9901 ( .C1(n8627), .C2(n8505), .A(n8403), .B(n8402), .ZN(P2_U3221) );
  INV_X1 U9902 ( .A(n8404), .ZN(n8408) );
  OAI222_X1 U9903 ( .A1(n9755), .A2(n8406), .B1(n9752), .B2(n8408), .C1(n8405), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  INV_X1 U9904 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10097) );
  OAI222_X1 U9905 ( .A1(n9125), .A2(n10097), .B1(n7807), .B2(n8408), .C1(n8407), .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9906 ( .A(n9597), .ZN(n9298) );
  NAND2_X1 U9907 ( .A1(n8409), .A2(n9298), .ZN(n8410) );
  NAND2_X1 U9908 ( .A1(n9709), .A2(n9297), .ZN(n8412) );
  AND2_X1 U9909 ( .A1(n9705), .A2(n9296), .ZN(n8414) );
  NOR2_X1 U9910 ( .A1(n9569), .A2(n9541), .ZN(n8415) );
  NAND2_X1 U9911 ( .A1(n9569), .A2(n9541), .ZN(n8416) );
  NAND2_X1 U9912 ( .A1(n9681), .A2(n9523), .ZN(n8417) );
  AND2_X1 U9913 ( .A1(n9676), .A2(n9508), .ZN(n8418) );
  INV_X1 U9914 ( .A(n9672), .ZN(n9478) );
  NAND2_X1 U9915 ( .A1(n9667), .A2(n9481), .ZN(n8419) );
  NAND2_X1 U9916 ( .A1(n8420), .A2(n8419), .ZN(n9449) );
  NAND2_X1 U9917 ( .A1(n9454), .A2(n9179), .ZN(n8421) );
  NAND2_X1 U9918 ( .A1(n9661), .A2(n9465), .ZN(n8422) );
  OR2_X1 U9919 ( .A1(n9656), .A2(n9456), .ZN(n8423) );
  OR2_X1 U9920 ( .A1(n9646), .A2(n9428), .ZN(n8426) );
  OR2_X1 U9921 ( .A1(n9642), .A2(n9415), .ZN(n8428) );
  AND2_X1 U9922 ( .A1(n9642), .A2(n9415), .ZN(n8427) );
  NAND2_X1 U9923 ( .A1(n9360), .A2(n9363), .ZN(n9359) );
  NAND2_X1 U9924 ( .A1(n9359), .A2(n5120), .ZN(n8429) );
  INV_X1 U9925 ( .A(n9656), .ZN(n9439) );
  INV_X1 U9926 ( .A(n9681), .ZN(n9512) );
  AND2_X2 U9927 ( .A1(n9529), .A2(n9512), .ZN(n9510) );
  INV_X1 U9928 ( .A(n9676), .ZN(n9493) );
  NAND2_X1 U9929 ( .A1(n9510), .A2(n9493), .ZN(n9488) );
  NOR2_X1 U9930 ( .A1(n9616), .A2(n10220), .ZN(n9485) );
  AOI22_X1 U9931 ( .A1(n8431), .A2(n10213), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9616), .ZN(n8432) );
  OAI21_X1 U9932 ( .B1(n8433), .B2(n9609), .A(n8432), .ZN(n8469) );
  INV_X1 U9933 ( .A(n8434), .ZN(n8436) );
  INV_X1 U9934 ( .A(n9577), .ZN(n8439) );
  INV_X1 U9935 ( .A(n8443), .ZN(n8444) );
  NOR2_X1 U9936 ( .A1(n8446), .A2(n8444), .ZN(n8445) );
  INV_X1 U9937 ( .A(n8446), .ZN(n8450) );
  INV_X1 U9938 ( .A(n8447), .ZN(n8448) );
  AOI21_X1 U9939 ( .B1(n8450), .B2(n8449), .A(n8448), .ZN(n8451) );
  INV_X1 U9940 ( .A(n9376), .ZN(n9293) );
  AOI21_X1 U9941 ( .B1(n8467), .B2(P1_B_REG_SCAN_IN), .A(n9927), .ZN(n9351) );
  OAI222_X1 U9942 ( .A1(n9755), .A2(n8471), .B1(n9752), .B2(n8470), .C1(
        P1_U3084), .C2(n5879), .ZN(P1_U3328) );
  XNOR2_X1 U9943 ( .A(n8473), .B(n8472), .ZN(n8481) );
  INV_X1 U9944 ( .A(n8743), .ZN(n8475) );
  OAI22_X1 U9945 ( .A1(n8624), .A2(n8475), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8474), .ZN(n8479) );
  INV_X1 U9946 ( .A(n8740), .ZN(n8477) );
  OAI22_X1 U9947 ( .A1(n8477), .A2(n8583), .B1(n8584), .B2(n8476), .ZN(n8478)
         );
  AOI211_X1 U9948 ( .C1(n8992), .C2(n8638), .A(n8479), .B(n8478), .ZN(n8480)
         );
  OAI21_X1 U9949 ( .B1(n8481), .B2(n8627), .A(n8480), .ZN(P2_U3216) );
  NOR3_X1 U9950 ( .A1(n8608), .A2(n8484), .A3(n8483), .ZN(n8485) );
  AOI21_X1 U9951 ( .B1(n4886), .B2(n8631), .A(n8485), .ZN(n8494) );
  AOI22_X1 U9952 ( .A1(n8637), .A2(n8649), .B1(n8636), .B2(n8913), .ZN(n8487)
         );
  OAI211_X1 U9953 ( .C1(n8624), .C2(n8488), .A(n8487), .B(n8486), .ZN(n8491)
         );
  NOR2_X1 U9954 ( .A1(n8489), .A2(n8627), .ZN(n8490) );
  AOI211_X1 U9955 ( .C1(n9061), .C2(n8638), .A(n8491), .B(n8490), .ZN(n8492)
         );
  OAI21_X1 U9956 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(P2_U3217) );
  NOR2_X1 U9957 ( .A1(n8496), .A2(n8495), .ZN(n8554) );
  AOI22_X1 U9958 ( .A1(n8497), .A2(n8631), .B1(n8629), .B2(n8645), .ZN(n8503)
         );
  INV_X1 U9959 ( .A(n8799), .ZN(n8499) );
  OAI22_X1 U9960 ( .A1(n8624), .A2(n8499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8498), .ZN(n8501) );
  OAI22_X1 U9961 ( .A1(n8512), .A2(n8584), .B1(n8583), .B2(n8557), .ZN(n8500)
         );
  AOI211_X1 U9962 ( .C1(n9012), .C2(n8638), .A(n8501), .B(n8500), .ZN(n8502)
         );
  OAI21_X1 U9963 ( .B1(n8554), .B2(n8503), .A(n8502), .ZN(P2_U3218) );
  NAND2_X1 U9964 ( .A1(n8505), .A2(n8504), .ZN(n8568) );
  OR2_X1 U9965 ( .A1(n8568), .A2(n8569), .ZN(n8566) );
  AOI21_X1 U9966 ( .B1(n8566), .B2(n8506), .A(n8627), .ZN(n8511) );
  NOR3_X1 U9967 ( .A1(n8507), .A2(n8513), .A3(n8608), .ZN(n8510) );
  AND2_X1 U9968 ( .A1(n8509), .A2(n8508), .ZN(n8576) );
  OAI21_X1 U9969 ( .B1(n8511), .B2(n8510), .A(n8576), .ZN(n8517) );
  NOR2_X1 U9970 ( .A1(n8624), .A2(n8833), .ZN(n8515) );
  OAI22_X1 U9971 ( .A1(n8513), .A2(n8584), .B1(n8583), .B2(n8512), .ZN(n8514)
         );
  AOI211_X1 U9972 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3152), .A(n8515), 
        .B(n8514), .ZN(n8516) );
  OAI211_X1 U9973 ( .C1(n8518), .C2(n8617), .A(n8517), .B(n8516), .ZN(P2_U3225) );
  INV_X1 U9974 ( .A(n8519), .ZN(n8763) );
  NAND2_X1 U9975 ( .A1(n8733), .A2(n8914), .ZN(n8521) );
  NAND2_X1 U9976 ( .A1(n5099), .A2(n8912), .ZN(n8520) );
  NAND2_X1 U9977 ( .A1(n8521), .A2(n8520), .ZN(n8767) );
  AOI22_X1 U9978 ( .A1(n8622), .A2(n8767), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8522) );
  OAI21_X1 U9979 ( .B1(n8763), .B2(n8624), .A(n8522), .ZN(n8528) );
  NAND3_X1 U9980 ( .A1(n8524), .A2(n8629), .A3(n8644), .ZN(n8525) );
  OAI21_X1 U9981 ( .B1(n8526), .B2(n8627), .A(n8525), .ZN(n8527) );
  XNOR2_X1 U9982 ( .A(n8530), .B(n8529), .ZN(n8632) );
  AOI22_X1 U9983 ( .A1(n8632), .A2(n8630), .B1(n8531), .B2(n8530), .ZN(n8535)
         );
  XNOR2_X1 U9984 ( .A(n8533), .B(n8532), .ZN(n8534) );
  XNOR2_X1 U9985 ( .A(n8535), .B(n8534), .ZN(n8541) );
  OAI22_X1 U9986 ( .A1(n8624), .A2(n8922), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8536), .ZN(n8539) );
  OAI22_X1 U9987 ( .A1(n8537), .A2(n8584), .B1(n8583), .B2(n8612), .ZN(n8538)
         );
  AOI211_X1 U9988 ( .C1(n9050), .C2(n8638), .A(n8539), .B(n8538), .ZN(n8540)
         );
  OAI21_X1 U9989 ( .B1(n8541), .B2(n8627), .A(n8540), .ZN(P2_U3228) );
  AOI21_X1 U9990 ( .B1(n8543), .B2(n8542), .A(n8627), .ZN(n8545) );
  NAND2_X1 U9991 ( .A1(n8545), .A2(n8544), .ZN(n8552) );
  OAI22_X1 U9992 ( .A1(n8546), .A2(n8934), .B1(n8935), .B2(n8932), .ZN(n8898)
         );
  INV_X1 U9993 ( .A(n8898), .ZN(n8548) );
  OAI22_X1 U9994 ( .A1(n8549), .A2(n8548), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8547), .ZN(n8550) );
  AOI21_X1 U9995 ( .B1(n8904), .B2(n8635), .A(n8550), .ZN(n8551) );
  OAI211_X1 U9996 ( .C1(n8906), .C2(n8617), .A(n8552), .B(n8551), .ZN(P2_U3230) );
  NOR2_X1 U9997 ( .A1(n8554), .A2(n8553), .ZN(n8556) );
  XNOR2_X1 U9998 ( .A(n8556), .B(n8555), .ZN(n8560) );
  OAI22_X1 U9999 ( .A1(n8560), .A2(n8627), .B1(n8557), .B2(n8608), .ZN(n8558)
         );
  OAI21_X1 U10000 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8565) );
  NOR2_X1 U10001 ( .A1(n8561), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8563) );
  OAI22_X1 U10002 ( .A1(n8810), .A2(n8584), .B1(n8583), .B2(n8779), .ZN(n8562)
         );
  AOI211_X1 U10003 ( .C1(n8635), .C2(n8785), .A(n8563), .B(n8562), .ZN(n8564)
         );
  OAI211_X1 U10004 ( .C1(n8782), .C2(n8617), .A(n8565), .B(n8564), .ZN(
        P2_U3231) );
  INV_X1 U10005 ( .A(n8566), .ZN(n8567) );
  AOI211_X1 U10006 ( .C1(n8569), .C2(n8568), .A(n8627), .B(n8567), .ZN(n8573)
         );
  AOI22_X1 U10007 ( .A1(n8635), .A2(n8850), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8571) );
  AOI22_X1 U10008 ( .A1(n8637), .A2(n8846), .B1(n8636), .B2(n8847), .ZN(n8570)
         );
  OAI211_X1 U10009 ( .C1(n8855), .C2(n8617), .A(n8571), .B(n8570), .ZN(n8572)
         );
  OR2_X1 U10010 ( .A1(n8573), .A2(n8572), .ZN(P2_U3235) );
  INV_X1 U10011 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U10012 ( .A1(n8576), .A2(n8575), .ZN(n8578) );
  XNOR2_X1 U10013 ( .A(n8578), .B(n8577), .ZN(n8580) );
  NAND3_X1 U10014 ( .A1(n8580), .A2(n8631), .A3(n8579), .ZN(n8589) );
  INV_X1 U10015 ( .A(n8580), .ZN(n8581) );
  NAND3_X1 U10016 ( .A1(n8581), .A2(n8629), .A3(n8831), .ZN(n8588) );
  OAI22_X1 U10017 ( .A1(n8624), .A2(n8816), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8582), .ZN(n8586) );
  OAI22_X1 U10018 ( .A1(n8809), .A2(n8584), .B1(n8583), .B2(n8810), .ZN(n8585)
         );
  AOI211_X1 U10019 ( .C1(n9019), .C2(n8638), .A(n8586), .B(n8585), .ZN(n8587)
         );
  NAND3_X1 U10020 ( .A1(n8589), .A2(n8588), .A3(n8587), .ZN(P2_U3237) );
  XNOR2_X1 U10021 ( .A(n8591), .B(n8590), .ZN(n8601) );
  AOI21_X1 U10022 ( .B1(n8598), .B2(n8593), .A(n8592), .ZN(n8594) );
  NOR3_X1 U10023 ( .A1(n8627), .A2(n8601), .A3(n8594), .ZN(n8595) );
  AOI21_X1 U10024 ( .B1(n8962), .B2(n8638), .A(n8595), .ZN(n8605) );
  AOI22_X1 U10025 ( .A1(n8622), .A2(n8597), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8596), .ZN(n8604) );
  OAI22_X1 U10026 ( .A1(n8599), .A2(n8608), .B1(n8627), .B2(n8598), .ZN(n8602)
         );
  NAND3_X1 U10027 ( .A1(n8602), .A2(n8601), .A3(n8600), .ZN(n8603) );
  NAND3_X1 U10028 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(P2_U3239) );
  INV_X1 U10029 ( .A(n8606), .ZN(n8607) );
  AOI21_X1 U10030 ( .B1(n8544), .B2(n8607), .A(n8627), .ZN(n8611) );
  NOR3_X1 U10031 ( .A1(n8609), .A2(n8612), .A3(n8608), .ZN(n8610) );
  OAI21_X1 U10032 ( .B1(n8611), .B2(n8610), .A(n4707), .ZN(n8616) );
  OAI22_X1 U10033 ( .A1(n8613), .A2(n8934), .B1(n8612), .B2(n8932), .ZN(n8883)
         );
  AND2_X1 U10034 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8690) );
  NOR2_X1 U10035 ( .A1(n8624), .A2(n8885), .ZN(n8614) );
  AOI211_X1 U10036 ( .C1(n8622), .C2(n8883), .A(n8690), .B(n8614), .ZN(n8615)
         );
  OAI211_X1 U10037 ( .C1(n4846), .C2(n8617), .A(n8616), .B(n8615), .ZN(
        P2_U3240) );
  XNOR2_X1 U10038 ( .A(n8619), .B(n8618), .ZN(n8628) );
  NAND2_X1 U10039 ( .A1(n8719), .A2(n8914), .ZN(n8621) );
  NAND2_X1 U10040 ( .A1(n8644), .A2(n8912), .ZN(n8620) );
  NAND2_X1 U10041 ( .A1(n8621), .A2(n8620), .ZN(n8754) );
  AOI22_X1 U10042 ( .A1(n8754), .A2(n8622), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8623) );
  OAI21_X1 U10043 ( .B1(n8758), .B2(n8624), .A(n8623), .ZN(n8625) );
  AOI21_X1 U10044 ( .B1(n8998), .B2(n8638), .A(n8625), .ZN(n8626) );
  OAI21_X1 U10045 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(P2_U3242) );
  NAND2_X1 U10046 ( .A1(n8629), .A2(n8913), .ZN(n8634) );
  NAND2_X1 U10047 ( .A1(n8631), .A2(n8630), .ZN(n8633) );
  MUX2_X1 U10048 ( .A(n8634), .B(n8633), .S(n8632), .Z(n8642) );
  AOI22_X1 U10049 ( .A1(n8635), .A2(n8945), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8641) );
  AOI22_X1 U10050 ( .A1(n8637), .A2(n8648), .B1(n8636), .B2(n8647), .ZN(n8640)
         );
  NAND2_X1 U10051 ( .A1(n9056), .A2(n8638), .ZN(n8639) );
  NAND4_X1 U10052 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), .ZN(
        P2_U3243) );
  MUX2_X1 U10053 ( .A(n8643), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8661), .Z(
        P2_U3582) );
  MUX2_X1 U10054 ( .A(n8740), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8661), .Z(
        P2_U3580) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8719), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10056 ( .A(n8733), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8661), .Z(
        P2_U3578) );
  MUX2_X1 U10057 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8644), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10058 ( .A(n5099), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8661), .Z(
        P2_U3576) );
  MUX2_X1 U10059 ( .A(n8645), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8661), .Z(
        P2_U3575) );
  MUX2_X1 U10060 ( .A(n8831), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8661), .Z(
        P2_U3574) );
  MUX2_X1 U10061 ( .A(n8847), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8661), .Z(
        P2_U3573) );
  MUX2_X1 U10062 ( .A(n8830), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8661), .Z(
        P2_U3572) );
  MUX2_X1 U10063 ( .A(n8846), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8661), .Z(
        P2_U3571) );
  MUX2_X1 U10064 ( .A(n8646), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8661), .Z(
        P2_U3570) );
  MUX2_X1 U10065 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8915), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10066 ( .A(n8647), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8661), .Z(
        P2_U3568) );
  MUX2_X1 U10067 ( .A(n8913), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8661), .Z(
        P2_U3567) );
  MUX2_X1 U10068 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8648), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10069 ( .A(n8649), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8661), .Z(
        P2_U3565) );
  MUX2_X1 U10070 ( .A(n8650), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8661), .Z(
        P2_U3564) );
  MUX2_X1 U10071 ( .A(n8651), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8661), .Z(
        P2_U3563) );
  MUX2_X1 U10072 ( .A(n8652), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8661), .Z(
        P2_U3562) );
  MUX2_X1 U10073 ( .A(n8653), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8661), .Z(
        P2_U3561) );
  MUX2_X1 U10074 ( .A(n8654), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8661), .Z(
        P2_U3560) );
  MUX2_X1 U10075 ( .A(n8655), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8661), .Z(
        P2_U3559) );
  MUX2_X1 U10076 ( .A(n8656), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8661), .Z(
        P2_U3558) );
  MUX2_X1 U10077 ( .A(n8657), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8661), .Z(
        P2_U3557) );
  MUX2_X1 U10078 ( .A(n8658), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8661), .Z(
        P2_U3556) );
  MUX2_X1 U10079 ( .A(n8659), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8661), .Z(
        P2_U3555) );
  MUX2_X1 U10080 ( .A(n6468), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8661), .Z(
        P2_U3554) );
  MUX2_X1 U10081 ( .A(n8660), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8661), .Z(
        P2_U3553) );
  MUX2_X1 U10082 ( .A(n6469), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8661), .Z(
        P2_U3552) );
  INV_X1 U10083 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10135) );
  AOI21_X1 U10084 ( .B1(n8663), .B2(n10135), .A(n8662), .ZN(n8665) );
  XNOR2_X1 U10085 ( .A(n8684), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U10086 ( .A1(n8664), .A2(n8665), .ZN(n8683) );
  OAI211_X1 U10087 ( .C1(n8665), .C2(n8664), .A(n9973), .B(n8683), .ZN(n8676)
         );
  NAND2_X1 U10088 ( .A1(n8678), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8668) );
  OAI21_X1 U10089 ( .B1(n8678), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8668), .ZN(
        n8669) );
  AOI211_X1 U10090 ( .C1(n8670), .C2(n8669), .A(n8677), .B(n9976), .ZN(n8674)
         );
  AND2_X1 U10091 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8671) );
  AOI21_X1 U10092 ( .B1(n9975), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8671), .ZN(
        n8672) );
  OAI21_X1 U10093 ( .B1(n9977), .B2(n8684), .A(n8672), .ZN(n8673) );
  NOR2_X1 U10094 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  NAND2_X1 U10095 ( .A1(n8676), .A2(n8675), .ZN(P2_U3262) );
  INV_X1 U10096 ( .A(n8681), .ZN(n8693) );
  NOR2_X1 U10097 ( .A1(n6272), .A2(n8679), .ZN(n8698) );
  AOI211_X1 U10098 ( .C1(n6272), .C2(n8679), .A(n8698), .B(n9976), .ZN(n8680)
         );
  INV_X1 U10099 ( .A(n8680), .ZN(n8692) );
  OR2_X1 U10100 ( .A1(n8681), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U10101 ( .A1(n8681), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U10102 ( .A1(n8694), .A2(n8682), .ZN(n8687) );
  OAI21_X1 U10103 ( .B1(n8685), .B2(n8684), .A(n8683), .ZN(n8686) );
  OR2_X1 U10104 ( .A1(n8687), .A2(n8686), .ZN(n8695) );
  NAND2_X1 U10105 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  AOI21_X1 U10106 ( .B1(n8695), .B2(n8688), .A(n9978), .ZN(n8689) );
  AOI211_X1 U10107 ( .C1(n9975), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8690), .B(
        n8689), .ZN(n8691) );
  OAI211_X1 U10108 ( .C1(n9977), .C2(n8693), .A(n8692), .B(n8691), .ZN(
        P2_U3263) );
  NAND2_X1 U10109 ( .A1(n8695), .A2(n8694), .ZN(n8696) );
  XNOR2_X1 U10110 ( .A(n8696), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8699) );
  INV_X1 U10111 ( .A(n8699), .ZN(n8700) );
  NAND2_X1 U10112 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8701) );
  INV_X1 U10113 ( .A(n8978), .ZN(n8708) );
  XNOR2_X1 U10114 ( .A(n8707), .B(n8977), .ZN(n8975) );
  NAND2_X1 U10115 ( .A1(n8975), .A2(n8944), .ZN(n8706) );
  NAND2_X1 U10116 ( .A1(n8704), .A2(n8703), .ZN(n8980) );
  NOR2_X1 U10117 ( .A1(n9998), .A2(n8980), .ZN(n8710) );
  AOI21_X1 U10118 ( .B1(n9998), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8710), .ZN(
        n8705) );
  OAI211_X1 U10119 ( .C1(n8948), .C2(n8977), .A(n8706), .B(n8705), .ZN(
        P2_U3265) );
  OAI21_X1 U10120 ( .B1(n4271), .B2(n8708), .A(n8707), .ZN(n8981) );
  NOR2_X1 U10121 ( .A1(n9996), .A2(n8709), .ZN(n8711) );
  AOI211_X1 U10122 ( .C1(n8978), .C2(n8963), .A(n8711), .B(n8710), .ZN(n8712)
         );
  OAI21_X1 U10123 ( .B1(n8981), .B2(n8713), .A(n8712), .ZN(P2_U3266) );
  XNOR2_X1 U10124 ( .A(n8715), .B(n8714), .ZN(n8991) );
  OAI211_X1 U10125 ( .C1(n8718), .C2(n8717), .A(n8716), .B(n8917), .ZN(n8721)
         );
  NAND2_X1 U10126 ( .A1(n8719), .A2(n8912), .ZN(n8720) );
  OAI211_X1 U10127 ( .C1(n8722), .C2(n8934), .A(n8721), .B(n8720), .ZN(n8987)
         );
  INV_X1 U10128 ( .A(n8741), .ZN(n8725) );
  INV_X1 U10129 ( .A(n8723), .ZN(n8724) );
  AOI21_X1 U10130 ( .B1(n4855), .B2(n8725), .A(n8724), .ZN(n8988) );
  NAND2_X1 U10131 ( .A1(n8988), .A2(n8944), .ZN(n8728) );
  AOI22_X1 U10132 ( .A1(n9998), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8726), .B2(
        n8955), .ZN(n8727) );
  OAI211_X1 U10133 ( .C1(n8729), .C2(n8948), .A(n8728), .B(n8727), .ZN(n8730)
         );
  AOI21_X1 U10134 ( .B1(n8987), .B2(n9996), .A(n8730), .ZN(n8731) );
  OAI21_X1 U10135 ( .B1(n8991), .B2(n8890), .A(n8731), .ZN(P2_U3268) );
  XNOR2_X1 U10136 ( .A(n8732), .B(n8737), .ZN(n8996) );
  INV_X1 U10137 ( .A(n8766), .ZN(n8735) );
  NAND2_X1 U10138 ( .A1(n8735), .A2(n8734), .ZN(n8769) );
  NAND2_X1 U10139 ( .A1(n8769), .A2(n8736), .ZN(n8751) );
  OR2_X1 U10140 ( .A1(n8995), .A2(n9998), .ZN(n8748) );
  INV_X1 U10141 ( .A(n8756), .ZN(n8742) );
  AOI21_X1 U10142 ( .B1(n8992), .B2(n8742), .A(n8741), .ZN(n8993) );
  AOI22_X1 U10143 ( .A1(n9998), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8743), .B2(
        n8955), .ZN(n8744) );
  OAI21_X1 U10144 ( .B1(n8745), .B2(n8948), .A(n8744), .ZN(n8746) );
  AOI21_X1 U10145 ( .B1(n8993), .B2(n8944), .A(n8746), .ZN(n8747) );
  OAI211_X1 U10146 ( .C1(n8996), .C2(n8890), .A(n8748), .B(n8747), .ZN(
        P2_U3269) );
  XNOR2_X1 U10147 ( .A(n8749), .B(n8752), .ZN(n9001) );
  AND2_X1 U10148 ( .A1(n8769), .A2(n8750), .ZN(n8753) );
  OAI21_X1 U10149 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8755) );
  AOI21_X1 U10150 ( .B1(n8755), .B2(n8917), .A(n8754), .ZN(n9000) );
  AOI211_X1 U10151 ( .C1(n8998), .C2(n8770), .A(n10022), .B(n8756), .ZN(n8997)
         );
  NAND2_X1 U10152 ( .A1(n8997), .A2(n6532), .ZN(n8757) );
  OAI211_X1 U10153 ( .C1(n9990), .C2(n8758), .A(n9000), .B(n8757), .ZN(n8759)
         );
  NAND2_X1 U10154 ( .A1(n8759), .A2(n9996), .ZN(n8761) );
  AOI22_X1 U10155 ( .A1(n8998), .A2(n8963), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n9998), .ZN(n8760) );
  OAI211_X1 U10156 ( .C1(n9001), .C2(n8890), .A(n8761), .B(n8760), .ZN(
        P2_U3270) );
  XNOR2_X1 U10157 ( .A(n8762), .B(n8765), .ZN(n9006) );
  OAI22_X1 U10158 ( .A1(n9996), .A2(n8764), .B1(n8763), .B2(n9990), .ZN(n8774)
         );
  AOI21_X1 U10159 ( .B1(n8766), .B2(n8765), .A(n8930), .ZN(n8768) );
  AOI21_X1 U10160 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(n9005) );
  INV_X1 U10161 ( .A(n8770), .ZN(n8771) );
  AOI211_X1 U10162 ( .C1(n9003), .C2(n8784), .A(n10022), .B(n8771), .ZN(n9002)
         );
  NAND2_X1 U10163 ( .A1(n9002), .A2(n6532), .ZN(n8772) );
  AOI21_X1 U10164 ( .B1(n9005), .B2(n8772), .A(n9998), .ZN(n8773) );
  AOI211_X1 U10165 ( .C1(n8963), .C2(n9003), .A(n8774), .B(n8773), .ZN(n8775)
         );
  OAI21_X1 U10166 ( .B1(n9006), .B2(n8890), .A(n8775), .ZN(P2_U3271) );
  AOI211_X1 U10167 ( .C1(n8778), .C2(n8777), .A(n8930), .B(n8776), .ZN(n8781)
         );
  OAI22_X1 U10168 ( .A1(n8779), .A2(n8934), .B1(n8810), .B2(n8932), .ZN(n8780)
         );
  NOR2_X1 U10169 ( .A1(n8781), .A2(n8780), .ZN(n9010) );
  OR2_X1 U10170 ( .A1(n4260), .A2(n8782), .ZN(n8783) );
  AND2_X1 U10171 ( .A1(n8784), .A2(n8783), .ZN(n9008) );
  NAND2_X1 U10172 ( .A1(n9007), .A2(n8963), .ZN(n8787) );
  NAND2_X1 U10173 ( .A1(n8785), .A2(n8955), .ZN(n8786) );
  OAI211_X1 U10174 ( .C1(n9996), .C2(n8788), .A(n8787), .B(n8786), .ZN(n8793)
         );
  AOI21_X1 U10175 ( .B1(n8791), .B2(n8790), .A(n8789), .ZN(n9011) );
  NOR2_X1 U10176 ( .A1(n9011), .A2(n8890), .ZN(n8792) );
  AOI211_X1 U10177 ( .C1(n9008), .C2(n8944), .A(n8793), .B(n8792), .ZN(n8794)
         );
  OAI21_X1 U10178 ( .B1(n9998), .B2(n9010), .A(n8794), .ZN(P2_U3272) );
  OAI21_X1 U10179 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8798) );
  AOI222_X1 U10180 ( .A1(n8917), .A2(n8798), .B1(n5099), .B2(n8914), .C1(n8831), .C2(n8912), .ZN(n9018) );
  AOI21_X1 U10181 ( .B1(n9012), .B2(n8814), .A(n4260), .ZN(n9013) );
  AOI22_X1 U10182 ( .A1(n9998), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8799), .B2(
        n8955), .ZN(n8800) );
  OAI21_X1 U10183 ( .B1(n8801), .B2(n8948), .A(n8800), .ZN(n8802) );
  AOI21_X1 U10184 ( .B1(n9013), .B2(n8944), .A(n8802), .ZN(n8806) );
  OR2_X1 U10185 ( .A1(n8804), .A2(n8803), .ZN(n9015) );
  NAND3_X1 U10186 ( .A1(n9015), .A2(n9014), .A3(n8965), .ZN(n8805) );
  OAI211_X1 U10187 ( .C1(n9018), .C2(n9998), .A(n8806), .B(n8805), .ZN(
        P2_U3273) );
  OR2_X1 U10188 ( .A1(n8825), .A2(n8826), .ZN(n8827) );
  NAND2_X1 U10189 ( .A1(n8827), .A2(n8807), .ZN(n8808) );
  XOR2_X1 U10190 ( .A(n8819), .B(n8808), .Z(n8812) );
  OAI22_X1 U10191 ( .A1(n8810), .A2(n8934), .B1(n8809), .B2(n8932), .ZN(n8811)
         );
  AOI21_X1 U10192 ( .B1(n8812), .B2(n8917), .A(n8811), .ZN(n9022) );
  INV_X1 U10193 ( .A(n8814), .ZN(n8815) );
  AOI21_X1 U10194 ( .B1(n9019), .B2(n8837), .A(n8815), .ZN(n9020) );
  INV_X1 U10195 ( .A(n8816), .ZN(n8817) );
  AOI22_X1 U10196 ( .A1(n9998), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8817), .B2(
        n8955), .ZN(n8818) );
  OAI21_X1 U10197 ( .B1(n8355), .B2(n8948), .A(n8818), .ZN(n8822) );
  XOR2_X1 U10198 ( .A(n8820), .B(n8819), .Z(n9023) );
  NOR2_X1 U10199 ( .A1(n9023), .A2(n8890), .ZN(n8821) );
  AOI211_X1 U10200 ( .C1(n9020), .C2(n8944), .A(n8822), .B(n8821), .ZN(n8823)
         );
  OAI21_X1 U10201 ( .B1(n9998), .B2(n9022), .A(n8823), .ZN(P2_U3274) );
  XNOR2_X1 U10202 ( .A(n8824), .B(n8826), .ZN(n9028) );
  INV_X1 U10203 ( .A(n8825), .ZN(n8829) );
  INV_X1 U10204 ( .A(n8826), .ZN(n8828) );
  OAI21_X1 U10205 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8832) );
  AOI222_X1 U10206 ( .A1(n8917), .A2(n8832), .B1(n8831), .B2(n8914), .C1(n8830), .C2(n8912), .ZN(n9027) );
  OAI22_X1 U10207 ( .A1(n9996), .A2(n8834), .B1(n8833), .B2(n9990), .ZN(n8835)
         );
  AOI21_X1 U10208 ( .B1(n9024), .B2(n8963), .A(n8835), .ZN(n8839) );
  NAND2_X1 U10209 ( .A1(n8857), .A2(n9024), .ZN(n8836) );
  AND2_X1 U10210 ( .A1(n8837), .A2(n8836), .ZN(n9025) );
  NAND2_X1 U10211 ( .A1(n9025), .A2(n8944), .ZN(n8838) );
  OAI211_X1 U10212 ( .C1(n9027), .C2(n9998), .A(n8839), .B(n8838), .ZN(n8840)
         );
  INV_X1 U10213 ( .A(n8840), .ZN(n8841) );
  OAI21_X1 U10214 ( .B1(n9028), .B2(n8890), .A(n8841), .ZN(P2_U3275) );
  XNOR2_X1 U10215 ( .A(n8842), .B(n8844), .ZN(n9033) );
  OAI211_X1 U10216 ( .C1(n8845), .C2(n8844), .A(n8843), .B(n8917), .ZN(n8849)
         );
  AOI22_X1 U10217 ( .A1(n8847), .A2(n8914), .B1(n8912), .B2(n8846), .ZN(n8848)
         );
  INV_X1 U10218 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8852) );
  INV_X1 U10219 ( .A(n8850), .ZN(n8851) );
  OAI22_X1 U10220 ( .A1(n9996), .A2(n8852), .B1(n8851), .B2(n9990), .ZN(n8853)
         );
  AOI21_X1 U10221 ( .B1(n9029), .B2(n8963), .A(n8853), .ZN(n8859) );
  OR2_X1 U10222 ( .A1(n8855), .A2(n8854), .ZN(n8856) );
  AND2_X1 U10223 ( .A1(n8857), .A2(n8856), .ZN(n9030) );
  NAND2_X1 U10224 ( .A1(n9030), .A2(n8944), .ZN(n8858) );
  OAI211_X1 U10225 ( .C1(n9032), .C2(n9998), .A(n8859), .B(n8858), .ZN(n8860)
         );
  INV_X1 U10226 ( .A(n8860), .ZN(n8861) );
  OAI21_X1 U10227 ( .B1(n8890), .B2(n9033), .A(n8861), .ZN(P2_U3276) );
  XOR2_X1 U10228 ( .A(n8864), .B(n8862), .Z(n9037) );
  INV_X1 U10229 ( .A(n8863), .ZN(n8877) );
  XOR2_X1 U10230 ( .A(n8865), .B(n8864), .Z(n8867) );
  OAI21_X1 U10231 ( .B1(n8867), .B2(n8930), .A(n8866), .ZN(n8871) );
  XNOR2_X1 U10232 ( .A(n4316), .B(n9034), .ZN(n8868) );
  AOI21_X1 U10233 ( .B1(n9091), .B2(n8868), .A(n8871), .ZN(n9036) );
  OAI21_X1 U10234 ( .B1(n9037), .B2(n8869), .A(n9036), .ZN(n8870) );
  OAI211_X1 U10235 ( .C1(n6532), .C2(n8871), .A(n8870), .B(n9996), .ZN(n8876)
         );
  OAI22_X1 U10236 ( .A1(n9996), .A2(n8873), .B1(n8872), .B2(n9990), .ZN(n8874)
         );
  AOI21_X1 U10237 ( .B1(n9034), .B2(n8963), .A(n8874), .ZN(n8875) );
  OAI211_X1 U10238 ( .C1(n9037), .C2(n8877), .A(n8876), .B(n8875), .ZN(
        P2_U3277) );
  NAND2_X1 U10239 ( .A1(n8911), .A2(n8926), .ZN(n8910) );
  NAND2_X1 U10240 ( .A1(n8910), .A2(n8878), .ZN(n8897) );
  NOR2_X1 U10241 ( .A1(n8897), .A2(n8902), .ZN(n8896) );
  NAND2_X1 U10242 ( .A1(n4437), .A2(n8879), .ZN(n8882) );
  OAI21_X1 U10243 ( .B1(n8896), .B2(n8880), .A(n8889), .ZN(n8881) );
  OAI21_X1 U10244 ( .B1(n8896), .B2(n8882), .A(n8881), .ZN(n8884) );
  AOI21_X1 U10245 ( .B1(n8884), .B2(n8917), .A(n8883), .ZN(n9041) );
  AOI211_X1 U10246 ( .C1(n9039), .C2(n8894), .A(n10022), .B(n4316), .ZN(n9038)
         );
  INV_X1 U10247 ( .A(n8885), .ZN(n8886) );
  AOI22_X1 U10248 ( .A1(n9998), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8886), .B2(
        n8955), .ZN(n8887) );
  OAI21_X1 U10249 ( .B1(n4846), .B2(n8948), .A(n8887), .ZN(n8892) );
  XOR2_X1 U10250 ( .A(n8889), .B(n8888), .Z(n9042) );
  NOR2_X1 U10251 ( .A1(n9042), .A2(n8890), .ZN(n8891) );
  AOI211_X1 U10252 ( .C1(n9038), .C2(n8969), .A(n8892), .B(n8891), .ZN(n8893)
         );
  OAI21_X1 U10253 ( .B1(n9041), .B2(n9998), .A(n8893), .ZN(P2_U3278) );
  INV_X1 U10254 ( .A(n8894), .ZN(n8895) );
  AOI211_X1 U10255 ( .C1(n9045), .C2(n8918), .A(n10022), .B(n8895), .ZN(n9044)
         );
  AOI211_X1 U10256 ( .C1(n8902), .C2(n8897), .A(n8930), .B(n8896), .ZN(n8899)
         );
  NOR2_X1 U10257 ( .A1(n8899), .A2(n8898), .ZN(n9047) );
  INV_X1 U10258 ( .A(n9047), .ZN(n8900) );
  AOI21_X1 U10259 ( .B1(n9044), .B2(n6532), .A(n8900), .ZN(n8909) );
  OAI21_X1 U10260 ( .B1(n8903), .B2(n8902), .A(n8901), .ZN(n9043) );
  AOI22_X1 U10261 ( .A1(n9998), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8904), .B2(
        n8955), .ZN(n8905) );
  OAI21_X1 U10262 ( .B1(n8906), .B2(n8948), .A(n8905), .ZN(n8907) );
  AOI21_X1 U10263 ( .B1(n9043), .B2(n8965), .A(n8907), .ZN(n8908) );
  OAI21_X1 U10264 ( .B1(n8909), .B2(n9998), .A(n8908), .ZN(P2_U3279) );
  OAI21_X1 U10265 ( .B1(n8926), .B2(n8911), .A(n8910), .ZN(n8916) );
  AOI222_X1 U10266 ( .A1(n8917), .A2(n8916), .B1(n8915), .B2(n8914), .C1(n8913), .C2(n8912), .ZN(n9053) );
  INV_X1 U10267 ( .A(n8942), .ZN(n8920) );
  INV_X1 U10268 ( .A(n8918), .ZN(n8919) );
  AOI21_X1 U10269 ( .B1(n9050), .B2(n8920), .A(n8919), .ZN(n9051) );
  NOR2_X1 U10270 ( .A1(n8921), .A2(n8948), .ZN(n8924) );
  OAI22_X1 U10271 ( .A1(n9996), .A2(n10063), .B1(n8922), .B2(n9990), .ZN(n8923) );
  AOI211_X1 U10272 ( .C1(n9051), .C2(n8944), .A(n8924), .B(n8923), .ZN(n8928)
         );
  AOI21_X1 U10273 ( .B1(n8926), .B2(n8925), .A(n4323), .ZN(n9049) );
  NAND2_X1 U10274 ( .A1(n9049), .A2(n8965), .ZN(n8927) );
  OAI211_X1 U10275 ( .C1(n9053), .C2(n9998), .A(n8928), .B(n8927), .ZN(
        P2_U3280) );
  AOI211_X1 U10276 ( .C1(n8931), .C2(n8939), .A(n8930), .B(n8929), .ZN(n8937)
         );
  OAI22_X1 U10277 ( .A1(n8935), .A2(n8934), .B1(n8933), .B2(n8932), .ZN(n8936)
         );
  NOR2_X1 U10278 ( .A1(n8937), .A2(n8936), .ZN(n9059) );
  OAI21_X1 U10279 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n9055) );
  INV_X1 U10280 ( .A(n8941), .ZN(n8943) );
  AOI21_X1 U10281 ( .B1(n9056), .B2(n8943), .A(n8942), .ZN(n9057) );
  NAND2_X1 U10282 ( .A1(n9057), .A2(n8944), .ZN(n8947) );
  AOI22_X1 U10283 ( .A1(n9998), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8945), .B2(
        n8955), .ZN(n8946) );
  OAI211_X1 U10284 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8950)
         );
  AOI21_X1 U10285 ( .B1(n8965), .B2(n9055), .A(n8950), .ZN(n8951) );
  OAI21_X1 U10286 ( .B1(n9059), .B2(n9998), .A(n8951), .ZN(P2_U3281) );
  AOI22_X1 U10287 ( .A1(n8965), .A2(n8953), .B1(n8963), .B2(n8952), .ZN(n8961)
         );
  AOI22_X1 U10288 ( .A1(n8969), .A2(n8956), .B1(n8955), .B2(n8954), .ZN(n8960)
         );
  MUX2_X1 U10289 ( .A(n8958), .B(n8957), .S(n9996), .Z(n8959) );
  NAND3_X1 U10290 ( .A1(n8961), .A2(n8960), .A3(n8959), .ZN(P2_U3293) );
  AOI22_X1 U10291 ( .A1(n8965), .A2(n8964), .B1(n8963), .B2(n8962), .ZN(n8974)
         );
  NOR2_X1 U10292 ( .A1(n9990), .A2(n8966), .ZN(n8967) );
  AOI21_X1 U10293 ( .B1(n8969), .B2(n8968), .A(n8967), .ZN(n8973) );
  MUX2_X1 U10294 ( .A(n8971), .B(n8970), .S(n9996), .Z(n8972) );
  NAND3_X1 U10295 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(P2_U3294) );
  NAND2_X1 U10296 ( .A1(n8975), .A2(n9091), .ZN(n8976) );
  OAI211_X1 U10297 ( .C1(n8977), .C2(n10020), .A(n8976), .B(n8980), .ZN(n9097)
         );
  MUX2_X1 U10298 ( .A(n9097), .B(P2_REG1_REG_31__SCAN_IN), .S(n4315), .Z(
        P2_U3551) );
  NAND2_X1 U10299 ( .A1(n8978), .A2(n9090), .ZN(n8979) );
  OAI211_X1 U10300 ( .C1(n8981), .C2(n10022), .A(n8980), .B(n8979), .ZN(n9098)
         );
  MUX2_X1 U10301 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9098), .S(n4333), .Z(
        P2_U3550) );
  AOI22_X1 U10302 ( .A1(n8983), .A2(n9091), .B1(n9090), .B2(n8982), .ZN(n8984)
         );
  INV_X1 U10303 ( .A(n8987), .ZN(n8990) );
  AOI22_X1 U10304 ( .A1(n8988), .A2(n9091), .B1(n9090), .B2(n4855), .ZN(n8989)
         );
  OAI211_X1 U10305 ( .C1(n8991), .C2(n9081), .A(n8990), .B(n8989), .ZN(n9099)
         );
  MUX2_X1 U10306 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9099), .S(n4333), .Z(
        P2_U3548) );
  AOI22_X1 U10307 ( .A1(n8993), .A2(n9091), .B1(n9090), .B2(n8992), .ZN(n8994)
         );
  MUX2_X1 U10308 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9100), .S(n4333), .Z(
        P2_U3547) );
  AOI21_X1 U10309 ( .B1(n9090), .B2(n8998), .A(n8997), .ZN(n8999) );
  OAI211_X1 U10310 ( .C1(n9001), .C2(n9081), .A(n9000), .B(n8999), .ZN(n9101)
         );
  MUX2_X1 U10311 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9101), .S(n4333), .Z(
        P2_U3546) );
  AOI21_X1 U10312 ( .B1(n9090), .B2(n9003), .A(n9002), .ZN(n9004) );
  OAI211_X1 U10313 ( .C1(n9006), .C2(n9081), .A(n9005), .B(n9004), .ZN(n9102)
         );
  MUX2_X1 U10314 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9102), .S(n4333), .Z(
        P2_U3545) );
  AOI22_X1 U10315 ( .A1(n9008), .A2(n9091), .B1(n9090), .B2(n9007), .ZN(n9009)
         );
  OAI211_X1 U10316 ( .C1(n9081), .C2(n9011), .A(n9010), .B(n9009), .ZN(n9103)
         );
  MUX2_X1 U10317 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9103), .S(n4333), .Z(
        P2_U3544) );
  AOI22_X1 U10318 ( .A1(n9013), .A2(n9091), .B1(n9090), .B2(n9012), .ZN(n9017)
         );
  NAND3_X1 U10319 ( .A1(n9015), .A2(n9014), .A3(n10028), .ZN(n9016) );
  NAND3_X1 U10320 ( .A1(n9018), .A2(n9017), .A3(n9016), .ZN(n9104) );
  MUX2_X1 U10321 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9104), .S(n4333), .Z(
        P2_U3543) );
  AOI22_X1 U10322 ( .A1(n9020), .A2(n9091), .B1(n9090), .B2(n9019), .ZN(n9021)
         );
  OAI211_X1 U10323 ( .C1(n9081), .C2(n9023), .A(n9022), .B(n9021), .ZN(n9105)
         );
  MUX2_X1 U10324 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9105), .S(n4333), .Z(
        P2_U3542) );
  AOI22_X1 U10325 ( .A1(n9025), .A2(n9091), .B1(n9090), .B2(n9024), .ZN(n9026)
         );
  OAI211_X1 U10326 ( .C1(n9081), .C2(n9028), .A(n9027), .B(n9026), .ZN(n9106)
         );
  MUX2_X1 U10327 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9106), .S(n4333), .Z(
        P2_U3541) );
  AOI22_X1 U10328 ( .A1(n9030), .A2(n9091), .B1(n9090), .B2(n9029), .ZN(n9031)
         );
  OAI211_X1 U10329 ( .C1(n9081), .C2(n9033), .A(n9032), .B(n9031), .ZN(n9107)
         );
  MUX2_X1 U10330 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9107), .S(n4333), .Z(
        P2_U3540) );
  NAND2_X1 U10331 ( .A1(n9034), .A2(n9090), .ZN(n9035) );
  OAI211_X1 U10332 ( .C1(n9081), .C2(n9037), .A(n9036), .B(n9035), .ZN(n9108)
         );
  MUX2_X1 U10333 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9108), .S(n4333), .Z(
        P2_U3539) );
  AOI21_X1 U10334 ( .B1(n9090), .B2(n9039), .A(n9038), .ZN(n9040) );
  OAI211_X1 U10335 ( .C1(n9081), .C2(n9042), .A(n9041), .B(n9040), .ZN(n9109)
         );
  MUX2_X1 U10336 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9109), .S(n4333), .Z(
        P2_U3538) );
  INV_X1 U10337 ( .A(n9043), .ZN(n9048) );
  AOI21_X1 U10338 ( .B1(n9090), .B2(n9045), .A(n9044), .ZN(n9046) );
  OAI211_X1 U10339 ( .C1(n9081), .C2(n9048), .A(n9047), .B(n9046), .ZN(n9110)
         );
  MUX2_X1 U10340 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9110), .S(n4333), .Z(
        P2_U3537) );
  INV_X1 U10341 ( .A(n9049), .ZN(n9054) );
  AOI22_X1 U10342 ( .A1(n9051), .A2(n9091), .B1(n9090), .B2(n9050), .ZN(n9052)
         );
  OAI211_X1 U10343 ( .C1(n9081), .C2(n9054), .A(n9053), .B(n9052), .ZN(n9111)
         );
  MUX2_X1 U10344 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9111), .S(n4333), .Z(
        P2_U3536) );
  INV_X1 U10345 ( .A(n9055), .ZN(n9060) );
  AOI22_X1 U10346 ( .A1(n9057), .A2(n9091), .B1(n9090), .B2(n9056), .ZN(n9058)
         );
  OAI211_X1 U10347 ( .C1(n9081), .C2(n9060), .A(n9059), .B(n9058), .ZN(n9112)
         );
  MUX2_X1 U10348 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9112), .S(n4333), .Z(
        P2_U3535) );
  AOI22_X1 U10349 ( .A1(n9062), .A2(n9091), .B1(n9090), .B2(n9061), .ZN(n9063)
         );
  OAI211_X1 U10350 ( .C1(n9081), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9113)
         );
  MUX2_X1 U10351 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9113), .S(n4333), .Z(
        P2_U3534) );
  AOI22_X1 U10352 ( .A1(n9067), .A2(n9091), .B1(n9090), .B2(n9066), .ZN(n9068)
         );
  OAI211_X1 U10353 ( .C1(n9081), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9114)
         );
  MUX2_X1 U10354 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9114), .S(n4333), .Z(
        P2_U3533) );
  AOI21_X1 U10355 ( .B1(n9090), .B2(n9072), .A(n9071), .ZN(n9073) );
  OAI211_X1 U10356 ( .C1(n9081), .C2(n9075), .A(n9074), .B(n9073), .ZN(n9115)
         );
  MUX2_X1 U10357 ( .A(n9115), .B(P2_REG1_REG_11__SCAN_IN), .S(n4315), .Z(
        P2_U3531) );
  AOI21_X1 U10358 ( .B1(n9090), .B2(n9077), .A(n9076), .ZN(n9078) );
  OAI211_X1 U10359 ( .C1(n9081), .C2(n9080), .A(n9079), .B(n9078), .ZN(n9116)
         );
  MUX2_X1 U10360 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9116), .S(n4333), .Z(
        P2_U3530) );
  INV_X1 U10361 ( .A(n9082), .ZN(n9087) );
  AOI22_X1 U10362 ( .A1(n9084), .A2(n9091), .B1(n9090), .B2(n9083), .ZN(n9085)
         );
  OAI211_X1 U10363 ( .C1(n9096), .C2(n9087), .A(n9086), .B(n9085), .ZN(n9117)
         );
  MUX2_X1 U10364 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9117), .S(n4333), .Z(
        P2_U3529) );
  INV_X1 U10365 ( .A(n9088), .ZN(n9095) );
  AOI22_X1 U10366 ( .A1(n9092), .A2(n9091), .B1(n9090), .B2(n9089), .ZN(n9093)
         );
  OAI211_X1 U10367 ( .C1(n9096), .C2(n9095), .A(n9094), .B(n9093), .ZN(n9118)
         );
  MUX2_X1 U10368 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9118), .S(n4333), .Z(
        P2_U3528) );
  MUX2_X1 U10369 ( .A(n9097), .B(P2_REG0_REG_31__SCAN_IN), .S(n4455), .Z(
        P2_U3519) );
  MUX2_X1 U10370 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9098), .S(n10030), .Z(
        P2_U3518) );
  MUX2_X1 U10371 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9099), .S(n10030), .Z(
        P2_U3516) );
  MUX2_X1 U10372 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9100), .S(n10030), .Z(
        P2_U3515) );
  MUX2_X1 U10373 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9101), .S(n10030), .Z(
        P2_U3514) );
  MUX2_X1 U10374 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9102), .S(n10030), .Z(
        P2_U3513) );
  MUX2_X1 U10375 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9103), .S(n10030), .Z(
        P2_U3512) );
  MUX2_X1 U10376 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9104), .S(n10030), .Z(
        P2_U3511) );
  MUX2_X1 U10377 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9105), .S(n10030), .Z(
        P2_U3510) );
  MUX2_X1 U10378 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9106), .S(n10030), .Z(
        P2_U3509) );
  MUX2_X1 U10379 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9107), .S(n10030), .Z(
        P2_U3508) );
  MUX2_X1 U10380 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9108), .S(n10030), .Z(
        P2_U3507) );
  MUX2_X1 U10381 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9109), .S(n10030), .Z(
        P2_U3505) );
  MUX2_X1 U10382 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9110), .S(n10030), .Z(
        P2_U3502) );
  MUX2_X1 U10383 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9111), .S(n10030), .Z(
        P2_U3499) );
  MUX2_X1 U10384 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9112), .S(n10030), .Z(
        P2_U3496) );
  MUX2_X1 U10385 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9113), .S(n10030), .Z(
        P2_U3493) );
  MUX2_X1 U10386 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9114), .S(n10030), .Z(
        P2_U3490) );
  MUX2_X1 U10387 ( .A(n9115), .B(P2_REG0_REG_11__SCAN_IN), .S(n4455), .Z(
        P2_U3484) );
  MUX2_X1 U10388 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9116), .S(n10030), .Z(
        P2_U3481) );
  MUX2_X1 U10389 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9117), .S(n10030), .Z(
        P2_U3478) );
  MUX2_X1 U10390 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n9118), .S(n10030), .Z(
        P2_U3475) );
  INV_X1 U10391 ( .A(n9119), .ZN(n9750) );
  NOR4_X1 U10392 ( .A1(n9121), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9120), .A4(
        P2_U3152), .ZN(n9122) );
  AOI21_X1 U10393 ( .B1(n9127), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9122), .ZN(
        n9123) );
  OAI21_X1 U10394 ( .B1(n9750), .B2(n7807), .A(n9123), .ZN(P2_U3327) );
  INV_X1 U10395 ( .A(n9124), .ZN(n9751) );
  OAI222_X1 U10396 ( .A1(P2_U3152), .A2(n4235), .B1(n7807), .B2(n9751), .C1(
        n9126), .C2(n9125), .ZN(P2_U3329) );
  NAND2_X1 U10397 ( .A1(n9127), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9128) );
  OAI211_X1 U10398 ( .C1(n9130), .C2(n7807), .A(n9129), .B(n9128), .ZN(
        P2_U3330) );
  MUX2_X1 U10399 ( .A(n9131), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10400 ( .A(n9134), .B(n9133), .ZN(n9135) );
  XNOR2_X1 U10401 ( .A(n9132), .B(n9135), .ZN(n9140) );
  OAI22_X1 U10402 ( .A1(n9382), .A2(n9286), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10075), .ZN(n9136) );
  AOI21_X1 U10403 ( .B1(n9272), .B2(n9415), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10404 ( .B1(n9376), .B2(n9275), .A(n9137), .ZN(n9138) );
  AOI21_X1 U10405 ( .B1(n9634), .B2(n9288), .A(n9138), .ZN(n9139) );
  OAI21_X1 U10406 ( .B1(n9140), .B2(n9278), .A(n9139), .ZN(P1_U3212) );
  NAND2_X1 U10407 ( .A1(n9141), .A2(n9142), .ZN(n9143) );
  XOR2_X1 U10408 ( .A(n9144), .B(n9143), .Z(n9150) );
  NAND2_X1 U10409 ( .A1(n9272), .A2(n9297), .ZN(n9146) );
  OAI211_X1 U10410 ( .C1(n9580), .C2(n9275), .A(n9146), .B(n9145), .ZN(n9148)
         );
  NOR2_X1 U10411 ( .A1(n9584), .A2(n9235), .ZN(n9147) );
  AOI211_X1 U10412 ( .C1(n9587), .C2(n9271), .A(n9148), .B(n9147), .ZN(n9149)
         );
  OAI21_X1 U10413 ( .B1(n9150), .B2(n9278), .A(n9149), .ZN(P1_U3213) );
  INV_X1 U10414 ( .A(n9151), .ZN(n9153) );
  NAND2_X1 U10415 ( .A1(n9153), .A2(n9152), .ZN(n9216) );
  NAND2_X1 U10416 ( .A1(n9151), .A2(n9154), .ZN(n9185) );
  NAND2_X1 U10417 ( .A1(n9216), .A2(n9185), .ZN(n9156) );
  XNOR2_X1 U10418 ( .A(n9156), .B(n9155), .ZN(n9162) );
  OAI22_X1 U10419 ( .A1(n9179), .A2(n9282), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9157), .ZN(n9158) );
  AOI21_X1 U10420 ( .B1(n9444), .B2(n9284), .A(n9158), .ZN(n9159) );
  OAI21_X1 U10421 ( .B1(n9286), .B2(n9436), .A(n9159), .ZN(n9160) );
  AOI21_X1 U10422 ( .B1(n9656), .B2(n9288), .A(n9160), .ZN(n9161) );
  OAI21_X1 U10423 ( .B1(n9162), .B2(n9278), .A(n9161), .ZN(P1_U3214) );
  OR2_X1 U10424 ( .A1(n9163), .A2(n9225), .ZN(n9167) );
  NOR2_X1 U10425 ( .A1(n4255), .A2(n9165), .ZN(n9256) );
  INV_X1 U10426 ( .A(n9164), .ZN(n9259) );
  NAND2_X1 U10427 ( .A1(n4255), .A2(n9165), .ZN(n9257) );
  OAI21_X1 U10428 ( .B1(n9256), .B2(n9259), .A(n9257), .ZN(n9166) );
  NOR2_X1 U10429 ( .A1(n9166), .A2(n9167), .ZN(n9226) );
  AOI21_X1 U10430 ( .B1(n9167), .B2(n9166), .A(n9226), .ZN(n9173) );
  NAND2_X1 U10431 ( .A1(n9272), .A2(n9523), .ZN(n9168) );
  NAND2_X1 U10432 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9346) );
  OAI211_X1 U10433 ( .C1(n9169), .C2(n9275), .A(n9168), .B(n9346), .ZN(n9171)
         );
  NOR2_X1 U10434 ( .A1(n9493), .A2(n9235), .ZN(n9170) );
  AOI211_X1 U10435 ( .C1(n9491), .C2(n9271), .A(n9171), .B(n9170), .ZN(n9172)
         );
  OAI21_X1 U10436 ( .B1(n9173), .B2(n9278), .A(n9172), .ZN(P1_U3217) );
  OAI21_X1 U10437 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9177) );
  NAND2_X1 U10438 ( .A1(n9177), .A2(n5905), .ZN(n9183) );
  NOR2_X1 U10439 ( .A1(n9286), .A2(n9470), .ZN(n9181) );
  OAI22_X1 U10440 ( .A1(n9179), .A2(n9275), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9178), .ZN(n9180) );
  AOI211_X1 U10441 ( .C1(n9272), .C2(n9496), .A(n9181), .B(n9180), .ZN(n9182)
         );
  OAI211_X1 U10442 ( .C1(n5015), .C2(n9235), .A(n9183), .B(n9182), .ZN(
        P1_U3221) );
  INV_X1 U10443 ( .A(n9646), .ZN(n9412) );
  NAND2_X1 U10444 ( .A1(n9185), .A2(n9184), .ZN(n9217) );
  AND2_X1 U10445 ( .A1(n9188), .A2(n9186), .ZN(n9215) );
  NAND3_X1 U10446 ( .A1(n9217), .A2(n9216), .A3(n9215), .ZN(n9214) );
  NAND3_X1 U10447 ( .A1(n9214), .A2(n9188), .A3(n9187), .ZN(n9190) );
  OAI22_X1 U10448 ( .A1(n9192), .A2(n9282), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9191), .ZN(n9194) );
  NOR2_X1 U10449 ( .A1(n9375), .A2(n9275), .ZN(n9193) );
  AOI211_X1 U10450 ( .C1(n9410), .C2(n9271), .A(n9194), .B(n9193), .ZN(n9195)
         );
  NAND2_X1 U10451 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  XNOR2_X1 U10452 ( .A(n4264), .B(n9198), .ZN(n9204) );
  OAI22_X1 U10453 ( .A1(n9275), .A2(n9199), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4701), .ZN(n9200) );
  AOI21_X1 U10454 ( .B1(n9272), .B2(n9541), .A(n9200), .ZN(n9201) );
  OAI21_X1 U10455 ( .B1(n9286), .B2(n9547), .A(n9201), .ZN(n9202) );
  AOI21_X1 U10456 ( .B1(n9693), .B2(n9288), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10457 ( .B1(n9204), .B2(n9278), .A(n9203), .ZN(P1_U3224) );
  OAI21_X1 U10458 ( .B1(n9207), .B2(n9205), .A(n9206), .ZN(n9208) );
  NAND2_X1 U10459 ( .A1(n9208), .A2(n5905), .ZN(n9213) );
  NOR2_X1 U10460 ( .A1(n9209), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9838) );
  AOI21_X1 U10461 ( .B1(n9284), .B2(n9523), .A(n9838), .ZN(n9210) );
  OAI21_X1 U10462 ( .B1(n9558), .B2(n9282), .A(n9210), .ZN(n9211) );
  AOI21_X1 U10463 ( .B1(n9530), .B2(n9271), .A(n9211), .ZN(n9212) );
  OAI211_X1 U10464 ( .C1(n5004), .C2(n9235), .A(n9213), .B(n9212), .ZN(
        P1_U3226) );
  INV_X1 U10465 ( .A(n9214), .ZN(n9219) );
  AOI21_X1 U10466 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9218) );
  OAI21_X1 U10467 ( .B1(n9219), .B2(n9218), .A(n5905), .ZN(n9223) );
  AOI22_X1 U10468 ( .A1(n9456), .A2(n9272), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9220) );
  OAI21_X1 U10469 ( .B1(n9286), .B2(n9423), .A(n9220), .ZN(n9221) );
  AOI21_X1 U10470 ( .B1(n9428), .B2(n9284), .A(n9221), .ZN(n9222) );
  OAI211_X1 U10471 ( .C1(n4698), .C2(n9235), .A(n9223), .B(n9222), .ZN(
        P1_U3227) );
  NOR3_X1 U10472 ( .A1(n9226), .A2(n9225), .A3(n5685), .ZN(n9229) );
  INV_X1 U10473 ( .A(n9227), .ZN(n9228) );
  OAI21_X1 U10474 ( .B1(n9229), .B2(n9228), .A(n5905), .ZN(n9234) );
  INV_X1 U10475 ( .A(n9230), .ZN(n9476) );
  AOI22_X1 U10476 ( .A1(n9481), .A2(n9284), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9231) );
  OAI21_X1 U10477 ( .B1(n9261), .B2(n9282), .A(n9231), .ZN(n9232) );
  AOI21_X1 U10478 ( .B1(n9476), .B2(n9271), .A(n9232), .ZN(n9233) );
  OAI211_X1 U10479 ( .C1(n9478), .C2(n9235), .A(n9234), .B(n9233), .ZN(
        P1_U3231) );
  XNOR2_X1 U10480 ( .A(n9237), .B(n9236), .ZN(n9238) );
  XNOR2_X1 U10481 ( .A(n9239), .B(n9238), .ZN(n9245) );
  AOI21_X1 U10482 ( .B1(n9272), .B2(n9298), .A(n9240), .ZN(n9242) );
  NAND2_X1 U10483 ( .A1(n9271), .A2(n9607), .ZN(n9241) );
  OAI211_X1 U10484 ( .C1(n9598), .C2(n9275), .A(n9242), .B(n9241), .ZN(n9243)
         );
  AOI21_X1 U10485 ( .B1(n9709), .B2(n9288), .A(n9243), .ZN(n9244) );
  OAI21_X1 U10486 ( .B1(n9245), .B2(n9278), .A(n9244), .ZN(P1_U3232) );
  NAND2_X1 U10487 ( .A1(n9246), .A2(n9247), .ZN(n9249) );
  XNOR2_X1 U10488 ( .A(n9249), .B(n9248), .ZN(n9255) );
  AOI22_X1 U10489 ( .A1(n9481), .A2(n9272), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9251) );
  NAND2_X1 U10490 ( .A1(n9452), .A2(n9271), .ZN(n9250) );
  OAI211_X1 U10491 ( .C1(n9252), .C2(n9275), .A(n9251), .B(n9250), .ZN(n9253)
         );
  AOI21_X1 U10492 ( .B1(n9661), .B2(n9288), .A(n9253), .ZN(n9254) );
  OAI21_X1 U10493 ( .B1(n9255), .B2(n9278), .A(n9254), .ZN(P1_U3233) );
  INV_X1 U10494 ( .A(n9256), .ZN(n9258) );
  NAND2_X1 U10495 ( .A1(n9258), .A2(n9257), .ZN(n9260) );
  XNOR2_X1 U10496 ( .A(n9260), .B(n9259), .ZN(n9266) );
  NAND2_X1 U10497 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9846) );
  OAI21_X1 U10498 ( .B1(n9275), .B2(n9261), .A(n9846), .ZN(n9262) );
  AOI21_X1 U10499 ( .B1(n9272), .B2(n9543), .A(n9262), .ZN(n9263) );
  OAI21_X1 U10500 ( .B1(n9286), .B2(n9513), .A(n9263), .ZN(n9264) );
  AOI21_X1 U10501 ( .B1(n9681), .B2(n9288), .A(n9264), .ZN(n9265) );
  OAI21_X1 U10502 ( .B1(n9266), .B2(n9278), .A(n9265), .ZN(P1_U3236) );
  NAND2_X1 U10503 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  XNOR2_X1 U10504 ( .A(n9267), .B(n9270), .ZN(n9279) );
  AOI22_X1 U10505 ( .A1(n9393), .A2(n9271), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9274) );
  NAND2_X1 U10506 ( .A1(n9428), .A2(n9272), .ZN(n9273) );
  OAI211_X1 U10507 ( .C1(n9294), .C2(n9275), .A(n9274), .B(n9273), .ZN(n9276)
         );
  AOI21_X1 U10508 ( .B1(n9642), .B2(n9288), .A(n9276), .ZN(n9277) );
  OAI21_X1 U10509 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(P1_U3238) );
  XOR2_X1 U10510 ( .A(n9281), .B(n9280), .Z(n9290) );
  NAND2_X1 U10511 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9312) );
  OAI21_X1 U10512 ( .B1(n9282), .B2(n9598), .A(n9312), .ZN(n9283) );
  AOI21_X1 U10513 ( .B1(n9284), .B2(n9522), .A(n9283), .ZN(n9285) );
  OAI21_X1 U10514 ( .B1(n9286), .B2(n9567), .A(n9285), .ZN(n9287) );
  AOI21_X1 U10515 ( .B1(n9569), .B2(n9288), .A(n9287), .ZN(n9289) );
  OAI21_X1 U10516 ( .B1(n9290), .B2(n9278), .A(n9289), .ZN(P1_U3239) );
  MUX2_X1 U10517 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9350), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10518 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9291), .S(P1_U4006), .Z(
        P1_U3585) );
  INV_X1 U10519 ( .A(n9292), .ZN(n9365) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9365), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10521 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9293), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10522 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9398), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10523 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9415), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9428), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9444), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9456), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9465), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9481), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10529 ( .A(n9496), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9295), .Z(
        P1_U3575) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9508), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9523), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9543), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10533 ( .A(n9522), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9295), .Z(
        P1_U3571) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9541), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9296), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9297), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9298), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9299), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9300), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9301), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9302), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9303), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9304), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9305), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9307), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9308), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7362), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9309), .S(P1_U4006), .Z(
        P1_U3556) );
  XOR2_X1 U10549 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9334), .Z(n9322) );
  INV_X1 U10550 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U10551 ( .A1(n9853), .A2(n9333), .ZN(n9313) );
  OAI211_X1 U10552 ( .C1(n9862), .C2(n9314), .A(n9313), .B(n9312), .ZN(n9321)
         );
  INV_X1 U10553 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9319) );
  OAI21_X1 U10554 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9325) );
  XNOR2_X1 U10555 ( .A(n9325), .B(n9333), .ZN(n9318) );
  NOR2_X1 U10556 ( .A1(n9318), .A2(n9319), .ZN(n9324) );
  AOI211_X1 U10557 ( .C1(n9319), .C2(n9318), .A(n9847), .B(n9324), .ZN(n9320)
         );
  AOI211_X1 U10558 ( .C1(n9841), .C2(n9322), .A(n9321), .B(n9320), .ZN(n9323)
         );
  INV_X1 U10559 ( .A(n9323), .ZN(P1_U3256) );
  NAND2_X1 U10560 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9828), .ZN(n9326) );
  OAI21_X1 U10561 ( .B1(n9828), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9326), .ZN(
        n9824) );
  NAND2_X1 U10562 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9839), .ZN(n9327) );
  OAI21_X1 U10563 ( .B1(n9839), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9327), .ZN(
        n9835) );
  INV_X1 U10564 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9328) );
  MUX2_X1 U10565 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9328), .S(n9854), .Z(n9329) );
  INV_X1 U10566 ( .A(n9329), .ZN(n9850) );
  XNOR2_X1 U10567 ( .A(n9854), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9857) );
  INV_X1 U10568 ( .A(n9839), .ZN(n9338) );
  XOR2_X1 U10569 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9839), .Z(n9842) );
  INV_X1 U10570 ( .A(n9331), .ZN(n9332) );
  AOI22_X1 U10571 ( .A1(n9334), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9333), .B2(
        n9332), .ZN(n9829) );
  XNOR2_X1 U10572 ( .A(n9828), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9830) );
  INV_X1 U10573 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9335) );
  OAI22_X1 U10574 ( .A1(n9829), .A2(n9830), .B1(n9336), .B2(n9335), .ZN(n9843)
         );
  NAND2_X1 U10575 ( .A1(n9842), .A2(n9843), .ZN(n9840) );
  OAI21_X1 U10576 ( .B1(n9338), .B2(n9337), .A(n9840), .ZN(n9856) );
  OAI22_X1 U10577 ( .A1(n9344), .A2(n9847), .B1(n9343), .B2(n9858), .ZN(n9345)
         );
  OAI21_X1 U10578 ( .B1(n9862), .B2(n9347), .A(n9346), .ZN(n9348) );
  NAND2_X1 U10579 ( .A1(n9355), .A2(n9623), .ZN(n9349) );
  XNOR2_X1 U10580 ( .A(n9349), .B(n9619), .ZN(n9617) );
  NAND2_X1 U10581 ( .A1(n9617), .A2(n9614), .ZN(n9353) );
  NAND2_X1 U10582 ( .A1(n9351), .A2(n9350), .ZN(n9621) );
  NOR2_X1 U10583 ( .A1(n10210), .A2(n9621), .ZN(n9356) );
  AOI21_X1 U10584 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(n9616), .A(n9356), .ZN(
        n9352) );
  OAI211_X1 U10585 ( .C1(n9619), .C2(n9609), .A(n9353), .B(n9352), .ZN(
        P1_U3261) );
  XNOR2_X1 U10586 ( .A(n9355), .B(n9354), .ZN(n9620) );
  NAND2_X1 U10587 ( .A1(n9620), .A2(n9614), .ZN(n9358) );
  AOI21_X1 U10588 ( .B1(n9616), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9356), .ZN(
        n9357) );
  OAI211_X1 U10589 ( .C1(n9623), .C2(n9609), .A(n9358), .B(n9357), .ZN(
        P1_U3262) );
  OAI21_X1 U10590 ( .B1(n9360), .B2(n9363), .A(n9359), .ZN(n9632) );
  AOI21_X1 U10591 ( .B1(n9628), .B2(n9380), .A(n4287), .ZN(n9629) );
  AOI22_X1 U10592 ( .A1(n9361), .A2(n10213), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n9616), .ZN(n9362) );
  OAI21_X1 U10593 ( .B1(n4998), .B2(n9609), .A(n9362), .ZN(n9370) );
  XNOR2_X1 U10594 ( .A(n9364), .B(n9363), .ZN(n9369) );
  XNOR2_X1 U10595 ( .A(n9372), .B(n9371), .ZN(n9633) );
  INV_X1 U10596 ( .A(n9633), .ZN(n9389) );
  XNOR2_X1 U10597 ( .A(n9373), .B(n4680), .ZN(n9374) );
  NAND2_X1 U10598 ( .A1(n9374), .A2(n9603), .ZN(n9379) );
  OAI22_X1 U10599 ( .A1(n9376), .A2(n9927), .B1(n9375), .B2(n9925), .ZN(n9377)
         );
  INV_X1 U10600 ( .A(n9377), .ZN(n9378) );
  NAND2_X1 U10601 ( .A1(n9379), .A2(n9378), .ZN(n9638) );
  OAI211_X1 U10602 ( .C1(n9391), .C2(n9385), .A(n4997), .B(n9380), .ZN(n9636)
         );
  INV_X1 U10603 ( .A(n9485), .ZN(n9381) );
  NOR2_X1 U10604 ( .A1(n9636), .A2(n9381), .ZN(n9387) );
  INV_X1 U10605 ( .A(n9382), .ZN(n9383) );
  AOI22_X1 U10606 ( .A1(n9383), .A2(n10213), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9616), .ZN(n9384) );
  OAI21_X1 U10607 ( .B1(n9385), .B2(n9609), .A(n9384), .ZN(n9386) );
  AOI211_X1 U10608 ( .C1(n9638), .C2(n10221), .A(n9387), .B(n9386), .ZN(n9388)
         );
  OAI21_X1 U10609 ( .B1(n9389), .B2(n9595), .A(n9388), .ZN(P1_U3264) );
  XOR2_X1 U10610 ( .A(n9397), .B(n9390), .Z(n9645) );
  INV_X1 U10611 ( .A(n9409), .ZN(n9392) );
  AOI211_X1 U10612 ( .C1(n9642), .C2(n9392), .A(n9949), .B(n9391), .ZN(n9641)
         );
  AOI22_X1 U10613 ( .A1(n9393), .A2(n10213), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9616), .ZN(n9394) );
  OAI21_X1 U10614 ( .B1(n9395), .B2(n9609), .A(n9394), .ZN(n9404) );
  XOR2_X1 U10615 ( .A(n9397), .B(n9396), .Z(n9402) );
  NAND2_X1 U10616 ( .A1(n9428), .A2(n9540), .ZN(n9399) );
  AOI211_X1 U10617 ( .C1(n9641), .C2(n9485), .A(n9404), .B(n9403), .ZN(n9405)
         );
  OAI21_X1 U10618 ( .B1(n9595), .B2(n9645), .A(n9405), .ZN(P1_U3265) );
  OAI21_X1 U10619 ( .B1(n9407), .B2(n9414), .A(n9406), .ZN(n9408) );
  INV_X1 U10620 ( .A(n9408), .ZN(n9650) );
  AOI21_X1 U10621 ( .B1(n9646), .B2(n9421), .A(n9409), .ZN(n9647) );
  AOI22_X1 U10622 ( .A1(n9410), .A2(n10213), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9616), .ZN(n9411) );
  OAI21_X1 U10623 ( .B1(n9412), .B2(n9609), .A(n9411), .ZN(n9418) );
  XOR2_X1 U10624 ( .A(n9414), .B(n9413), .Z(n9416) );
  AOI222_X1 U10625 ( .A1(n9603), .A2(n9416), .B1(n9415), .B2(n9542), .C1(n9444), .C2(n9540), .ZN(n9649) );
  NOR2_X1 U10626 ( .A1(n9649), .A2(n10210), .ZN(n9417) );
  AOI211_X1 U10627 ( .C1(n9647), .C2(n9614), .A(n9418), .B(n9417), .ZN(n9419)
         );
  OAI21_X1 U10628 ( .B1(n9650), .B2(n9595), .A(n9419), .ZN(P1_U3266) );
  XNOR2_X1 U10629 ( .A(n9420), .B(n9427), .ZN(n9655) );
  INV_X1 U10630 ( .A(n9421), .ZN(n9422) );
  AOI211_X1 U10631 ( .C1(n9652), .C2(n9434), .A(n9949), .B(n9422), .ZN(n9651)
         );
  INV_X1 U10632 ( .A(n9423), .ZN(n9424) );
  AOI22_X1 U10633 ( .A1(n9424), .A2(n10213), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9616), .ZN(n9425) );
  OAI21_X1 U10634 ( .B1(n4698), .B2(n9609), .A(n9425), .ZN(n9431) );
  XNOR2_X1 U10635 ( .A(n9426), .B(n9427), .ZN(n9429) );
  AOI222_X1 U10636 ( .A1(n9603), .A2(n9429), .B1(n9428), .B2(n9542), .C1(n9456), .C2(n9540), .ZN(n9654) );
  NOR2_X1 U10637 ( .A1(n9654), .A2(n10210), .ZN(n9430) );
  AOI211_X1 U10638 ( .C1(n9651), .C2(n9485), .A(n9431), .B(n9430), .ZN(n9432)
         );
  OAI21_X1 U10639 ( .B1(n9595), .B2(n9655), .A(n9432), .ZN(P1_U3267) );
  XNOR2_X1 U10640 ( .A(n9433), .B(n9442), .ZN(n9660) );
  INV_X1 U10641 ( .A(n9450), .ZN(n9435) );
  AOI21_X1 U10642 ( .B1(n9656), .B2(n9435), .A(n5011), .ZN(n9657) );
  INV_X1 U10643 ( .A(n9436), .ZN(n9437) );
  AOI22_X1 U10644 ( .A1(n9437), .A2(n10213), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9616), .ZN(n9438) );
  OAI21_X1 U10645 ( .B1(n9439), .B2(n9609), .A(n9438), .ZN(n9447) );
  NAND2_X1 U10646 ( .A1(n9441), .A2(n9440), .ZN(n9443) );
  XNOR2_X1 U10647 ( .A(n9443), .B(n9442), .ZN(n9445) );
  AOI222_X1 U10648 ( .A1(n9603), .A2(n9445), .B1(n9444), .B2(n9542), .C1(n9465), .C2(n9540), .ZN(n9659) );
  NOR2_X1 U10649 ( .A1(n9659), .A2(n10210), .ZN(n9446) );
  AOI211_X1 U10650 ( .C1(n9657), .C2(n9614), .A(n9447), .B(n9446), .ZN(n9448)
         );
  OAI21_X1 U10651 ( .B1(n9595), .B2(n9660), .A(n9448), .ZN(P1_U3268) );
  XNOR2_X1 U10652 ( .A(n9449), .B(n9455), .ZN(n9665) );
  INV_X1 U10653 ( .A(n9467), .ZN(n9451) );
  AOI21_X1 U10654 ( .B1(n9661), .B2(n9451), .A(n9450), .ZN(n9662) );
  AOI22_X1 U10655 ( .A1(n9452), .A2(n10213), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n9616), .ZN(n9453) );
  OAI21_X1 U10656 ( .B1(n9454), .B2(n9609), .A(n9453), .ZN(n9459) );
  AOI222_X1 U10657 ( .A1(n9603), .A2(n9457), .B1(n9456), .B2(n9542), .C1(n9481), .C2(n9540), .ZN(n9664) );
  NOR2_X1 U10658 ( .A1(n9664), .A2(n10210), .ZN(n9458) );
  AOI211_X1 U10659 ( .C1(n9662), .C2(n9614), .A(n9459), .B(n9458), .ZN(n9460)
         );
  OAI21_X1 U10660 ( .B1(n9595), .B2(n9665), .A(n9460), .ZN(P1_U3269) );
  XNOR2_X1 U10661 ( .A(n9462), .B(n9461), .ZN(n9670) );
  XNOR2_X1 U10662 ( .A(n9463), .B(n9464), .ZN(n9466) );
  AOI222_X1 U10663 ( .A1(n9603), .A2(n9466), .B1(n9496), .B2(n9540), .C1(n9465), .C2(n9542), .ZN(n9669) );
  AOI211_X1 U10664 ( .C1(n9667), .C2(n9475), .A(n9949), .B(n9467), .ZN(n9666)
         );
  NAND2_X1 U10665 ( .A1(n9666), .A2(n9468), .ZN(n9469) );
  OAI211_X1 U10666 ( .C1(n9566), .C2(n9470), .A(n9669), .B(n9469), .ZN(n9471)
         );
  NAND2_X1 U10667 ( .A1(n9471), .A2(n10221), .ZN(n9473) );
  AOI22_X1 U10668 ( .A1(n9667), .A2(n9588), .B1(n9616), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9472) );
  OAI211_X1 U10669 ( .C1(n9670), .C2(n9595), .A(n9473), .B(n9472), .ZN(
        P1_U3270) );
  XNOR2_X1 U10670 ( .A(n9474), .B(n9480), .ZN(n9675) );
  AOI211_X1 U10671 ( .C1(n9672), .C2(n9488), .A(n9949), .B(n5010), .ZN(n9671)
         );
  AOI22_X1 U10672 ( .A1(n9476), .A2(n10213), .B1(n9616), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9477) );
  OAI21_X1 U10673 ( .B1(n9478), .B2(n9609), .A(n9477), .ZN(n9484) );
  XNOR2_X1 U10674 ( .A(n9479), .B(n9480), .ZN(n9482) );
  AOI222_X1 U10675 ( .A1(n9603), .A2(n9482), .B1(n9481), .B2(n9542), .C1(n9508), .C2(n9540), .ZN(n9674) );
  NOR2_X1 U10676 ( .A1(n9674), .A2(n10210), .ZN(n9483) );
  AOI211_X1 U10677 ( .C1(n9671), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9486)
         );
  OAI21_X1 U10678 ( .B1(n9675), .B2(n9595), .A(n9486), .ZN(P1_U3271) );
  XOR2_X1 U10679 ( .A(n9494), .B(n9487), .Z(n9680) );
  INV_X1 U10680 ( .A(n9510), .ZN(n9490) );
  INV_X1 U10681 ( .A(n9488), .ZN(n9489) );
  AOI21_X1 U10682 ( .B1(n9676), .B2(n9490), .A(n9489), .ZN(n9677) );
  AOI22_X1 U10683 ( .A1(n9616), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9491), .B2(
        n10213), .ZN(n9492) );
  OAI21_X1 U10684 ( .B1(n9493), .B2(n9609), .A(n9492), .ZN(n9499) );
  XNOR2_X1 U10685 ( .A(n9495), .B(n9494), .ZN(n9497) );
  AOI222_X1 U10686 ( .A1(n9603), .A2(n9497), .B1(n9496), .B2(n9542), .C1(n9523), .C2(n9540), .ZN(n9679) );
  NOR2_X1 U10687 ( .A1(n9679), .A2(n9616), .ZN(n9498) );
  AOI211_X1 U10688 ( .C1(n9677), .C2(n9614), .A(n9499), .B(n9498), .ZN(n9500)
         );
  OAI21_X1 U10689 ( .B1(n9595), .B2(n9680), .A(n9500), .ZN(P1_U3272) );
  NAND2_X1 U10690 ( .A1(n9502), .A2(n9501), .ZN(n9539) );
  NAND2_X1 U10691 ( .A1(n9539), .A2(n9503), .ZN(n9521) );
  INV_X1 U10692 ( .A(n9504), .ZN(n9506) );
  OAI21_X1 U10693 ( .B1(n9521), .B2(n9506), .A(n9505), .ZN(n9507) );
  XOR2_X1 U10694 ( .A(n9507), .B(n9517), .Z(n9509) );
  AOI222_X1 U10695 ( .A1(n9603), .A2(n9509), .B1(n9508), .B2(n9542), .C1(n9543), .C2(n9540), .ZN(n9686) );
  INV_X1 U10696 ( .A(n9529), .ZN(n9511) );
  AOI21_X1 U10697 ( .B1(n9681), .B2(n9511), .A(n9510), .ZN(n9682) );
  NOR2_X1 U10698 ( .A1(n9512), .A2(n9609), .ZN(n9515) );
  OAI22_X1 U10699 ( .A1(n10221), .A2(n9328), .B1(n9513), .B2(n9566), .ZN(n9514) );
  AOI211_X1 U10700 ( .C1(n9682), .C2(n9614), .A(n9515), .B(n9514), .ZN(n9520)
         );
  NAND2_X1 U10701 ( .A1(n9518), .A2(n9517), .ZN(n9683) );
  NAND3_X1 U10702 ( .A1(n9516), .A2(n9683), .A3(n9573), .ZN(n9519) );
  OAI211_X1 U10703 ( .C1(n9686), .C2(n9616), .A(n9520), .B(n9519), .ZN(
        P1_U3273) );
  XNOR2_X1 U10704 ( .A(n9521), .B(n9525), .ZN(n9524) );
  AOI222_X1 U10705 ( .A1(n9603), .A2(n9524), .B1(n9523), .B2(n9542), .C1(n9522), .C2(n9540), .ZN(n9690) );
  INV_X1 U10706 ( .A(n9525), .ZN(n9526) );
  XNOR2_X1 U10707 ( .A(n9527), .B(n9526), .ZN(n9691) );
  INV_X1 U10708 ( .A(n9691), .ZN(n9534) );
  AND2_X1 U10709 ( .A1(n9545), .A2(n9687), .ZN(n9528) );
  NOR2_X1 U10710 ( .A1(n9529), .A2(n9528), .ZN(n9688) );
  NAND2_X1 U10711 ( .A1(n9688), .A2(n9614), .ZN(n9532) );
  AOI22_X1 U10712 ( .A1(n10210), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9530), 
        .B2(n10213), .ZN(n9531) );
  OAI211_X1 U10713 ( .C1(n5004), .C2(n9609), .A(n9532), .B(n9531), .ZN(n9533)
         );
  AOI21_X1 U10714 ( .B1(n9534), .B2(n9573), .A(n9533), .ZN(n9535) );
  OAI21_X1 U10715 ( .B1(n9690), .B2(n9616), .A(n9535), .ZN(P1_U3274) );
  NAND3_X1 U10716 ( .A1(n9537), .A2(n9550), .A3(n9536), .ZN(n9538) );
  NAND2_X1 U10717 ( .A1(n9539), .A2(n9538), .ZN(n9544) );
  AOI222_X1 U10718 ( .A1(n9603), .A2(n9544), .B1(n9543), .B2(n9542), .C1(n9541), .C2(n9540), .ZN(n9695) );
  INV_X1 U10719 ( .A(n9545), .ZN(n9546) );
  AOI211_X1 U10720 ( .C1(n9693), .C2(n9565), .A(n9949), .B(n9546), .ZN(n9692)
         );
  INV_X1 U10721 ( .A(n9547), .ZN(n9548) );
  AOI22_X1 U10722 ( .A1(n9616), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9548), .B2(
        n10213), .ZN(n9549) );
  OAI21_X1 U10723 ( .B1(n5007), .B2(n9609), .A(n9549), .ZN(n9553) );
  XNOR2_X1 U10724 ( .A(n9551), .B(n9550), .ZN(n9696) );
  NOR2_X1 U10725 ( .A1(n9696), .A2(n9595), .ZN(n9552) );
  AOI211_X1 U10726 ( .C1(n9692), .C2(n9554), .A(n9553), .B(n9552), .ZN(n9555)
         );
  OAI21_X1 U10727 ( .B1(n9695), .B2(n10210), .A(n9555), .ZN(P1_U3275) );
  XNOR2_X1 U10728 ( .A(n9556), .B(n9562), .ZN(n9557) );
  NAND2_X1 U10729 ( .A1(n9557), .A2(n9603), .ZN(n9561) );
  OAI22_X1 U10730 ( .A1(n9558), .A2(n9927), .B1(n9598), .B2(n9925), .ZN(n9559)
         );
  INV_X1 U10731 ( .A(n9559), .ZN(n9560) );
  NAND2_X1 U10732 ( .A1(n9561), .A2(n9560), .ZN(n9701) );
  INV_X1 U10733 ( .A(n9701), .ZN(n9575) );
  XNOR2_X1 U10734 ( .A(n9563), .B(n9562), .ZN(n9697) );
  OR2_X1 U10735 ( .A1(n9586), .A2(n9698), .ZN(n9564) );
  NAND2_X1 U10736 ( .A1(n9565), .A2(n9564), .ZN(n9699) );
  OAI22_X1 U10737 ( .A1(n10221), .A2(n9319), .B1(n9567), .B2(n9566), .ZN(n9568) );
  AOI21_X1 U10738 ( .B1(n9569), .B2(n9588), .A(n9568), .ZN(n9570) );
  OAI21_X1 U10739 ( .B1(n9699), .B2(n9571), .A(n9570), .ZN(n9572) );
  AOI21_X1 U10740 ( .B1(n9697), .B2(n9573), .A(n9572), .ZN(n9574) );
  OAI21_X1 U10741 ( .B1(n9575), .B2(n9616), .A(n9574), .ZN(P1_U3276) );
  XNOR2_X1 U10742 ( .A(n9576), .B(n9577), .ZN(n9708) );
  AOI21_X1 U10743 ( .B1(n9578), .B2(n9577), .A(n9923), .ZN(n9583) );
  OAI22_X1 U10744 ( .A1(n9580), .A2(n9927), .B1(n9579), .B2(n9925), .ZN(n9581)
         );
  AOI21_X1 U10745 ( .B1(n9583), .B2(n9582), .A(n9581), .ZN(n9707) );
  INV_X1 U10746 ( .A(n9707), .ZN(n9593) );
  OAI21_X1 U10747 ( .B1(n9605), .B2(n9584), .A(n4997), .ZN(n9585) );
  OR2_X1 U10748 ( .A1(n9586), .A2(n9585), .ZN(n9703) );
  AOI22_X1 U10749 ( .A1(n9616), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9587), .B2(
        n10213), .ZN(n9590) );
  NAND2_X1 U10750 ( .A1(n9705), .A2(n9588), .ZN(n9589) );
  OAI211_X1 U10751 ( .C1(n9703), .C2(n9591), .A(n9590), .B(n9589), .ZN(n9592)
         );
  AOI21_X1 U10752 ( .B1(n9593), .B2(n10221), .A(n9592), .ZN(n9594) );
  OAI21_X1 U10753 ( .B1(n9708), .B2(n9595), .A(n9594), .ZN(P1_U3277) );
  XNOR2_X1 U10754 ( .A(n9596), .B(n9599), .ZN(n9604) );
  OAI22_X1 U10755 ( .A1(n9598), .A2(n9927), .B1(n9597), .B2(n9925), .ZN(n9602)
         );
  XOR2_X1 U10756 ( .A(n9600), .B(n9599), .Z(n9713) );
  NOR2_X1 U10757 ( .A1(n9713), .A2(n9897), .ZN(n9601) );
  AOI211_X1 U10758 ( .C1(n9604), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9712)
         );
  AOI21_X1 U10759 ( .B1(n9709), .B2(n9606), .A(n9605), .ZN(n9710) );
  AOI22_X1 U10760 ( .A1(n9616), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9607), .B2(
        n10213), .ZN(n9608) );
  OAI21_X1 U10761 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(n9613) );
  NOR2_X1 U10762 ( .A1(n9713), .A2(n9611), .ZN(n9612) );
  AOI211_X1 U10763 ( .C1(n9710), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9615)
         );
  OAI21_X1 U10764 ( .B1(n9712), .B2(n9616), .A(n9615), .ZN(P1_U3278) );
  NAND2_X1 U10765 ( .A1(n9617), .A2(n4997), .ZN(n9618) );
  OAI211_X1 U10766 ( .C1(n9619), .C2(n9947), .A(n9618), .B(n9621), .ZN(n9726)
         );
  MUX2_X1 U10767 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9726), .S(n9972), .Z(
        P1_U3554) );
  NAND2_X1 U10768 ( .A1(n9620), .A2(n4997), .ZN(n9622) );
  OAI211_X1 U10769 ( .C1(n9623), .C2(n9947), .A(n9622), .B(n9621), .ZN(n9727)
         );
  MUX2_X1 U10770 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9727), .S(n9972), .Z(
        P1_U3553) );
  AOI21_X1 U10771 ( .B1(n9893), .B2(n9625), .A(n9624), .ZN(n9626) );
  AOI22_X1 U10772 ( .A1(n9629), .A2(n4997), .B1(n9893), .B2(n9628), .ZN(n9630)
         );
  OAI211_X1 U10773 ( .C1(n9632), .C2(n9719), .A(n9631), .B(n9630), .ZN(n9728)
         );
  MUX2_X1 U10774 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9728), .S(n9972), .Z(
        P1_U3551) );
  NAND2_X1 U10775 ( .A1(n9633), .A2(n9952), .ZN(n9640) );
  NAND2_X1 U10776 ( .A1(n9634), .A2(n9893), .ZN(n9635) );
  NAND2_X1 U10777 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NOR2_X1 U10778 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NAND2_X1 U10779 ( .A1(n9640), .A2(n9639), .ZN(n9729) );
  MUX2_X1 U10780 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9729), .S(n9972), .Z(
        P1_U3550) );
  AOI21_X1 U10781 ( .B1(n9893), .B2(n9642), .A(n9641), .ZN(n9643) );
  OAI211_X1 U10782 ( .C1(n9645), .C2(n9719), .A(n9644), .B(n9643), .ZN(n9730)
         );
  MUX2_X1 U10783 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9730), .S(n9972), .Z(
        P1_U3549) );
  AOI22_X1 U10784 ( .A1(n9647), .A2(n4997), .B1(n9893), .B2(n9646), .ZN(n9648)
         );
  OAI211_X1 U10785 ( .C1(n9650), .C2(n9719), .A(n9649), .B(n9648), .ZN(n9731)
         );
  MUX2_X1 U10786 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9731), .S(n9972), .Z(
        P1_U3548) );
  AOI21_X1 U10787 ( .B1(n9893), .B2(n9652), .A(n9651), .ZN(n9653) );
  OAI211_X1 U10788 ( .C1(n9655), .C2(n9719), .A(n9654), .B(n9653), .ZN(n9732)
         );
  MUX2_X1 U10789 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9732), .S(n9972), .Z(
        P1_U3547) );
  AOI22_X1 U10790 ( .A1(n9657), .A2(n4997), .B1(n9893), .B2(n9656), .ZN(n9658)
         );
  OAI211_X1 U10791 ( .C1(n9660), .C2(n9719), .A(n9659), .B(n9658), .ZN(n9733)
         );
  MUX2_X1 U10792 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9733), .S(n9972), .Z(
        P1_U3546) );
  AOI22_X1 U10793 ( .A1(n9662), .A2(n4997), .B1(n9893), .B2(n9661), .ZN(n9663)
         );
  OAI211_X1 U10794 ( .C1(n9719), .C2(n9665), .A(n9664), .B(n9663), .ZN(n9734)
         );
  MUX2_X1 U10795 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9734), .S(n9972), .Z(
        P1_U3545) );
  AOI21_X1 U10796 ( .B1(n9893), .B2(n9667), .A(n9666), .ZN(n9668) );
  OAI211_X1 U10797 ( .C1(n9670), .C2(n9719), .A(n9669), .B(n9668), .ZN(n9735)
         );
  MUX2_X1 U10798 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9735), .S(n9972), .Z(
        P1_U3544) );
  AOI21_X1 U10799 ( .B1(n9893), .B2(n9672), .A(n9671), .ZN(n9673) );
  OAI211_X1 U10800 ( .C1(n9675), .C2(n9719), .A(n9674), .B(n9673), .ZN(n9736)
         );
  MUX2_X1 U10801 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9736), .S(n9972), .Z(
        P1_U3543) );
  AOI22_X1 U10802 ( .A1(n9677), .A2(n4997), .B1(n9893), .B2(n9676), .ZN(n9678)
         );
  OAI211_X1 U10803 ( .C1(n9680), .C2(n9719), .A(n9679), .B(n9678), .ZN(n9737)
         );
  MUX2_X1 U10804 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9737), .S(n9972), .Z(
        P1_U3542) );
  AOI22_X1 U10805 ( .A1(n9682), .A2(n4997), .B1(n9893), .B2(n9681), .ZN(n9685)
         );
  NAND3_X1 U10806 ( .A1(n9516), .A2(n9683), .A3(n9952), .ZN(n9684) );
  NAND3_X1 U10807 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n9738) );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9738), .S(n9972), .Z(
        P1_U3541) );
  AOI22_X1 U10809 ( .A1(n9688), .A2(n4997), .B1(n9893), .B2(n9687), .ZN(n9689)
         );
  OAI211_X1 U10810 ( .C1(n9719), .C2(n9691), .A(n9690), .B(n9689), .ZN(n9739)
         );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9739), .S(n9972), .Z(
        P1_U3540) );
  AOI21_X1 U10812 ( .B1(n9893), .B2(n9693), .A(n9692), .ZN(n9694) );
  OAI211_X1 U10813 ( .C1(n9719), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9740)
         );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9740), .S(n9972), .Z(
        P1_U3539) );
  AND2_X1 U10815 ( .A1(n9697), .A2(n9952), .ZN(n9702) );
  OAI22_X1 U10816 ( .A1(n9699), .A2(n9949), .B1(n9698), .B2(n9947), .ZN(n9700)
         );
  MUX2_X1 U10817 ( .A(n9741), .B(P1_REG1_REG_15__SCAN_IN), .S(n9969), .Z(
        P1_U3538) );
  INV_X1 U10818 ( .A(n9703), .ZN(n9704) );
  AOI21_X1 U10819 ( .B1(n9893), .B2(n9705), .A(n9704), .ZN(n9706) );
  OAI211_X1 U10820 ( .C1(n9719), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9742)
         );
  MUX2_X1 U10821 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9742), .S(n9972), .Z(
        P1_U3537) );
  AOI22_X1 U10822 ( .A1(n9710), .A2(n4997), .B1(n9893), .B2(n9709), .ZN(n9711)
         );
  OAI211_X1 U10823 ( .C1(n9896), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9743)
         );
  MUX2_X1 U10824 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9743), .S(n9972), .Z(
        P1_U3536) );
  AOI21_X1 U10825 ( .B1(n9893), .B2(n9715), .A(n9714), .ZN(n9716) );
  OAI211_X1 U10826 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9744)
         );
  MUX2_X1 U10827 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9744), .S(n9972), .Z(
        P1_U3533) );
  AOI22_X1 U10828 ( .A1(n9721), .A2(n4997), .B1(n9893), .B2(n9720), .ZN(n9722)
         );
  OAI211_X1 U10829 ( .C1(n9896), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9745)
         );
  MUX2_X1 U10830 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9745), .S(n9972), .Z(
        P1_U3532) );
  MUX2_X1 U10831 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9725), .S(n9972), .Z(
        P1_U3523) );
  MUX2_X1 U10832 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9726), .S(n9958), .Z(
        P1_U3522) );
  MUX2_X1 U10833 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9727), .S(n9958), .Z(
        P1_U3521) );
  MUX2_X1 U10834 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9728), .S(n9958), .Z(
        P1_U3519) );
  MUX2_X1 U10835 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9729), .S(n9958), .Z(
        P1_U3518) );
  MUX2_X1 U10836 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9730), .S(n9958), .Z(
        P1_U3517) );
  MUX2_X1 U10837 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9731), .S(n9958), .Z(
        P1_U3516) );
  MUX2_X1 U10838 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9732), .S(n9958), .Z(
        P1_U3515) );
  MUX2_X1 U10839 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9733), .S(n9958), .Z(
        P1_U3514) );
  MUX2_X1 U10840 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9734), .S(n9958), .Z(
        P1_U3513) );
  MUX2_X1 U10841 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9735), .S(n9958), .Z(
        P1_U3512) );
  MUX2_X1 U10842 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9736), .S(n9958), .Z(
        P1_U3511) );
  MUX2_X1 U10843 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9737), .S(n9958), .Z(
        P1_U3510) );
  MUX2_X1 U10844 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9738), .S(n9958), .Z(
        P1_U3508) );
  MUX2_X1 U10845 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9739), .S(n9958), .Z(
        P1_U3505) );
  MUX2_X1 U10846 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9740), .S(n9958), .Z(
        P1_U3502) );
  MUX2_X1 U10847 ( .A(n9741), .B(P1_REG0_REG_15__SCAN_IN), .S(n9956), .Z(
        P1_U3499) );
  MUX2_X1 U10848 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9742), .S(n9958), .Z(
        P1_U3496) );
  MUX2_X1 U10849 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9743), .S(n9958), .Z(
        P1_U3493) );
  MUX2_X1 U10850 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9744), .S(n9958), .Z(
        P1_U3484) );
  MUX2_X1 U10851 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n9745), .S(n9958), .Z(
        P1_U3481) );
  NOR4_X1 U10852 ( .A1(n9746), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4609), .A4(
        P1_U3084), .ZN(n9747) );
  AOI21_X1 U10853 ( .B1(n9748), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9747), .ZN(
        n9749) );
  OAI21_X1 U10854 ( .B1(n9750), .B2(n9752), .A(n9749), .ZN(P1_U3322) );
  OAI222_X1 U10855 ( .A1(n9755), .A2(n9754), .B1(P1_U3084), .B2(n9753), .C1(
        n9752), .C2(n9751), .ZN(P1_U3324) );
  MUX2_X1 U10856 ( .A(n9756), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10857 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U10858 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9757) );
  AOI21_X1 U10859 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9757), .ZN(n10041) );
  NOR2_X1 U10860 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9758) );
  AOI21_X1 U10861 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9758), .ZN(n10044) );
  NOR2_X1 U10862 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9759) );
  AOI21_X1 U10863 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9759), .ZN(n10047) );
  NOR2_X1 U10864 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9760) );
  AOI21_X1 U10865 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9760), .ZN(n10050) );
  NOR2_X1 U10866 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9761) );
  AOI21_X1 U10867 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9761), .ZN(n10053) );
  NOR2_X1 U10868 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9767) );
  XNOR2_X1 U10869 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10244) );
  NAND2_X1 U10870 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9765) );
  XOR2_X1 U10871 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10242) );
  NAND2_X1 U10872 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9763) );
  AOI21_X1 U10873 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10035) );
  NAND3_X1 U10874 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U10875 ( .A1(n9765), .A2(n9764), .ZN(n10243) );
  NOR2_X1 U10876 ( .A1(n10244), .A2(n10243), .ZN(n9766) );
  NOR2_X1 U10877 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  NOR2_X1 U10878 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9768), .ZN(n10227) );
  NAND2_X1 U10879 ( .A1(n9769), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U10880 ( .A1(n10226), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U10881 ( .A1(n9771), .A2(n9770), .ZN(n9772) );
  NAND2_X1 U10882 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9772), .ZN(n9773) );
  NAND2_X1 U10883 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9774), .ZN(n9776) );
  NAND2_X1 U10884 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10237), .ZN(n9775) );
  AND2_X1 U10885 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9777), .ZN(n9778) );
  NAND2_X1 U10886 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9779) );
  OAI21_X1 U10887 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9779), .ZN(n10061) );
  NOR2_X1 U10888 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  AOI21_X1 U10889 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10060), .ZN(n10059) );
  NAND2_X1 U10890 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9780) );
  OAI21_X1 U10891 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9780), .ZN(n10058) );
  NOR2_X1 U10892 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  NOR2_X1 U10893 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9781) );
  AOI21_X1 U10894 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9781), .ZN(n10055) );
  NAND2_X1 U10895 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  NAND2_X1 U10896 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  NAND2_X1 U10897 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  OAI21_X1 U10898 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10042), .ZN(n10040) );
  XOR2_X1 U10899 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9782) );
  XNOR2_X1 U10900 ( .A(n9783), .B(n9782), .ZN(ADD_1071_U4) );
  XNOR2_X1 U10901 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10902 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10903 ( .B1(n4239), .B2(n4621), .A(n9784), .ZN(n9786) );
  XNOR2_X1 U10904 ( .A(n9786), .B(n9785), .ZN(n9787) );
  AOI22_X1 U10905 ( .A1(n9789), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9788), .B2(
        n9787), .ZN(n9790) );
  OAI21_X1 U10906 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9791), .A(n9790), .ZN(
        P1_U3241) );
  INV_X1 U10907 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9792) );
  OR2_X1 U10908 ( .A1(n9862), .A2(n9792), .ZN(n9801) );
  NAND2_X1 U10909 ( .A1(n9853), .A2(n9793), .ZN(n9800) );
  NAND2_X1 U10910 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U10911 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9794) );
  NAND2_X1 U10912 ( .A1(n9795), .A2(n9794), .ZN(n9796) );
  NAND3_X1 U10913 ( .A1(n9841), .A2(n9797), .A3(n9796), .ZN(n9798) );
  AND4_X1 U10914 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n9798), .ZN(n9806)
         );
  OAI211_X1 U10915 ( .C1(n9804), .C2(n6765), .A(n9817), .B(n9803), .ZN(n9805)
         );
  NAND2_X1 U10916 ( .A1(n9806), .A2(n9805), .ZN(P1_U3242) );
  INV_X1 U10917 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9813) );
  OAI211_X1 U10918 ( .C1(n9809), .C2(n9808), .A(n9841), .B(n9807), .ZN(n9812)
         );
  NAND2_X1 U10919 ( .A1(n9853), .A2(n9810), .ZN(n9811) );
  OAI211_X1 U10920 ( .C1(n9813), .C2(n9862), .A(n9812), .B(n9811), .ZN(n9814)
         );
  NOR2_X1 U10921 ( .A1(n9815), .A2(n9814), .ZN(n9821) );
  OAI211_X1 U10922 ( .C1(n9819), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9820)
         );
  OAI211_X1 U10923 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9822), .A(n9821), .B(
        n9820), .ZN(P1_U3243) );
  INV_X1 U10924 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U10925 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n4701), .ZN(n9827) );
  AOI211_X1 U10926 ( .C1(n9825), .C2(n9824), .A(n9847), .B(n9823), .ZN(n9826)
         );
  AOI211_X1 U10927 ( .C1(n9853), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9833)
         );
  XOR2_X1 U10928 ( .A(n9830), .B(n9829), .Z(n9831) );
  NAND2_X1 U10929 ( .A1(n9831), .A2(n9841), .ZN(n9832) );
  OAI211_X1 U10930 ( .C1(n9834), .C2(n9862), .A(n9833), .B(n9832), .ZN(
        P1_U3257) );
  AOI211_X1 U10931 ( .C1(n9836), .C2(n9835), .A(n4312), .B(n9847), .ZN(n9837)
         );
  AOI211_X1 U10932 ( .C1(n9853), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9845)
         );
  OAI211_X1 U10933 ( .C1(n9843), .C2(n9842), .A(n9841), .B(n9840), .ZN(n9844)
         );
  OAI211_X1 U10934 ( .C1(n4522), .C2(n9862), .A(n9845), .B(n9844), .ZN(
        P1_U3258) );
  INV_X1 U10935 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9863) );
  INV_X1 U10936 ( .A(n9846), .ZN(n9852) );
  AOI211_X1 U10937 ( .C1(n9850), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9851)
         );
  AOI211_X1 U10938 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9861)
         );
  AOI21_X1 U10939 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9859) );
  OR2_X1 U10940 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  OAI211_X1 U10941 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9860), .ZN(
        P1_U3259) );
  INV_X1 U10942 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9864) );
  NOR2_X1 U10943 ( .A1(n9891), .A2(n9864), .ZN(P1_U3292) );
  INV_X1 U10944 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9865) );
  NOR2_X1 U10945 ( .A1(n9891), .A2(n9865), .ZN(P1_U3293) );
  INV_X1 U10946 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10155) );
  NOR2_X1 U10947 ( .A1(n9891), .A2(n10155), .ZN(P1_U3294) );
  INV_X1 U10948 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U10949 ( .A1(n9875), .A2(n9866), .ZN(P1_U3295) );
  INV_X1 U10950 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9867) );
  NOR2_X1 U10951 ( .A1(n9875), .A2(n9867), .ZN(P1_U3296) );
  INV_X1 U10952 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9868) );
  NOR2_X1 U10953 ( .A1(n9875), .A2(n9868), .ZN(P1_U3297) );
  INV_X1 U10954 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9869) );
  NOR2_X1 U10955 ( .A1(n9875), .A2(n9869), .ZN(P1_U3298) );
  INV_X1 U10956 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U10957 ( .A1(n9875), .A2(n9870), .ZN(P1_U3299) );
  INV_X1 U10958 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10176) );
  NOR2_X1 U10959 ( .A1(n9875), .A2(n10176), .ZN(P1_U3300) );
  INV_X1 U10960 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U10961 ( .A1(n9875), .A2(n9871), .ZN(P1_U3301) );
  INV_X1 U10962 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9872) );
  NOR2_X1 U10963 ( .A1(n9875), .A2(n9872), .ZN(P1_U3302) );
  INV_X1 U10964 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9873) );
  NOR2_X1 U10965 ( .A1(n9875), .A2(n9873), .ZN(P1_U3303) );
  INV_X1 U10966 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U10967 ( .A1(n9875), .A2(n9874), .ZN(P1_U3304) );
  INV_X1 U10968 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9876) );
  NOR2_X1 U10969 ( .A1(n9891), .A2(n9876), .ZN(P1_U3305) );
  INV_X1 U10970 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9877) );
  NOR2_X1 U10971 ( .A1(n9891), .A2(n9877), .ZN(P1_U3306) );
  INV_X1 U10972 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9878) );
  NOR2_X1 U10973 ( .A1(n9891), .A2(n9878), .ZN(P1_U3307) );
  INV_X1 U10974 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9879) );
  NOR2_X1 U10975 ( .A1(n9891), .A2(n9879), .ZN(P1_U3308) );
  INV_X1 U10976 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9880) );
  NOR2_X1 U10977 ( .A1(n9891), .A2(n9880), .ZN(P1_U3309) );
  INV_X1 U10978 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9881) );
  NOR2_X1 U10979 ( .A1(n9891), .A2(n9881), .ZN(P1_U3310) );
  INV_X1 U10980 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9882) );
  NOR2_X1 U10981 ( .A1(n9891), .A2(n9882), .ZN(P1_U3311) );
  INV_X1 U10982 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U10983 ( .A1(n9891), .A2(n9883), .ZN(P1_U3312) );
  INV_X1 U10984 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U10985 ( .A1(n9891), .A2(n10119), .ZN(P1_U3313) );
  INV_X1 U10986 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9884) );
  NOR2_X1 U10987 ( .A1(n9891), .A2(n9884), .ZN(P1_U3314) );
  INV_X1 U10988 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9885) );
  NOR2_X1 U10989 ( .A1(n9891), .A2(n9885), .ZN(P1_U3315) );
  INV_X1 U10990 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9886) );
  NOR2_X1 U10991 ( .A1(n9891), .A2(n9886), .ZN(P1_U3316) );
  INV_X1 U10992 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9887) );
  NOR2_X1 U10993 ( .A1(n9891), .A2(n9887), .ZN(P1_U3317) );
  INV_X1 U10994 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U10995 ( .A1(n9891), .A2(n9888), .ZN(P1_U3318) );
  INV_X1 U10996 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9889) );
  NOR2_X1 U10997 ( .A1(n9891), .A2(n9889), .ZN(P1_U3319) );
  INV_X1 U10998 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U10999 ( .A1(n9891), .A2(n9890), .ZN(P1_U3320) );
  INV_X1 U11000 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10152) );
  NOR2_X1 U11001 ( .A1(n9891), .A2(n10152), .ZN(P1_U3321) );
  NAND2_X1 U11002 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  OAI211_X1 U11003 ( .C1(n9898), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9900)
         );
  NOR2_X1 U11004 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  NOR3_X1 U11005 ( .A1(n9901), .A2(n9900), .A3(n9899), .ZN(n9959) );
  AOI22_X1 U11006 ( .A1(n9958), .A2(n9959), .B1(n5209), .B2(n9956), .ZN(
        P1_U3457) );
  INV_X1 U11007 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U11008 ( .A1(n9958), .A2(n9902), .B1(n10166), .B2(n9956), .ZN(
        P1_U3460) );
  INV_X1 U11009 ( .A(n9903), .ZN(n9908) );
  OAI22_X1 U11010 ( .A1(n9904), .A2(n9949), .B1(n4989), .B2(n9947), .ZN(n9907)
         );
  INV_X1 U11011 ( .A(n9905), .ZN(n9906) );
  AOI211_X1 U11012 ( .C1(n9912), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9961)
         );
  INV_X1 U11013 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U11014 ( .A1(n9958), .A2(n9961), .B1(n10132), .B2(n9956), .ZN(
        P1_U3463) );
  OAI22_X1 U11015 ( .A1(n9910), .A2(n9949), .B1(n9909), .B2(n9947), .ZN(n9911)
         );
  AOI21_X1 U11016 ( .B1(n9913), .B2(n9912), .A(n9911), .ZN(n9914) );
  AND2_X1 U11017 ( .A1(n9915), .A2(n9914), .ZN(n9963) );
  INV_X1 U11018 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U11019 ( .A1(n9958), .A2(n9963), .B1(n9916), .B2(n9956), .ZN(
        P1_U3466) );
  INV_X1 U11020 ( .A(n9917), .ZN(n9921) );
  AOI21_X1 U11021 ( .B1(n9919), .B2(n9918), .A(n7472), .ZN(n9920) );
  NOR2_X1 U11022 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  OAI222_X1 U11023 ( .A1(n9927), .A2(n9926), .B1(n9925), .B2(n9924), .C1(n9923), .C2(n9922), .ZN(n10223) );
  NAND2_X1 U11024 ( .A1(n7475), .A2(n7472), .ZN(n10215) );
  NAND3_X1 U11025 ( .A1(n10216), .A2(n10215), .A3(n9952), .ZN(n9930) );
  OAI211_X1 U11026 ( .C1(n9929), .C2(n10209), .A(n4997), .B(n9928), .ZN(n10219) );
  OAI211_X1 U11027 ( .C1(n10209), .C2(n9947), .A(n9930), .B(n10219), .ZN(n9931) );
  NOR2_X1 U11028 ( .A1(n10223), .A2(n9931), .ZN(n9965) );
  INV_X1 U11029 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U11030 ( .A1(n9958), .A2(n9965), .B1(n9932), .B2(n9956), .ZN(
        P1_U3469) );
  OAI22_X1 U11031 ( .A1(n9934), .A2(n9949), .B1(n9933), .B2(n9947), .ZN(n9936)
         );
  AOI211_X1 U11032 ( .C1(n9937), .C2(n9952), .A(n9936), .B(n9935), .ZN(n9966)
         );
  INV_X1 U11033 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U11034 ( .A1(n9958), .A2(n9966), .B1(n9938), .B2(n9956), .ZN(
        P1_U3472) );
  AND2_X1 U11035 ( .A1(n9939), .A2(n9952), .ZN(n9943) );
  OAI21_X1 U11036 ( .B1(n9941), .B2(n9947), .A(n9940), .ZN(n9942) );
  NOR3_X1 U11037 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9968) );
  INV_X1 U11038 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9945) );
  AOI22_X1 U11039 ( .A1(n9958), .A2(n9968), .B1(n9945), .B2(n9956), .ZN(
        P1_U3475) );
  INV_X1 U11040 ( .A(n9946), .ZN(n9953) );
  OAI22_X1 U11041 ( .A1(n9950), .A2(n9949), .B1(n9948), .B2(n9947), .ZN(n9951)
         );
  AOI21_X1 U11042 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9954) );
  AND2_X1 U11043 ( .A1(n9955), .A2(n9954), .ZN(n9971) );
  INV_X1 U11044 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11045 ( .A1(n9958), .A2(n9971), .B1(n9957), .B2(n9956), .ZN(
        P1_U3478) );
  AOI22_X1 U11046 ( .A1(n9972), .A2(n9959), .B1(n6782), .B2(n9969), .ZN(
        P1_U3524) );
  INV_X1 U11047 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11048 ( .A1(n9972), .A2(n9961), .B1(n9960), .B2(n9969), .ZN(
        P1_U3526) );
  AOI22_X1 U11049 ( .A1(n9972), .A2(n9963), .B1(n9962), .B2(n9969), .ZN(
        P1_U3527) );
  INV_X1 U11050 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11051 ( .A1(n9972), .A2(n9965), .B1(n9964), .B2(n9969), .ZN(
        P1_U3528) );
  AOI22_X1 U11052 ( .A1(n9972), .A2(n9966), .B1(n4389), .B2(n9969), .ZN(
        P1_U3529) );
  INV_X1 U11053 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9967) );
  AOI22_X1 U11054 ( .A1(n9972), .A2(n9968), .B1(n9967), .B2(n9969), .ZN(
        P1_U3530) );
  AOI22_X1 U11055 ( .A1(n9972), .A2(n9971), .B1(n9970), .B2(n9969), .ZN(
        P1_U3531) );
  AOI22_X1 U11056 ( .A1(n9974), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n9973), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11057 ( .A1(n9975), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9982) );
  NOR2_X1 U11058 ( .A1(n9976), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9980) );
  OAI21_X1 U11059 ( .B1(n9978), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9977), .ZN(
        n9979) );
  OAI21_X1 U11060 ( .B1(n9980), .B2(n9979), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9981) );
  OAI211_X1 U11061 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9983), .A(n9982), .B(
        n9981), .ZN(P2_U3245) );
  NAND2_X1 U11062 ( .A1(n9984), .A2(n6532), .ZN(n9988) );
  NAND2_X1 U11063 ( .A1(n9986), .A2(n9985), .ZN(n9987) );
  OAI211_X1 U11064 ( .C1(n9990), .C2(n9989), .A(n9988), .B(n9987), .ZN(n9993)
         );
  INV_X1 U11065 ( .A(n9991), .ZN(n9992) );
  AOI211_X1 U11066 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(n9997)
         );
  AOI22_X1 U11067 ( .A1(n9998), .A2(n6952), .B1(n9997), .B2(n9996), .ZN(
        P2_U3291) );
  AND2_X1 U11068 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10004), .ZN(P2_U3297) );
  AND2_X1 U11069 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10004), .ZN(P2_U3298) );
  AND2_X1 U11070 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10004), .ZN(P2_U3299) );
  AND2_X1 U11071 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10004), .ZN(P2_U3300) );
  AND2_X1 U11072 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10004), .ZN(P2_U3301) );
  AND2_X1 U11073 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10004), .ZN(P2_U3302) );
  AND2_X1 U11074 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10004), .ZN(P2_U3303) );
  AND2_X1 U11075 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10004), .ZN(P2_U3304) );
  AND2_X1 U11076 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10004), .ZN(P2_U3305) );
  AND2_X1 U11077 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10004), .ZN(P2_U3306) );
  AND2_X1 U11078 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10004), .ZN(P2_U3307) );
  AND2_X1 U11079 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10004), .ZN(P2_U3308) );
  AND2_X1 U11080 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10004), .ZN(P2_U3309) );
  INV_X1 U11081 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U11082 ( .A1(n10001), .A2(n10109), .ZN(P2_U3310) );
  AND2_X1 U11083 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10004), .ZN(P2_U3311) );
  AND2_X1 U11084 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10004), .ZN(P2_U3312) );
  AND2_X1 U11085 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10004), .ZN(P2_U3313) );
  AND2_X1 U11086 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10004), .ZN(P2_U3314) );
  INV_X1 U11087 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U11088 ( .A1(n10001), .A2(n10191), .ZN(P2_U3315) );
  AND2_X1 U11089 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10004), .ZN(P2_U3316) );
  AND2_X1 U11090 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10004), .ZN(P2_U3317) );
  AND2_X1 U11091 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10004), .ZN(P2_U3318) );
  INV_X1 U11092 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U11093 ( .A1(n10001), .A2(n10149), .ZN(P2_U3319) );
  AND2_X1 U11094 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10004), .ZN(P2_U3320) );
  INV_X1 U11095 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U11096 ( .A1(n10001), .A2(n10163), .ZN(P2_U3321) );
  AND2_X1 U11097 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10004), .ZN(P2_U3322) );
  AND2_X1 U11098 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10004), .ZN(P2_U3323) );
  AND2_X1 U11099 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10004), .ZN(P2_U3324) );
  AND2_X1 U11100 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10004), .ZN(P2_U3325) );
  AND2_X1 U11101 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10004), .ZN(P2_U3326) );
  AOI22_X1 U11102 ( .A1(n10007), .A2(n10003), .B1(n10002), .B2(n10004), .ZN(
        P2_U3437) );
  AOI22_X1 U11103 ( .A1(n10007), .A2(n10006), .B1(n10005), .B2(n10004), .ZN(
        P2_U3438) );
  OAI21_X1 U11104 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10011) );
  AOI21_X1 U11105 ( .B1(n10028), .B2(n10012), .A(n10011), .ZN(n10031) );
  INV_X1 U11106 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10013) );
  AOI22_X1 U11107 ( .A1(n10030), .A2(n10031), .B1(n10013), .B2(n4455), .ZN(
        P2_U3451) );
  INV_X1 U11108 ( .A(n10014), .ZN(n10016) );
  OAI22_X1 U11109 ( .A1(n10016), .A2(n10022), .B1(n10015), .B2(n10020), .ZN(
        n10017) );
  AOI211_X1 U11110 ( .C1(n10028), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10033) );
  AOI22_X1 U11111 ( .A1(n10030), .A2(n10033), .B1(n6043), .B2(n4455), .ZN(
        P2_U3463) );
  OAI22_X1 U11112 ( .A1(n10023), .A2(n10022), .B1(n10021), .B2(n10020), .ZN(
        n10026) );
  INV_X1 U11113 ( .A(n10024), .ZN(n10025) );
  AOI211_X1 U11114 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10034) );
  INV_X1 U11115 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U11116 ( .A1(n10030), .A2(n10034), .B1(n10029), .B2(n4455), .ZN(
        P2_U3469) );
  AOI22_X1 U11117 ( .A1(n4333), .A2(n10031), .B1(n6913), .B2(n4315), .ZN(
        P2_U3520) );
  AOI22_X1 U11118 ( .A1(n4333), .A2(n10033), .B1(n10032), .B2(n4315), .ZN(
        P2_U3524) );
  AOI22_X1 U11119 ( .A1(n4333), .A2(n10034), .B1(n6974), .B2(n4315), .ZN(
        P2_U3526) );
  INV_X1 U11120 ( .A(n10035), .ZN(n10036) );
  NAND2_X1 U11121 ( .A1(n10037), .A2(n10036), .ZN(n10038) );
  XNOR2_X1 U11122 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10038), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11123 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11124 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(ADD_1071_U56) );
  OAI21_X1 U11125 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(ADD_1071_U57) );
  OAI21_X1 U11126 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(ADD_1071_U58) );
  OAI21_X1 U11127 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(ADD_1071_U59) );
  OAI21_X1 U11128 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(ADD_1071_U60) );
  OAI21_X1 U11129 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(ADD_1071_U61) );
  AOI21_X1 U11130 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(ADD_1071_U62) );
  AOI21_X1 U11131 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(ADD_1071_U63) );
  INV_X1 U11132 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10179) );
  NOR4_X1 U11133 ( .A1(SI_25_), .A2(P2_REG3_REG_19__SCAN_IN), .A3(n10182), 
        .A4(n10179), .ZN(n10074) );
  NOR4_X1 U11134 ( .A1(n10138), .A2(P1_DATAO_REG_11__SCAN_IN), .A3(
        P1_DATAO_REG_4__SCAN_IN), .A4(P2_DATAO_REG_8__SCAN_IN), .ZN(n10073) );
  AND4_X1 U11135 ( .A1(n10063), .A2(P1_DATAO_REG_26__SCAN_IN), .A3(SI_27_), 
        .A4(P1_DATAO_REG_31__SCAN_IN), .ZN(n10072) );
  NOR3_X1 U11136 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P2_REG1_REG_16__SCAN_IN), 
        .A3(P2_REG2_REG_8__SCAN_IN), .ZN(n10067) );
  NOR4_X1 U11137 ( .A1(P1_REG0_REG_3__SCAN_IN), .A2(P2_REG2_REG_25__SCAN_IN), 
        .A3(P2_REG0_REG_15__SCAN_IN), .A4(n6974), .ZN(n10066) );
  NOR3_X1 U11138 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(n10064), .ZN(n10065) );
  NAND4_X1 U11139 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(n10067), .A3(n10066), .A4(
        n10065), .ZN(n10068) );
  OR4_X1 U11140 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(n10120), .A3(P2_B_REG_SCAN_IN), .A4(n10068), .ZN(n10070) );
  NAND4_X1 U11141 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(P2_DATAO_REG_9__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n10069) );
  NOR4_X1 U11142 ( .A1(n10070), .A2(P1_D_REG_10__SCAN_IN), .A3(n10176), .A4(
        n10069), .ZN(n10071) );
  AND4_X1 U11143 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10207) );
  NOR4_X1 U11144 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), 
        .A3(P2_REG0_REG_20__SCAN_IN), .A4(n10075), .ZN(n10087) );
  NAND4_X1 U11145 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_16__SCAN_IN), .A3(P2_D_REG_18__SCAN_IN), .A4(
        P2_REG3_REG_6__SCAN_IN), .ZN(n10078) );
  NAND4_X1 U11146 ( .A1(n10163), .A2(n10076), .A3(P2_ADDR_REG_13__SCAN_IN), 
        .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n10077) );
  NOR2_X1 U11147 ( .A1(n10078), .A2(n10077), .ZN(n10086) );
  NOR2_X1 U11148 ( .A1(P2_RD_REG_SCAN_IN), .A2(SI_31_), .ZN(n10080) );
  NOR4_X1 U11149 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), 
        .A3(P2_REG2_REG_23__SCAN_IN), .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n10079) );
  AND4_X1 U11150 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(P2_REG3_REG_1__SCAN_IN), 
        .A3(n10080), .A4(n10079), .ZN(n10081) );
  NAND4_X1 U11151 ( .A1(n10082), .A2(n10105), .A3(P1_ADDR_REG_19__SCAN_IN), 
        .A4(n10081), .ZN(n10084) );
  NAND4_X1 U11152 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(SI_21_), .A3(
        P2_REG3_REG_7__SCAN_IN), .A4(P1_DATAO_REG_30__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U11153 ( .A1(n10084), .A2(n10083), .ZN(n10085) );
  AND4_X1 U11154 ( .A1(n10087), .A2(n10091), .A3(n10086), .A4(n10085), .ZN(
        n10089) );
  NOR4_X1 U11155 ( .A1(P1_D_REG_29__SCAN_IN), .A2(SI_22_), .A3(
        P2_DATAO_REG_21__SCAN_IN), .A4(n10152), .ZN(n10088) );
  AND2_X1 U11156 ( .A1(n10089), .A2(n10088), .ZN(n10206) );
  INV_X1 U11157 ( .A(SI_21_), .ZN(n10092) );
  AOI22_X1 U11158 ( .A1(n10092), .A2(keyinput17), .B1(n10091), .B2(keyinput2), 
        .ZN(n10090) );
  OAI221_X1 U11159 ( .B1(n10092), .B2(keyinput17), .C1(n10091), .C2(keyinput2), 
        .A(n10090), .ZN(n10103) );
  INV_X1 U11160 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10095) );
  INV_X1 U11161 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11162 ( .A1(n10095), .A2(keyinput59), .B1(n10094), .B2(keyinput29), 
        .ZN(n10093) );
  OAI221_X1 U11163 ( .B1(n10095), .B2(keyinput59), .C1(n10094), .C2(keyinput29), .A(n10093), .ZN(n10102) );
  AOI22_X1 U11164 ( .A1(n6092), .A2(keyinput56), .B1(keyinput48), .B2(n10097), 
        .ZN(n10096) );
  OAI221_X1 U11165 ( .B1(n6092), .B2(keyinput56), .C1(n10097), .C2(keyinput48), 
        .A(n10096), .ZN(n10101) );
  XOR2_X1 U11166 ( .A(n6523), .B(keyinput43), .Z(n10099) );
  XNOR2_X1 U11167 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput41), .ZN(n10098) );
  NAND2_X1 U11168 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NOR4_X1 U11169 ( .A1(n10103), .A2(n10102), .A3(n10101), .A4(n10100), .ZN(
        n10146) );
  AOI22_X1 U11170 ( .A1(n10105), .A2(keyinput20), .B1(keyinput52), .B2(n6976), 
        .ZN(n10104) );
  OAI221_X1 U11171 ( .B1(n10105), .B2(keyinput20), .C1(n6976), .C2(keyinput52), 
        .A(n10104), .ZN(n10117) );
  AOI22_X1 U11172 ( .A1(n10108), .A2(keyinput53), .B1(n10107), .B2(keyinput31), 
        .ZN(n10106) );
  OAI221_X1 U11173 ( .B1(n10108), .B2(keyinput53), .C1(n10107), .C2(keyinput31), .A(n10106), .ZN(n10116) );
  XNOR2_X1 U11174 ( .A(n10109), .B(keyinput30), .ZN(n10115) );
  XOR2_X1 U11175 ( .A(n10110), .B(keyinput33), .Z(n10113) );
  XNOR2_X1 U11176 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput39), .ZN(n10112)
         );
  XNOR2_X1 U11177 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput47), .ZN(n10111) );
  NAND3_X1 U11178 ( .A1(n10113), .A2(n10112), .A3(n10111), .ZN(n10114) );
  NOR4_X1 U11179 ( .A1(n10117), .A2(n10116), .A3(n10115), .A4(n10114), .ZN(
        n10145) );
  AOI22_X1 U11180 ( .A1(n6169), .A2(keyinput5), .B1(n10119), .B2(keyinput57), 
        .ZN(n10118) );
  OAI221_X1 U11181 ( .B1(n6169), .B2(keyinput5), .C1(n10119), .C2(keyinput57), 
        .A(n10118), .ZN(n10129) );
  XNOR2_X1 U11182 ( .A(n10120), .B(keyinput26), .ZN(n10128) );
  XNOR2_X1 U11183 ( .A(keyinput54), .B(n10121), .ZN(n10127) );
  XNOR2_X1 U11184 ( .A(P2_B_REG_SCAN_IN), .B(keyinput63), .ZN(n10125) );
  XNOR2_X1 U11185 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput12), .ZN(n10124)
         );
  XNOR2_X1 U11186 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput1), .ZN(n10123) );
  XNOR2_X1 U11187 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput18), .ZN(n10122)
         );
  NAND4_X1 U11188 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10126) );
  NOR4_X1 U11189 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        n10144) );
  AOI22_X1 U11190 ( .A1(n6974), .A2(keyinput7), .B1(n8764), .B2(keyinput14), 
        .ZN(n10130) );
  OAI221_X1 U11191 ( .B1(n6974), .B2(keyinput7), .C1(n8764), .C2(keyinput14), 
        .A(n10130), .ZN(n10142) );
  INV_X1 U11192 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11193 ( .A1(n10133), .A2(keyinput3), .B1(n10132), .B2(keyinput36), 
        .ZN(n10131) );
  OAI221_X1 U11194 ( .B1(n10133), .B2(keyinput3), .C1(n10132), .C2(keyinput36), 
        .A(n10131), .ZN(n10141) );
  AOI22_X1 U11195 ( .A1(n10136), .A2(keyinput51), .B1(keyinput60), .B2(n10135), 
        .ZN(n10134) );
  OAI221_X1 U11196 ( .B1(n10136), .B2(keyinput51), .C1(n10135), .C2(keyinput60), .A(n10134), .ZN(n10140) );
  AOI22_X1 U11197 ( .A1(n7644), .A2(keyinput11), .B1(n10138), .B2(keyinput24), 
        .ZN(n10137) );
  OAI221_X1 U11198 ( .B1(n7644), .B2(keyinput11), .C1(n10138), .C2(keyinput24), 
        .A(n10137), .ZN(n10139) );
  NOR4_X1 U11199 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10143) );
  NAND4_X1 U11200 ( .A1(n10146), .A2(n10145), .A3(n10144), .A4(n10143), .ZN(
        n10205) );
  AOI22_X1 U11201 ( .A1(n10149), .A2(keyinput37), .B1(keyinput10), .B2(n10148), 
        .ZN(n10147) );
  OAI221_X1 U11202 ( .B1(n10149), .B2(keyinput37), .C1(n10148), .C2(keyinput10), .A(n10147), .ZN(n10161) );
  AOI22_X1 U11203 ( .A1(n10152), .A2(keyinput27), .B1(keyinput58), .B2(n10151), 
        .ZN(n10150) );
  OAI221_X1 U11204 ( .B1(n10152), .B2(keyinput27), .C1(n10151), .C2(keyinput58), .A(n10150), .ZN(n10160) );
  AOI22_X1 U11205 ( .A1(n10155), .A2(keyinput34), .B1(keyinput40), .B2(n10154), 
        .ZN(n10153) );
  OAI221_X1 U11206 ( .B1(n10155), .B2(keyinput34), .C1(n10154), .C2(keyinput40), .A(n10153), .ZN(n10159) );
  XNOR2_X1 U11207 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput46), .ZN(n10157)
         );
  XNOR2_X1 U11208 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput38), .ZN(n10156)
         );
  NAND2_X1 U11209 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NOR4_X1 U11210 ( .A1(n10161), .A2(n10160), .A3(n10159), .A4(n10158), .ZN(
        n10203) );
  AOI22_X1 U11211 ( .A1(n10163), .A2(keyinput61), .B1(keyinput9), .B2(n7756), 
        .ZN(n10162) );
  OAI221_X1 U11212 ( .B1(n10163), .B2(keyinput61), .C1(n7756), .C2(keyinput9), 
        .A(n10162), .ZN(n10173) );
  AOI22_X1 U11213 ( .A1(n6341), .A2(keyinput45), .B1(keyinput21), .B2(n10165), 
        .ZN(n10164) );
  OAI221_X1 U11214 ( .B1(n6341), .B2(keyinput45), .C1(n10165), .C2(keyinput21), 
        .A(n10164), .ZN(n10172) );
  XOR2_X1 U11215 ( .A(n10166), .B(keyinput32), .Z(n10170) );
  XNOR2_X1 U11216 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput0), .ZN(n10169) );
  XNOR2_X1 U11217 ( .A(SI_12_), .B(keyinput62), .ZN(n10168) );
  XNOR2_X1 U11218 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput42), .ZN(n10167)
         );
  NAND4_X1 U11219 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10171) );
  NOR3_X1 U11220 ( .A1(n10173), .A2(n10172), .A3(n10171), .ZN(n10202) );
  AOI22_X1 U11221 ( .A1(n10176), .A2(keyinput22), .B1(keyinput19), .B2(n10175), 
        .ZN(n10174) );
  OAI221_X1 U11222 ( .B1(n10176), .B2(keyinput22), .C1(n10175), .C2(keyinput19), .A(n10174), .ZN(n10188) );
  AOI22_X1 U11223 ( .A1(n10179), .A2(keyinput4), .B1(n10178), .B2(keyinput49), 
        .ZN(n10177) );
  OAI221_X1 U11224 ( .B1(n10179), .B2(keyinput4), .C1(n10178), .C2(keyinput49), 
        .A(n10177), .ZN(n10187) );
  AOI22_X1 U11225 ( .A1(n10182), .A2(keyinput50), .B1(n10181), .B2(keyinput6), 
        .ZN(n10180) );
  OAI221_X1 U11226 ( .B1(n10182), .B2(keyinput50), .C1(n10181), .C2(keyinput6), 
        .A(n10180), .ZN(n10186) );
  XNOR2_X1 U11227 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput28), .ZN(n10184)
         );
  XNOR2_X1 U11228 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput23), .ZN(n10183) );
  NAND2_X1 U11229 ( .A1(n10184), .A2(n10183), .ZN(n10185) );
  NOR4_X1 U11230 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10201) );
  AOI22_X1 U11231 ( .A1(n10191), .A2(keyinput8), .B1(n10190), .B2(keyinput35), 
        .ZN(n10189) );
  OAI221_X1 U11232 ( .B1(n10191), .B2(keyinput8), .C1(n10190), .C2(keyinput35), 
        .A(n10189), .ZN(n10199) );
  XOR2_X1 U11233 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput44), .Z(n10198) );
  XNOR2_X1 U11234 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(keyinput13), .ZN(n10195)
         );
  XNOR2_X1 U11235 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput55), .ZN(n10194)
         );
  XNOR2_X1 U11236 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(keyinput25), .ZN(n10193)
         );
  XNOR2_X1 U11237 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput16), .ZN(n10192)
         );
  NAND4_X1 U11238 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10197) );
  XNOR2_X1 U11239 ( .A(keyinput15), .B(n10063), .ZN(n10196) );
  NOR4_X1 U11240 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NAND4_X1 U11241 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  AOI211_X1 U11242 ( .C1(n10207), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        n10225) );
  NOR2_X1 U11243 ( .A1(n10209), .A2(n10208), .ZN(n10211) );
  AOI211_X1 U11244 ( .C1(n10213), .C2(n10212), .A(n10211), .B(n10210), .ZN(
        n10218) );
  NAND3_X1 U11245 ( .A1(n10216), .A2(n10215), .A3(n10214), .ZN(n10217) );
  OAI211_X1 U11246 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        n10222) );
  OAI22_X1 U11247 ( .A1(n10223), .A2(n10222), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n10221), .ZN(n10224) );
  XNOR2_X1 U11248 ( .A(n10225), .B(n10224), .ZN(P1_U3286) );
  XOR2_X1 U11249 ( .A(n10226), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11250 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  XNOR2_X1 U11251 ( .A(n10229), .B(n4526), .ZN(ADD_1071_U51) );
  OAI21_X1 U11252 ( .B1(n10232), .B2(n10231), .A(n10230), .ZN(n10233) );
  XNOR2_X1 U11253 ( .A(n10233), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11254 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(ADD_1071_U47) );
  XOR2_X1 U11255 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10237), .Z(ADD_1071_U48) );
  XOR2_X1 U11256 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10238), .Z(ADD_1071_U49) );
  XOR2_X1 U11257 ( .A(n10240), .B(n10239), .Z(ADD_1071_U54) );
  XOR2_X1 U11258 ( .A(n10242), .B(n10241), .Z(ADD_1071_U53) );
  XNOR2_X1 U11259 ( .A(n10244), .B(n10243), .ZN(ADD_1071_U52) );
  NAND2_X1 U8005 ( .A1(n6368), .A2(n6367), .ZN(n8998) );
  CLKBUF_X1 U4752 ( .A(n4303), .Z(n4633) );
  AND2_X1 U4757 ( .A1(n6910), .A2(n5270), .ZN(n6040) );
  CLKBUF_X2 U4782 ( .A(n6037), .Z(n6249) );
  NOR2_X2 U4799 ( .A1(n8770), .A2(n8998), .ZN(n8756) );
  CLKBUF_X2 U4913 ( .A(n5368), .Z(n4626) );
  AND2_X1 U6124 ( .A1(n9406), .A2(n8426), .ZN(n9390) );
  XNOR2_X1 U6549 ( .A(n5538), .B(n5533), .ZN(n6829) );
endmodule

