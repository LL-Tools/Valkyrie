

module b20_C_AntiSAT_k_256_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691;

  AOI211_X1 U5017 ( .C1(n10612), .C2(n9482), .A(n9481), .B(n9480), .ZN(n9485)
         );
  NAND2_X1 U5018 ( .A1(n5049), .A2(n5046), .ZN(n4693) );
  AOI21_X1 U5019 ( .B1(n5031), .B2(n5030), .A(n5029), .ZN(n8209) );
  NAND2_X2 U5020 ( .A1(n5836), .A2(n5835), .ZN(n10275) );
  XNOR2_X1 U5021 ( .A(n5566), .B(n5565), .ZN(n7523) );
  INV_X1 U5022 ( .A(n5333), .ZN(n5555) );
  CLKBUF_X2 U5023 ( .A(n5340), .Z(n4522) );
  AND2_X1 U5024 ( .A1(n5276), .A2(n9802), .ZN(n8442) );
  BUF_X1 U5025 ( .A(n6296), .Z(n6479) );
  NAND2_X1 U5026 ( .A1(n4989), .A2(n5947), .ZN(n10477) );
  INV_X1 U5027 ( .A(n8530), .ZN(n6049) );
  INV_X2 U5028 ( .A(n5147), .ZN(n5788) );
  CLKBUF_X3 U5029 ( .A(n5788), .Z(n4517) );
  CLKBUF_X2 U5030 ( .A(n8442), .Z(n4520) );
  AND2_X1 U5031 ( .A1(n8118), .A2(n8117), .ZN(n8159) );
  AOI21_X2 U5032 ( .B1(n9587), .B2(n8402), .A(n8401), .ZN(n9576) );
  NAND2_X1 U5033 ( .A1(n8285), .A2(n8280), .ZN(n6861) );
  AND2_X1 U5034 ( .A1(n6478), .A2(n6477), .ZN(n9880) );
  XNOR2_X1 U5035 ( .A(n8159), .B(n8177), .ZN(n8120) );
  INV_X1 U5036 ( .A(n8521), .ZN(n9521) );
  AND2_X1 U5037 ( .A1(n5049), .A2(n5048), .ZN(n9885) );
  AND4_X1 U5038 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n6932)
         );
  AND2_X1 U5039 ( .A1(n6185), .A2(n8701), .ZN(n8765) );
  XNOR2_X1 U5040 ( .A(n5413), .B(n5412), .ZN(n6630) );
  INV_X1 U5041 ( .A(n6166), .ZN(n8816) );
  AND4_X2 U5042 ( .A1(n4683), .A2(n4684), .A3(n5066), .A4(n5778), .ZN(n4511)
         );
  INV_X1 U5043 ( .A(n8453), .ZN(n8448) );
  AND3_X2 U5045 ( .A1(n4912), .A2(n9519), .A3(n4913), .ZN(n9520) );
  AOI21_X2 U5046 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9475), .A(n9474), .ZN(
        n9488) );
  NAND2_X2 U5047 ( .A1(n5297), .A2(n5296), .ZN(n5150) );
  NAND2_X2 U5048 ( .A1(n5146), .A2(n5145), .ZN(n5297) );
  NAND2_X2 U5049 ( .A1(n8132), .A2(n8131), .ZN(n8165) );
  BUF_X4 U5050 ( .A(n5908), .Z(n8537) );
  BUF_X1 U5051 ( .A(n6979), .Z(n4512) );
  BUF_X2 U5052 ( .A(n6979), .Z(n4513) );
  NAND3_X1 U5053 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(n6979) );
  OR2_X2 U5054 ( .A1(n10486), .A2(n7640), .ZN(n8658) );
  AOI211_X1 U5055 ( .C1(n8834), .C2(n8833), .A(n8832), .B(n8831), .ZN(n8836)
         );
  OR2_X2 U5057 ( .A1(n9467), .A2(n4613), .ZN(n4912) );
  AND2_X4 U5058 ( .A1(n6274), .A2(n6272), .ZN(n6354) );
  INV_X2 U5059 ( .A(n7692), .ZN(n7341) );
  OAI21_X2 U5060 ( .B1(n6616), .B2(n5913), .A(n5916), .ZN(n7692) );
  NOR2_X2 U5061 ( .A1(n7550), .A2(n7549), .ZN(n7551) );
  OAI22_X2 U5062 ( .A1(n7269), .A2(n4856), .B1(n4583), .B2(n7160), .ZN(n7550)
         );
  AND2_X2 U5063 ( .A1(n4905), .A2(n4621), .ZN(n9506) );
  NAND4_X2 U5064 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n9387)
         );
  XNOR2_X2 U5065 ( .A(n5337), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10549) );
  XNOR2_X2 U5066 ( .A(n5264), .B(n5271), .ZN(n5668) );
  OAI21_X1 U5067 ( .B1(n9634), .B2(n9374), .A(n9626), .ZN(n9614) );
  AOI21_X1 U5068 ( .B1(n8057), .B2(n8763), .A(n6045), .ZN(n8144) );
  OAI22_X1 U5069 ( .A1(n7594), .A2(n5449), .B1(n7780), .B2(n8011), .ZN(n7656)
         );
  NAND2_X1 U5070 ( .A1(n5935), .A2(n5934), .ZN(n10442) );
  NAND2_X2 U5071 ( .A1(n6978), .A2(n7099), .ZN(n8285) );
  AND2_X1 U5072 ( .A1(n8293), .A2(n8292), .ZN(n8281) );
  NAND2_X2 U5073 ( .A1(n6514), .A2(n6517), .ZN(n6296) );
  INV_X1 U5074 ( .A(n9725), .ZN(n7099) );
  INV_X2 U5075 ( .A(n6514), .ZN(n6327) );
  INV_X2 U5076 ( .A(n4512), .ZN(n8244) );
  INV_X4 U5077 ( .A(n6517), .ZN(n4514) );
  CLKBUF_X2 U5079 ( .A(n5339), .Z(n4525) );
  BUF_X2 U5080 ( .A(n5340), .Z(n4523) );
  AND2_X1 U5081 ( .A1(n5276), .A2(n5277), .ZN(n5340) );
  BUF_X4 U5082 ( .A(n5339), .Z(n4515) );
  NOR2_X1 U5083 ( .A1(n5819), .A2(n5043), .ZN(n5038) );
  CLKBUF_X3 U5084 ( .A(n5788), .Z(n4516) );
  MUX2_X1 U5085 ( .A(n10294), .B(n10293), .S(n10523), .Z(n10295) );
  MUX2_X1 U5086 ( .A(n10224), .B(n10293), .S(n10537), .Z(n10225) );
  NOR2_X1 U5087 ( .A1(n10057), .A2(n4618), .ZN(n6558) );
  NAND2_X1 U5088 ( .A1(n4739), .A2(n4737), .ZN(n4935) );
  NAND2_X1 U5089 ( .A1(n10068), .A2(n10069), .ZN(n10067) );
  NAND2_X1 U5090 ( .A1(n5064), .A2(n5063), .ZN(n5062) );
  OR2_X1 U5091 ( .A1(n4770), .A2(n4740), .ZN(n4739) );
  NAND2_X1 U5092 ( .A1(n10088), .A2(n10092), .ZN(n6194) );
  NAND2_X1 U5093 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5094 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  OR2_X1 U5095 ( .A1(n8907), .A2(n8908), .ZN(n8909) );
  NOR2_X1 U5096 ( .A1(n9545), .A2(n5699), .ZN(n9666) );
  OAI21_X1 U5097 ( .B1(n5678), .B2(n9642), .A(n5677), .ZN(n9545) );
  NAND2_X1 U5098 ( .A1(n10169), .A2(n8697), .ZN(n10149) );
  OAI21_X1 U5099 ( .B1(n6259), .B2(n9642), .A(n6258), .ZN(n9553) );
  AOI21_X1 U5100 ( .B1(n10175), .B2(n6072), .A(n5020), .ZN(n10155) );
  OR2_X1 U5101 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  OAI21_X1 U5102 ( .B1(n6255), .B2(n5692), .A(n8415), .ZN(n5747) );
  AOI21_X1 U5103 ( .B1(n4870), .B2(n4531), .A(n4608), .ZN(n4674) );
  XNOR2_X1 U5104 ( .A(n9506), .B(n9507), .ZN(n9467) );
  AND2_X1 U5105 ( .A1(n4906), .A2(n4616), .ZN(n4621) );
  NAND2_X1 U5106 ( .A1(n6186), .A2(n6185), .ZN(n8201) );
  NAND2_X1 U5107 ( .A1(n5028), .A2(n6058), .ZN(n10206) );
  AND2_X1 U5108 ( .A1(n8415), .A2(n5693), .ZN(n8507) );
  NAND2_X1 U5109 ( .A1(n9655), .A2(n9654), .ZN(n9653) );
  NAND2_X1 U5110 ( .A1(n4976), .A2(n4975), .ZN(n8151) );
  OR2_X1 U5111 ( .A1(n8218), .A2(n8500), .ZN(n8220) );
  INV_X1 U5112 ( .A(n8059), .ZN(n4976) );
  OAI21_X1 U5113 ( .B1(n4627), .B2(n4625), .A(n4622), .ZN(n8218) );
  AOI21_X1 U5114 ( .B1(n4992), .B2(n8208), .A(n8699), .ZN(n4990) );
  NAND2_X1 U5115 ( .A1(n6119), .A2(n6118), .ZN(n10095) );
  CLKBUF_X1 U5116 ( .A(n6190), .Z(n10142) );
  OR2_X1 U5117 ( .A1(n6190), .A2(n9886), .ZN(n8615) );
  NOR2_X1 U5118 ( .A1(n10205), .A2(n4993), .ZN(n4992) );
  OR2_X1 U5119 ( .A1(n10124), .A2(n9834), .ZN(n10102) );
  NAND2_X1 U5120 ( .A1(n4669), .A2(n4536), .ZN(n7930) );
  AOI21_X1 U5121 ( .B1(n4533), .B2(n5089), .A(n4588), .ZN(n5088) );
  NAND2_X1 U5122 ( .A1(n6063), .A2(n6062), .ZN(n10177) );
  XNOR2_X1 U5123 ( .A(n5584), .B(n5585), .ZN(n7778) );
  AND2_X1 U5124 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  INV_X1 U5125 ( .A(n8703), .ZN(n6185) );
  NAND2_X1 U5126 ( .A1(n5557), .A2(n5556), .ZN(n9652) );
  OAI21_X1 U5127 ( .B1(n5566), .B2(n5223), .A(n5222), .ZN(n5576) );
  AND2_X1 U5128 ( .A1(n8150), .A2(n9945), .ZN(n8703) );
  NAND2_X1 U5129 ( .A1(n5286), .A2(n5285), .ZN(n9634) );
  AND2_X1 U5130 ( .A1(n5537), .A2(n5536), .ZN(n9790) );
  NAND2_X1 U5131 ( .A1(n6037), .A2(n6036), .ZN(n9848) );
  NAND2_X1 U5132 ( .A1(n7307), .A2(n5396), .ZN(n7584) );
  NAND2_X1 U5133 ( .A1(n7473), .A2(n7470), .ZN(n7845) );
  AOI21_X1 U5134 ( .B1(n5054), .B2(n5052), .A(n5051), .ZN(n5050) );
  NAND2_X1 U5135 ( .A1(n5525), .A2(n5524), .ZN(n8250) );
  NAND2_X1 U5136 ( .A1(n6870), .A2(n5061), .ZN(n7227) );
  AND2_X1 U5137 ( .A1(n5497), .A2(n5496), .ZN(n9717) );
  NAND2_X1 U5138 ( .A1(n7457), .A2(n7458), .ZN(n7473) );
  NAND2_X1 U5139 ( .A1(n6024), .A2(n6023), .ZN(n10281) );
  NOR2_X1 U5140 ( .A1(n6180), .A2(n6172), .ZN(n8834) );
  AND2_X1 U5141 ( .A1(n8682), .A2(n8837), .ZN(n10430) );
  AND2_X1 U5142 ( .A1(n8655), .A2(n8663), .ZN(n8756) );
  NAND2_X1 U5143 ( .A1(n5468), .A2(n5467), .ZN(n8349) );
  NAND2_X1 U5144 ( .A1(n5999), .A2(n5998), .ZN(n10432) );
  NAND2_X1 U5145 ( .A1(n5842), .A2(n5841), .ZN(n7768) );
  NAND2_X1 U5146 ( .A1(n4918), .A2(n4917), .ZN(n7753) );
  NAND2_X1 U5147 ( .A1(n7021), .A2(n8526), .ZN(n9355) );
  AND2_X1 U5148 ( .A1(n5973), .A2(n5972), .ZN(n10494) );
  OR2_X1 U5149 ( .A1(n10578), .A2(n7552), .ZN(n7554) );
  OAI21_X1 U5150 ( .B1(n5439), .B2(n5438), .A(n5176), .ZN(n5451) );
  OAI21_X1 U5151 ( .B1(n5425), .B2(n5167), .A(n5170), .ZN(n5439) );
  INV_X2 U5152 ( .A(n6750), .ZN(n6915) );
  NAND2_X1 U5153 ( .A1(n4934), .A2(n4932), .ZN(n5409) );
  AND4_X1 U5154 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n7641)
         );
  AND4_X1 U5155 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n7134)
         );
  NAND2_X1 U5156 ( .A1(n4662), .A2(n4661), .ZN(n4934) );
  CLKBUF_X3 U5157 ( .A(n5961), .Z(n6154) );
  OAI211_X1 U5158 ( .C1(n5901), .C2(n9996), .A(n5890), .B(n5889), .ZN(n5891)
         );
  NAND4_X1 U5159 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n9726)
         );
  AND3_X1 U5160 ( .A1(n5316), .A2(n5315), .A3(n5314), .ZN(n7108) );
  NAND2_X1 U5161 ( .A1(n5670), .A2(n8448), .ZN(n9644) );
  AND2_X1 U5162 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  NAND2_X1 U5163 ( .A1(n6266), .A2(n6265), .ZN(n6268) );
  NAND2_X1 U5164 ( .A1(n6196), .A2(n6195), .ZN(n10427) );
  INV_X2 U5165 ( .A(n5913), .ZN(n8529) );
  AND3_X1 U5166 ( .A1(n5328), .A2(n5327), .A3(n5326), .ZN(n10623) );
  AND2_X1 U5167 ( .A1(n5812), .A2(n8883), .ZN(n5907) );
  AND2_X1 U5168 ( .A1(n5714), .A2(n5713), .ZN(n6965) );
  NAND2_X2 U5169 ( .A1(n5901), .A2(n4518), .ZN(n8530) );
  NAND2_X1 U5170 ( .A1(n5901), .A2(n4517), .ZN(n5913) );
  NAND2_X1 U5171 ( .A1(n6165), .A2(n6223), .ZN(n6265) );
  NAND2_X1 U5172 ( .A1(n5808), .A2(n10341), .ZN(n8883) );
  NAND2_X2 U5173 ( .A1(n8142), .A2(n6197), .ZN(n5901) );
  INV_X2 U5174 ( .A(n5336), .ZN(n8438) );
  OR2_X1 U5175 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  CLKBUF_X1 U5176 ( .A(n6968), .Z(n8513) );
  AND2_X1 U5177 ( .A1(n6239), .A2(n7957), .ZN(n6221) );
  NAND2_X1 U5178 ( .A1(n4687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U5179 ( .A1(n4765), .A2(n4762), .ZN(n8142) );
  XNOR2_X1 U5180 ( .A(n5662), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U5181 ( .A1(n6602), .A2(n4518), .ZN(n5336) );
  NAND2_X1 U5182 ( .A1(n7073), .A2(n7145), .ZN(n7291) );
  XNOR2_X1 U5183 ( .A(n5705), .B(n5263), .ZN(n8070) );
  INV_X2 U5184 ( .A(n6602), .ZN(n5554) );
  NAND2_X1 U5185 ( .A1(n10557), .A2(n7072), .ZN(n7073) );
  NOR2_X1 U5186 ( .A1(n5038), .A2(n5039), .ZN(n5037) );
  XNOR2_X1 U5187 ( .A(n5139), .B(SI_2_), .ZN(n5322) );
  NAND2_X1 U5188 ( .A1(n5661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5662) );
  OAI21_X1 U5189 ( .B1(n4516), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5138), .ZN(
        n5139) );
  XNOR2_X1 U5190 ( .A(n5273), .B(n4819), .ZN(n8897) );
  NAND2_X1 U5191 ( .A1(n10558), .A2(n10559), .ZN(n10557) );
  XNOR2_X1 U5192 ( .A(n5151), .B(SI_5_), .ZN(n5360) );
  NAND2_X1 U5193 ( .A1(n9793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  AND2_X1 U5194 ( .A1(n4511), .A2(n5781), .ZN(n6208) );
  AND2_X1 U5195 ( .A1(n5658), .A2(n5114), .ZN(n5663) );
  NAND2_X1 U5196 ( .A1(n4904), .A2(n4903), .ZN(n10559) );
  NOR2_X2 U5197 ( .A1(n4645), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U5198 ( .A1(n4640), .A2(n4639), .ZN(n4645) );
  INV_X1 U5199 ( .A(n5898), .ZN(n4684) );
  NOR2_X1 U5200 ( .A1(n5508), .A2(n5257), .ZN(n5258) );
  AND2_X1 U5201 ( .A1(n5778), .A2(n5777), .ZN(n4682) );
  NAND2_X1 U5202 ( .A1(n5931), .A2(n4675), .ZN(n5837) );
  AND3_X1 U5203 ( .A1(n5774), .A2(n5773), .A3(n6007), .ZN(n5777) );
  AND3_X1 U5204 ( .A1(n4642), .A2(n4643), .A3(n4641), .ZN(n4640) );
  AND2_X1 U5205 ( .A1(n4919), .A2(n4644), .ZN(n4639) );
  AND4_X1 U5206 ( .A1(n5772), .A2(n5771), .A3(n6019), .A4(n5770), .ZN(n5778)
         );
  NAND2_X1 U5207 ( .A1(n10347), .A2(n5128), .ZN(n5131) );
  INV_X1 U5208 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5931) );
  INV_X1 U5209 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4643) );
  INV_X1 U5210 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5779) );
  INV_X1 U5211 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4675) );
  INV_X1 U5212 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6224) );
  NOR2_X1 U5213 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5259) );
  NOR2_X1 U5214 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5261) );
  NOR2_X1 U5215 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5260) );
  INV_X1 U5216 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6160) );
  AND2_X1 U5217 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10347) );
  INV_X4 U5218 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5219 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4819) );
  INV_X1 U5220 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4919) );
  NOR2_X1 U5221 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5035) );
  INV_X4 U5222 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5223 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5774) );
  BUF_X4 U5224 ( .A(n5147), .Z(n4518) );
  AND2_X2 U5225 ( .A1(n5130), .A2(n5131), .ZN(n5147) );
  XNOR2_X2 U5226 ( .A(n9671), .B(n9366), .ZN(n8474) );
  NAND2_X2 U5227 ( .A1(n8561), .A2(n8560), .ZN(n8559) );
  AOI22_X2 U5228 ( .A1(n8238), .A2(n8237), .B1(n8236), .B2(n8235), .ZN(n8561)
         );
  AOI21_X2 U5229 ( .B1(n4658), .B2(n5117), .A(n4655), .ZN(n7594) );
  AOI211_X1 U5230 ( .C1(n7692), .C2(n5127), .A(n10502), .B(n7128), .ZN(n7690)
         );
  BUF_X4 U5231 ( .A(n5341), .Z(n4519) );
  NAND2_X1 U5232 ( .A1(n6514), .A2(n6517), .ZN(n4521) );
  NAND3_X1 U5233 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(n4524) );
  INV_X4 U5234 ( .A(n8244), .ZN(n8600) );
  AND2_X1 U5235 ( .A1(n8897), .A2(n5277), .ZN(n5339) );
  INV_X2 U5237 ( .A(n6354), .ZN(n4527) );
  INV_X1 U5238 ( .A(n4946), .ZN(n4945) );
  OAI21_X1 U5239 ( .B1(n5598), .B2(n4947), .A(n5610), .ZN(n4946) );
  INV_X1 U5240 ( .A(n8897), .ZN(n5276) );
  OAI21_X1 U5241 ( .B1(n4531), .B2(n4867), .A(n4866), .ZN(n4865) );
  NOR2_X1 U5242 ( .A1(n4570), .A2(n4871), .ZN(n4866) );
  XNOR2_X1 U5243 ( .A(n4524), .B(n6978), .ZN(n6980) );
  INV_X1 U5244 ( .A(n7531), .ZN(n4917) );
  INV_X1 U5245 ( .A(n5062), .ZN(n6563) );
  NAND2_X1 U5246 ( .A1(n4726), .A2(n8641), .ZN(n8642) );
  AND3_X1 U5247 ( .A1(n4724), .A2(n8638), .A3(n8748), .ZN(n4723) );
  AND2_X1 U5248 ( .A1(n4742), .A2(n4773), .ZN(n8662) );
  NAND2_X1 U5249 ( .A1(n4772), .A2(n4775), .ZN(n4742) );
  NOR2_X1 U5250 ( .A1(n4776), .A2(n8737), .ZN(n4774) );
  INV_X1 U5251 ( .A(n8360), .ZN(n4825) );
  NAND2_X1 U5252 ( .A1(n8670), .A2(n8669), .ZN(n8684) );
  INV_X1 U5253 ( .A(n8723), .ZN(n4794) );
  OR2_X1 U5254 ( .A1(n8418), .A2(n4832), .ZN(n8452) );
  NAND2_X1 U5255 ( .A1(n4833), .A2(n4538), .ZN(n4832) );
  NAND2_X1 U5256 ( .A1(n8452), .A2(n4830), .ZN(n8461) );
  NAND2_X1 U5257 ( .A1(n4831), .A2(n4833), .ZN(n4830) );
  INV_X1 U5258 ( .A(n8451), .ZN(n4831) );
  NAND2_X1 U5259 ( .A1(n7289), .A2(n7155), .ZN(n7156) );
  NOR2_X1 U5260 ( .A1(n4806), .A2(n8507), .ZN(n4804) );
  OR2_X1 U5261 ( .A1(n8601), .A2(n9367), .ZN(n8415) );
  OR2_X1 U5262 ( .A1(n9580), .A2(n9594), .ZN(n8397) );
  OR2_X1 U5263 ( .A1(n9634), .A2(n9647), .ZN(n8381) );
  NAND2_X1 U5264 ( .A1(n4586), .A2(n5533), .ZN(n4880) );
  OR2_X1 U5265 ( .A1(n9652), .A2(n9630), .ZN(n8371) );
  OR2_X1 U5266 ( .A1(n8261), .A2(n9645), .ZN(n8370) );
  NAND2_X1 U5267 ( .A1(n7930), .A2(n5489), .ZN(n7920) );
  INV_X1 U5268 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4641) );
  NOR2_X1 U5269 ( .A1(n5703), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5084) );
  INV_X1 U5270 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5265) );
  AND2_X1 U5271 ( .A1(n4936), .A2(n4738), .ZN(n4737) );
  AOI22_X1 U5272 ( .A1(n4542), .A2(n4767), .B1(n4937), .B2(n4530), .ZN(n4738)
         );
  INV_X1 U5273 ( .A(n8883), .ZN(n5811) );
  INV_X1 U5274 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6159) );
  AND2_X1 U5275 ( .A1(n10094), .A2(n4886), .ZN(n8533) );
  NOR2_X1 U5276 ( .A1(n4887), .A2(n10053), .ZN(n4886) );
  INV_X1 U5277 ( .A(n4888), .ZN(n4887) );
  NAND2_X1 U5278 ( .A1(n5015), .A2(n5014), .ZN(n5013) );
  INV_X1 U5279 ( .A(n5016), .ZN(n5014) );
  INV_X1 U5280 ( .A(n5001), .ZN(n4998) );
  OR2_X1 U5281 ( .A1(n10432), .A2(n9949), .ZN(n5004) );
  INV_X1 U5282 ( .A(n8660), .ZN(n8653) );
  XNOR2_X1 U5283 ( .A(n8422), .B(n8421), .ZN(n8420) );
  NOR2_X1 U5284 ( .A1(n4760), .A2(n4759), .ZN(n5781) );
  NOR2_X1 U5285 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4761) );
  AND2_X1 U5286 ( .A1(n5243), .A2(n5242), .ZN(n5610) );
  NAND2_X1 U5287 ( .A1(n5233), .A2(n5232), .ZN(n5599) );
  AOI21_X1 U5288 ( .B1(n4969), .B2(n4967), .A(n4966), .ZN(n4965) );
  NOR2_X1 U5289 ( .A1(n5398), .A2(n4933), .ZN(n4932) );
  INV_X1 U5290 ( .A(n5157), .ZN(n4933) );
  AND2_X1 U5291 ( .A1(n5072), .A2(n5074), .ZN(n5071) );
  NAND2_X1 U5292 ( .A1(n6966), .A2(n6965), .ZN(n6974) );
  NOR2_X1 U5293 ( .A1(n6980), .A2(n9725), .ZN(n6982) );
  INV_X1 U5294 ( .A(n4519), .ZN(n5638) );
  AND4_X1 U5295 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n7468)
         );
  NAND2_X1 U5296 ( .A1(n5341), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5331) );
  NOR2_X1 U5297 ( .A1(n10581), .A2(n7535), .ZN(n10580) );
  OR2_X1 U5298 ( .A1(n7987), .A2(n7986), .ZN(n7991) );
  NAND2_X1 U5299 ( .A1(n7753), .A2(n7752), .ZN(n7967) );
  NAND2_X1 U5300 ( .A1(n9491), .A2(n4853), .ZN(n4852) );
  INV_X1 U5301 ( .A(n4865), .ZN(n4864) );
  NOR2_X1 U5302 ( .A1(n4604), .A2(n4608), .ZN(n4872) );
  NAND2_X1 U5303 ( .A1(n9592), .A2(n4874), .ZN(n4870) );
  INV_X1 U5304 ( .A(n9368), .ZN(n9571) );
  INV_X1 U5305 ( .A(n9369), .ZN(n9583) );
  AOI21_X1 U5306 ( .B1(n9606), .B2(n8388), .A(n5691), .ZN(n9596) );
  NAND2_X1 U5307 ( .A1(n8220), .A2(n8370), .ZN(n9655) );
  NAND2_X1 U5308 ( .A1(n4818), .A2(n8352), .ZN(n7919) );
  INV_X1 U5309 ( .A(n9730), .ZN(n9642) );
  XNOR2_X1 U5310 ( .A(n5275), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5277) );
  INV_X1 U5311 ( .A(n5270), .ZN(n5272) );
  OR2_X1 U5312 ( .A1(n8530), .A2(n4826), .ZN(n5856) );
  AND2_X1 U5313 ( .A1(n9804), .A2(n5047), .ZN(n5046) );
  NOR2_X1 U5314 ( .A1(n9860), .A2(n9883), .ZN(n5047) );
  NAND2_X1 U5315 ( .A1(n5795), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6052) );
  INV_X1 U5316 ( .A(n6041), .ZN(n5795) );
  AND2_X1 U5317 ( .A1(n6635), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6598) );
  AND2_X1 U5318 ( .A1(n5811), .A2(n5812), .ZN(n5961) );
  AND2_X1 U5319 ( .A1(n5777), .A2(n5775), .ZN(n4683) );
  NAND2_X1 U5320 ( .A1(n4982), .A2(n7620), .ZN(n7623) );
  NAND2_X1 U5321 ( .A1(n7621), .A2(n8663), .ZN(n4982) );
  NAND2_X1 U5322 ( .A1(n6137), .A2(n6136), .ZN(n6548) );
  INV_X1 U5323 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5128) );
  NOR2_X1 U5324 ( .A1(n6560), .A2(n6559), .ZN(n5063) );
  OAI21_X1 U5325 ( .B1(n4528), .B2(n4535), .A(n4577), .ZN(n4778) );
  NOR2_X1 U5326 ( .A1(n8631), .A2(n4528), .ZN(n4780) );
  OAI21_X1 U5327 ( .B1(n8643), .B2(n4776), .A(n8651), .ZN(n4772) );
  NAND2_X1 U5328 ( .A1(n8632), .A2(n8748), .ZN(n8633) );
  NAND2_X1 U5329 ( .A1(n4779), .A2(n4777), .ZN(n8632) );
  NAND2_X1 U5330 ( .A1(n4781), .A2(n4780), .ZN(n4779) );
  INV_X1 U5331 ( .A(n4778), .ZN(n4777) );
  INV_X1 U5332 ( .A(n8650), .ZN(n4775) );
  OAI21_X1 U5333 ( .B1(n4717), .B2(n8350), .A(n4715), .ZN(n4714) );
  NAND2_X1 U5334 ( .A1(n8351), .A2(n4718), .ZN(n4715) );
  NOR2_X1 U5335 ( .A1(n8348), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U5336 ( .A1(n4712), .A2(n4711), .ZN(n4710) );
  NOR2_X1 U5337 ( .A1(n4716), .A2(n8492), .ZN(n4711) );
  OR2_X1 U5338 ( .A1(n8344), .A2(n8448), .ZN(n4712) );
  NOR2_X1 U5339 ( .A1(n8351), .A2(n4719), .ZN(n4716) );
  AOI21_X1 U5340 ( .B1(n8662), .B2(n8652), .A(n8832), .ZN(n8654) );
  AOI21_X1 U5341 ( .B1(n8361), .B2(n4823), .A(n4822), .ZN(n4821) );
  NAND2_X1 U5342 ( .A1(n8365), .A2(n8364), .ZN(n4822) );
  NOR2_X1 U5343 ( .A1(n4825), .A2(n4824), .ZN(n4823) );
  NAND2_X1 U5344 ( .A1(n4699), .A2(n4698), .ZN(n4697) );
  AOI21_X1 U5345 ( .B1(n4704), .B2(n8381), .A(n4702), .ZN(n4698) );
  NAND2_X1 U5346 ( .A1(n4558), .A2(n8381), .ZN(n4699) );
  NAND2_X1 U5347 ( .A1(n4703), .A2(n4701), .ZN(n4700) );
  NOR2_X1 U5348 ( .A1(n4704), .A2(n4702), .ZN(n4701) );
  INV_X1 U5349 ( .A(n4820), .ZN(n4703) );
  NAND2_X1 U5350 ( .A1(n8678), .A2(n8677), .ZN(n8681) );
  OAI21_X1 U5351 ( .B1(n4835), .B2(n4834), .A(n8393), .ZN(n8403) );
  NOR2_X1 U5352 ( .A1(n8386), .A2(n8453), .ZN(n4835) );
  OAI21_X1 U5353 ( .B1(n8387), .B2(n8448), .A(n8476), .ZN(n4834) );
  OR2_X1 U5354 ( .A1(n4567), .A2(n4734), .ZN(n4731) );
  OAI21_X1 U5355 ( .B1(n8721), .B2(n8789), .A(n4794), .ZN(n4784) );
  AND2_X1 U5356 ( .A1(n4792), .A2(n8710), .ZN(n4730) );
  NOR2_X1 U5357 ( .A1(n4732), .A2(n4728), .ZN(n4727) );
  AND2_X1 U5358 ( .A1(n4792), .A2(n4733), .ZN(n4732) );
  INV_X1 U5359 ( .A(n8716), .ZN(n4733) );
  NAND2_X1 U5360 ( .A1(n4791), .A2(n4785), .ZN(n4789) );
  OAI211_X1 U5361 ( .C1(n4791), .C2(n4790), .A(n4782), .B(n4785), .ZN(n4788)
         );
  NAND2_X1 U5362 ( .A1(n4792), .A2(n8789), .ZN(n4782) );
  OR2_X1 U5363 ( .A1(n9842), .A2(n5060), .ZN(n5059) );
  INV_X1 U5364 ( .A(n6426), .ZN(n5060) );
  NAND2_X1 U5365 ( .A1(n4771), .A2(n8739), .ZN(n4770) );
  AND2_X1 U5366 ( .A1(n5775), .A2(n5818), .ZN(n4681) );
  INV_X1 U5367 ( .A(SI_17_), .ZN(n5198) );
  OR2_X1 U5368 ( .A1(n9353), .A2(n5111), .ZN(n5110) );
  NOR2_X1 U5369 ( .A1(n5105), .A2(n9353), .ZN(n5104) );
  INV_X1 U5370 ( .A(n5107), .ZN(n5105) );
  INV_X1 U5371 ( .A(n9353), .ZN(n5102) );
  INV_X1 U5372 ( .A(n4924), .ZN(n4923) );
  OAI21_X1 U5373 ( .B1(n7291), .B2(n4925), .A(n7166), .ZN(n4924) );
  NAND2_X1 U5374 ( .A1(n9407), .A2(n9406), .ZN(n9411) );
  AND2_X1 U5375 ( .A1(n8389), .A2(n8388), .ZN(n8476) );
  OR2_X1 U5376 ( .A1(n8936), .A2(n9631), .ZN(n8384) );
  AND2_X1 U5377 ( .A1(n4878), .A2(n4667), .ZN(n4666) );
  INV_X1 U5378 ( .A(n9654), .ZN(n4667) );
  INV_X1 U5379 ( .A(n8345), .ZN(n4651) );
  NAND2_X1 U5380 ( .A1(n4673), .A2(n4564), .ZN(n8321) );
  NAND2_X1 U5381 ( .A1(n5304), .A2(n5303), .ZN(n8302) );
  AND2_X1 U5382 ( .A1(n7305), .A2(n5384), .ZN(n4875) );
  OR2_X1 U5383 ( .A1(n6584), .A2(n6577), .ZN(n6953) );
  INV_X1 U5384 ( .A(n9938), .ZN(n6500) );
  INV_X1 U5385 ( .A(n4988), .ZN(n4987) );
  OAI21_X1 U5386 ( .B1(n10069), .B2(n8794), .A(n8799), .ZN(n4988) );
  NAND2_X1 U5387 ( .A1(n10304), .A2(n6500), .ZN(n5018) );
  NOR2_X1 U5388 ( .A1(n10142), .A2(n10159), .ZN(n4882) );
  AND2_X1 U5389 ( .A1(n5000), .A2(n6033), .ZN(n4999) );
  NOR2_X1 U5390 ( .A1(n4898), .A2(n10432), .ZN(n4897) );
  INV_X1 U5391 ( .A(n4899), .ZN(n4898) );
  INV_X1 U5392 ( .A(n5987), .ZN(n5793) );
  INV_X1 U5393 ( .A(n8756), .ZN(n5994) );
  OR2_X1 U5394 ( .A1(n10442), .A2(n7641), .ZN(n8749) );
  NAND2_X1 U5395 ( .A1(n4529), .A2(n4892), .ZN(n4891) );
  NOR2_X1 U5396 ( .A1(n8624), .A2(n8623), .ZN(n8631) );
  AND2_X1 U5397 ( .A1(n6523), .A2(n6522), .ZN(n7409) );
  XNOR2_X1 U5398 ( .A(n6277), .B(n9963), .ZN(n7480) );
  OR2_X1 U5399 ( .A1(n7873), .A2(n10281), .ZN(n5126) );
  NOR2_X1 U5400 ( .A1(n7491), .A2(n5879), .ZN(n6901) );
  NAND2_X1 U5401 ( .A1(n5753), .A2(n5752), .ZN(n8422) );
  NOR2_X1 U5402 ( .A1(n4539), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U5403 ( .A1(n4943), .A2(n4941), .ZN(n5625) );
  AOI21_X1 U5404 ( .B1(n4945), .B2(n4947), .A(n4942), .ZN(n4941) );
  INV_X1 U5405 ( .A(n5243), .ZN(n4942) );
  AND2_X1 U5406 ( .A1(n5546), .A2(n5211), .ZN(n5212) );
  NAND2_X1 U5407 ( .A1(n4957), .A2(n5191), .ZN(n4956) );
  INV_X1 U5408 ( .A(n5506), .ZN(n4957) );
  INV_X1 U5409 ( .A(n4955), .ZN(n4954) );
  OAI21_X1 U5410 ( .B1(n4958), .B2(n4956), .A(n5197), .ZN(n4955) );
  NOR2_X1 U5411 ( .A1(n5192), .A2(n4959), .ZN(n4958) );
  INV_X1 U5412 ( .A(n5188), .ZN(n4959) );
  INV_X1 U5413 ( .A(n5490), .ZN(n5192) );
  AOI21_X1 U5414 ( .B1(n4929), .B2(n5155), .A(n5391), .ZN(n4661) );
  NAND2_X1 U5415 ( .A1(n5150), .A2(n4930), .ZN(n4663) );
  AOI22_X1 U5416 ( .A1(n8549), .A2(n5093), .B1(n4590), .B2(n5094), .ZN(n5092)
         );
  INV_X1 U5417 ( .A(n8242), .ZN(n5093) );
  AOI21_X1 U5418 ( .B1(n5078), .B2(n4574), .A(n5075), .ZN(n5074) );
  INV_X1 U5419 ( .A(n8015), .ZN(n5075) );
  NAND2_X1 U5420 ( .A1(n5080), .A2(n5079), .ZN(n8582) );
  AOI21_X1 U5421 ( .B1(n5081), .B2(n5083), .A(n4561), .ZN(n5079) );
  INV_X1 U5422 ( .A(n4551), .ZN(n5089) );
  AND2_X1 U5423 ( .A1(n8940), .A2(n5108), .ZN(n5107) );
  OR2_X1 U5424 ( .A1(n9315), .A2(n5109), .ZN(n5108) );
  INV_X1 U5425 ( .A(n8594), .ZN(n5109) );
  AND2_X1 U5426 ( .A1(n8470), .A2(n8513), .ZN(n4817) );
  OR2_X1 U5427 ( .A1(n9746), .A2(n9665), .ZN(n8469) );
  AND2_X1 U5428 ( .A1(n8515), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U5429 ( .A1(n4587), .A2(n8513), .ZN(n4816) );
  OAI21_X1 U5430 ( .B1(n4721), .B2(n8454), .A(n8465), .ZN(n4720) );
  INV_X1 U5431 ( .A(n8464), .ZN(n8465) );
  OAI21_X1 U5432 ( .B1(n8458), .B2(n8457), .A(n4722), .ZN(n4721) );
  OAI21_X1 U5433 ( .B1(n5085), .B2(n4746), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5266) );
  NAND2_X1 U5434 ( .A1(n4745), .A2(n5362), .ZN(n4746) );
  AND2_X1 U5435 ( .A1(n5249), .A2(n5248), .ZN(n4745) );
  AND2_X1 U5436 ( .A1(n4748), .A2(n4747), .ZN(n7053) );
  NAND2_X1 U5437 ( .A1(n7050), .A2(n7071), .ZN(n4747) );
  INV_X1 U5438 ( .A(n10560), .ZN(n4748) );
  NAND2_X1 U5439 ( .A1(n7053), .A2(n7052), .ZN(n7144) );
  NAND2_X1 U5440 ( .A1(n7074), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7292) );
  OR2_X1 U5441 ( .A1(n7156), .A2(n7279), .ZN(n7157) );
  NAND2_X1 U5442 ( .A1(n7554), .A2(n7553), .ZN(n7738) );
  INV_X1 U5443 ( .A(n7555), .ZN(n7553) );
  XNOR2_X1 U5444 ( .A(n7967), .B(n7977), .ZN(n7754) );
  OR2_X1 U5445 ( .A1(n5426), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U5446 ( .A1(n7991), .A2(n7990), .ZN(n8118) );
  NOR2_X1 U5447 ( .A1(n7577), .A2(n7754), .ZN(n7969) );
  OR2_X1 U5448 ( .A1(n8171), .A2(n8170), .ZN(n9407) );
  XNOR2_X1 U5449 ( .A(n9411), .B(n9410), .ZN(n10601) );
  NAND2_X1 U5450 ( .A1(n9458), .A2(n4907), .ZN(n4906) );
  INV_X1 U5451 ( .A(n9459), .ZN(n4907) );
  OR2_X1 U5452 ( .A1(n9423), .A2(n4908), .ZN(n4905) );
  OR2_X1 U5453 ( .A1(n9459), .A2(n9424), .ZN(n4908) );
  NOR2_X1 U5454 ( .A1(n10597), .A2(n10404), .ZN(n4757) );
  AOI21_X1 U5455 ( .B1(n9490), .B2(n4855), .A(n9517), .ZN(n4854) );
  AOI21_X1 U5456 ( .B1(n4804), .B2(n4801), .A(n4589), .ZN(n4800) );
  INV_X1 U5457 ( .A(n4556), .ZN(n4801) );
  INV_X1 U5458 ( .A(n4804), .ZN(n4802) );
  INV_X1 U5459 ( .A(n4870), .ZN(n4863) );
  OR2_X1 U5460 ( .A1(n8410), .A2(n8411), .ZN(n9563) );
  OR2_X1 U5461 ( .A1(n9572), .A2(n9583), .ZN(n8404) );
  NAND2_X1 U5462 ( .A1(n4874), .A2(n5597), .ZN(n4869) );
  AND2_X1 U5463 ( .A1(n8399), .A2(n8404), .ZN(n9575) );
  NAND2_X1 U5464 ( .A1(n8920), .A2(n9371), .ZN(n4874) );
  AOI22_X1 U5465 ( .A1(n9614), .A2(n9619), .B1(n9631), .B2(n9777), .ZN(n9602)
         );
  OAI21_X1 U5466 ( .B1(n9618), .B2(n8375), .A(n8384), .ZN(n9606) );
  AND3_X1 U5467 ( .A1(n5291), .A2(n5290), .A3(n5289), .ZN(n9647) );
  INV_X1 U5468 ( .A(n4879), .ZN(n4878) );
  OAI22_X1 U5469 ( .A1(n8498), .A2(n4880), .B1(n9376), .B2(n8261), .ZN(n4879)
         );
  OR2_X1 U5470 ( .A1(n8084), .A2(n4880), .ZN(n4668) );
  AND2_X1 U5471 ( .A1(n4668), .A2(n4666), .ZN(n9641) );
  AND2_X1 U5472 ( .A1(n8371), .A2(n8379), .ZN(n9654) );
  AOI21_X1 U5473 ( .B1(n4632), .B2(n4630), .A(n4629), .ZN(n4628) );
  INV_X1 U5474 ( .A(n8358), .ZN(n4630) );
  INV_X1 U5475 ( .A(n8363), .ZN(n4629) );
  INV_X1 U5476 ( .A(n7919), .ZN(n4627) );
  NAND2_X1 U5477 ( .A1(n7656), .A2(n8492), .ZN(n4876) );
  AND4_X1 U5478 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n8236)
         );
  NAND2_X1 U5479 ( .A1(n7596), .A2(n5686), .ZN(n7654) );
  AND4_X1 U5480 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n7892)
         );
  NAND2_X1 U5481 ( .A1(n7498), .A2(n8485), .ZN(n5683) );
  NAND2_X1 U5482 ( .A1(n7009), .A2(n8302), .ZN(n7086) );
  OR2_X1 U5483 ( .A1(n10623), .A2(n9387), .ZN(n8292) );
  AND2_X1 U5484 ( .A1(n5395), .A2(n5394), .ZN(n7331) );
  AND2_X1 U5485 ( .A1(n5382), .A2(n5381), .ZN(n7316) );
  AND3_X1 U5486 ( .A1(n5366), .A2(n5365), .A3(n5364), .ZN(n7320) );
  NAND2_X1 U5487 ( .A1(n5667), .A2(n5666), .ZN(n9730) );
  AND2_X1 U5488 ( .A1(n6965), .A2(n5715), .ZN(n5719) );
  INV_X1 U5489 ( .A(n5085), .ZN(n4813) );
  XNOR2_X1 U5490 ( .A(n5665), .B(n5664), .ZN(n6967) );
  OR2_X1 U5491 ( .A1(n5663), .A2(n9792), .ZN(n5665) );
  OR2_X1 U5492 ( .A1(n5428), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5452) );
  XNOR2_X1 U5493 ( .A(n6280), .B(n4514), .ZN(n6281) );
  AND2_X1 U5494 ( .A1(n6270), .A2(n6269), .ZN(n6282) );
  INV_X1 U5495 ( .A(n9860), .ZN(n5044) );
  OR2_X1 U5496 ( .A1(n6039), .A2(n6038), .ZN(n6041) );
  NOR2_X1 U5497 ( .A1(n9860), .A2(n9861), .ZN(n5045) );
  NAND2_X1 U5498 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U5499 ( .A1(n6370), .A2(n6369), .ZN(n5055) );
  NAND2_X1 U5500 ( .A1(n6075), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U5501 ( .A(n6299), .B(n4514), .ZN(n6305) );
  AND2_X1 U5502 ( .A1(n6127), .A2(n6126), .ZN(n9835) );
  AND2_X1 U5503 ( .A1(n6057), .A2(n6056), .ZN(n9815) );
  INV_X1 U5504 ( .A(n6154), .ZN(n6111) );
  NAND2_X1 U5505 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(n5042), .ZN(n5041) );
  NAND2_X1 U5506 ( .A1(n5801), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5040) );
  AND2_X1 U5507 ( .A1(n6158), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U5508 ( .A1(n6160), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5043) );
  OAI21_X1 U5509 ( .B1(n8732), .B2(n4987), .A(n4985), .ZN(n4984) );
  OAI21_X1 U5510 ( .B1(n8732), .B2(n8735), .A(n4987), .ZN(n4985) );
  OR2_X1 U5511 ( .A1(n8807), .A2(n8893), .ZN(n9887) );
  AND2_X1 U5512 ( .A1(n10049), .A2(n6142), .ZN(n10059) );
  AND2_X1 U5513 ( .A1(n5018), .A2(n6106), .ZN(n5016) );
  OR2_X1 U5514 ( .A1(n6109), .A2(n9836), .ZN(n6120) );
  NOR2_X1 U5515 ( .A1(n10177), .A2(n5021), .ZN(n5020) );
  NAND2_X1 U5516 ( .A1(n6061), .A2(n5025), .ZN(n10188) );
  OR2_X1 U5517 ( .A1(n10208), .A2(n6059), .ZN(n5025) );
  NAND2_X1 U5518 ( .A1(n8151), .A2(n6184), .ZN(n6186) );
  OR2_X1 U5519 ( .A1(n8201), .A2(n8208), .ZN(n8203) );
  AND2_X1 U5520 ( .A1(n10275), .A2(n9945), .ZN(n5029) );
  NAND2_X1 U5521 ( .A1(n8150), .A2(n8205), .ZN(n5030) );
  INV_X1 U5522 ( .A(n8144), .ZN(n5031) );
  AND2_X1 U5523 ( .A1(n4554), .A2(n5004), .ZN(n5000) );
  NAND2_X1 U5524 ( .A1(n5002), .A2(n4554), .ZN(n5001) );
  INV_X1 U5525 ( .A(n5003), .ZN(n5002) );
  AOI21_X1 U5526 ( .B1(n10430), .B2(n5004), .A(n4582), .ZN(n5003) );
  INV_X1 U5527 ( .A(n8758), .ZN(n7620) );
  NAND2_X1 U5528 ( .A1(n7602), .A2(n7603), .ZN(n5027) );
  NAND2_X1 U5529 ( .A1(n7604), .A2(n8653), .ZN(n4617) );
  NAND2_X1 U5530 ( .A1(n7247), .A2(n5943), .ZN(n5009) );
  INV_X1 U5531 ( .A(n10427), .ZN(n10203) );
  NAND2_X1 U5532 ( .A1(n6051), .A2(n6050), .ZN(n8212) );
  NAND2_X1 U5533 ( .A1(n6627), .A2(n8529), .ZN(n4989) );
  AND2_X1 U5534 ( .A1(n6240), .A2(n10336), .ZN(n7407) );
  AND3_X1 U5535 ( .A1(n6521), .A2(n6236), .A3(n6522), .ZN(n6250) );
  NAND2_X1 U5536 ( .A1(n6265), .A2(n8742), .ZN(n7436) );
  XNOR2_X1 U5537 ( .A(n5810), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U5538 ( .A1(n5809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5810) );
  XNOR2_X1 U5539 ( .A(n5749), .B(n5748), .ZN(n8190) );
  INV_X1 U5540 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5541 ( .A1(n4511), .A2(n5033), .ZN(n5786) );
  NOR2_X1 U5542 ( .A1(n5787), .A2(n4766), .ZN(n4763) );
  NAND2_X1 U5543 ( .A1(n4944), .A2(n5238), .ZN(n5611) );
  OR2_X1 U5544 ( .A1(n6208), .A2(n6214), .ZN(n6215) );
  NOR2_X1 U5545 ( .A1(n5575), .A2(n4972), .ZN(n4971) );
  INV_X1 U5546 ( .A(n5222), .ZN(n4972) );
  AND2_X1 U5547 ( .A1(n5232), .A2(n5231), .ZN(n5585) );
  AOI21_X1 U5548 ( .B1(n4971), .B2(n5223), .A(n4970), .ZN(n4969) );
  INV_X1 U5549 ( .A(n5227), .ZN(n4970) );
  XNOR2_X1 U5550 ( .A(n6225), .B(n6224), .ZN(n6635) );
  NAND2_X1 U5551 ( .A1(n6223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6225) );
  AND2_X1 U5552 ( .A1(n5609), .A2(n5608), .ZN(n9594) );
  AND3_X1 U5553 ( .A1(n5543), .A2(n5542), .A3(n5541), .ZN(n9645) );
  NOR2_X1 U5554 ( .A1(n6982), .A2(n6981), .ZN(n7024) );
  NAND2_X1 U5555 ( .A1(n5601), .A2(n5600), .ZN(n9580) );
  AND3_X1 U5556 ( .A1(n5563), .A2(n5562), .A3(n5561), .ZN(n9630) );
  NAND2_X1 U5557 ( .A1(n5578), .A2(n5577), .ZN(n9607) );
  AND4_X1 U5558 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n8259)
         );
  NAND2_X1 U5559 ( .A1(n5282), .A2(n5281), .ZN(n9368) );
  NAND2_X1 U5560 ( .A1(n5622), .A2(n5621), .ZN(n9369) );
  AND4_X1 U5561 ( .A1(n5519), .A2(n5518), .A3(n5517), .A4(n5516), .ZN(n8563)
         );
  OR2_X1 U5562 ( .A1(n7057), .A2(n6600), .ZN(n9500) );
  NAND2_X1 U5563 ( .A1(n10573), .A2(n10572), .ZN(n10571) );
  NAND2_X1 U5564 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  NOR2_X1 U5565 ( .A1(n7263), .A2(n4749), .ZN(n7151) );
  NOR2_X1 U5566 ( .A1(n4750), .A2(n7148), .ZN(n4749) );
  INV_X1 U5567 ( .A(n7149), .ZN(n4750) );
  NAND2_X1 U5568 ( .A1(n7151), .A2(n7150), .ZN(n7539) );
  NAND2_X1 U5569 ( .A1(n10591), .A2(n10592), .ZN(n10590) );
  OR2_X1 U5570 ( .A1(n10580), .A2(n7529), .ZN(n4918) );
  XNOR2_X1 U5571 ( .A(n5399), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7751) );
  NOR2_X1 U5572 ( .A1(n7740), .A2(n7739), .ZN(n7986) );
  OR2_X1 U5573 ( .A1(n7975), .A2(n7974), .ZN(n8132) );
  OR2_X1 U5574 ( .A1(n9423), .A2(n9424), .ZN(n4911) );
  AND2_X1 U5575 ( .A1(P2_U3893), .A2(n5668), .ZN(n10612) );
  XOR2_X1 U5576 ( .A(n9455), .B(n9446), .Z(n9423) );
  INV_X1 U5577 ( .A(n10566), .ZN(n10615) );
  NAND2_X1 U5578 ( .A1(n5755), .A2(n5754), .ZN(n8904) );
  INV_X1 U5579 ( .A(n9671), .ZN(n9548) );
  NOR2_X1 U5580 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  NAND2_X1 U5581 ( .A1(n9744), .A2(n9739), .ZN(n9715) );
  OR2_X1 U5582 ( .A1(n9904), .A2(n9905), .ZN(n5065) );
  OR2_X1 U5583 ( .A1(n8813), .A2(n6166), .ZN(n8814) );
  INV_X1 U5584 ( .A(n6532), .ZN(n8871) );
  AND4_X1 U5585 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n9950)
         );
  NAND2_X1 U5586 ( .A1(n8534), .A2(n10435), .ZN(n8884) );
  OR2_X1 U5587 ( .A1(n6529), .A2(n8875), .ZN(n10190) );
  NAND2_X1 U5588 ( .A1(n6149), .A2(n6148), .ZN(n10053) );
  NAND2_X1 U5589 ( .A1(n8884), .A2(n10216), .ZN(n10287) );
  INV_X1 U5590 ( .A(n10063), .ZN(n4619) );
  NAND2_X1 U5591 ( .A1(n10058), .A2(n10520), .ZN(n4620) );
  NAND2_X1 U5592 ( .A1(n10523), .A2(n10282), .ZN(n10329) );
  INV_X1 U5593 ( .A(n5807), .ZN(n10341) );
  XNOR2_X1 U5594 ( .A(n8437), .B(n8436), .ZN(n10344) );
  OAI21_X1 U5595 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8437) );
  INV_X1 U5596 ( .A(n8640), .ZN(n4781) );
  AND3_X1 U5597 ( .A1(n4707), .A2(n8321), .A3(n4705), .ZN(n8329) );
  NAND2_X1 U5598 ( .A1(n4706), .A2(n8453), .ZN(n4705) );
  OR2_X1 U5599 ( .A1(n8320), .A2(n8453), .ZN(n4707) );
  NAND2_X1 U5600 ( .A1(n8326), .A2(n8325), .ZN(n4706) );
  INV_X1 U5601 ( .A(n5942), .ZN(n4776) );
  INV_X1 U5602 ( .A(n8496), .ZN(n4824) );
  NAND2_X1 U5603 ( .A1(n4541), .A2(n4713), .ZN(n4708) );
  NAND2_X1 U5604 ( .A1(n4710), .A2(n4713), .ZN(n4709) );
  INV_X1 U5605 ( .A(n4714), .ZN(n4713) );
  OAI21_X1 U5606 ( .B1(n4821), .B2(n4700), .A(n4697), .ZN(n4696) );
  OAI21_X1 U5607 ( .B1(n8704), .B2(n8703), .A(n8850), .ZN(n4744) );
  NAND2_X1 U5608 ( .A1(n8403), .A2(n8475), .ZN(n8395) );
  AOI21_X1 U5609 ( .B1(n4585), .B2(n4791), .A(n4784), .ZN(n4783) );
  NAND2_X1 U5610 ( .A1(n4731), .A2(n8716), .ZN(n8717) );
  NAND2_X1 U5611 ( .A1(n8711), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U5612 ( .A1(n8738), .A2(n8737), .ZN(n4769) );
  INV_X1 U5613 ( .A(n4872), .ZN(n4867) );
  NOR2_X1 U5614 ( .A1(n4939), .A2(n4768), .ZN(n4767) );
  NOR2_X1 U5615 ( .A1(n10043), .A2(n8737), .ZN(n4768) );
  NAND2_X1 U5616 ( .A1(n4940), .A2(n9933), .ZN(n4939) );
  AND2_X1 U5617 ( .A1(n8740), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U5618 ( .A1(n10043), .A2(n8737), .ZN(n4938) );
  NOR2_X1 U5619 ( .A1(n4767), .A2(n4937), .ZN(n4740) );
  INV_X1 U5620 ( .A(n5238), .ZN(n4947) );
  NOR2_X1 U5621 ( .A1(n4968), .A2(n4963), .ZN(n4962) );
  INV_X1 U5622 ( .A(n5218), .ZN(n4963) );
  INV_X1 U5623 ( .A(n4969), .ZN(n4968) );
  INV_X1 U5624 ( .A(n4971), .ZN(n4967) );
  INV_X1 U5625 ( .A(n5585), .ZN(n4966) );
  AOI21_X1 U5626 ( .B1(n4954), .B2(n4956), .A(n4952), .ZN(n4951) );
  INV_X1 U5627 ( .A(n5520), .ZN(n4952) );
  NAND2_X1 U5628 ( .A1(n4954), .A2(n5476), .ZN(n4949) );
  INV_X1 U5629 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6007) );
  AND2_X1 U5630 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  INV_X1 U5631 ( .A(SI_20_), .ZN(n8947) );
  INV_X1 U5632 ( .A(SI_14_), .ZN(n9262) );
  INV_X1 U5633 ( .A(n7844), .ZN(n5076) );
  INV_X1 U5634 ( .A(n5082), .ZN(n5081) );
  OAI21_X1 U5635 ( .B1(n8575), .B2(n5083), .A(n8931), .ZN(n5082) );
  INV_X1 U5636 ( .A(n8579), .ZN(n5083) );
  NOR2_X1 U5637 ( .A1(n8452), .A2(n8451), .ZN(n8456) );
  AOI21_X1 U5638 ( .B1(n8456), .B2(n8455), .A(n8473), .ZN(n4722) );
  AOI21_X1 U5639 ( .B1(n4829), .B2(n4828), .A(n8463), .ZN(n8464) );
  NOR2_X1 U5640 ( .A1(n8459), .A2(n8460), .ZN(n4828) );
  NAND2_X1 U5641 ( .A1(n8461), .A2(n9548), .ZN(n4829) );
  XNOR2_X1 U5642 ( .A(n7049), .B(n4751), .ZN(n10544) );
  NOR2_X1 U5643 ( .A1(n10544), .A2(n10543), .ZN(n10542) );
  INV_X1 U5644 ( .A(n5324), .ZN(n7061) );
  NAND2_X1 U5645 ( .A1(n7290), .A2(n7279), .ZN(n4921) );
  NAND2_X1 U5646 ( .A1(n7976), .A2(n4603), .ZN(n8122) );
  INV_X1 U5647 ( .A(n8164), .ZN(n4845) );
  XNOR2_X1 U5648 ( .A(n9390), .B(n9409), .ZN(n10604) );
  OR2_X1 U5649 ( .A1(n8904), .A2(n8607), .ZN(n8467) );
  NOR2_X1 U5650 ( .A1(n4867), .A2(n4861), .ZN(n4860) );
  INV_X1 U5651 ( .A(n4874), .ZN(n4861) );
  INV_X1 U5652 ( .A(n8404), .ZN(n4809) );
  OR2_X1 U5653 ( .A1(n8920), .A2(n9604), .ZN(n8475) );
  AND2_X1 U5654 ( .A1(n5559), .A2(n5287), .ZN(n5570) );
  INV_X1 U5655 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U5656 ( .A1(n5527), .A2(n5526), .ZN(n5540) );
  AND2_X1 U5657 ( .A1(n5514), .A2(n9192), .ZN(n5527) );
  NOR2_X1 U5658 ( .A1(n5456), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5470) );
  OR2_X1 U5659 ( .A1(n5443), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U5660 ( .A1(n7579), .A2(n7843), .ZN(n8326) );
  NAND2_X1 U5661 ( .A1(n8266), .A2(n7468), .ZN(n8325) );
  NOR2_X1 U5662 ( .A1(n6645), .A2(n5734), .ZN(n6577) );
  NAND2_X1 U5663 ( .A1(n8285), .A2(n4637), .ZN(n9732) );
  NAND2_X1 U5664 ( .A1(n4638), .A2(n8280), .ZN(n4637) );
  INV_X1 U5665 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5737) );
  INV_X1 U5666 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5255) );
  INV_X1 U5667 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5254) );
  NOR2_X1 U5668 ( .A1(n5452), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U5669 ( .A1(n5057), .A2(n5056), .ZN(n6450) );
  AOI21_X1 U5670 ( .B1(n4534), .B2(n5060), .A(n4579), .ZN(n5056) );
  INV_X1 U5671 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5772) );
  INV_X1 U5672 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5770) );
  AND2_X1 U5673 ( .A1(n5776), .A2(n5769), .ZN(n5066) );
  NOR2_X1 U5674 ( .A1(n10080), .A2(n6548), .ZN(n4888) );
  AND2_X1 U5675 ( .A1(n10296), .A2(n9936), .ZN(n8785) );
  INV_X1 U5676 ( .A(n8700), .ZN(n8712) );
  NOR2_X1 U5677 ( .A1(n10275), .A2(n8212), .ZN(n4885) );
  INV_X1 U5678 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U5679 ( .A1(n5794), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6039) );
  NOR2_X1 U5680 ( .A1(n4981), .A2(n4979), .ZN(n4978) );
  INV_X1 U5681 ( .A(n8663), .ZN(n4979) );
  INV_X1 U5682 ( .A(n8838), .ZN(n4981) );
  NAND2_X1 U5683 ( .A1(n8758), .A2(n8838), .ZN(n4980) );
  NOR2_X1 U5684 ( .A1(n6001), .A2(n7190), .ZN(n6000) );
  NOR2_X1 U5685 ( .A1(n7916), .A2(n7768), .ZN(n4899) );
  AND2_X1 U5686 ( .A1(n6174), .A2(n8824), .ZN(n8744) );
  INV_X1 U5687 ( .A(n10334), .ZN(n6238) );
  AND2_X1 U5688 ( .A1(n5644), .A2(n5630), .ZN(n5642) );
  AND2_X1 U5689 ( .A1(n5626), .A2(n5247), .ZN(n5624) );
  AND2_X1 U5690 ( .A1(n5238), .A2(n5237), .ZN(n5598) );
  NAND2_X1 U5691 ( .A1(n4685), .A2(n4576), .ZN(n4687) );
  AOI21_X1 U5692 ( .B1(n5409), .B2(n5166), .A(n5165), .ZN(n5425) );
  INV_X1 U5693 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5769) );
  OAI21_X1 U5694 ( .B1(n4518), .B2(n4826), .A(n4736), .ZN(n5135) );
  NAND2_X1 U5695 ( .A1(n4518), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4736) );
  XNOR2_X1 U5696 ( .A(n5135), .B(n4735), .ZN(n5134) );
  INV_X1 U5697 ( .A(SI_1_), .ZN(n4735) );
  INV_X1 U5698 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5129) );
  NAND2_X1 U5699 ( .A1(n5103), .A2(n5100), .ZN(n8907) );
  AND2_X1 U5700 ( .A1(n4610), .A2(n5101), .ZN(n5100) );
  OR2_X1 U5701 ( .A1(n5617), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U5702 ( .A1(n7845), .A2(n7844), .ZN(n8010) );
  XNOR2_X1 U5703 ( .A(n7108), .B(n4512), .ZN(n6997) );
  OAI21_X1 U5704 ( .B1(n5096), .B2(n7318), .A(n5095), .ZN(n9304) );
  NOR2_X1 U5705 ( .A1(n5097), .A2(n7001), .ZN(n5096) );
  INV_X1 U5706 ( .A(n6998), .ZN(n5097) );
  NAND2_X1 U5707 ( .A1(n8576), .A2(n8575), .ZN(n9321) );
  NOR2_X1 U5708 ( .A1(n5498), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U5709 ( .A1(n4813), .A2(n4812), .ZN(n5270) );
  AND2_X1 U5710 ( .A1(n5086), .A2(n4560), .ZN(n4812) );
  NAND2_X1 U5711 ( .A1(n4525), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U5712 ( .A1(n4920), .A2(n4919), .ZN(n5324) );
  NAND2_X1 U5713 ( .A1(n10570), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5714 ( .A1(n7292), .A2(n7291), .ZN(n4922) );
  NAND2_X1 U5715 ( .A1(n7144), .A2(n4563), .ZN(n7281) );
  NOR2_X1 U5716 ( .A1(n7281), .A2(n7282), .ZN(n7280) );
  OR2_X1 U5717 ( .A1(n7269), .A2(n7268), .ZN(n4857) );
  OR2_X1 U5718 ( .A1(n7160), .A2(n7268), .ZN(n4856) );
  NOR2_X1 U5719 ( .A1(n5377), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U5720 ( .A1(n7743), .A2(n7744), .ZN(n7745) );
  NAND2_X1 U5721 ( .A1(n7745), .A2(n7746), .ZN(n7976) );
  XNOR2_X1 U5722 ( .A(n8122), .B(n8121), .ZN(n7979) );
  XNOR2_X1 U5723 ( .A(n8165), .B(n8133), .ZN(n8134) );
  NOR2_X1 U5724 ( .A1(n8134), .A2(n8135), .ZN(n8167) );
  NOR2_X1 U5725 ( .A1(n9412), .A2(n10600), .ZN(n9415) );
  INV_X1 U5726 ( .A(n9411), .ZN(n9408) );
  AOI21_X1 U5727 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9433), .A(n9422), .ZN(
        n9455) );
  INV_X1 U5728 ( .A(n9522), .ZN(n4853) );
  NAND2_X1 U5729 ( .A1(n9508), .A2(n4914), .ZN(n4913) );
  INV_X1 U5730 ( .A(n9510), .ZN(n4914) );
  AOI21_X1 U5731 ( .B1(n4799), .B2(n4798), .A(n4797), .ZN(n8468) );
  NOR2_X1 U5732 ( .A1(n4802), .A2(n8604), .ZN(n4798) );
  OAI21_X1 U5733 ( .B1(n4800), .B2(n8604), .A(n4584), .ZN(n4797) );
  NOR2_X1 U5734 ( .A1(n9562), .A2(n9644), .ZN(n5676) );
  NAND2_X1 U5735 ( .A1(n4807), .A2(n8409), .ZN(n4806) );
  OR2_X1 U5736 ( .A1(n8410), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U5737 ( .A1(n8396), .A2(n8404), .ZN(n4808) );
  OR2_X1 U5738 ( .A1(n5588), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5602) );
  NOR2_X1 U5739 ( .A1(n5602), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5615) );
  NOR2_X1 U5740 ( .A1(n9633), .A2(n5690), .ZN(n9618) );
  AOI21_X1 U5741 ( .B1(n9621), .B2(n4523), .A(n5574), .ZN(n9631) );
  AOI21_X1 U5742 ( .B1(n8084), .B2(n4666), .A(n4664), .ZN(n9627) );
  INV_X1 U5743 ( .A(n4665), .ZN(n4664) );
  AOI21_X1 U5744 ( .B1(n4666), .B2(n4880), .A(n5564), .ZN(n4665) );
  NAND2_X1 U5745 ( .A1(n9627), .A2(n9632), .ZN(n9626) );
  NAND2_X1 U5746 ( .A1(n9653), .A2(n8371), .ZN(n9633) );
  OR2_X1 U5747 ( .A1(n5540), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5558) );
  AOI21_X1 U5748 ( .B1(n4624), .B2(n4631), .A(n4623), .ZN(n4622) );
  INV_X1 U5749 ( .A(n8278), .ZN(n4623) );
  OAI21_X1 U5750 ( .B1(n7596), .B2(n4552), .A(n4649), .ZN(n7934) );
  INV_X1 U5751 ( .A(n4650), .ZN(n4649) );
  OAI21_X1 U5752 ( .B1(n5686), .B2(n4552), .A(n5687), .ZN(n4650) );
  OR2_X1 U5753 ( .A1(n5483), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5754 ( .A1(n4876), .A2(n4569), .ZN(n4669) );
  INV_X1 U5755 ( .A(n5461), .ZN(n4670) );
  AOI21_X1 U5756 ( .B1(n7585), .B2(n8490), .A(n4548), .ZN(n4655) );
  INV_X1 U5757 ( .A(n7584), .ZN(n4658) );
  OAI21_X1 U5758 ( .B1(n7589), .B2(n5685), .A(n8334), .ZN(n7597) );
  AND2_X1 U5759 ( .A1(n8339), .A2(n8336), .ZN(n8477) );
  NAND2_X1 U5760 ( .A1(n4657), .A2(n4656), .ZN(n7585) );
  INV_X1 U5761 ( .A(n5122), .ZN(n4656) );
  INV_X1 U5762 ( .A(n7566), .ZN(n4657) );
  INV_X1 U5763 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5417) );
  INV_X1 U5764 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7460) );
  AND2_X1 U5765 ( .A1(n5402), .A2(n7460), .ZN(n5418) );
  AOI21_X1 U5766 ( .B1(n8487), .B2(n4648), .A(n4647), .ZN(n4646) );
  INV_X1 U5767 ( .A(n8319), .ZN(n4647) );
  NOR2_X1 U5768 ( .A1(n5385), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5402) );
  OR2_X1 U5769 ( .A1(n5369), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5385) );
  OR2_X1 U5770 ( .A1(n9386), .A2(n7320), .ZN(n8303) );
  AND4_X1 U5771 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n7321)
         );
  OAI21_X1 U5772 ( .B1(n5681), .B2(n4636), .A(n4634), .ZN(n7009) );
  INV_X1 U5773 ( .A(n4635), .ZN(n4634) );
  NAND2_X1 U5774 ( .A1(n8309), .A2(n8301), .ZN(n6887) );
  NAND2_X1 U5775 ( .A1(n7036), .A2(n5384), .ZN(n7309) );
  INV_X1 U5776 ( .A(n4654), .ZN(n4858) );
  OAI22_X1 U5777 ( .A1(n5336), .A2(n5855), .B1(n10549), .B2(n6602), .ZN(n4654)
         );
  OR2_X1 U5778 ( .A1(n8453), .A2(n6575), .ZN(n6842) );
  NOR2_X1 U5779 ( .A1(n6953), .A2(n5740), .ZN(n6988) );
  INV_X1 U5780 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5720) );
  INV_X1 U5781 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5657) );
  OR2_X1 U5782 ( .A1(n5974), .A2(n7820), .ZN(n5987) );
  NAND2_X1 U5783 ( .A1(n8038), .A2(n6410), .ZN(n6417) );
  OR2_X1 U5784 ( .A1(n6087), .A2(n9808), .ZN(n6099) );
  OAI21_X1 U5785 ( .B1(n9885), .B2(n9880), .A(n9804), .ZN(n9862) );
  NAND2_X1 U5786 ( .A1(n9880), .A2(n4553), .ZN(n4695) );
  AND2_X1 U5787 ( .A1(n7761), .A2(n7359), .ZN(n4678) );
  INV_X1 U5788 ( .A(n7761), .ZN(n4676) );
  INV_X1 U5789 ( .A(n6369), .ZN(n5052) );
  INV_X1 U5790 ( .A(n6385), .ZN(n5051) );
  OR2_X1 U5791 ( .A1(n7700), .A2(n6370), .ZN(n5053) );
  INV_X1 U5792 ( .A(n6805), .ZN(n6293) );
  OR2_X1 U5793 ( .A1(n8875), .A2(n6535), .ZN(n7406) );
  OR2_X1 U5794 ( .A1(n8807), .A2(n6665), .ZN(n9908) );
  INV_X1 U5795 ( .A(n9887), .ZN(n9910) );
  NAND2_X1 U5796 ( .A1(n9919), .A2(n9921), .ZN(n9920) );
  NOR2_X1 U5797 ( .A1(n6525), .A2(n6524), .ZN(n6531) );
  INV_X1 U5798 ( .A(n4935), .ZN(n8780) );
  NAND2_X1 U5799 ( .A1(n4935), .A2(n4573), .ZN(n8783) );
  OR2_X1 U5800 ( .A1(n4940), .A2(n8804), .ZN(n8866) );
  AND2_X1 U5801 ( .A1(n6105), .A2(n6104), .ZN(n9834) );
  AND2_X1 U5802 ( .A1(n6083), .A2(n6082), .ZN(n9827) );
  AND3_X1 U5803 ( .A1(n5833), .A2(n5832), .A3(n5831), .ZN(n8205) );
  AND3_X1 U5804 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n8153) );
  INV_X1 U5805 ( .A(n5907), .ZN(n8540) );
  AND4_X1 U5806 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n7868)
         );
  AND4_X1 U5807 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n7640)
         );
  AND4_X1 U5808 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n7678)
         );
  AND4_X1 U5809 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n7362)
         );
  NAND2_X1 U5810 ( .A1(n5015), .A2(n4600), .ZN(n5011) );
  NAND2_X1 U5811 ( .A1(n4543), .A2(n4600), .ZN(n5010) );
  NAND2_X1 U5812 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  NAND2_X1 U5813 ( .A1(n10094), .A2(n10296), .ZN(n10077) );
  NAND2_X1 U5814 ( .A1(n10156), .A2(n4578), .ZN(n10110) );
  NOR2_X1 U5815 ( .A1(n10110), .A2(n10095), .ZN(n10094) );
  NAND2_X1 U5816 ( .A1(n10156), .A2(n4882), .ZN(n10140) );
  INV_X1 U5817 ( .A(n8616), .ZN(n10154) );
  NAND2_X1 U5818 ( .A1(n10156), .A2(n6206), .ZN(n10157) );
  AND2_X1 U5819 ( .A1(n10197), .A2(n9943), .ZN(n5022) );
  NAND2_X1 U5820 ( .A1(n10322), .A2(n9826), .ZN(n5023) );
  INV_X1 U5821 ( .A(n10188), .ZN(n5024) );
  XNOR2_X1 U5822 ( .A(n10177), .B(n9888), .ZN(n10174) );
  NAND2_X1 U5823 ( .A1(n8145), .A2(n4883), .ZN(n10193) );
  AND2_X1 U5824 ( .A1(n4540), .A2(n10322), .ZN(n4883) );
  NOR2_X1 U5825 ( .A1(n10193), .A2(n10177), .ZN(n10156) );
  NAND2_X1 U5826 ( .A1(n5798), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6065) );
  OR2_X1 U5827 ( .A1(n8212), .A2(n9944), .ZN(n6058) );
  NAND2_X1 U5828 ( .A1(n8209), .A2(n4571), .ZN(n5028) );
  NAND2_X1 U5829 ( .A1(n8145), .A2(n4885), .ZN(n10207) );
  NOR2_X1 U5830 ( .A1(n5126), .A2(n9848), .ZN(n8145) );
  NAND2_X1 U5831 ( .A1(n8145), .A2(n8150), .ZN(n8211) );
  INV_X1 U5832 ( .A(n8763), .ZN(n4975) );
  NAND2_X1 U5833 ( .A1(n4996), .A2(n4995), .ZN(n8057) );
  AOI21_X1 U5834 ( .B1(n4998), .B2(n6033), .A(n4580), .ZN(n4996) );
  NOR2_X1 U5835 ( .A1(n7874), .A2(n4896), .ZN(n4895) );
  INV_X1 U5836 ( .A(n4897), .ZN(n4896) );
  AND2_X1 U5837 ( .A1(n8683), .A2(n8671), .ZN(n8760) );
  NAND2_X1 U5838 ( .A1(n7867), .A2(n8760), .ZN(n7866) );
  OR2_X1 U5839 ( .A1(n5989), .A2(n6821), .ZN(n6001) );
  NAND2_X1 U5840 ( .A1(n7610), .A2(n4899), .ZN(n10433) );
  NAND2_X1 U5841 ( .A1(n7610), .A2(n10501), .ZN(n7627) );
  AND2_X1 U5842 ( .A1(n5994), .A2(n5981), .ZN(n5026) );
  AND2_X1 U5843 ( .A1(n7681), .A2(n10494), .ZN(n7610) );
  NOR2_X1 U5844 ( .A1(n5118), .A2(n10486), .ZN(n7681) );
  AND2_X1 U5845 ( .A1(n5980), .A2(n8653), .ZN(n8755) );
  NAND2_X1 U5846 ( .A1(n4974), .A2(n8834), .ZN(n4973) );
  INV_X1 U5847 ( .A(n7377), .ZN(n4974) );
  NOR2_X1 U5848 ( .A1(n6936), .A2(n10442), .ZN(n4889) );
  INV_X1 U5849 ( .A(n4891), .ZN(n4890) );
  NOR2_X1 U5850 ( .A1(n4891), .A2(n6936), .ZN(n7373) );
  NAND2_X1 U5851 ( .A1(n4893), .A2(n4529), .ZN(n7248) );
  NAND2_X1 U5852 ( .A1(n4893), .A2(n7449), .ZN(n5127) );
  INV_X1 U5853 ( .A(n8627), .ZN(n8746) );
  OAI211_X1 U5854 ( .C1(n6271), .C2(n6266), .A(n8873), .B(n7436), .ZN(n7871)
         );
  NAND2_X1 U5855 ( .A1(n7485), .A2(n6173), .ZN(n8624) );
  INV_X1 U5856 ( .A(n7480), .ZN(n4994) );
  NAND2_X1 U5857 ( .A1(n7486), .A2(n7480), .ZN(n7485) );
  NOR2_X1 U5858 ( .A1(n10502), .A2(n8816), .ZN(n6528) );
  OR2_X1 U5859 ( .A1(n8737), .A2(n8871), .ZN(n10499) );
  INV_X1 U5860 ( .A(n10502), .ZN(n10435) );
  OR2_X1 U5861 ( .A1(n7436), .A2(n6266), .ZN(n10517) );
  NAND2_X1 U5862 ( .A1(n7871), .A2(n10499), .ZN(n10520) );
  NAND2_X1 U5863 ( .A1(n8424), .A2(n8423), .ZN(n8434) );
  OR2_X1 U5864 ( .A1(n8422), .A2(n8421), .ZN(n8423) );
  OR2_X1 U5865 ( .A1(n8420), .A2(n8419), .ZN(n8424) );
  XNOR2_X1 U5866 ( .A(n8434), .B(n8433), .ZN(n8544) );
  XNOR2_X1 U5867 ( .A(n8420), .B(SI_29_), .ZN(n8881) );
  INV_X1 U5868 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U5869 ( .A(n5643), .B(n5642), .ZN(n8091) );
  XNOR2_X1 U5870 ( .A(n6219), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6239) );
  INV_X1 U5871 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6163) );
  AOI21_X1 U5872 ( .B1(n5545), .B2(n5214), .A(n4601), .ZN(n5284) );
  AND2_X1 U5873 ( .A1(n5218), .A2(n5217), .ZN(n5283) );
  XNOR2_X1 U5874 ( .A(n5549), .B(n5548), .ZN(n7432) );
  NAND2_X1 U5875 ( .A1(n6046), .A2(n6160), .ZN(n6048) );
  NAND2_X1 U5876 ( .A1(n5819), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U5877 ( .A1(n4950), .A2(n4954), .ZN(n5521) );
  OR2_X1 U5878 ( .A1(n4960), .A2(n4956), .ZN(n4950) );
  NAND2_X1 U5879 ( .A1(n4953), .A2(n5191), .ZN(n5507) );
  NAND2_X1 U5880 ( .A1(n5409), .A2(n5408), .ZN(n5413) );
  NAND2_X1 U5881 ( .A1(n4934), .A2(n5157), .ZN(n5397) );
  NAND2_X1 U5882 ( .A1(n4660), .A2(n5155), .ZN(n5392) );
  NAND2_X1 U5883 ( .A1(n4663), .A2(n4928), .ZN(n4660) );
  INV_X1 U5884 ( .A(n5360), .ZN(n4927) );
  AND2_X1 U5885 ( .A1(n5069), .A2(n5077), .ZN(n5068) );
  NAND2_X1 U5886 ( .A1(n7845), .A2(n5071), .ZN(n5070) );
  OR2_X1 U5887 ( .A1(n8027), .A2(n9379), .ZN(n5077) );
  INV_X1 U5888 ( .A(n9381), .ZN(n8011) );
  XNOR2_X1 U5889 ( .A(n6997), .B(n9726), .ZN(n6993) );
  NAND2_X1 U5890 ( .A1(n6992), .A2(n5098), .ZN(n6999) );
  NAND2_X1 U5891 ( .A1(n8289), .A2(n6977), .ZN(n7023) );
  NAND2_X1 U5892 ( .A1(n4513), .A2(n7044), .ZN(n6977) );
  NAND2_X1 U5893 ( .A1(n9321), .A2(n8579), .ZN(n8932) );
  NAND2_X1 U5894 ( .A1(n5568), .A2(n5567), .ZN(n8936) );
  NAND2_X1 U5895 ( .A1(n5106), .A2(n8594), .ZN(n8939) );
  NAND2_X1 U5896 ( .A1(n5091), .A2(n4551), .ZN(n5090) );
  INV_X1 U5897 ( .A(n8559), .ZN(n5091) );
  AND2_X1 U5898 ( .A1(n6999), .A2(n5096), .ZN(n7319) );
  NAND2_X1 U5899 ( .A1(n6999), .A2(n6998), .ZN(n7002) );
  AND2_X1 U5900 ( .A1(n6960), .A2(n6961), .ZN(n9346) );
  NAND2_X1 U5901 ( .A1(n5088), .A2(n5087), .ZN(n8572) );
  NAND2_X1 U5902 ( .A1(n8559), .A2(n4533), .ZN(n5087) );
  NOR2_X1 U5903 ( .A1(n4537), .A2(n8596), .ZN(n9352) );
  XNOR2_X1 U5904 ( .A(n8597), .B(n9368), .ZN(n9353) );
  NAND2_X1 U5905 ( .A1(n5268), .A2(n5267), .ZN(n9361) );
  NAND2_X1 U5906 ( .A1(n6957), .A2(n8222), .ZN(n9360) );
  INV_X1 U5907 ( .A(n9346), .ZN(n9358) );
  NAND2_X1 U5908 ( .A1(n4720), .A2(n6967), .ZN(n8519) );
  XNOR2_X1 U5909 ( .A(n5660), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8523) );
  AND4_X1 U5910 ( .A1(n8446), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8449)
         );
  INV_X1 U5911 ( .A(n9645), .ZN(n9376) );
  INV_X1 U5912 ( .A(n7321), .ZN(n9386) );
  NAND2_X1 U5913 ( .A1(n4515), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U5914 ( .A1(n4515), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5329) );
  NOR2_X1 U5915 ( .A1(n7207), .A2(n4920), .ZN(n10543) );
  NAND2_X1 U5916 ( .A1(n4846), .A2(n7285), .ZN(n7065) );
  NAND2_X1 U5917 ( .A1(n4922), .A2(n7290), .ZN(n7294) );
  NAND2_X1 U5918 ( .A1(n7539), .A2(n7540), .ZN(n10591) );
  XNOR2_X1 U5919 ( .A(n7983), .B(n7977), .ZN(n7740) );
  AND2_X1 U5920 ( .A1(n5429), .A2(n5452), .ZN(n7997) );
  INV_X1 U5921 ( .A(n7991), .ZN(n7993) );
  INV_X1 U5922 ( .A(n7967), .ZN(n7968) );
  NOR2_X1 U5923 ( .A1(n8177), .A2(n8159), .ZN(n8160) );
  INV_X1 U5924 ( .A(n4839), .ZN(n9443) );
  OR2_X1 U5925 ( .A1(n9435), .A2(n9434), .ZN(n4839) );
  INV_X1 U5926 ( .A(n9444), .ZN(n4838) );
  NAND2_X1 U5927 ( .A1(n4906), .A2(n4905), .ZN(n9466) );
  NAND2_X1 U5928 ( .A1(n4840), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4837) );
  NAND2_X1 U5929 ( .A1(n9444), .A2(n4840), .ZN(n4836) );
  INV_X1 U5930 ( .A(n9445), .ZN(n4840) );
  INV_X1 U5931 ( .A(n4755), .ZN(n4754) );
  NOR2_X1 U5932 ( .A1(n4757), .A2(n9504), .ZN(n4756) );
  NAND2_X1 U5933 ( .A1(n9513), .A2(n9514), .ZN(n4752) );
  NAND2_X1 U5934 ( .A1(n9505), .A2(n10612), .ZN(n4753) );
  NAND2_X1 U5935 ( .A1(n4854), .A2(n4853), .ZN(n4851) );
  OAI21_X1 U5936 ( .B1(n9576), .B2(n4802), .A(n4800), .ZN(n5763) );
  AOI21_X1 U5937 ( .B1(n9366), .B2(n6257), .A(n6256), .ZN(n6258) );
  NOR2_X1 U5938 ( .A1(n9571), .A2(n9644), .ZN(n6256) );
  XNOR2_X1 U5939 ( .A(n4653), .B(n4652), .ZN(n9557) );
  INV_X1 U5940 ( .A(n8507), .ZN(n4652) );
  NAND2_X1 U5941 ( .A1(n4805), .A2(n4803), .ZN(n4653) );
  INV_X1 U5942 ( .A(n4806), .ZN(n4803) );
  OAI22_X1 U5943 ( .A1(n4863), .A2(n4862), .B1(n4872), .B2(n4871), .ZN(n9560)
         );
  NAND2_X1 U5944 ( .A1(n4531), .A2(n4873), .ZN(n4862) );
  OAI21_X1 U5945 ( .B1(n9576), .B2(n8396), .A(n8404), .ZN(n9564) );
  XNOR2_X1 U5946 ( .A(n4674), .B(n9575), .ZN(n9570) );
  NAND2_X1 U5947 ( .A1(n5613), .A2(n5612), .ZN(n9572) );
  NAND2_X1 U5948 ( .A1(n4868), .A2(n4874), .ZN(n9581) );
  NAND2_X1 U5949 ( .A1(n4668), .A2(n4878), .ZN(n9643) );
  NAND2_X1 U5950 ( .A1(n8084), .A2(n8498), .ZN(n4877) );
  INV_X1 U5951 ( .A(n9790), .ZN(n8261) );
  NAND2_X1 U5952 ( .A1(n4626), .A2(n4628), .ZN(n8086) );
  NAND2_X1 U5953 ( .A1(n4627), .A2(n4632), .ZN(n4626) );
  NAND2_X1 U5954 ( .A1(n7654), .A2(n8345), .ZN(n7827) );
  NAND2_X1 U5955 ( .A1(n4876), .A2(n5461), .ZN(n7828) );
  NAND2_X1 U5956 ( .A1(n5682), .A2(n8313), .ZN(n7306) );
  OR2_X1 U5957 ( .A1(n5333), .A2(n6609), .ZN(n5302) );
  OR2_X1 U5958 ( .A1(n5336), .A2(n6610), .ZN(n5301) );
  INV_X1 U5959 ( .A(n10628), .ZN(n8222) );
  INV_X1 U5960 ( .A(n9651), .ZN(n9637) );
  NAND2_X1 U5961 ( .A1(n6844), .A2(n8222), .ZN(n10629) );
  AND2_X1 U5962 ( .A1(n8441), .A2(n8440), .ZN(n9662) );
  NAND2_X1 U5963 ( .A1(n5648), .A2(n5647), .ZN(n9671) );
  INV_X1 U5964 ( .A(n9662), .ZN(n9746) );
  INV_X1 U5965 ( .A(n9361), .ZN(n9757) );
  NAND2_X1 U5966 ( .A1(n4673), .A2(n5416), .ZN(n7579) );
  NAND2_X1 U5967 ( .A1(n5718), .A2(n5717), .ZN(n6640) );
  AND2_X1 U5968 ( .A1(n7057), .A2(n7020), .ZN(n6952) );
  AND2_X1 U5969 ( .A1(n7055), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7020) );
  AND2_X1 U5970 ( .A1(n5086), .A2(n4811), .ZN(n4810) );
  AND2_X1 U5971 ( .A1(n4560), .A2(n5067), .ZN(n4811) );
  NOR2_X1 U5972 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5067) );
  INV_X1 U5973 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9792) );
  INV_X1 U5974 ( .A(n5277), .ZN(n9802) );
  INV_X1 U5975 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8964) );
  XNOR2_X1 U5976 ( .A(n5702), .B(n5701), .ZN(n8009) );
  INV_X1 U5977 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5978 ( .A1(n5722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5702) );
  INV_X1 U5979 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7886) );
  INV_X1 U5980 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7777) );
  INV_X1 U5981 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7814) );
  INV_X1 U5982 ( .A(n8523), .ZN(n7816) );
  INV_X1 U5983 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7562) );
  INV_X1 U5984 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9197) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7315) );
  INV_X1 U5986 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7259) );
  INV_X1 U5987 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7215) );
  INV_X1 U5988 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7097) );
  INV_X1 U5989 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9278) );
  INV_X1 U5990 ( .A(n9419), .ZN(n9433) );
  INV_X1 U5991 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8970) );
  INV_X1 U5992 ( .A(n7997), .ZN(n7988) );
  INV_X1 U5993 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6632) );
  INV_X1 U5994 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9206) );
  INV_X1 U5995 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9234) );
  NOR2_X1 U5997 ( .A1(n4555), .A2(n9833), .ZN(n4689) );
  AND2_X1 U5998 ( .A1(n4553), .A2(n4694), .ZN(n4690) );
  NAND2_X1 U5999 ( .A1(n5058), .A2(n6426), .ZN(n9851) );
  NAND2_X1 U6000 ( .A1(n9841), .A2(n9842), .ZN(n5058) );
  NAND2_X1 U6001 ( .A1(n4691), .A2(n4695), .ZN(n9864) );
  AND2_X1 U6002 ( .A1(n4693), .A2(n4692), .ZN(n4691) );
  INV_X1 U6003 ( .A(n5045), .ZN(n4692) );
  AND2_X1 U6004 ( .A1(n6531), .A2(n6266), .ZN(n9916) );
  NAND2_X1 U6005 ( .A1(n6274), .A2(n6598), .ZN(n8875) );
  OR2_X1 U6006 ( .A1(n10109), .A2(n6111), .ZN(n6116) );
  INV_X1 U6007 ( .A(n9834), .ZN(n9939) );
  INV_X1 U6008 ( .A(n9827), .ZN(n9941) );
  OR2_X1 U6009 ( .A1(n6599), .A2(n6274), .ZN(n9942) );
  INV_X1 U6010 ( .A(n8205), .ZN(n9945) );
  AND4_X1 U6011 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n9952)
         );
  NAND2_X1 U6012 ( .A1(n5870), .A2(n5125), .ZN(n9962) );
  AND3_X1 U6013 ( .A1(n5869), .A2(n5868), .A3(n5867), .ZN(n5125) );
  NAND2_X2 U6014 ( .A1(n5851), .A2(n5852), .ZN(n9963) );
  AND3_X1 U6015 ( .A1(n5850), .A2(n5849), .A3(n5848), .ZN(n5851) );
  OR2_X1 U6016 ( .A1(n6739), .A2(n6665), .ZN(n10007) );
  NAND2_X1 U6017 ( .A1(n5819), .A2(n5042), .ZN(n5036) );
  NAND2_X1 U6018 ( .A1(n5041), .A2(n5040), .ZN(n5039) );
  AOI211_X1 U6019 ( .C1(n10043), .C2(n10042), .A(n10502), .B(n10041), .ZN(
        n10218) );
  NAND2_X1 U6020 ( .A1(n8732), .A2(n8735), .ZN(n4986) );
  NAND2_X1 U6021 ( .A1(n5012), .A2(n5015), .ZN(n10093) );
  NAND2_X1 U6022 ( .A1(n8203), .A2(n8702), .ZN(n10200) );
  INV_X1 U6023 ( .A(n10281), .ZN(n6032) );
  NAND2_X1 U6024 ( .A1(n4997), .A2(n5001), .ZN(n7854) );
  NAND2_X1 U6025 ( .A1(n10431), .A2(n5000), .ZN(n4997) );
  NAND2_X1 U6026 ( .A1(n7623), .A2(n8838), .ZN(n10425) );
  INV_X1 U6027 ( .A(n5116), .ZN(n5007) );
  INV_X1 U6028 ( .A(n10190), .ZN(n10452) );
  INV_X1 U6029 ( .A(n10194), .ZN(n10450) );
  INV_X1 U6030 ( .A(n8822), .ZN(n6205) );
  OR2_X1 U6031 ( .A1(n10215), .A2(n7412), .ZN(n10456) );
  INV_X1 U6032 ( .A(n10456), .ZN(n10441) );
  INV_X1 U6033 ( .A(n10095), .ZN(n10300) );
  INV_X1 U6034 ( .A(n10142), .ZN(n10311) );
  INV_X1 U6035 ( .A(n8212), .ZN(n10330) );
  AND2_X1 U6036 ( .A1(n10334), .A2(n10333), .ZN(n10469) );
  INV_X1 U6037 ( .A(n5812), .ZN(n8545) );
  NAND2_X1 U6038 ( .A1(n5805), .A2(n5804), .ZN(n5808) );
  NAND2_X1 U6039 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  AOI21_X1 U6040 ( .B1(n6219), .B2(n4764), .A(n4763), .ZN(n4762) );
  OR2_X1 U6041 ( .A1(n6219), .A2(n4766), .ZN(n4765) );
  AND2_X1 U6042 ( .A1(n5787), .A2(n4766), .ZN(n4764) );
  INV_X1 U6043 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9258) );
  XNOR2_X1 U6044 ( .A(n6210), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7957) );
  INV_X1 U6045 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U6046 ( .A1(n5566), .A2(n4971), .ZN(n4964) );
  INV_X1 U6047 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9285) );
  INV_X1 U6048 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7813) );
  INV_X1 U6049 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7524) );
  INV_X1 U6050 ( .A(n4526), .ZN(n8742) );
  INV_X1 U6051 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7405) );
  INV_X1 U6052 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7338) );
  INV_X1 U6053 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7261) );
  INV_X1 U6054 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7214) );
  INV_X1 U6055 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7043) );
  INV_X1 U6056 ( .A(n7713), .ZN(n7723) );
  INV_X1 U6057 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6745) );
  INV_X1 U6058 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6735) );
  INV_X1 U6059 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6639) );
  INV_X1 U6060 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U6061 ( .A1(n5150), .A2(n5149), .ZN(n5361) );
  XNOR2_X1 U6062 ( .A(n5297), .B(n5296), .ZN(n6610) );
  INV_X1 U6063 ( .A(n4918), .ZN(n7532) );
  OAI21_X1 U6064 ( .B1(n6588), .B2(n9715), .A(n6587), .ZN(n6589) );
  NOR2_X1 U6065 ( .A1(n5115), .A2(n5766), .ZN(n5767) );
  OAI21_X1 U6066 ( .B1(n10296), .B2(n9931), .A(n6571), .ZN(n6572) );
  NAND2_X1 U6067 ( .A1(n5062), .A2(n4602), .ZN(n6553) );
  OAI21_X1 U6068 ( .B1(n6558), .B2(n10534), .A(n6557), .ZN(P1_U3550) );
  NOR2_X1 U6069 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  OAI21_X1 U6070 ( .B1(n10287), .B2(n6596), .A(n4894), .ZN(n10288) );
  OR2_X1 U6071 ( .A1(n10523), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n4894) );
  INV_X1 U6072 ( .A(n6594), .ZN(n6595) );
  OAI22_X1 U6073 ( .A1(n6593), .A2(n10329), .B1(n10523), .B2(n6592), .ZN(n6594) );
  INV_X1 U6074 ( .A(n6253), .ZN(n6254) );
  NAND2_X1 U6075 ( .A1(n8638), .A2(n8637), .ZN(n4528) );
  AND2_X1 U6076 ( .A1(n7341), .A2(n7449), .ZN(n4529) );
  NAND2_X1 U6077 ( .A1(n4769), .A2(n4741), .ZN(n4530) );
  AND2_X1 U6078 ( .A1(n4869), .A2(n9589), .ZN(n4531) );
  OR2_X1 U6079 ( .A1(n6167), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4532) );
  AOI21_X1 U6080 ( .B1(n10344), .B2(n8529), .A(n8528), .ZN(n10289) );
  INV_X1 U6081 ( .A(n10289), .ZN(n4940) );
  AND2_X1 U6082 ( .A1(n5092), .A2(n4562), .ZN(n4533) );
  INV_X1 U6083 ( .A(n9833), .ZN(n4694) );
  AND2_X1 U6084 ( .A1(n9852), .A2(n5059), .ZN(n4534) );
  INV_X1 U6085 ( .A(n8721), .ZN(n4785) );
  INV_X1 U6086 ( .A(n8347), .ZN(n4718) );
  INV_X1 U6087 ( .A(n10177), .ZN(n10318) );
  AND2_X1 U6088 ( .A1(n8635), .A2(n8825), .ZN(n4535) );
  AND2_X1 U6089 ( .A1(n4671), .A2(n8348), .ZN(n4536) );
  AND2_X1 U6090 ( .A1(n5099), .A2(n5107), .ZN(n4537) );
  OR2_X1 U6091 ( .A1(n8417), .A2(n8416), .ZN(n4538) );
  NAND2_X1 U6092 ( .A1(n4766), .A2(n5783), .ZN(n4539) );
  AND2_X1 U6093 ( .A1(n4885), .A2(n4884), .ZN(n4540) );
  NOR2_X1 U6094 ( .A1(n8343), .A2(n8453), .ZN(n4541) );
  INV_X1 U6095 ( .A(n8920), .ZN(n9769) );
  NAND2_X1 U6096 ( .A1(n5587), .A2(n5586), .ZN(n8920) );
  NAND2_X1 U6097 ( .A1(n10043), .A2(n4769), .ZN(n4542) );
  NAND2_X1 U6098 ( .A1(n4591), .A2(n5018), .ZN(n5015) );
  NAND2_X1 U6099 ( .A1(n5013), .A2(n6128), .ZN(n4543) );
  AND2_X1 U6100 ( .A1(n4882), .A2(n4881), .ZN(n4544) );
  AND4_X1 U6101 ( .A1(n5423), .A2(n5422), .A3(n5421), .A4(n5420), .ZN(n7843)
         );
  INV_X1 U6102 ( .A(n7843), .ZN(n4672) );
  OR2_X1 U6103 ( .A1(n10477), .A2(n9956), .ZN(n4545) );
  INV_X2 U6104 ( .A(n8066), .ZN(n10215) );
  INV_X1 U6105 ( .A(n8737), .ZN(n8629) );
  NAND2_X1 U6106 ( .A1(n8816), .A2(n6532), .ZN(n6264) );
  INV_X1 U6107 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4920) );
  INV_X1 U6108 ( .A(n4520), .ZN(n5592) );
  AND2_X1 U6109 ( .A1(n9746), .A2(n8447), .ZN(n4546) );
  NAND4_X1 U6110 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n9725)
         );
  AND2_X1 U6111 ( .A1(n5152), .A2(SI_5_), .ZN(n4547) );
  NOR2_X1 U6112 ( .A1(n7851), .A2(n9382), .ZN(n4548) );
  NAND2_X1 U6113 ( .A1(n5037), .A2(n5036), .ZN(n6166) );
  OR2_X1 U6114 ( .A1(n6478), .A2(n6477), .ZN(n5049) );
  NOR2_X1 U6115 ( .A1(n5377), .A2(n5550), .ZN(n5658) );
  OR2_X1 U6116 ( .A1(n9906), .A2(n5065), .ZN(n5064) );
  NAND2_X1 U6117 ( .A1(n8719), .A2(n8629), .ZN(n4549) );
  AND2_X1 U6118 ( .A1(n10094), .A2(n4888), .ZN(n4550) );
  OR2_X1 U6119 ( .A1(n8549), .A2(n5094), .ZN(n4551) );
  OR2_X1 U6120 ( .A1(n4651), .A2(n5688), .ZN(n4552) );
  NAND2_X1 U6121 ( .A1(n6222), .A2(n6221), .ZN(n6274) );
  NAND2_X1 U6122 ( .A1(n8718), .A2(n4549), .ZN(n4793) );
  NAND2_X1 U6123 ( .A1(n5086), .A2(n5249), .ZN(n5377) );
  INV_X1 U6124 ( .A(n8313), .ZN(n4648) );
  XNOR2_X1 U6125 ( .A(n5313), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7051) );
  AND2_X1 U6126 ( .A1(n5044), .A2(n9804), .ZN(n4553) );
  OR2_X1 U6127 ( .A1(n7874), .A2(n9948), .ZN(n4554) );
  NOR2_X1 U6128 ( .A1(n5045), .A2(n6497), .ZN(n4555) );
  NOR2_X1 U6129 ( .A1(n8410), .A2(n4809), .ZN(n4556) );
  NAND2_X1 U6130 ( .A1(n9895), .A2(n9813), .ZN(n4557) );
  AND2_X1 U6131 ( .A1(n8373), .A2(n8374), .ZN(n4558) );
  INV_X1 U6132 ( .A(n8702), .ZN(n4993) );
  AND2_X1 U6133 ( .A1(n4877), .A2(n5533), .ZN(n4559) );
  NAND2_X1 U6134 ( .A1(n5338), .A2(n4858), .ZN(n6862) );
  INV_X1 U6135 ( .A(n6862), .ZN(n6978) );
  NAND2_X1 U6136 ( .A1(n4964), .A2(n4969), .ZN(n5584) );
  NAND2_X1 U6137 ( .A1(n8802), .A2(n8800), .ZN(n8732) );
  XNOR2_X1 U6138 ( .A(n5599), .B(n5598), .ZN(n6094) );
  AND2_X1 U6139 ( .A1(n5249), .A2(n5265), .ZN(n4560) );
  AND2_X1 U6140 ( .A1(n8581), .A2(n9631), .ZN(n4561) );
  NAND2_X1 U6141 ( .A1(n8749), .A2(n7636), .ZN(n7376) );
  OR2_X1 U6142 ( .A1(n8253), .A2(n8259), .ZN(n4562) );
  OR2_X1 U6143 ( .A1(n7146), .A2(n7145), .ZN(n4563) );
  AND2_X1 U6144 ( .A1(n4672), .A2(n5416), .ZN(n4564) );
  AND3_X1 U6145 ( .A1(n5878), .A2(n5877), .A3(n5876), .ZN(n7417) );
  OR2_X1 U6146 ( .A1(n10501), .A2(n9952), .ZN(n4565) );
  INV_X1 U6147 ( .A(n10275), .ZN(n8150) );
  AND3_X1 U6148 ( .A1(n4695), .A2(n4693), .A3(n4555), .ZN(n4566) );
  AND2_X1 U6149 ( .A1(n8709), .A2(n8737), .ZN(n4567) );
  AND3_X1 U6150 ( .A1(n4754), .A2(n4753), .A3(n4752), .ZN(n4568) );
  INV_X1 U6151 ( .A(n10080), .ZN(n10296) );
  NAND2_X1 U6152 ( .A1(n6130), .A2(n6129), .ZN(n10080) );
  NOR2_X1 U6153 ( .A1(n8351), .A2(n4670), .ZN(n4569) );
  INV_X1 U6154 ( .A(n7874), .ZN(n8044) );
  NAND2_X1 U6155 ( .A1(n6011), .A2(n6010), .ZN(n7874) );
  AND2_X1 U6156 ( .A1(n6108), .A2(n6107), .ZN(n10304) );
  NOR2_X1 U6157 ( .A1(n9368), .A2(n9361), .ZN(n4570) );
  OR2_X1 U6158 ( .A1(n10330), .A2(n9815), .ZN(n4571) );
  AND2_X1 U6159 ( .A1(n4980), .A2(n10430), .ZN(n4572) );
  NAND2_X1 U6160 ( .A1(n8808), .A2(n8629), .ZN(n4573) );
  OR2_X1 U6161 ( .A1(n7890), .A2(n5076), .ZN(n4574) );
  AND2_X1 U6162 ( .A1(n4912), .A2(n4913), .ZN(n4575) );
  AND2_X1 U6163 ( .A1(n5780), .A2(n4686), .ZN(n4576) );
  INV_X1 U6164 ( .A(n4632), .ZN(n4631) );
  INV_X1 U6165 ( .A(n8351), .ZN(n4827) );
  AND2_X1 U6166 ( .A1(n8634), .A2(n8641), .ZN(n4577) );
  INV_X1 U6167 ( .A(n4725), .ZN(n8826) );
  NAND2_X1 U6168 ( .A1(n8634), .A2(n8635), .ZN(n4725) );
  OR2_X1 U6169 ( .A1(n9726), .A2(n7108), .ZN(n8309) );
  INV_X1 U6170 ( .A(n8309), .ZN(n4636) );
  NAND2_X1 U6171 ( .A1(n6281), .A2(n6282), .ZN(n6295) );
  AND2_X1 U6172 ( .A1(n4544), .A2(n10304), .ZN(n4578) );
  NAND2_X1 U6173 ( .A1(n7738), .A2(n7737), .ZN(n7983) );
  AND2_X1 U6174 ( .A1(n6433), .A2(n6432), .ZN(n4579) );
  NOR2_X1 U6175 ( .A1(n6032), .A2(n8675), .ZN(n4580) );
  OR2_X1 U6176 ( .A1(n5704), .A2(n5703), .ZN(n4581) );
  AND2_X1 U6177 ( .A1(n7874), .A2(n9948), .ZN(n4582) );
  AND2_X1 U6178 ( .A1(n5055), .A2(n6380), .ZN(n5054) );
  INV_X1 U6179 ( .A(n8379), .ZN(n4704) );
  NAND2_X1 U6180 ( .A1(n7156), .A2(n7279), .ZN(n4583) );
  INV_X1 U6181 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U6182 ( .A1(n9548), .A2(n9366), .ZN(n4584) );
  INV_X1 U6183 ( .A(n8350), .ZN(n4719) );
  AND2_X1 U6184 ( .A1(n4793), .A2(n4785), .ZN(n4585) );
  INV_X1 U6185 ( .A(n4625), .ZN(n4624) );
  NAND2_X1 U6186 ( .A1(n4628), .A2(n8275), .ZN(n4625) );
  OR2_X1 U6187 ( .A1(n9790), .A2(n9645), .ZN(n4586) );
  OR2_X1 U6188 ( .A1(n4546), .A2(n8472), .ZN(n4587) );
  NOR2_X1 U6189 ( .A1(n8254), .A2(n9377), .ZN(n4588) );
  NAND2_X1 U6190 ( .A1(n4795), .A2(n4549), .ZN(n4791) );
  INV_X1 U6191 ( .A(n4791), .ZN(n4728) );
  NOR2_X1 U6192 ( .A1(n9562), .A2(n8601), .ZN(n4589) );
  INV_X1 U6193 ( .A(n10117), .ZN(n4796) );
  INV_X1 U6194 ( .A(n4793), .ZN(n4792) );
  NAND2_X1 U6195 ( .A1(n8243), .A2(n8242), .ZN(n4590) );
  NAND2_X1 U6196 ( .A1(n6117), .A2(n5017), .ZN(n4591) );
  INV_X1 U6197 ( .A(n5669), .ZN(n8521) );
  XNOR2_X1 U6198 ( .A(n5266), .B(n5265), .ZN(n5669) );
  NOR2_X1 U6199 ( .A1(n10442), .A2(n9957), .ZN(n4592) );
  NOR2_X1 U6200 ( .A1(n8708), .A2(n8707), .ZN(n4593) );
  AND2_X1 U6201 ( .A1(n4951), .A2(n4949), .ZN(n4594) );
  NAND2_X1 U6202 ( .A1(n8532), .A2(n8531), .ZN(n10043) );
  INV_X1 U6203 ( .A(n10043), .ZN(n4741) );
  INV_X1 U6204 ( .A(n7305), .ZN(n8487) );
  INV_X1 U6205 ( .A(n10197), .ZN(n10322) );
  NAND2_X1 U6206 ( .A1(n5790), .A2(n5789), .ZN(n10197) );
  AND2_X1 U6207 ( .A1(n4987), .A2(n8777), .ZN(n4595) );
  AND2_X1 U6208 ( .A1(n4916), .A2(n4915), .ZN(n4596) );
  AND2_X1 U6209 ( .A1(n4911), .A2(n4910), .ZN(n4597) );
  INV_X1 U6210 ( .A(n5956), .ZN(n5006) );
  INV_X1 U6211 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6158) );
  INV_X1 U6212 ( .A(n8808), .ZN(n4936) );
  INV_X1 U6213 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4644) );
  INV_X1 U6214 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5818) );
  INV_X1 U6215 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4642) );
  INV_X1 U6216 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U6217 ( .A1(n5053), .A2(n6369), .ZN(n7817) );
  INV_X1 U6218 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4826) );
  INV_X1 U6219 ( .A(n10549), .ZN(n4751) );
  AND2_X1 U6220 ( .A1(n8145), .A2(n4540), .ZN(n4598) );
  AND2_X1 U6221 ( .A1(n10156), .A2(n4544), .ZN(n4599) );
  NAND2_X1 U6222 ( .A1(n10095), .A2(n9937), .ZN(n4600) );
  NOR2_X1 U6223 ( .A1(n5213), .A2(n5212), .ZN(n4601) );
  NAND2_X1 U6224 ( .A1(n9920), .A2(n6418), .ZN(n9841) );
  AND3_X1 U6225 ( .A1(n6545), .A2(n9922), .A3(n6544), .ZN(n4602) );
  NAND2_X1 U6226 ( .A1(n8559), .A2(n8242), .ZN(n8548) );
  NAND2_X1 U6227 ( .A1(n5090), .A2(n5092), .ZN(n8255) );
  NAND2_X1 U6228 ( .A1(n8467), .A2(n8431), .ZN(n8508) );
  INV_X1 U6229 ( .A(n8508), .ZN(n4833) );
  INV_X1 U6230 ( .A(n9617), .ZN(n4702) );
  INV_X1 U6231 ( .A(n8789), .ZN(n4790) );
  NAND2_X1 U6232 ( .A1(n6096), .A2(n6095), .ZN(n10124) );
  INV_X1 U6233 ( .A(n10124), .ZN(n4881) );
  OR2_X1 U6234 ( .A1(n5679), .A2(n7044), .ZN(n8289) );
  INV_X1 U6235 ( .A(n8289), .ZN(n4638) );
  XNOR2_X1 U6236 ( .A(n6417), .B(n6415), .ZN(n9919) );
  INV_X1 U6237 ( .A(n9371), .ZN(n9604) );
  OR2_X1 U6238 ( .A1(n7978), .A2(n7977), .ZN(n4603) );
  AND2_X1 U6239 ( .A1(n9572), .A2(n9369), .ZN(n4604) );
  AND2_X1 U6240 ( .A1(n6071), .A2(n6070), .ZN(n9888) );
  INV_X1 U6241 ( .A(n9888), .ZN(n5021) );
  NAND2_X1 U6242 ( .A1(n5633), .A2(n5632), .ZN(n8601) );
  INV_X1 U6243 ( .A(n9883), .ZN(n5048) );
  AND2_X1 U6244 ( .A1(n4839), .A2(n4838), .ZN(n4605) );
  INV_X1 U6245 ( .A(n4873), .ZN(n4871) );
  NAND2_X1 U6246 ( .A1(n9761), .A2(n9583), .ZN(n4873) );
  AND2_X1 U6247 ( .A1(n4669), .A2(n8348), .ZN(n4606) );
  NAND2_X1 U6248 ( .A1(n9872), .A2(n9871), .ZN(n4607) );
  AND2_X1 U6249 ( .A1(n9370), .A2(n9580), .ZN(n4608) );
  AND2_X1 U6250 ( .A1(n4724), .A2(n8638), .ZN(n4609) );
  AND2_X1 U6251 ( .A1(n5110), .A2(n8599), .ZN(n4610) );
  INV_X1 U6252 ( .A(n5019), .ZN(n5017) );
  AND2_X1 U6253 ( .A1(n10124), .A2(n9939), .ZN(n5019) );
  INV_X1 U6254 ( .A(n10462), .ZN(n8066) );
  AOI21_X1 U6255 ( .B1(n6217), .B2(n6216), .A(n6215), .ZN(n6222) );
  NAND2_X1 U6256 ( .A1(n5821), .A2(n5820), .ZN(n10208) );
  INV_X1 U6257 ( .A(n10208), .ZN(n4884) );
  NAND2_X1 U6258 ( .A1(n6353), .A2(n7359), .ZN(n7700) );
  NAND2_X1 U6259 ( .A1(n5735), .A2(n8070), .ZN(n6975) );
  AND2_X1 U6260 ( .A1(n10418), .A2(n6346), .ZN(n7360) );
  NAND2_X1 U6261 ( .A1(n5050), .A2(n4680), .ZN(n7760) );
  OAI21_X1 U6262 ( .B1(n5700), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6263 ( .A1(n5073), .A2(n5074), .ZN(n8029) );
  NAND2_X1 U6264 ( .A1(n5383), .A2(n8482), .ZN(n7036) );
  NAND2_X1 U6265 ( .A1(n6870), .A2(n6316), .ZN(n7226) );
  INV_X1 U6266 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U6267 ( .A1(n5027), .A2(n5981), .ZN(n7506) );
  NAND2_X1 U6268 ( .A1(n7610), .A2(n4897), .ZN(n4900) );
  AND2_X1 U6269 ( .A1(n8353), .A2(n8352), .ZN(n8495) );
  INV_X1 U6270 ( .A(n8495), .ZN(n4671) );
  NOR2_X1 U6271 ( .A1(n8161), .A2(n8160), .ZN(n4611) );
  AND2_X1 U6272 ( .A1(n5009), .A2(n5007), .ZN(n4612) );
  NAND4_X1 U6273 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n5305)
         );
  NAND2_X1 U6274 ( .A1(n6861), .A2(n5349), .ZN(n6863) );
  NAND2_X1 U6275 ( .A1(n5681), .A2(n8478), .ZN(n6884) );
  NOR2_X1 U6276 ( .A1(n6265), .A2(n6166), .ZN(n6271) );
  NAND2_X1 U6277 ( .A1(n7206), .A2(n9521), .ZN(n10606) );
  INV_X1 U6278 ( .A(n9463), .ZN(n9475) );
  INV_X1 U6279 ( .A(n6936), .ZN(n4893) );
  NAND2_X1 U6280 ( .A1(n5922), .A2(n5921), .ZN(n10449) );
  INV_X1 U6281 ( .A(n10449), .ZN(n4892) );
  INV_X1 U6282 ( .A(n9491), .ZN(n4855) );
  OR2_X1 U6283 ( .A1(n9510), .A2(n9468), .ZN(n4613) );
  AND2_X1 U6284 ( .A1(n4855), .A2(n9522), .ZN(n4614) );
  AND2_X1 U6285 ( .A1(n4857), .A2(n4583), .ZN(n4615) );
  OR2_X1 U6286 ( .A1(n9463), .A2(n4909), .ZN(n4616) );
  NAND2_X1 U6287 ( .A1(n4847), .A2(n7145), .ZN(n7285) );
  INV_X1 U6288 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5256) );
  INV_X1 U6289 ( .A(n6967), .ZN(n8516) );
  INV_X1 U6290 ( .A(n7290), .ZN(n4925) );
  INV_X1 U6291 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n4909) );
  NOR2_X1 U6292 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10346) );
  XNOR2_X1 U6293 ( .A(n7528), .B(n10585), .ZN(n10581) );
  NAND2_X1 U6294 ( .A1(n5764), .A2(n9711), .ZN(n5765) );
  AOI21_X1 U6295 ( .B1(n9557), .B2(n9711), .A(n9553), .ZN(n9674) );
  AND2_X1 U6296 ( .A1(n9550), .A2(n9711), .ZN(n5699) );
  AOI211_X2 U6297 ( .C1(n10223), .C2(n10520), .A(n10222), .B(n10221), .ZN(
        n10293) );
  INV_X1 U6298 ( .A(n5149), .ZN(n4931) );
  OAI21_X1 U6299 ( .B1(n9435), .B2(n4837), .A(n4836), .ZN(n9474) );
  NAND2_X1 U6300 ( .A1(n4843), .A2(n4844), .ZN(n9389) );
  NOR2_X1 U6301 ( .A1(n9391), .A2(n10603), .ZN(n9393) );
  NOR2_X1 U6302 ( .A1(n9492), .A2(n9491), .ZN(n9518) );
  OAI21_X1 U6303 ( .B1(n9515), .B2(n10606), .A(n4756), .ZN(n4755) );
  AOI21_X1 U6304 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9433), .A(n9432), .ZN(
        n9442) );
  NAND3_X1 U6305 ( .A1(n7051), .A2(n10571), .A3(n7064), .ZN(n4846) );
  NAND2_X2 U6306 ( .A1(n4617), .A2(n8756), .ZN(n7621) );
  NOR2_X1 U6307 ( .A1(n9964), .A2(n7492), .ZN(n7486) );
  NAND2_X2 U6308 ( .A1(n6194), .A2(n8818), .ZN(n10068) );
  NOR2_X1 U6309 ( .A1(n8167), .A2(n8168), .ZN(n8171) );
  NAND2_X1 U6310 ( .A1(n4596), .A2(n9510), .ZN(n9511) );
  NOR2_X1 U6311 ( .A1(n7969), .A2(n7970), .ZN(n7975) );
  NOR2_X1 U6312 ( .A1(n7175), .A2(n7174), .ZN(n7527) );
  INV_X1 U6313 ( .A(n9512), .ZN(n4758) );
  XNOR2_X1 U6314 ( .A(n7551), .B(n10585), .ZN(n10579) );
  NAND2_X1 U6315 ( .A1(n4758), .A2(n4568), .ZN(P2_U3200) );
  OAI21_X1 U6316 ( .B1(n7919), .B2(n8357), .A(n8358), .ZN(n8050) );
  AOI21_X1 U6317 ( .B1(n8357), .B2(n8358), .A(n4633), .ZN(n4632) );
  INV_X1 U6318 ( .A(n8362), .ZN(n4633) );
  OAI21_X1 U6319 ( .B1(n8478), .B2(n4636), .A(n8299), .ZN(n4635) );
  INV_X1 U6320 ( .A(n8281), .ZN(n5680) );
  NAND2_X1 U6321 ( .A1(n9732), .A2(n8281), .ZN(n6885) );
  NAND2_X1 U6322 ( .A1(n6862), .A2(n9725), .ZN(n8280) );
  NAND4_X1 U6323 ( .A1(n4643), .A2(n4644), .A3(n4919), .A4(n4642), .ZN(n5298)
         );
  INV_X1 U6324 ( .A(n4645), .ZN(n5362) );
  OAI21_X1 U6325 ( .B1(n5682), .B2(n7305), .A(n4646), .ZN(n7498) );
  NAND2_X1 U6326 ( .A1(n7934), .A2(n8353), .ZN(n4818) );
  NAND2_X2 U6327 ( .A1(n5668), .A2(n5669), .ZN(n6602) );
  AND2_X1 U6328 ( .A1(n4930), .A2(n5155), .ZN(n4659) );
  NAND2_X1 U6329 ( .A1(n5150), .A2(n4659), .ZN(n4662) );
  NAND2_X1 U6330 ( .A1(n6630), .A2(n8438), .ZN(n4673) );
  OR2_X1 U6331 ( .A1(n5050), .A2(n4676), .ZN(n4679) );
  NAND3_X1 U6332 ( .A1(n4679), .A2(n6393), .A3(n4677), .ZN(n7835) );
  NAND3_X1 U6333 ( .A1(n5054), .A2(n6353), .A3(n4678), .ZN(n4677) );
  NAND3_X1 U6334 ( .A1(n5054), .A2(n6353), .A3(n7359), .ZN(n4680) );
  NAND4_X1 U6335 ( .A1(n4684), .A2(n4682), .A3(n4681), .A4(n5066), .ZN(n6157)
         );
  INV_X1 U6336 ( .A(n6157), .ZN(n6162) );
  INV_X1 U6337 ( .A(n6167), .ZN(n4685) );
  INV_X1 U6338 ( .A(n4687), .ZN(n6213) );
  INV_X1 U6341 ( .A(n4696), .ZN(n8385) );
  OAI21_X1 U6342 ( .B1(n4821), .B2(n4820), .A(n4558), .ZN(n8380) );
  NAND3_X1 U6343 ( .A1(n4709), .A2(n8495), .A3(n4708), .ZN(n8356) );
  NAND3_X1 U6344 ( .A1(n8634), .A2(n8635), .A3(n8639), .ZN(n4724) );
  OAI21_X1 U6345 ( .B1(n4725), .B2(n8640), .A(n4723), .ZN(n4726) );
  OAI21_X1 U6346 ( .B1(n4567), .B2(n4729), .A(n4727), .ZN(n8724) );
  NAND2_X1 U6347 ( .A1(n8711), .A2(n8710), .ZN(n4734) );
  INV_X1 U6348 ( .A(n5134), .ZN(n5334) );
  NAND2_X1 U6349 ( .A1(n4743), .A2(n4593), .ZN(n8709) );
  NAND2_X1 U6350 ( .A1(n4744), .A2(n8851), .ZN(n4743) );
  NAND2_X1 U6351 ( .A1(n8695), .A2(n8701), .ZN(n8704) );
  XNOR2_X1 U6352 ( .A(n5361), .B(n5360), .ZN(n6616) );
  NAND2_X1 U6353 ( .A1(n5258), .A2(n5084), .ZN(n5085) );
  INV_X1 U6354 ( .A(n5086), .ZN(n5375) );
  MUX2_X1 U6355 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n8521), .Z(n7207) );
  MUX2_X1 U6356 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n8521), .Z(n7049) );
  NAND4_X1 U6357 ( .A1(n5779), .A2(n5780), .A3(n4686), .A4(n5818), .ZN(n4759)
         );
  NAND4_X1 U6358 ( .A1(n4761), .A2(n6158), .A3(n6224), .A4(n6160), .ZN(n4760)
         );
  OAI21_X1 U6359 ( .B1(n8733), .B2(n8732), .A(n5121), .ZN(n4771) );
  NAND3_X1 U6360 ( .A1(n4775), .A2(n8633), .A3(n4774), .ZN(n4773) );
  OAI21_X1 U6361 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8640) );
  NAND2_X1 U6362 ( .A1(n8717), .A2(n4783), .ZN(n4787) );
  NAND3_X1 U6363 ( .A1(n4787), .A2(n8725), .A3(n4786), .ZN(n8722) );
  NAND3_X1 U6364 ( .A1(n4788), .A2(n4794), .A3(n4789), .ZN(n4786) );
  NAND2_X1 U6365 ( .A1(n8720), .A2(n4796), .ZN(n4795) );
  INV_X1 U6366 ( .A(n9576), .ZN(n4799) );
  NAND2_X1 U6367 ( .A1(n9576), .A2(n4556), .ZN(n4805) );
  NAND2_X1 U6368 ( .A1(n4810), .A2(n4813), .ZN(n9793) );
  NAND2_X1 U6369 ( .A1(n4814), .A2(n4815), .ZN(n8517) );
  NAND3_X1 U6370 ( .A1(n8471), .A2(n8469), .A3(n4817), .ZN(n4814) );
  NAND3_X1 U6371 ( .A1(n8366), .A2(n8370), .A3(n8369), .ZN(n4820) );
  XNOR2_X1 U6372 ( .A(n9442), .B(n9456), .ZN(n9435) );
  INV_X1 U6373 ( .A(n4841), .ZN(n4844) );
  OAI21_X1 U6374 ( .B1(n8160), .B2(P2_REG1_REG_11__SCAN_IN), .A(n4845), .ZN(
        n4841) );
  NAND2_X1 U6375 ( .A1(n4842), .A2(n8120), .ZN(n4843) );
  INV_X1 U6376 ( .A(n8160), .ZN(n4842) );
  NOR2_X1 U6377 ( .A1(n8120), .A2(n8119), .ZN(n8161) );
  NAND2_X1 U6378 ( .A1(n7287), .A2(n7285), .ZN(n7154) );
  NAND3_X1 U6379 ( .A1(n7285), .A2(n4846), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n7287) );
  NAND2_X1 U6380 ( .A1(n10571), .A2(n7064), .ZN(n4847) );
  OAI211_X1 U6381 ( .C1(n9489), .C2(n4851), .A(n4849), .B(n4848), .ZN(n9537)
         );
  NAND2_X1 U6382 ( .A1(n9489), .A2(n4614), .ZN(n4848) );
  OAI21_X1 U6383 ( .B1(n4854), .B2(n9522), .A(n4850), .ZN(n4849) );
  NAND2_X1 U6384 ( .A1(n4854), .A2(n4852), .ZN(n4850) );
  NOR2_X1 U6385 ( .A1(n9489), .A2(n9490), .ZN(n9492) );
  INV_X1 U6386 ( .A(n4857), .ZN(n7267) );
  NAND4_X1 U6387 ( .A1(n5262), .A2(n5260), .A3(n5261), .A4(n5259), .ZN(n5703)
         );
  NAND2_X1 U6388 ( .A1(n9592), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U6389 ( .A1(n4859), .A2(n4864), .ZN(n5623) );
  OR2_X1 U6390 ( .A1(n9592), .A2(n5597), .ZN(n4868) );
  NAND2_X1 U6391 ( .A1(n7036), .A2(n4875), .ZN(n7307) );
  NAND2_X1 U6392 ( .A1(n5352), .A2(n7011), .ZN(n7090) );
  AOI21_X1 U6393 ( .B1(n5762), .B2(n9730), .A(n5761), .ZN(n8906) );
  OAI22_X2 U6394 ( .A1(n8048), .A2(n8496), .B1(n8563), .B2(n8200), .ZN(n8084)
         );
  OAI21_X1 U6395 ( .B1(n9757), .B2(n9571), .A(n5623), .ZN(n6255) );
  OAI21_X1 U6396 ( .B1(n7090), .B2(n7321), .A(n7320), .ZN(n5368) );
  OAI22_X2 U6397 ( .A1(n9602), .A2(n8476), .B1(n9372), .B2(n9607), .ZN(n9592)
         );
  NAND2_X1 U6398 ( .A1(n6888), .A2(n5351), .ZN(n7011) );
  OAI22_X1 U6399 ( .A1(n5747), .A2(n5746), .B1(n8912), .B2(n9548), .ZN(n5756)
         );
  AOI22_X2 U6400 ( .A1(n7920), .A2(n5505), .B1(n8240), .B2(n7927), .ZN(n8048)
         );
  INV_X1 U6401 ( .A(n7116), .ZN(n5303) );
  AND3_X2 U6402 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n7116) );
  INV_X1 U6403 ( .A(n8483), .ZN(n8299) );
  NAND2_X1 U6404 ( .A1(n4890), .A2(n4889), .ZN(n7647) );
  NAND2_X1 U6405 ( .A1(n7610), .A2(n4895), .ZN(n7873) );
  INV_X1 U6406 ( .A(n4900), .ZN(n10434) );
  NAND2_X1 U6407 ( .A1(n9536), .A2(n4901), .ZN(P2_U3201) );
  NAND2_X1 U6408 ( .A1(n4902), .A2(n10575), .ZN(n4901) );
  INV_X1 U6409 ( .A(n9537), .ZN(n4902) );
  OR2_X1 U6410 ( .A1(n10570), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4904) );
  XNOR2_X2 U6411 ( .A(n5325), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10570) );
  INV_X1 U6412 ( .A(n4911), .ZN(n9457) );
  INV_X1 U6413 ( .A(n9458), .ZN(n4910) );
  INV_X1 U6414 ( .A(n9508), .ZN(n4915) );
  OR2_X1 U6415 ( .A1(n9467), .A2(n9468), .ZN(n4916) );
  INV_X1 U6416 ( .A(n4916), .ZN(n9509) );
  OAI21_X1 U6417 ( .B1(n7292), .B2(n4925), .A(n4923), .ZN(n7167) );
  OAI22_X1 U6418 ( .A1(n7292), .A2(n4921), .B1(n4923), .B2(n7148), .ZN(n7170)
         );
  OAI21_X1 U6419 ( .B1(n5150), .B2(n4927), .A(n4926), .ZN(n5380) );
  AOI21_X1 U6420 ( .B1(n4931), .B2(n5360), .A(n4547), .ZN(n4926) );
  INV_X1 U6421 ( .A(n4929), .ZN(n4928) );
  OAI21_X1 U6422 ( .B1(n5360), .B2(n4547), .A(n5153), .ZN(n4929) );
  NOR2_X1 U6423 ( .A1(n4547), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U6424 ( .A1(n5599), .A2(n4945), .ZN(n4943) );
  NAND2_X1 U6425 ( .A1(n5599), .A2(n5598), .ZN(n4944) );
  OR2_X1 U6426 ( .A1(n5477), .A2(n5476), .ZN(n4960) );
  NAND2_X1 U6427 ( .A1(n4948), .A2(n4594), .ZN(n5203) );
  NAND2_X1 U6428 ( .A1(n5477), .A2(n4954), .ZN(n4948) );
  NAND2_X1 U6429 ( .A1(n4960), .A2(n4958), .ZN(n4953) );
  NAND2_X1 U6430 ( .A1(n4960), .A2(n5188), .ZN(n5491) );
  NAND2_X1 U6431 ( .A1(n5219), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U6432 ( .A1(n4961), .A2(n4965), .ZN(n5233) );
  NAND2_X1 U6433 ( .A1(n7605), .A2(n8755), .ZN(n7604) );
  AND2_X1 U6434 ( .A1(n4973), .A2(n8830), .ZN(n7605) );
  OAI21_X2 U6435 ( .B1(n7855), .B2(n8762), .A(n8687), .ZN(n8059) );
  NAND2_X1 U6436 ( .A1(n7621), .A2(n4978), .ZN(n4977) );
  NAND2_X1 U6437 ( .A1(n4977), .A2(n4572), .ZN(n6181) );
  NAND2_X1 U6438 ( .A1(n10068), .A2(n4595), .ZN(n4983) );
  OAI211_X1 U6439 ( .C1(n10068), .C2(n4986), .A(n4984), .B(n4983), .ZN(n6204)
         );
  XNOR2_X1 U6440 ( .A(n5397), .B(n5398), .ZN(n6627) );
  NAND2_X1 U6441 ( .A1(n8201), .A2(n4992), .ZN(n4991) );
  NAND2_X2 U6442 ( .A1(n4991), .A2(n4990), .ZN(n10185) );
  NAND2_X1 U6443 ( .A1(n10185), .A2(n10189), .ZN(n6188) );
  NAND2_X1 U6444 ( .A1(n4994), .A2(n7481), .ZN(n7484) );
  NAND2_X1 U6445 ( .A1(n10431), .A2(n4999), .ZN(n4995) );
  OAI21_X1 U6446 ( .B1(n10431), .B2(n10430), .A(n5004), .ZN(n7865) );
  OAI211_X1 U6447 ( .C1(n5006), .C2(n5008), .A(n5005), .B(n4545), .ZN(n7672)
         );
  NAND3_X1 U6448 ( .A1(n7247), .A2(n5943), .A3(n5956), .ZN(n5005) );
  NOR2_X1 U6449 ( .A1(n5116), .A2(n4592), .ZN(n5008) );
  NAND2_X1 U6450 ( .A1(n5009), .A2(n5008), .ZN(n7634) );
  OAI21_X1 U6451 ( .B1(n10123), .B2(n5011), .A(n5010), .ZN(n10076) );
  NAND2_X1 U6452 ( .A1(n10123), .A2(n5016), .ZN(n5012) );
  AOI21_X1 U6453 ( .B1(n10123), .B2(n6106), .A(n5019), .ZN(n10107) );
  AOI21_X2 U6454 ( .B1(n5024), .B2(n5023), .A(n5022), .ZN(n10175) );
  NAND2_X1 U6455 ( .A1(n5027), .A2(n5026), .ZN(n7505) );
  AND2_X1 U6456 ( .A1(n5781), .A2(n5034), .ZN(n5032) );
  AND2_X1 U6457 ( .A1(n5781), .A2(n5782), .ZN(n5033) );
  NAND2_X1 U6458 ( .A1(n4511), .A2(n5032), .ZN(n5800) );
  NOR2_X2 U6459 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5871) );
  NAND2_X1 U6460 ( .A1(n5871), .A2(n5035), .ZN(n5898) );
  INV_X1 U6461 ( .A(n5049), .ZN(n9881) );
  NAND2_X1 U6462 ( .A1(n9841), .A2(n4534), .ZN(n5057) );
  AND2_X1 U6463 ( .A1(n6321), .A2(n6316), .ZN(n5061) );
  NAND2_X2 U6464 ( .A1(n6871), .A2(n6872), .ZN(n6870) );
  NAND2_X1 U6465 ( .A1(n4684), .A2(n5769), .ZN(n5914) );
  NAND3_X1 U6466 ( .A1(n6334), .A2(n6345), .A3(n7343), .ZN(n10418) );
  NAND2_X1 U6467 ( .A1(n6334), .A2(n7343), .ZN(n10415) );
  NAND3_X1 U6468 ( .A1(n6455), .A2(n4607), .A3(n6454), .ZN(n9822) );
  NAND2_X1 U6469 ( .A1(n6455), .A2(n6454), .ZN(n9870) );
  NAND2_X1 U6470 ( .A1(n9822), .A2(n6467), .ZN(n6471) );
  NAND2_X1 U6471 ( .A1(n5272), .A2(n5271), .ZN(n5274) );
  INV_X1 U6472 ( .A(n8028), .ZN(n5072) );
  OR2_X1 U6473 ( .A1(n7845), .A2(n7899), .ZN(n5073) );
  NAND2_X1 U6474 ( .A1(n5070), .A2(n5068), .ZN(n8238) );
  NAND3_X1 U6475 ( .A1(n5072), .A2(n5074), .A3(n7899), .ZN(n5069) );
  INV_X1 U6476 ( .A(n7899), .ZN(n5078) );
  NAND2_X1 U6477 ( .A1(n8576), .A2(n5081), .ZN(n5080) );
  NAND3_X1 U6478 ( .A1(n4919), .A2(n4642), .A3(n4644), .ZN(n5312) );
  INV_X1 U6479 ( .A(n5258), .ZN(n5550) );
  INV_X1 U6480 ( .A(n8563), .ZN(n5094) );
  NAND3_X1 U6481 ( .A1(n6992), .A2(n5098), .A3(n7317), .ZN(n5095) );
  AND2_X1 U6482 ( .A1(n6993), .A2(n6991), .ZN(n5098) );
  OR2_X1 U6483 ( .A1(n9314), .A2(n5109), .ZN(n5099) );
  NAND2_X1 U6484 ( .A1(n9314), .A2(n5104), .ZN(n5103) );
  NAND2_X1 U6485 ( .A1(n9314), .A2(n9315), .ZN(n5106) );
  NAND3_X1 U6486 ( .A1(n5102), .A2(n5107), .A3(n5109), .ZN(n5101) );
  INV_X1 U6487 ( .A(n8596), .ZN(n5111) );
  NAND2_X1 U6488 ( .A1(n5880), .A2(n5879), .ZN(n6174) );
  AND2_X1 U6489 ( .A1(n5317), .A2(n7010), .ZN(n5352) );
  NAND2_X1 U6490 ( .A1(n6889), .A2(n6890), .ZN(n6888) );
  NAND2_X1 U6491 ( .A1(n5680), .A2(n5350), .ZN(n6889) );
  NAND2_X1 U6492 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  OR2_X1 U6493 ( .A1(n8299), .A2(n7012), .ZN(n7010) );
  NAND2_X1 U6494 ( .A1(n10287), .A2(n10537), .ZN(n8887) );
  NAND2_X1 U6495 ( .A1(n6157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U6496 ( .A1(n5908), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5850) );
  AND2_X2 U6497 ( .A1(n8883), .A2(n8545), .ZN(n5908) );
  NAND2_X1 U6498 ( .A1(n8536), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5870) );
  INV_X1 U6499 ( .A(n8536), .ZN(n6152) );
  CLKBUF_X1 U6500 ( .A(n7480), .Z(n8741) );
  INV_X1 U6501 ( .A(n6271), .ZN(n6276) );
  AND2_X2 U6502 ( .A1(n8897), .A2(n9802), .ZN(n5341) );
  NAND2_X1 U6503 ( .A1(n5786), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U6504 ( .A1(n7125), .A2(n5919), .ZN(n7247) );
  AND2_X1 U6505 ( .A1(n6980), .A2(n9725), .ZN(n6981) );
  INV_X1 U6506 ( .A(n5305), .ZN(n5304) );
  INV_X1 U6507 ( .A(n10094), .ZN(n10079) );
  NAND2_X2 U6508 ( .A1(n5960), .A2(n5959), .ZN(n10486) );
  AND2_X1 U6509 ( .A1(n6681), .A2(n8142), .ZN(n10033) );
  CLKBUF_X1 U6510 ( .A(n6197), .Z(n8893) );
  OR2_X1 U6511 ( .A1(n10652), .A2(n9716), .ZN(n9789) );
  INV_X1 U6512 ( .A(n9789), .ZN(n6261) );
  INV_X2 U6513 ( .A(n10652), .ZN(n10649) );
  AND3_X2 U6514 ( .A1(n6840), .A2(n6585), .A3(n6584), .ZN(n9744) );
  AND2_X1 U6515 ( .A1(n5456), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5112) );
  NOR2_X1 U6516 ( .A1(n5550), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5113) );
  AND2_X1 U6517 ( .A1(n5657), .A2(n5656), .ZN(n5114) );
  INV_X1 U6518 ( .A(n9646), .ZN(n6257) );
  INV_X2 U6519 ( .A(n10629), .ZN(n10632) );
  AND4_X1 U6520 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n7856)
         );
  AND4_X1 U6521 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n8554)
         );
  INV_X1 U6522 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5803) );
  OR2_X1 U6523 ( .A1(n6031), .A2(n6030), .ZN(n9947) );
  INV_X1 U6524 ( .A(n9947), .ZN(n8675) );
  INV_X1 U6525 ( .A(n6971), .ZN(n5698) );
  AND2_X1 U6526 ( .A1(n10652), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5115) );
  NOR2_X1 U6527 ( .A1(n5942), .A2(n7370), .ZN(n5116) );
  NOR2_X1 U6528 ( .A1(n7583), .A2(n4548), .ZN(n5117) );
  INV_X1 U6529 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5656) );
  AND2_X1 U6530 ( .A1(n5829), .A2(n5828), .ZN(n6441) );
  INV_X1 U6531 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5469) );
  OR2_X1 U6532 ( .A1(n7647), .A2(n10477), .ZN(n5118) );
  AND2_X1 U6533 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5119) );
  AND2_X2 U6534 ( .A1(n6250), .A2(n7407), .ZN(n10537) );
  AND2_X1 U6535 ( .A1(n10053), .A2(n8889), .ZN(n5120) );
  OR2_X1 U6536 ( .A1(n8802), .A2(n8737), .ZN(n5121) );
  NOR2_X1 U6537 ( .A1(n7579), .A2(n4672), .ZN(n5122) );
  NAND2_X1 U6538 ( .A1(n8713), .A2(n8712), .ZN(n5123) );
  AND2_X1 U6539 ( .A1(n5744), .A2(n5743), .ZN(n5124) );
  XNOR2_X1 U6540 ( .A(n6245), .B(n8774), .ZN(n10058) );
  AND2_X1 U6541 ( .A1(n7031), .A2(n9737), .ZN(n9718) );
  NAND2_X1 U6542 ( .A1(n8625), .A2(n8629), .ZN(n8626) );
  AND2_X1 U6543 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  NAND2_X1 U6544 ( .A1(n8642), .A2(n8737), .ZN(n8643) );
  NOR2_X1 U6545 ( .A1(n8659), .A2(n8832), .ZN(n8661) );
  AOI21_X1 U6546 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8665) );
  NAND2_X1 U6547 ( .A1(n8668), .A2(n8629), .ZN(n8669) );
  NAND2_X1 U6548 ( .A1(n8692), .A2(n8629), .ZN(n8693) );
  INV_X1 U6549 ( .A(n8714), .ZN(n8715) );
  NAND2_X1 U6550 ( .A1(n5123), .A2(n8715), .ZN(n8716) );
  INV_X1 U6551 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5773) );
  INV_X1 U6552 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5248) );
  INV_X1 U6553 ( .A(n6174), .ZN(n8623) );
  INV_X1 U6554 ( .A(n6972), .ZN(n6973) );
  NAND2_X1 U6555 ( .A1(n7891), .A2(n9382), .ZN(n7888) );
  INV_X1 U6556 ( .A(n8165), .ZN(n8166) );
  AND2_X1 U6557 ( .A1(n9652), .A2(n9375), .ZN(n5564) );
  INV_X1 U6558 ( .A(n6441), .ZN(n6059) );
  INV_X1 U6559 ( .A(n7417), .ZN(n5879) );
  AND3_X1 U6560 ( .A1(n6160), .A2(n6159), .A3(n6158), .ZN(n6161) );
  INV_X1 U6561 ( .A(n8554), .ZN(n8240) );
  NAND2_X1 U6562 ( .A1(n8514), .A2(n6970), .ZN(n8515) );
  INV_X1 U6563 ( .A(n9409), .ZN(n9410) );
  INV_X1 U6564 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9192) );
  OR2_X1 U6565 ( .A1(n5432), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5443) );
  INV_X1 U6566 ( .A(n6887), .ZN(n8478) );
  AND2_X1 U6567 ( .A1(n5792), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5948) );
  INV_X1 U6568 ( .A(n7229), .ZN(n6321) );
  OR2_X1 U6569 ( .A1(n4527), .A2(n7492), .ZN(n6284) );
  INV_X1 U6570 ( .A(n6077), .ZN(n6075) );
  OR2_X1 U6571 ( .A1(n6065), .A2(n6064), .ZN(n6077) );
  AND2_X1 U6572 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  NAND2_X1 U6573 ( .A1(n9962), .A2(n7417), .ZN(n8824) );
  INV_X1 U6574 ( .A(P1_B_REG_SCAN_IN), .ZN(n6211) );
  INV_X1 U6575 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5782) );
  AND2_X1 U6576 ( .A1(n5801), .A2(n5779), .ZN(n6214) );
  INV_X1 U6577 ( .A(SI_19_), .ZN(n5204) );
  INV_X1 U6578 ( .A(SI_16_), .ZN(n5193) );
  NOR2_X1 U6579 ( .A1(n5634), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U6580 ( .A1(n7842), .A2(n4672), .ZN(n7844) );
  NAND2_X1 U6581 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  INV_X1 U6582 ( .A(n9324), .ZN(n8575) );
  INV_X1 U6583 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5271) );
  OR2_X1 U6584 ( .A1(n5579), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U6585 ( .A1(n5570), .A2(n5569), .ZN(n5579) );
  INV_X1 U6586 ( .A(n7554), .ZN(n7556) );
  INV_X1 U6587 ( .A(n7992), .ZN(n7990) );
  NAND2_X1 U6588 ( .A1(n9477), .A2(n9476), .ZN(n9478) );
  XNOR2_X1 U6589 ( .A(n9507), .B(n9488), .ZN(n9477) );
  NAND2_X1 U6590 ( .A1(n5470), .A2(n5469), .ZN(n5483) );
  INV_X1 U6591 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5354) );
  INV_X1 U6592 ( .A(n8901), .ZN(n5764) );
  NAND2_X1 U6593 ( .A1(n8305), .A2(n8313), .ZN(n8482) );
  AND2_X1 U6594 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  OR2_X1 U6595 ( .A1(n6120), .A2(n9913), .ZN(n6141) );
  AND2_X1 U6596 ( .A1(n6141), .A2(n6121), .ZN(n10096) );
  INV_X1 U6597 ( .A(n10159), .ZN(n6206) );
  NOR2_X1 U6598 ( .A1(n10061), .A2(n10273), .ZN(n6555) );
  OR2_X1 U6599 ( .A1(n10080), .A2(n9936), .ZN(n6135) );
  OR2_X1 U6600 ( .A1(n7957), .A2(n6211), .ZN(n6218) );
  AND2_X1 U6601 ( .A1(n5544), .A2(n5210), .ZN(n5214) );
  OR3_X1 U6602 ( .A1(n5971), .A2(P1_IR_REG_11__SCAN_IN), .A3(
        P1_IR_REG_10__SCAN_IN), .ZN(n5995) );
  INV_X1 U6603 ( .A(n5410), .ZN(n5165) );
  NAND2_X1 U6604 ( .A1(n5788), .A2(n6608), .ZN(n5138) );
  AND2_X1 U6605 ( .A1(n7471), .A2(n7472), .ZN(n7470) );
  OR2_X1 U6606 ( .A1(n6962), .A2(n6961), .ZN(n9327) );
  NOR2_X1 U6607 ( .A1(n10597), .A2(n10400), .ZN(n9483) );
  INV_X1 U6608 ( .A(n9366), .ZN(n8912) );
  INV_X1 U6609 ( .A(n9367), .ZN(n9562) );
  INV_X1 U6610 ( .A(n8476), .ZN(n9605) );
  NOR2_X1 U6611 ( .A1(n5558), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5559) );
  AND2_X1 U6612 ( .A1(n8363), .A2(n8362), .ZN(n8496) );
  NAND2_X1 U6613 ( .A1(n5418), .A2(n5417), .ZN(n5432) );
  AND2_X1 U6614 ( .A1(n8320), .A2(n8325), .ZN(n8485) );
  OR2_X1 U6615 ( .A1(n9716), .A2(n5698), .ZN(n10622) );
  NAND2_X1 U6616 ( .A1(n6961), .A2(n8448), .ZN(n9646) );
  INV_X1 U6617 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5664) );
  INV_X1 U6618 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7820) );
  AND2_X1 U6619 ( .A1(n6510), .A2(n6509), .ZN(n6559) );
  AND2_X1 U6620 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5905) );
  AND2_X1 U6621 ( .A1(n5905), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5923) );
  INV_X1 U6622 ( .A(n8537), .ZN(n6124) );
  INV_X1 U6623 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6821) );
  INV_X1 U6624 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7190) );
  AND2_X1 U6625 ( .A1(n7802), .A2(n7728), .ZN(n7729) );
  INV_X1 U6626 ( .A(n8533), .ZN(n10042) );
  INV_X1 U6627 ( .A(n10156), .ZN(n10176) );
  AND2_X1 U6628 ( .A1(n8712), .A2(n6187), .ZN(n10189) );
  INV_X1 U6629 ( .A(n8766), .ZN(n8208) );
  AND2_X1 U6630 ( .A1(n9848), .A2(n9946), .ZN(n6045) );
  NAND2_X1 U6631 ( .A1(n6272), .A2(n6166), .ZN(n7493) );
  OR2_X1 U6632 ( .A1(n7436), .A2(n8871), .ZN(n10502) );
  INV_X1 U6633 ( .A(n8744), .ZN(n6852) );
  AND2_X1 U6634 ( .A1(n5202), .A2(n5201), .ZN(n5520) );
  OAI21_X1 U6635 ( .B1(n5451), .B2(n5180), .A(n5179), .ZN(n5463) );
  INV_X1 U6636 ( .A(n9327), .ZN(n9354) );
  AND4_X1 U6637 ( .A1(n8446), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n8607)
         );
  AOI21_X1 U6638 ( .B1(n9608), .B2(n4523), .A(n5583), .ZN(n9616) );
  AND4_X1 U6639 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n8074)
         );
  INV_X1 U6640 ( .A(n10597), .ZN(n7301) );
  INV_X1 U6641 ( .A(n10598), .ZN(n10586) );
  AND2_X1 U6642 ( .A1(n7206), .A2(n8521), .ZN(n10566) );
  AND2_X1 U6643 ( .A1(n8220), .A2(n8219), .ZN(n9712) );
  INV_X1 U6644 ( .A(n8900), .ZN(n9657) );
  AND2_X2 U6645 ( .A1(n6952), .A2(n6841), .ZN(n10628) );
  AND2_X1 U6646 ( .A1(n6952), .A2(n6578), .ZN(n6840) );
  NAND2_X1 U6647 ( .A1(n7816), .A2(n6970), .ZN(n9716) );
  INV_X1 U6648 ( .A(n9716), .ZN(n9739) );
  INV_X1 U6649 ( .A(n9718), .ZN(n9711) );
  OR3_X1 U6650 ( .A1(n8009), .A2(n5735), .A3(n8070), .ZN(n7057) );
  INV_X1 U6651 ( .A(n5719), .ZN(n6645) );
  INV_X1 U6652 ( .A(n6549), .ZN(n6550) );
  INV_X1 U6653 ( .A(n9908), .ZN(n9865) );
  INV_X1 U6654 ( .A(n9931), .ZN(n10421) );
  AND2_X1 U6655 ( .A1(n6531), .A2(n6526), .ZN(n9922) );
  AND2_X1 U6656 ( .A1(n5817), .A2(n5816), .ZN(n9826) );
  OR2_X1 U6657 ( .A1(n6739), .A2(n8874), .ZN(n7948) );
  INV_X1 U6658 ( .A(n7948), .ZN(n10025) );
  INV_X1 U6659 ( .A(n8893), .ZN(n6665) );
  NOR2_X1 U6660 ( .A1(n10537), .A2(n6241), .ZN(n6242) );
  NOR2_X1 U6661 ( .A1(n10534), .A2(n10517), .ZN(n8889) );
  OAI22_X1 U6662 ( .A1(n10061), .A2(n10329), .B1(n10523), .B2(n6252), .ZN(
        n6253) );
  NAND2_X1 U6663 ( .A1(n6220), .A2(n6239), .ZN(n10334) );
  NAND2_X1 U6664 ( .A1(n5137), .A2(n5136), .ZN(n5323) );
  INV_X1 U6665 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10381) );
  AND2_X1 U6666 ( .A1(n6990), .A2(n6989), .ZN(n9363) );
  NAND2_X1 U6667 ( .A1(n5641), .A2(n5640), .ZN(n9367) );
  INV_X1 U6668 ( .A(n9647), .ZN(n9374) );
  INV_X1 U6669 ( .A(n7892), .ZN(n9382) );
  OR2_X1 U6670 ( .A1(P2_U3150), .A2(n7058), .ZN(n10597) );
  AND2_X1 U6671 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  AND2_X1 U6672 ( .A1(n7088), .A2(n7087), .ZN(n7222) );
  AND2_X1 U6673 ( .A1(n7221), .A2(n7032), .ZN(n8900) );
  INV_X1 U6674 ( .A(n8601), .ZN(n9677) );
  INV_X1 U6675 ( .A(n9744), .ZN(n9743) );
  INV_X1 U6676 ( .A(n8936), .ZN(n9777) );
  AND2_X1 U6677 ( .A1(n5742), .A2(n5741), .ZN(n10652) );
  INV_X1 U6678 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9061) );
  INV_X1 U6679 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8272) );
  INV_X1 U6680 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6761) );
  INV_X1 U6681 ( .A(n7148), .ZN(n7279) );
  INV_X1 U6682 ( .A(n9916), .ZN(n10413) );
  INV_X1 U6683 ( .A(n9922), .ZN(n10416) );
  AND2_X1 U6684 ( .A1(n6530), .A2(n10190), .ZN(n9931) );
  INV_X1 U6685 ( .A(n9835), .ZN(n9937) );
  INV_X1 U6686 ( .A(n9826), .ZN(n9943) );
  INV_X1 U6687 ( .A(n10033), .ZN(n8109) );
  OR2_X1 U6688 ( .A1(n7413), .A2(n6166), .ZN(n10194) );
  INV_X1 U6689 ( .A(n10458), .ZN(n8158) );
  AND2_X1 U6690 ( .A1(n7413), .A2(n10190), .ZN(n10462) );
  NOR2_X1 U6691 ( .A1(n5120), .A2(n6242), .ZN(n6243) );
  INV_X1 U6692 ( .A(n8889), .ZN(n10273) );
  INV_X1 U6693 ( .A(n10537), .ZN(n10534) );
  INV_X1 U6694 ( .A(n10523), .ZN(n6596) );
  AND2_X1 U6695 ( .A1(n10484), .A2(n10483), .ZN(n10526) );
  AND2_X2 U6696 ( .A1(n6251), .A2(n6250), .ZN(n10523) );
  INV_X1 U6697 ( .A(n10469), .ZN(n10470) );
  INV_X1 U6698 ( .A(n6222), .ZN(n7885) );
  INV_X1 U6699 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7433) );
  INV_X1 U6700 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9269) );
  INV_X2 U6701 ( .A(n9500), .ZN(P2_U3893) );
  INV_X2 U6702 ( .A(n9942), .ZN(P1_U3973) );
  OAI21_X1 U6703 ( .B1(n6558), .B2(n6596), .A(n6254), .ZN(P1_U3518) );
  NAND2_X1 U6704 ( .A1(n10346), .A2(n5129), .ZN(n5130) );
  AND2_X1 U6705 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6706 ( .A1(n4518), .A2(n5132), .ZN(n5348) );
  AND2_X1 U6707 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6708 ( .A1(n4517), .A2(n5133), .ZN(n5864) );
  NAND2_X1 U6709 ( .A1(n5348), .A2(n5864), .ZN(n5335) );
  NAND2_X1 U6710 ( .A1(n5335), .A2(n5134), .ZN(n5137) );
  NAND2_X1 U6711 ( .A1(n5135), .A2(SI_1_), .ZN(n5136) );
  INV_X1 U6712 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6614) );
  INV_X1 U6713 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U6714 ( .A1(n5323), .A2(n5322), .ZN(n5142) );
  INV_X1 U6715 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6716 ( .A1(n5140), .A2(SI_2_), .ZN(n5141) );
  NAND2_X1 U6717 ( .A1(n5142), .A2(n5141), .ZN(n5311) );
  INV_X1 U6718 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6606) );
  INV_X1 U6719 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6611) );
  MUX2_X1 U6720 ( .A(n6606), .B(n6611), .S(n4518), .Z(n5143) );
  XNOR2_X1 U6721 ( .A(n5143), .B(SI_3_), .ZN(n5310) );
  NAND2_X1 U6722 ( .A1(n5311), .A2(n5310), .ZN(n5146) );
  INV_X1 U6723 ( .A(n5143), .ZN(n5144) );
  NAND2_X1 U6724 ( .A1(n5144), .A2(SI_3_), .ZN(n5145) );
  MUX2_X1 U6725 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5788), .Z(n5148) );
  INV_X1 U6726 ( .A(SI_4_), .ZN(n9195) );
  XNOR2_X1 U6727 ( .A(n5148), .B(n9195), .ZN(n5296) );
  NAND2_X1 U6728 ( .A1(n5148), .A2(SI_4_), .ZN(n5149) );
  INV_X1 U6729 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6615) );
  MUX2_X1 U6730 ( .A(n9234), .B(n6615), .S(n4517), .Z(n5151) );
  INV_X1 U6731 ( .A(n5151), .ZN(n5152) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4516), .Z(n5154) );
  XNOR2_X1 U6733 ( .A(n5154), .B(SI_6_), .ZN(n5379) );
  INV_X1 U6734 ( .A(n5379), .ZN(n5153) );
  NAND2_X1 U6735 ( .A1(n5154), .A2(SI_6_), .ZN(n5155) );
  MUX2_X1 U6736 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4517), .Z(n5156) );
  XNOR2_X1 U6737 ( .A(n5156), .B(SI_7_), .ZN(n5391) );
  NAND2_X1 U6738 ( .A1(n5156), .A2(SI_7_), .ZN(n5157) );
  INV_X1 U6739 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6628) );
  MUX2_X1 U6740 ( .A(n9206), .B(n6628), .S(n4516), .Z(n5159) );
  INV_X1 U6741 ( .A(SI_8_), .ZN(n5158) );
  NAND2_X1 U6742 ( .A1(n5159), .A2(n5158), .ZN(n5408) );
  INV_X1 U6743 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6744 ( .A1(n5160), .A2(SI_8_), .ZN(n5161) );
  NAND2_X1 U6745 ( .A1(n5408), .A2(n5161), .ZN(n5398) );
  MUX2_X1 U6746 ( .A(n6632), .B(n6631), .S(n4517), .Z(n5163) );
  INV_X1 U6747 ( .A(SI_9_), .ZN(n5162) );
  NAND2_X1 U6748 ( .A1(n5163), .A2(n5162), .ZN(n5411) );
  AND2_X1 U6749 ( .A1(n5408), .A2(n5411), .ZN(n5166) );
  INV_X1 U6750 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6751 ( .A1(n5164), .A2(SI_9_), .ZN(n5410) );
  MUX2_X1 U6752 ( .A(n8970), .B(n6639), .S(n4517), .Z(n5168) );
  XNOR2_X1 U6753 ( .A(n5168), .B(SI_10_), .ZN(n5424) );
  INV_X1 U6754 ( .A(n5424), .ZN(n5167) );
  INV_X1 U6755 ( .A(n5168), .ZN(n5169) );
  NAND2_X1 U6756 ( .A1(n5169), .A2(SI_10_), .ZN(n5170) );
  INV_X1 U6757 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5171) );
  MUX2_X1 U6758 ( .A(n5171), .B(n6735), .S(n4516), .Z(n5173) );
  INV_X1 U6759 ( .A(SI_11_), .ZN(n5172) );
  NAND2_X1 U6760 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
  INV_X1 U6761 ( .A(n5173), .ZN(n5174) );
  NAND2_X1 U6762 ( .A1(n5174), .A2(SI_11_), .ZN(n5175) );
  NAND2_X1 U6763 ( .A1(n5176), .A2(n5175), .ZN(n5438) );
  MUX2_X1 U6764 ( .A(n6761), .B(n6745), .S(n4517), .Z(n5177) );
  XNOR2_X1 U6765 ( .A(n5177), .B(SI_12_), .ZN(n5450) );
  INV_X1 U6766 ( .A(n5450), .ZN(n5180) );
  INV_X1 U6767 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6768 ( .A1(n5178), .A2(SI_12_), .ZN(n5179) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4516), .Z(n5182) );
  XNOR2_X1 U6770 ( .A(n5182), .B(SI_13_), .ZN(n5462) );
  INV_X1 U6771 ( .A(n5462), .ZN(n5181) );
  NAND2_X1 U6772 ( .A1(n5463), .A2(n5181), .ZN(n5184) );
  NAND2_X1 U6773 ( .A1(n5182), .A2(SI_13_), .ZN(n5183) );
  NAND2_X1 U6774 ( .A1(n5184), .A2(n5183), .ZN(n5477) );
  MUX2_X1 U6775 ( .A(n9278), .B(n9269), .S(n4516), .Z(n5185) );
  NAND2_X1 U6776 ( .A1(n5185), .A2(n9262), .ZN(n5188) );
  INV_X1 U6777 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6778 ( .A1(n5186), .A2(SI_14_), .ZN(n5187) );
  NAND2_X1 U6779 ( .A1(n5188), .A2(n5187), .ZN(n5476) );
  MUX2_X1 U6780 ( .A(n7097), .B(n7043), .S(n4516), .Z(n5189) );
  XNOR2_X1 U6781 ( .A(n5189), .B(SI_15_), .ZN(n5490) );
  INV_X1 U6782 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6783 ( .A1(n5190), .A2(SI_15_), .ZN(n5191) );
  MUX2_X1 U6784 ( .A(n7215), .B(n7214), .S(n4516), .Z(n5194) );
  NAND2_X1 U6785 ( .A1(n5194), .A2(n5193), .ZN(n5197) );
  INV_X1 U6786 ( .A(n5194), .ZN(n5195) );
  NAND2_X1 U6787 ( .A1(n5195), .A2(SI_16_), .ZN(n5196) );
  NAND2_X1 U6788 ( .A1(n5197), .A2(n5196), .ZN(n5506) );
  MUX2_X1 U6789 ( .A(n7259), .B(n7261), .S(n4517), .Z(n5199) );
  NAND2_X1 U6790 ( .A1(n5199), .A2(n5198), .ZN(n5202) );
  INV_X1 U6791 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6792 ( .A1(n5200), .A2(SI_17_), .ZN(n5201) );
  NAND2_X1 U6793 ( .A1(n5203), .A2(n5202), .ZN(n5534) );
  INV_X1 U6794 ( .A(n5534), .ZN(n5545) );
  MUX2_X1 U6795 ( .A(n7315), .B(n7338), .S(n4516), .Z(n5205) );
  XNOR2_X1 U6796 ( .A(n5205), .B(SI_18_), .ZN(n5544) );
  MUX2_X1 U6797 ( .A(n9197), .B(n7433), .S(n4517), .Z(n5207) );
  NAND2_X1 U6798 ( .A1(n5207), .A2(n5204), .ZN(n5210) );
  INV_X1 U6799 ( .A(n5210), .ZN(n5213) );
  INV_X1 U6800 ( .A(n5205), .ZN(n5206) );
  NAND2_X1 U6801 ( .A1(n5206), .A2(SI_18_), .ZN(n5546) );
  INV_X1 U6802 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U6803 ( .A1(n5208), .A2(SI_19_), .ZN(n5209) );
  NAND2_X1 U6804 ( .A1(n5210), .A2(n5209), .ZN(n5548) );
  INV_X1 U6805 ( .A(n5548), .ZN(n5211) );
  MUX2_X1 U6806 ( .A(n8272), .B(n7405), .S(n4517), .Z(n5215) );
  NAND2_X1 U6807 ( .A1(n5215), .A2(n8947), .ZN(n5218) );
  INV_X1 U6808 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6809 ( .A1(n5216), .A2(SI_20_), .ZN(n5217) );
  NAND2_X1 U6810 ( .A1(n5284), .A2(n5283), .ZN(n5219) );
  MUX2_X1 U6811 ( .A(n7562), .B(n7524), .S(n4517), .Z(n5220) );
  XNOR2_X1 U6812 ( .A(n5220), .B(SI_21_), .ZN(n5565) );
  INV_X1 U6813 ( .A(n5565), .ZN(n5223) );
  INV_X1 U6814 ( .A(n5220), .ZN(n5221) );
  NAND2_X1 U6815 ( .A1(n5221), .A2(SI_21_), .ZN(n5222) );
  MUX2_X1 U6816 ( .A(n7814), .B(n7813), .S(n4516), .Z(n5224) );
  INV_X1 U6817 ( .A(SI_22_), .ZN(n8959) );
  NAND2_X1 U6818 ( .A1(n5224), .A2(n8959), .ZN(n5227) );
  INV_X1 U6819 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6820 ( .A1(n5225), .A2(SI_22_), .ZN(n5226) );
  NAND2_X1 U6821 ( .A1(n5227), .A2(n5226), .ZN(n5575) );
  MUX2_X1 U6822 ( .A(n7777), .B(n9285), .S(n4516), .Z(n5229) );
  INV_X1 U6823 ( .A(SI_23_), .ZN(n5228) );
  NAND2_X1 U6824 ( .A1(n5229), .A2(n5228), .ZN(n5232) );
  INV_X1 U6825 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6826 ( .A1(n5230), .A2(SI_23_), .ZN(n5231) );
  MUX2_X1 U6827 ( .A(n7886), .B(n7884), .S(n4517), .Z(n5235) );
  INV_X1 U6828 ( .A(SI_24_), .ZN(n5234) );
  NAND2_X1 U6829 ( .A1(n5235), .A2(n5234), .ZN(n5238) );
  INV_X1 U6830 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6831 ( .A1(n5236), .A2(SI_24_), .ZN(n5237) );
  INV_X1 U6832 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7958) );
  MUX2_X1 U6833 ( .A(n8964), .B(n7958), .S(n4516), .Z(n5240) );
  INV_X1 U6834 ( .A(SI_25_), .ZN(n5239) );
  NAND2_X1 U6835 ( .A1(n5240), .A2(n5239), .ZN(n5243) );
  INV_X1 U6836 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6837 ( .A1(n5241), .A2(SI_25_), .ZN(n5242) );
  MUX2_X1 U6838 ( .A(n9061), .B(n9258), .S(n4517), .Z(n5245) );
  INV_X1 U6839 ( .A(SI_26_), .ZN(n5244) );
  NAND2_X1 U6840 ( .A1(n5245), .A2(n5244), .ZN(n5626) );
  INV_X1 U6841 ( .A(n5245), .ZN(n5246) );
  NAND2_X1 U6842 ( .A1(n5246), .A2(SI_26_), .ZN(n5247) );
  XNOR2_X1 U6843 ( .A(n5625), .B(n5624), .ZN(n8055) );
  INV_X1 U6844 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5249) );
  NOR2_X1 U6845 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5253) );
  NOR2_X1 U6846 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5252) );
  NOR2_X1 U6847 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5251) );
  NOR2_X1 U6848 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5250) );
  NAND4_X1 U6849 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n5508)
         );
  NAND3_X1 U6850 ( .A1(n5256), .A2(n5255), .A3(n5254), .ZN(n5257) );
  INV_X1 U6851 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5263) );
  NOR2_X1 U6852 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5262) );
  NAND2_X1 U6853 ( .A1(n5270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6854 ( .A1(n8055), .A2(n8438), .ZN(n5268) );
  NAND2_X2 U6855 ( .A1(n6602), .A2(n4517), .ZN(n5333) );
  OR2_X1 U6856 ( .A1(n5333), .A2(n9061), .ZN(n5267) );
  NOR2_X1 U6857 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5353) );
  NAND2_X1 U6858 ( .A1(n5353), .A2(n5354), .ZN(n5369) );
  INV_X1 U6859 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5287) );
  INV_X1 U6860 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5569) );
  INV_X1 U6861 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6862 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  NAND2_X1 U6863 ( .A1(n5617), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6864 ( .A1(n5634), .A2(n5269), .ZN(n9565) );
  NAND2_X1 U6865 ( .A1(n5274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6866 ( .A1(n9565), .A2(n4523), .ZN(n5282) );
  INV_X1 U6867 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U6868 ( .A1(n4520), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6869 ( .A1(n4515), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5278) );
  OAI211_X1 U6870 ( .C1(n5638), .C2(n9755), .A(n5279), .B(n5278), .ZN(n5280)
         );
  INV_X1 U6871 ( .A(n5280), .ZN(n5281) );
  XNOR2_X1 U6872 ( .A(n5284), .B(n5283), .ZN(n8271) );
  NAND2_X1 U6873 ( .A1(n8271), .A2(n8438), .ZN(n5286) );
  OR2_X1 U6874 ( .A1(n5333), .A2(n8272), .ZN(n5285) );
  NOR2_X1 U6875 ( .A1(n5559), .A2(n5287), .ZN(n5288) );
  OR2_X1 U6876 ( .A1(n5570), .A2(n5288), .ZN(n9635) );
  NAND2_X1 U6877 ( .A1(n9635), .A2(n4522), .ZN(n5291) );
  AOI22_X1 U6878 ( .A1(n4519), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n4515), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6879 ( .A1(n4520), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6880 ( .A1(n4519), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6881 ( .A1(n5119), .A2(n5353), .ZN(n7114) );
  NAND2_X1 U6882 ( .A1(n4522), .A2(n7114), .ZN(n5293) );
  NAND2_X1 U6883 ( .A1(n8442), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5292) );
  INV_X1 U6884 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U6885 ( .A1(n5298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5299) );
  XNOR2_X1 U6886 ( .A(n5299), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U6887 ( .A1(n5554), .A2(n7165), .ZN(n5300) );
  NAND2_X1 U6888 ( .A1(n5304), .A2(n7116), .ZN(n5317) );
  NAND2_X1 U6889 ( .A1(n5305), .A2(n7116), .ZN(n8311) );
  NAND2_X1 U6890 ( .A1(n8302), .A2(n8311), .ZN(n8483) );
  INV_X1 U6891 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U6892 ( .A1(n4522), .A2(n6958), .ZN(n5309) );
  NAND2_X1 U6893 ( .A1(n4525), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6894 ( .A1(n8442), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6895 ( .A1(n4519), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5306) );
  XNOR2_X1 U6896 ( .A(n5311), .B(n5310), .ZN(n6612) );
  OR2_X1 U6897 ( .A1(n5336), .A2(n6612), .ZN(n5316) );
  OR2_X1 U6898 ( .A1(n5333), .A2(n6611), .ZN(n5315) );
  NAND2_X1 U6899 ( .A1(n5312), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6900 ( .A1(n5554), .A2(n7051), .ZN(n5314) );
  INV_X1 U6901 ( .A(n7108), .ZN(n6964) );
  OR2_X1 U6902 ( .A1(n9726), .A2(n6964), .ZN(n7012) );
  NAND2_X1 U6903 ( .A1(n4523), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6904 ( .A1(n8442), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6905 ( .A1(n4519), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6906 ( .A1(n5333), .A2(n6614), .ZN(n5328) );
  XNOR2_X1 U6907 ( .A(n5323), .B(n5322), .ZN(n6613) );
  OR2_X1 U6908 ( .A1(n5336), .A2(n6613), .ZN(n5327) );
  NAND2_X1 U6909 ( .A1(n5554), .A2(n10570), .ZN(n5326) );
  NAND2_X1 U6910 ( .A1(n9387), .A2(n10623), .ZN(n8293) );
  NAND2_X1 U6911 ( .A1(n8442), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6912 ( .A1(n5340), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5330) );
  OR2_X1 U6913 ( .A1(n5333), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6914 ( .A(n5334), .B(n5335), .ZN(n5855) );
  NAND2_X1 U6915 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5337) );
  NAND2_X1 U6916 ( .A1(n4515), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6917 ( .A1(n4523), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6918 ( .A1(n4519), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6919 ( .A1(n8442), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5342) );
  NAND4_X1 U6920 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n5679)
         );
  INV_X1 U6921 ( .A(SI_0_), .ZN(n5863) );
  INV_X1 U6922 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U6923 ( .B1(n4516), .B2(n5863), .A(n5346), .ZN(n5347) );
  AND2_X1 U6924 ( .A1(n5348), .A2(n5347), .ZN(n9803) );
  MUX2_X1 U6925 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9803), .S(n6602), .Z(n6976) );
  NAND2_X1 U6926 ( .A1(n5679), .A2(n6976), .ZN(n5349) );
  NAND2_X1 U6927 ( .A1(n7099), .A2(n6862), .ZN(n9722) );
  NAND2_X1 U6928 ( .A1(n6863), .A2(n9722), .ZN(n5350) );
  INV_X1 U6929 ( .A(n10623), .ZN(n9738) );
  OR2_X1 U6930 ( .A1(n9387), .A2(n9738), .ZN(n6890) );
  NAND2_X1 U6931 ( .A1(n9726), .A2(n7108), .ZN(n8301) );
  AND2_X1 U6932 ( .A1(n6887), .A2(n8483), .ZN(n5351) );
  NAND2_X1 U6933 ( .A1(n4515), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6934 ( .A1(n4520), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5358) );
  OR2_X1 U6935 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6936 ( .A1(n5369), .A2(n5355), .ZN(n9309) );
  NAND2_X1 U6937 ( .A1(n4523), .A2(n9309), .ZN(n5357) );
  NAND2_X1 U6938 ( .A1(n4519), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6939 ( .A1(n5336), .A2(n6616), .ZN(n5366) );
  OR2_X1 U6940 ( .A1(n5333), .A2(n9234), .ZN(n5365) );
  OR2_X1 U6941 ( .A1(n5362), .A2(n9792), .ZN(n5363) );
  XNOR2_X1 U6942 ( .A(n5363), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U6943 ( .A1(n5554), .A2(n7148), .ZN(n5364) );
  NAND2_X1 U6944 ( .A1(n7090), .A2(n7321), .ZN(n5367) );
  NAND2_X1 U6945 ( .A1(n5368), .A2(n5367), .ZN(n7035) );
  INV_X1 U6946 ( .A(n7035), .ZN(n5383) );
  NAND2_X1 U6947 ( .A1(n4519), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6948 ( .A1(n4525), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6949 ( .A1(n5369), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6950 ( .A1(n5385), .A2(n5370), .ZN(n9347) );
  NAND2_X1 U6951 ( .A1(n4523), .A2(n9347), .ZN(n5372) );
  NAND2_X1 U6952 ( .A1(n4520), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5371) );
  NAND4_X1 U6953 ( .A1(n5374), .A2(n5373), .A3(n5372), .A4(n5371), .ZN(n9385)
         );
  NAND2_X1 U6954 ( .A1(n5375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5376) );
  MUX2_X1 U6955 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5376), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5378) );
  AND2_X1 U6956 ( .A1(n5378), .A2(n5377), .ZN(n7172) );
  AOI22_X1 U6957 ( .A1(n5555), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5554), .B2(
        n7172), .ZN(n5382) );
  XNOR2_X1 U6958 ( .A(n5380), .B(n5379), .ZN(n6617) );
  NAND2_X1 U6959 ( .A1(n6617), .A2(n8438), .ZN(n5381) );
  OR2_X1 U6960 ( .A1(n9385), .A2(n7316), .ZN(n8305) );
  NAND2_X1 U6961 ( .A1(n9385), .A2(n7316), .ZN(n8313) );
  INV_X1 U6962 ( .A(n7316), .ZN(n9345) );
  NAND2_X1 U6963 ( .A1(n9385), .A2(n9345), .ZN(n5384) );
  NAND2_X1 U6964 ( .A1(n4519), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6965 ( .A1(n4515), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5389) );
  AND2_X1 U6966 ( .A1(n5385), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6967 ( .A1(n5386), .A2(n5402), .ZN(n7353) );
  NAND2_X1 U6968 ( .A1(n4522), .A2(n7353), .ZN(n5388) );
  NAND2_X1 U6969 ( .A1(n4520), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5387) );
  NAND4_X1 U6970 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n9384)
         );
  XNOR2_X1 U6971 ( .A(n5392), .B(n5391), .ZN(n6623) );
  NAND2_X1 U6972 ( .A1(n6623), .A2(n8438), .ZN(n5395) );
  NAND2_X1 U6973 ( .A1(n5377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5393) );
  XNOR2_X1 U6974 ( .A(n5393), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U6975 ( .A1(n5555), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5554), .B2(
        n10585), .ZN(n5394) );
  OR2_X1 U6976 ( .A1(n9384), .A2(n7331), .ZN(n8324) );
  NAND2_X1 U6977 ( .A1(n7331), .A2(n9384), .ZN(n8319) );
  NAND2_X1 U6978 ( .A1(n8324), .A2(n8319), .ZN(n7305) );
  INV_X1 U6979 ( .A(n9384), .ZN(n7463) );
  NAND2_X1 U6980 ( .A1(n7463), .A2(n7331), .ZN(n5396) );
  NAND2_X1 U6981 ( .A1(n6627), .A2(n8438), .ZN(n5401) );
  OR2_X1 U6982 ( .A1(n5510), .A2(n9792), .ZN(n5399) );
  AOI22_X1 U6983 ( .A1(n5555), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5554), .B2(
        n7751), .ZN(n5400) );
  NAND2_X1 U6984 ( .A1(n5401), .A2(n5400), .ZN(n8266) );
  NAND2_X1 U6985 ( .A1(n4519), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6986 ( .A1(n4515), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5406) );
  NOR2_X1 U6987 ( .A1(n5402), .A2(n7460), .ZN(n5403) );
  OR2_X1 U6988 ( .A1(n5418), .A2(n5403), .ZN(n8265) );
  NAND2_X1 U6989 ( .A1(n4522), .A2(n8265), .ZN(n5405) );
  NAND2_X1 U6990 ( .A1(n4520), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5404) );
  OR2_X1 U6991 ( .A1(n8266), .A2(n7468), .ZN(n8320) );
  AND2_X1 U6992 ( .A1(n5411), .A2(n5410), .ZN(n5412) );
  INV_X1 U6993 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6994 ( .A1(n5510), .A2(n5414), .ZN(n5426) );
  NAND2_X1 U6995 ( .A1(n5426), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6996 ( .A(n5415), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7985) );
  AOI22_X1 U6997 ( .A1(n5555), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5554), .B2(
        n7985), .ZN(n5416) );
  NAND2_X1 U6998 ( .A1(n4515), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6999 ( .A1(n4520), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5422) );
  OR2_X1 U7000 ( .A1(n5418), .A2(n5417), .ZN(n5419) );
  NAND2_X1 U7001 ( .A1(n5432), .A2(n5419), .ZN(n7578) );
  NAND2_X1 U7002 ( .A1(n4522), .A2(n7578), .ZN(n5421) );
  NAND2_X1 U7003 ( .A1(n4519), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5420) );
  OR2_X1 U7004 ( .A1(n8485), .A2(n5122), .ZN(n7583) );
  XNOR2_X1 U7005 ( .A(n5425), .B(n5424), .ZN(n6638) );
  NAND2_X1 U7006 ( .A1(n6638), .A2(n8438), .ZN(n5431) );
  NAND2_X1 U7007 ( .A1(n5428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5427) );
  MUX2_X1 U7008 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5427), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5429) );
  AOI22_X1 U7009 ( .A1(n5555), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5554), .B2(
        n7997), .ZN(n5430) );
  NAND2_X1 U7010 ( .A1(n5431), .A2(n5430), .ZN(n7851) );
  NAND2_X1 U7011 ( .A1(n4515), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7012 ( .A1(n4520), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7013 ( .A1(n5432), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7014 ( .A1(n5443), .A2(n5433), .ZN(n7847) );
  NAND2_X1 U7015 ( .A1(n4523), .A2(n7847), .ZN(n5435) );
  NAND2_X1 U7016 ( .A1(n4519), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5434) );
  OR2_X1 U7017 ( .A1(n7851), .A2(n7892), .ZN(n8338) );
  NAND2_X1 U7018 ( .A1(n7851), .A2(n7892), .ZN(n8334) );
  NAND2_X1 U7019 ( .A1(n8338), .A2(n8334), .ZN(n8490) );
  NAND2_X1 U7020 ( .A1(n8321), .A2(n8326), .ZN(n7569) );
  INV_X1 U7021 ( .A(n7468), .ZN(n9383) );
  NAND2_X1 U7022 ( .A1(n8266), .A2(n9383), .ZN(n7565) );
  AND2_X1 U7023 ( .A1(n7569), .A2(n7565), .ZN(n7566) );
  XNOR2_X1 U7024 ( .A(n5439), .B(n5438), .ZN(n6732) );
  NAND2_X1 U7025 ( .A1(n6732), .A2(n8438), .ZN(n5442) );
  NAND2_X1 U7026 ( .A1(n5452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U7027 ( .A(n5440), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8177) );
  AOI22_X1 U7028 ( .A1(n5555), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5554), .B2(
        n8177), .ZN(n5441) );
  NAND2_X1 U7029 ( .A1(n5442), .A2(n5441), .ZN(n8082) );
  NAND2_X1 U7030 ( .A1(n4519), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7031 ( .A1(n4525), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7032 ( .A1(n5443), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7033 ( .A1(n5456), .A2(n5444), .ZN(n8071) );
  NAND2_X1 U7034 ( .A1(n4522), .A2(n8071), .ZN(n5446) );
  NAND2_X1 U7035 ( .A1(n4520), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5445) );
  NAND4_X1 U7036 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n9381)
         );
  NOR2_X1 U7037 ( .A1(n8082), .A2(n9381), .ZN(n5449) );
  INV_X1 U7038 ( .A(n8082), .ZN(n7780) );
  XNOR2_X1 U7039 ( .A(n5451), .B(n5450), .ZN(n6744) );
  NAND2_X1 U7040 ( .A1(n6744), .A2(n8438), .ZN(n5455) );
  OR2_X1 U7041 ( .A1(n5465), .A2(n9792), .ZN(n5453) );
  XNOR2_X1 U7042 ( .A(n5453), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8174) );
  AOI22_X1 U7043 ( .A1(n5555), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8174), .B2(
        n5554), .ZN(n5454) );
  NAND2_X1 U7044 ( .A1(n5455), .A2(n5454), .ZN(n8024) );
  NAND2_X1 U7045 ( .A1(n4519), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7046 ( .A1(n4515), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5459) );
  OR2_X1 U7047 ( .A1(n5112), .A2(n5470), .ZN(n8019) );
  NAND2_X1 U7048 ( .A1(n4523), .A2(n8019), .ZN(n5458) );
  NAND2_X1 U7049 ( .A1(n4520), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5457) );
  OR2_X1 U7050 ( .A1(n8024), .A2(n8074), .ZN(n8345) );
  NAND2_X1 U7051 ( .A1(n8024), .A2(n8074), .ZN(n8346) );
  NAND2_X1 U7052 ( .A1(n8345), .A2(n8346), .ZN(n8492) );
  INV_X1 U7053 ( .A(n8074), .ZN(n9380) );
  NAND2_X1 U7054 ( .A1(n8024), .A2(n9380), .ZN(n5461) );
  XNOR2_X1 U7055 ( .A(n5463), .B(n5462), .ZN(n6857) );
  NAND2_X1 U7056 ( .A1(n6857), .A2(n8438), .ZN(n5468) );
  INV_X1 U7057 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7058 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  NAND2_X1 U7059 ( .A1(n5466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U7060 ( .A(n5479), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9409) );
  AOI22_X1 U7061 ( .A1(n9409), .A2(n5554), .B1(n5555), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7062 ( .A1(n4519), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7063 ( .A1(n4525), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5474) );
  OR2_X1 U7064 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7065 ( .A1(n5483), .A2(n5471), .ZN(n7900) );
  NAND2_X1 U7066 ( .A1(n4523), .A2(n7900), .ZN(n5473) );
  NAND2_X1 U7067 ( .A1(n4520), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5472) );
  NAND4_X1 U7068 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9379)
         );
  AND2_X1 U7069 ( .A1(n8349), .A2(n9379), .ZN(n8351) );
  OR2_X1 U7070 ( .A1(n8349), .A2(n9379), .ZN(n8348) );
  XNOR2_X1 U7071 ( .A(n5477), .B(n5476), .ZN(n6897) );
  NAND2_X1 U7072 ( .A1(n6897), .A2(n8438), .ZN(n5482) );
  INV_X1 U7073 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7074 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  NAND2_X1 U7075 ( .A1(n5480), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5493) );
  XNOR2_X1 U7076 ( .A(n5493), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9419) );
  AOI22_X1 U7077 ( .A1(n9419), .A2(n5554), .B1(n5555), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7078 ( .A1(n5482), .A2(n5481), .ZN(n8034) );
  NAND2_X1 U7079 ( .A1(n4519), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7080 ( .A1(n4515), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7081 ( .A1(n5483), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7082 ( .A1(n5498), .A2(n5484), .ZN(n8030) );
  NAND2_X1 U7083 ( .A1(n4523), .A2(n8030), .ZN(n5486) );
  NAND2_X1 U7084 ( .A1(n4520), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5485) );
  OR2_X1 U7085 ( .A1(n8034), .A2(n8236), .ZN(n8353) );
  NAND2_X1 U7086 ( .A1(n8034), .A2(n8236), .ZN(n8352) );
  INV_X1 U7087 ( .A(n8236), .ZN(n9378) );
  NAND2_X1 U7088 ( .A1(n8034), .A2(n9378), .ZN(n5489) );
  XNOR2_X1 U7089 ( .A(n5491), .B(n5490), .ZN(n7042) );
  NAND2_X1 U7090 ( .A1(n7042), .A2(n8438), .ZN(n5497) );
  INV_X1 U7091 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7092 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  NAND2_X1 U7093 ( .A1(n5494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U7094 ( .A(n5495), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9456) );
  AOI22_X1 U7095 ( .A1(n9456), .A2(n5554), .B1(n5555), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7096 ( .A1(n4515), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7097 ( .A1(n4519), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5503) );
  INV_X1 U7098 ( .A(n5514), .ZN(n5500) );
  NAND2_X1 U7099 ( .A1(n5498), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7100 ( .A1(n5500), .A2(n5499), .ZN(n8565) );
  NAND2_X1 U7101 ( .A1(n4522), .A2(n8565), .ZN(n5502) );
  NAND2_X1 U7102 ( .A1(n4520), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7103 ( .A1(n9717), .A2(n8554), .ZN(n5505) );
  INV_X1 U7104 ( .A(n9717), .ZN(n7927) );
  XNOR2_X1 U7105 ( .A(n5507), .B(n5506), .ZN(n7213) );
  NAND2_X1 U7106 ( .A1(n7213), .A2(n8438), .ZN(n5513) );
  INV_X1 U7107 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7108 ( .A1(n5510), .A2(n5509), .ZN(n5522) );
  NAND2_X1 U7109 ( .A1(n5522), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5511) );
  XNOR2_X1 U7110 ( .A(n5511), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U7111 ( .A1(n5555), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5554), .B2(
        n9463), .ZN(n5512) );
  NAND2_X1 U7112 ( .A1(n5513), .A2(n5512), .ZN(n8556) );
  NAND2_X1 U7113 ( .A1(n4519), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7114 ( .A1(n4525), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5518) );
  NOR2_X1 U7115 ( .A1(n5514), .A2(n9192), .ZN(n5515) );
  OR2_X1 U7116 ( .A1(n5527), .A2(n5515), .ZN(n8551) );
  NAND2_X1 U7117 ( .A1(n4523), .A2(n8551), .ZN(n5517) );
  NAND2_X1 U7118 ( .A1(n4520), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5516) );
  OR2_X1 U7119 ( .A1(n8556), .A2(n8563), .ZN(n8363) );
  NAND2_X1 U7120 ( .A1(n8556), .A2(n8563), .ZN(n8362) );
  INV_X1 U7121 ( .A(n8556), .ZN(n8200) );
  XNOR2_X1 U7122 ( .A(n5521), .B(n5520), .ZN(n7258) );
  NAND2_X1 U7123 ( .A1(n7258), .A2(n8438), .ZN(n5525) );
  OAI21_X1 U7124 ( .B1(n5522), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5523) );
  XNOR2_X1 U7125 ( .A(n5523), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9507) );
  AOI22_X1 U7126 ( .A1(n5555), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5554), .B2(
        n9507), .ZN(n5524) );
  NAND2_X1 U7127 ( .A1(n4515), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7128 ( .A1(n4520), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5531) );
  OR2_X1 U7129 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  NAND2_X1 U7130 ( .A1(n5540), .A2(n5528), .ZN(n8246) );
  NAND2_X1 U7131 ( .A1(n4522), .A2(n8246), .ZN(n5530) );
  NAND2_X1 U7132 ( .A1(n4519), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5529) );
  OR2_X1 U7133 ( .A1(n8250), .A2(n8259), .ZN(n8275) );
  NAND2_X1 U7134 ( .A1(n8250), .A2(n8259), .ZN(n8278) );
  NAND2_X1 U7135 ( .A1(n8275), .A2(n8278), .ZN(n8498) );
  INV_X1 U7136 ( .A(n8259), .ZN(n9377) );
  NAND2_X1 U7137 ( .A1(n8250), .A2(n9377), .ZN(n5533) );
  XNOR2_X1 U7138 ( .A(n5534), .B(n5544), .ZN(n7314) );
  NAND2_X1 U7139 ( .A1(n7314), .A2(n8438), .ZN(n5537) );
  INV_X1 U7140 ( .A(n5658), .ZN(n5704) );
  NAND2_X1 U7141 ( .A1(n5704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5535) );
  XNOR2_X1 U7142 ( .A(n5535), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9514) );
  AOI22_X1 U7143 ( .A1(n5555), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5554), .B2(
        n9514), .ZN(n5536) );
  NAND2_X1 U7144 ( .A1(n4525), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7145 ( .A1(n4520), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5538) );
  AND2_X1 U7146 ( .A1(n5539), .A2(n5538), .ZN(n5543) );
  XNOR2_X1 U7147 ( .A(n5540), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U7148 ( .A1(n8256), .A2(n4522), .ZN(n5542) );
  NAND2_X1 U7149 ( .A1(n4519), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7150 ( .A1(n5545), .A2(n5544), .ZN(n5547) );
  NAND2_X1 U7151 ( .A1(n5547), .A2(n5546), .ZN(n5549) );
  NAND2_X1 U7152 ( .A1(n7432), .A2(n8438), .ZN(n5557) );
  INV_X1 U7153 ( .A(n5377), .ZN(n5551) );
  NAND2_X1 U7154 ( .A1(n5551), .A2(n5113), .ZN(n5552) );
  NAND2_X1 U7155 ( .A1(n5552), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5553) );
  XNOR2_X1 U7156 ( .A(n5553), .B(n5657), .ZN(n5694) );
  INV_X1 U7157 ( .A(n5694), .ZN(n5697) );
  AOI22_X1 U7158 ( .A1(n5555), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5697), .B2(
        n5554), .ZN(n5556) );
  AND2_X1 U7159 ( .A1(n5558), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5560) );
  OR2_X1 U7160 ( .A1(n5560), .A2(n5559), .ZN(n9650) );
  NAND2_X1 U7161 ( .A1(n9650), .A2(n4523), .ZN(n5563) );
  AOI22_X1 U7162 ( .A1(n4519), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n4515), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7163 ( .A1(n4520), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7164 ( .A1(n9652), .A2(n9630), .ZN(n8379) );
  INV_X1 U7165 ( .A(n9630), .ZN(n9375) );
  NAND2_X1 U7166 ( .A1(n9634), .A2(n9647), .ZN(n9617) );
  NAND2_X1 U7167 ( .A1(n8381), .A2(n9617), .ZN(n9632) );
  NAND2_X1 U7168 ( .A1(n7523), .A2(n8438), .ZN(n5568) );
  OR2_X1 U7169 ( .A1(n5333), .A2(n7562), .ZN(n5567) );
  OR2_X1 U7170 ( .A1(n5570), .A2(n5569), .ZN(n5571) );
  NAND2_X1 U7171 ( .A1(n5579), .A2(n5571), .ZN(n9621) );
  INV_X1 U7172 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U7173 ( .A1(n4520), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7174 ( .A1(n4515), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5572) );
  OAI211_X1 U7175 ( .C1(n5638), .C2(n9775), .A(n5573), .B(n5572), .ZN(n5574)
         );
  NAND2_X1 U7176 ( .A1(n8936), .A2(n9631), .ZN(n8382) );
  NAND2_X1 U7177 ( .A1(n8384), .A2(n8382), .ZN(n9619) );
  XNOR2_X1 U7178 ( .A(n5576), .B(n5575), .ZN(n7812) );
  NAND2_X1 U7179 ( .A1(n7812), .A2(n8438), .ZN(n5578) );
  OR2_X1 U7180 ( .A1(n5333), .A2(n7814), .ZN(n5577) );
  NAND2_X1 U7181 ( .A1(n5579), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7182 ( .A1(n5588), .A2(n5580), .ZN(n9608) );
  INV_X1 U7183 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9771) );
  NAND2_X1 U7184 ( .A1(n4520), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7185 ( .A1(n4525), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U7186 ( .C1(n5638), .C2(n9771), .A(n5582), .B(n5581), .ZN(n5583)
         );
  OR2_X1 U7187 ( .A1(n9607), .A2(n9616), .ZN(n8389) );
  NAND2_X1 U7188 ( .A1(n9607), .A2(n9616), .ZN(n8388) );
  INV_X1 U7189 ( .A(n9616), .ZN(n9372) );
  NAND2_X1 U7190 ( .A1(n7778), .A2(n8438), .ZN(n5587) );
  OR2_X1 U7191 ( .A1(n5333), .A2(n7777), .ZN(n5586) );
  NAND2_X1 U7192 ( .A1(n5588), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7193 ( .A1(n5602), .A2(n5589), .ZN(n9597) );
  NAND2_X1 U7194 ( .A1(n9597), .A2(n4522), .ZN(n5596) );
  INV_X1 U7195 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7196 ( .A1(n4515), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7197 ( .A1(n4519), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5590) );
  OAI211_X1 U7198 ( .C1(n5593), .C2(n5592), .A(n5591), .B(n5590), .ZN(n5594)
         );
  INV_X1 U7199 ( .A(n5594), .ZN(n5595) );
  NAND2_X1 U7200 ( .A1(n5596), .A2(n5595), .ZN(n9371) );
  NOR2_X1 U7201 ( .A1(n8920), .A2(n9371), .ZN(n5597) );
  NAND2_X1 U7202 ( .A1(n6094), .A2(n8438), .ZN(n5601) );
  OR2_X1 U7203 ( .A1(n5333), .A2(n7886), .ZN(n5600) );
  INV_X1 U7204 ( .A(n5615), .ZN(n5604) );
  NAND2_X1 U7205 ( .A1(n5602), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7206 ( .A1(n5604), .A2(n5603), .ZN(n9585) );
  NAND2_X1 U7207 ( .A1(n9585), .A2(n4522), .ZN(n5609) );
  INV_X1 U7208 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9763) );
  NAND2_X1 U7209 ( .A1(n4525), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7210 ( .A1(n4520), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5605) );
  OAI211_X1 U7211 ( .C1(n5638), .C2(n9763), .A(n5606), .B(n5605), .ZN(n5607)
         );
  INV_X1 U7212 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7213 ( .A1(n9580), .A2(n9594), .ZN(n8394) );
  NAND2_X1 U7214 ( .A1(n8397), .A2(n8394), .ZN(n9589) );
  INV_X1 U7215 ( .A(n9594), .ZN(n9370) );
  XNOR2_X1 U7216 ( .A(n5611), .B(n5610), .ZN(n7956) );
  NAND2_X1 U7217 ( .A1(n7956), .A2(n8438), .ZN(n5613) );
  OR2_X1 U7218 ( .A1(n5333), .A2(n8964), .ZN(n5612) );
  OR2_X1 U7219 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  NAND2_X1 U7220 ( .A1(n5617), .A2(n5616), .ZN(n9574) );
  NAND2_X1 U7221 ( .A1(n9574), .A2(n4523), .ZN(n5622) );
  INV_X1 U7222 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U7223 ( .A1(n4520), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7224 ( .A1(n4515), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5618) );
  OAI211_X1 U7225 ( .C1(n5638), .C2(n9759), .A(n5619), .B(n5618), .ZN(n5620)
         );
  INV_X1 U7226 ( .A(n5620), .ZN(n5621) );
  INV_X1 U7227 ( .A(n9572), .ZN(n9761) );
  NAND2_X1 U7228 ( .A1(n5625), .A2(n5624), .ZN(n5627) );
  NAND2_X1 U7229 ( .A1(n5627), .A2(n5626), .ZN(n5643) );
  INV_X1 U7230 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5631) );
  INV_X1 U7231 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8141) );
  MUX2_X1 U7232 ( .A(n5631), .B(n8141), .S(n4516), .Z(n5628) );
  INV_X1 U7233 ( .A(SI_27_), .ZN(n9059) );
  NAND2_X1 U7234 ( .A1(n5628), .A2(n9059), .ZN(n5644) );
  INV_X1 U7235 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7236 ( .A1(n5629), .A2(SI_27_), .ZN(n5630) );
  NAND2_X1 U7237 ( .A1(n8091), .A2(n8438), .ZN(n5633) );
  OR2_X1 U7238 ( .A1(n5333), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U7239 ( .A1(n5634), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5635) );
  INV_X1 U7240 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7241 ( .A1(n5635), .A2(n5650), .ZN(n9554) );
  NAND2_X1 U7242 ( .A1(n9554), .A2(n4523), .ZN(n5641) );
  INV_X1 U7243 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7244 ( .A1(n4520), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7245 ( .A1(n4515), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U7246 ( .C1(n5638), .C2(n6260), .A(n5637), .B(n5636), .ZN(n5639)
         );
  INV_X1 U7247 ( .A(n5639), .ZN(n5640) );
  AND2_X1 U7248 ( .A1(n8601), .A2(n9367), .ZN(n5692) );
  NAND2_X1 U7249 ( .A1(n5643), .A2(n5642), .ZN(n5645) );
  NAND2_X1 U7250 ( .A1(n5645), .A2(n5644), .ZN(n5749) );
  INV_X1 U7251 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5646) );
  INV_X1 U7252 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8892) );
  MUX2_X1 U7253 ( .A(n5646), .B(n8892), .S(n4517), .Z(n5751) );
  XNOR2_X1 U7254 ( .A(n5751), .B(SI_28_), .ZN(n5748) );
  NAND2_X1 U7255 ( .A1(n8190), .A2(n8438), .ZN(n5648) );
  OR2_X1 U7256 ( .A1(n5333), .A2(n5646), .ZN(n5647) );
  NAND2_X1 U7257 ( .A1(n4519), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7258 ( .A1(n4525), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7259 ( .A1(n8978), .A2(n5649), .ZN(n5671) );
  NAND2_X1 U7260 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n5650), .ZN(n5651) );
  NAND2_X1 U7261 ( .A1(n5671), .A2(n5651), .ZN(n9546) );
  NAND2_X1 U7262 ( .A1(n4522), .A2(n9546), .ZN(n5653) );
  NAND2_X1 U7263 ( .A1(n4520), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5652) );
  NAND4_X1 U7264 ( .A1(n5655), .A2(n5654), .A3(n5653), .A4(n5652), .ZN(n9366)
         );
  XNOR2_X1 U7265 ( .A(n5747), .B(n8474), .ZN(n5678) );
  NOR2_X1 U7266 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5659) );
  NAND2_X1 U7267 ( .A1(n5659), .A2(n5663), .ZN(n5700) );
  NAND2_X1 U7268 ( .A1(n5700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7269 ( .A1(n8523), .A2(n5697), .ZN(n5667) );
  NAND2_X1 U7270 ( .A1(n5663), .A2(n5664), .ZN(n5661) );
  NAND2_X1 U7271 ( .A1(n8513), .A2(n8516), .ZN(n5666) );
  INV_X1 U7272 ( .A(n5668), .ZN(n7047) );
  XNOR2_X1 U7273 ( .A(n7047), .B(n8521), .ZN(n6961) );
  INV_X1 U7274 ( .A(n6961), .ZN(n5670) );
  NAND2_X2 U7275 ( .A1(n8523), .A2(n8513), .ZN(n8453) );
  INV_X1 U7276 ( .A(n5671), .ZN(n8898) );
  NAND2_X1 U7277 ( .A1(n4522), .A2(n8898), .ZN(n8446) );
  NAND2_X1 U7278 ( .A1(n4515), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7279 ( .A1(n4520), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7280 ( .A1(n4519), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5672) );
  NOR2_X1 U7281 ( .A1(n8607), .A2(n9646), .ZN(n5675) );
  INV_X1 U7282 ( .A(n6976), .ZN(n7044) );
  NAND2_X1 U7283 ( .A1(n6885), .A2(n8292), .ZN(n5681) );
  NAND2_X1 U7284 ( .A1(n9386), .A2(n7320), .ZN(n8310) );
  NAND2_X1 U7285 ( .A1(n8303), .A2(n8310), .ZN(n8481) );
  INV_X1 U7286 ( .A(n8481), .ZN(n7089) );
  NAND2_X1 U7287 ( .A1(n7086), .A2(n7089), .ZN(n7088) );
  AND2_X1 U7288 ( .A1(n8303), .A2(n8305), .ZN(n8314) );
  NAND2_X1 U7289 ( .A1(n7088), .A2(n8314), .ZN(n5682) );
  NAND2_X1 U7290 ( .A1(n5683), .A2(n8320), .ZN(n7564) );
  INV_X1 U7291 ( .A(n7569), .ZN(n8486) );
  NAND2_X1 U7292 ( .A1(n7564), .A2(n8486), .ZN(n5684) );
  NAND2_X1 U7293 ( .A1(n5684), .A2(n8321), .ZN(n7589) );
  INV_X1 U7294 ( .A(n8338), .ZN(n5685) );
  OR2_X1 U7295 ( .A1(n8082), .A2(n8011), .ZN(n8339) );
  NAND2_X1 U7296 ( .A1(n8082), .A2(n8011), .ZN(n8336) );
  NAND2_X1 U7297 ( .A1(n7597), .A2(n8477), .ZN(n7596) );
  INV_X1 U7298 ( .A(n8336), .ZN(n8340) );
  NOR2_X1 U7299 ( .A1(n8492), .A2(n8340), .ZN(n5686) );
  INV_X1 U7300 ( .A(n9379), .ZN(n8022) );
  NOR2_X1 U7301 ( .A1(n8349), .A2(n8022), .ZN(n5688) );
  NAND2_X1 U7302 ( .A1(n8349), .A2(n8022), .ZN(n5687) );
  AND2_X1 U7303 ( .A1(n7927), .A2(n8554), .ZN(n8357) );
  NAND2_X1 U7304 ( .A1(n9717), .A2(n8240), .ZN(n8358) );
  INV_X1 U7305 ( .A(n8275), .ZN(n5689) );
  NAND2_X1 U7306 ( .A1(n8261), .A2(n9645), .ZN(n8276) );
  NAND2_X1 U7307 ( .A1(n8370), .A2(n8276), .ZN(n8500) );
  INV_X1 U7308 ( .A(n8381), .ZN(n5690) );
  NAND2_X1 U7309 ( .A1(n8382), .A2(n9617), .ZN(n8375) );
  INV_X1 U7310 ( .A(n8389), .ZN(n5691) );
  NAND2_X1 U7311 ( .A1(n9596), .A2(n8475), .ZN(n9587) );
  NAND2_X1 U7312 ( .A1(n8920), .A2(n9604), .ZN(n9586) );
  AND2_X1 U7313 ( .A1(n8394), .A2(n9586), .ZN(n8402) );
  INV_X1 U7314 ( .A(n8397), .ZN(n8401) );
  AND2_X1 U7315 ( .A1(n9572), .A2(n9583), .ZN(n8396) );
  NOR2_X1 U7316 ( .A1(n9361), .A2(n9571), .ZN(n8410) );
  NAND2_X1 U7317 ( .A1(n9361), .A2(n9571), .ZN(n8409) );
  INV_X1 U7318 ( .A(n5692), .ZN(n5693) );
  XOR2_X1 U7319 ( .A(n8474), .B(n5763), .Z(n9550) );
  NAND2_X1 U7320 ( .A1(n6967), .A2(n5694), .ZN(n6575) );
  NAND2_X1 U7321 ( .A1(n8523), .A2(n5694), .ZN(n5696) );
  OR2_X1 U7322 ( .A1(n6575), .A2(n6970), .ZN(n5695) );
  NAND2_X1 U7323 ( .A1(n5696), .A2(n5695), .ZN(n6579) );
  NAND2_X1 U7324 ( .A1(n6842), .A2(n6579), .ZN(n7031) );
  NAND2_X1 U7325 ( .A1(n5697), .A2(n6967), .ZN(n6971) );
  NAND2_X1 U7326 ( .A1(n7816), .A2(n5698), .ZN(n9737) );
  NAND2_X1 U7327 ( .A1(n5736), .A2(n5737), .ZN(n5712) );
  NAND2_X1 U7328 ( .A1(n5712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7329 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NAND2_X1 U7330 ( .A1(n4581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7331 ( .A1(n8009), .A2(n8070), .ZN(n5718) );
  INV_X1 U7332 ( .A(n5712), .ZN(n5710) );
  NOR2_X1 U7333 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5707) );
  INV_X1 U7334 ( .A(P2_B_REG_SCAN_IN), .ZN(n5706) );
  AOI22_X1 U7335 ( .A1(n5707), .A2(P2_B_REG_SCAN_IN), .B1(n5706), .B2(
        P2_IR_REG_24__SCAN_IN), .ZN(n5708) );
  INV_X1 U7336 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U7337 ( .A1(n5710), .A2(n5709), .ZN(n5714) );
  XNOR2_X1 U7338 ( .A(P2_IR_REG_24__SCAN_IN), .B(P2_B_REG_SCAN_IN), .ZN(n5711)
         );
  NAND3_X1 U7339 ( .A1(n5712), .A2(P2_IR_REG_25__SCAN_IN), .A3(n5711), .ZN(
        n5713) );
  INV_X1 U7340 ( .A(n8070), .ZN(n5715) );
  INV_X1 U7341 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7342 ( .A1(n5719), .A2(n5716), .ZN(n5717) );
  OR2_X1 U7343 ( .A1(n5721), .A2(n5720), .ZN(n5723) );
  NAND2_X1 U7344 ( .A1(n5723), .A2(n5722), .ZN(n5735) );
  OAI21_X1 U7345 ( .B1(n6645), .B2(P2_D_REG_0__SCAN_IN), .A(n6975), .ZN(n6583)
         );
  OR2_X1 U7346 ( .A1(n6640), .A2(n6583), .ZN(n6837) );
  NOR2_X1 U7347 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n5727) );
  NOR4_X1 U7348 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5726) );
  NOR4_X1 U7349 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5725) );
  NOR4_X1 U7350 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5724) );
  NAND4_X1 U7351 ( .A1(n5727), .A2(n5726), .A3(n5725), .A4(n5724), .ZN(n5733)
         );
  NOR4_X1 U7352 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U7353 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5730) );
  NOR4_X1 U7354 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5729) );
  NOR4_X1 U7355 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U7356 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n5732)
         );
  NOR2_X1 U7357 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  NOR2_X1 U7358 ( .A1(n6837), .A2(n6577), .ZN(n6946) );
  XNOR2_X1 U7359 ( .A(n5736), .B(n5737), .ZN(n7055) );
  NAND2_X1 U7360 ( .A1(n6946), .A2(n6952), .ZN(n6986) );
  AND3_X1 U7361 ( .A1(n6970), .A2(n8516), .A3(n5697), .ZN(n5738) );
  NAND2_X1 U7362 ( .A1(n5738), .A2(n8523), .ZN(n6947) );
  AND2_X1 U7363 ( .A1(n6842), .A2(n6947), .ZN(n5739) );
  OR2_X1 U7364 ( .A1(n6986), .A2(n5739), .ZN(n5742) );
  NAND2_X1 U7365 ( .A1(n6640), .A2(n6583), .ZN(n6584) );
  INV_X1 U7366 ( .A(n6952), .ZN(n5740) );
  NAND3_X1 U7367 ( .A1(n6947), .A2(n8453), .A3(n9716), .ZN(n6985) );
  NAND2_X1 U7368 ( .A1(n6985), .A2(n10622), .ZN(n6944) );
  NAND2_X1 U7369 ( .A1(n6988), .A2(n6944), .ZN(n5741) );
  OR2_X1 U7370 ( .A1(n9666), .A2(n10652), .ZN(n5745) );
  NAND2_X1 U7371 ( .A1(n9671), .A2(n6261), .ZN(n5744) );
  NAND2_X1 U7372 ( .A1(n10652), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7373 ( .A1(n5745), .A2(n5124), .ZN(P2_U3455) );
  NOR2_X1 U7374 ( .A1(n9671), .A2(n9366), .ZN(n5746) );
  NAND2_X1 U7375 ( .A1(n5749), .A2(n5748), .ZN(n5753) );
  INV_X1 U7376 ( .A(SI_28_), .ZN(n5750) );
  NAND2_X1 U7377 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  INV_X1 U7378 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9799) );
  INV_X1 U7379 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8882) );
  MUX2_X1 U7380 ( .A(n9799), .B(n8882), .S(n4516), .Z(n8421) );
  NAND2_X1 U7381 ( .A1(n8881), .A2(n8438), .ZN(n5755) );
  OR2_X1 U7382 ( .A1(n5333), .A2(n9799), .ZN(n5754) );
  NAND2_X1 U7383 ( .A1(n8904), .A2(n8607), .ZN(n8431) );
  XNOR2_X1 U7384 ( .A(n5756), .B(n4833), .ZN(n5762) );
  NAND2_X1 U7385 ( .A1(n4519), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7386 ( .A1(n4515), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7387 ( .A1(n4520), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5757) );
  AND2_X1 U7388 ( .A1(n6602), .A2(P2_B_REG_SCAN_IN), .ZN(n5760) );
  OR2_X1 U7389 ( .A1(n9646), .A2(n5760), .ZN(n9538) );
  OAI22_X1 U7390 ( .A1(n8449), .A2(n9538), .B1(n8912), .B2(n9644), .ZN(n5761)
         );
  XNOR2_X1 U7391 ( .A(n8468), .B(n8508), .ZN(n8901) );
  NAND2_X1 U7392 ( .A1(n8906), .A2(n5765), .ZN(n6586) );
  NAND2_X1 U7393 ( .A1(n6586), .A2(n10649), .ZN(n5768) );
  INV_X1 U7394 ( .A(n8904), .ZN(n6588) );
  NOR2_X1 U7395 ( .A1(n6588), .A2(n9789), .ZN(n5766) );
  NAND2_X1 U7396 ( .A1(n5768), .A2(n5767), .ZN(P2_U3456) );
  INV_X2 U7397 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5771) );
  NOR2_X1 U7398 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5776) );
  INV_X1 U7399 ( .A(n5837), .ZN(n5775) );
  INV_X1 U7400 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7401 ( .A1(n5800), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U7402 ( .A(n5785), .B(n5784), .ZN(n6197) );
  NAND2_X1 U7403 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5787) );
  NAND2_X1 U7404 ( .A1(n8271), .A2(n8529), .ZN(n5790) );
  OR2_X1 U7405 ( .A1(n8530), .A2(n7405), .ZN(n5789) );
  NAND2_X1 U7406 ( .A1(n5923), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5936) );
  INV_X1 U7407 ( .A(n5936), .ZN(n5791) );
  NAND2_X1 U7408 ( .A1(n5791), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5950) );
  INV_X1 U7409 ( .A(n5950), .ZN(n5792) );
  NAND2_X1 U7410 ( .A1(n5948), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7411 ( .A1(n5793), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7412 ( .A1(n6000), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6025) );
  INV_X1 U7413 ( .A(n6025), .ZN(n5794) );
  INV_X1 U7414 ( .A(n6052), .ZN(n5797) );
  AND2_X1 U7415 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5796) );
  INV_X1 U7416 ( .A(n5798), .ZN(n5823) );
  INV_X1 U7417 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U7418 ( .A1(n5823), .A2(n8952), .ZN(n5799) );
  NAND2_X1 U7419 ( .A1(n6065), .A2(n5799), .ZN(n10191) );
  NOR2_X2 U7420 ( .A1(n5800), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5806) );
  INV_X1 U7421 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5801) );
  OR2_X1 U7422 ( .A1(n5806), .A2(n5801), .ZN(n5802) );
  NAND2_X1 U7423 ( .A1(n5802), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7424 ( .A1(n5806), .A2(n5803), .ZN(n5809) );
  INV_X1 U7425 ( .A(n5809), .ZN(n5807) );
  OR2_X1 U7426 ( .A1(n10191), .A2(n6111), .ZN(n5817) );
  INV_X1 U7427 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10320) );
  AND2_X4 U7428 ( .A1(n8545), .A2(n5811), .ZN(n8536) );
  NAND2_X1 U7429 ( .A1(n8536), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7430 ( .A1(n6198), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5813) );
  OAI211_X1 U7431 ( .C1(n6124), .C2(n10320), .A(n5814), .B(n5813), .ZN(n5815)
         );
  INV_X1 U7432 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7433 ( .A1(n7432), .A2(n8529), .ZN(n5821) );
  NAND2_X1 U7434 ( .A1(n5834), .A2(n6159), .ZN(n5819) );
  INV_X2 U7435 ( .A(n5901), .ZN(n6634) );
  AOI22_X1 U7436 ( .A1(n6049), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6166), .B2(
        n6634), .ZN(n5820) );
  INV_X1 U7437 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9898) );
  INV_X1 U7438 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5822) );
  OAI21_X1 U7439 ( .B1(n6052), .B2(n9898), .A(n5822), .ZN(n5824) );
  AND2_X1 U7440 ( .A1(n5824), .A2(n5823), .ZN(n10209) );
  NAND2_X1 U7441 ( .A1(n10209), .A2(n6154), .ZN(n5829) );
  INV_X1 U7442 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U7443 ( .A1(n6198), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7444 ( .A1(n8537), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5825) );
  OAI211_X1 U7445 ( .C1(n10266), .C2(n6152), .A(n5826), .B(n5825), .ZN(n5827)
         );
  INV_X1 U7446 ( .A(n5827), .ZN(n5828) );
  INV_X1 U7447 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U7448 ( .A1(n6041), .A2(n9272), .ZN(n5830) );
  NAND2_X1 U7449 ( .A1(n6052), .A2(n5830), .ZN(n9856) );
  OR2_X1 U7450 ( .A1(n9856), .A2(n6111), .ZN(n5833) );
  AOI22_X1 U7451 ( .A1(n6198), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8537), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7452 ( .A1(n8536), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7453 ( .A1(n7258), .A2(n8529), .ZN(n5836) );
  XNOR2_X1 U7454 ( .A(n5834), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7937) );
  AOI22_X1 U7455 ( .A1(n6049), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6634), .B2(
        n7937), .ZN(n5835) );
  NAND2_X1 U7456 ( .A1(n6744), .A2(n8529), .ZN(n5842) );
  NOR2_X1 U7457 ( .A1(n5914), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5920) );
  NOR2_X1 U7458 ( .A1(n5837), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5838) );
  AND2_X1 U7459 ( .A1(n5920), .A2(n5838), .ZN(n5957) );
  INV_X1 U7460 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7461 ( .A1(n5957), .A2(n5839), .ZN(n5971) );
  NAND2_X1 U7462 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7463 ( .A(n5840), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7192) );
  AOI22_X1 U7464 ( .A1(n6049), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6634), .B2(
        n7192), .ZN(n5841) );
  INV_X1 U7465 ( .A(n7768), .ZN(n10511) );
  NAND2_X1 U7466 ( .A1(n8536), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7467 ( .A1(n5989), .A2(n6821), .ZN(n5843) );
  AND2_X1 U7468 ( .A1(n6001), .A2(n5843), .ZN(n7762) );
  NAND2_X1 U7469 ( .A1(n6154), .A2(n7762), .ZN(n5846) );
  NAND2_X1 U7470 ( .A1(n8537), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5845) );
  INV_X2 U7471 ( .A(n8540), .ZN(n6198) );
  NAND2_X1 U7472 ( .A1(n6198), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U7473 ( .A1(n8536), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7474 ( .A1(n5907), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7475 ( .A1(n5961), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5848) );
  INV_X1 U7476 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7477 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5853) );
  XNOR2_X1 U7478 ( .A(n5854), .B(n5853), .ZN(n9969) );
  INV_X1 U7479 ( .A(n5855), .ZN(n6622) );
  OR2_X1 U7480 ( .A1(n5913), .A2(n6622), .ZN(n5857) );
  OAI211_X1 U7481 ( .C1(n5901), .C2(n9969), .A(n5857), .B(n5856), .ZN(n6277)
         );
  NAND2_X1 U7482 ( .A1(n5961), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7483 ( .A1(n8536), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7484 ( .A1(n5908), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7485 ( .A1(n5907), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5858) );
  NAND4_X2 U7486 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n9964)
         );
  INV_X1 U7487 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6740) );
  INV_X1 U7488 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5862) );
  OAI21_X1 U7489 ( .B1(n4518), .B2(n5863), .A(n5862), .ZN(n5865) );
  NAND2_X1 U7490 ( .A1(n5865), .A2(n5864), .ZN(n6604) );
  MUX2_X1 U7491 ( .A(n6740), .B(n6604), .S(n5901), .Z(n7492) );
  INV_X1 U7492 ( .A(n7492), .ZN(n7435) );
  NAND2_X1 U7493 ( .A1(n9964), .A2(n7435), .ZN(n7481) );
  INV_X1 U7494 ( .A(n9963), .ZN(n8823) );
  NAND2_X1 U7495 ( .A1(n8823), .A2(n6205), .ZN(n5866) );
  NAND2_X1 U7496 ( .A1(n7484), .A2(n5866), .ZN(n6849) );
  NAND2_X1 U7497 ( .A1(n5908), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7498 ( .A1(n5961), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7499 ( .A1(n5907), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5867) );
  INV_X1 U7500 ( .A(n9962), .ZN(n5880) );
  OR2_X1 U7501 ( .A1(n5913), .A2(n6613), .ZN(n5878) );
  OR2_X1 U7502 ( .A1(n8530), .A2(n6608), .ZN(n5877) );
  NOR2_X1 U7503 ( .A1(n5871), .A2(n5801), .ZN(n5872) );
  NAND2_X1 U7504 ( .A1(n5872), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5875) );
  INV_X1 U7505 ( .A(n5872), .ZN(n5874) );
  INV_X1 U7506 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7507 ( .A1(n5874), .A2(n5873), .ZN(n5886) );
  AND2_X1 U7508 ( .A1(n5875), .A2(n5886), .ZN(n9983) );
  NAND2_X1 U7509 ( .A1(n6634), .A2(n9983), .ZN(n5876) );
  NAND2_X1 U7510 ( .A1(n6849), .A2(n6852), .ZN(n6848) );
  NAND2_X1 U7511 ( .A1(n5880), .A2(n7417), .ZN(n5881) );
  NAND2_X1 U7512 ( .A1(n6848), .A2(n5881), .ZN(n6900) );
  INV_X1 U7513 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U7514 ( .A1(n6154), .A2(n7423), .ZN(n5885) );
  NAND2_X1 U7515 ( .A1(n8536), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7516 ( .A1(n8537), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7517 ( .A1(n5907), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7518 ( .A1(n5886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5888) );
  INV_X1 U7519 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7520 ( .A(n5888), .B(n5887), .ZN(n9996) );
  OR2_X1 U7521 ( .A1(n5913), .A2(n6612), .ZN(n5890) );
  OR2_X1 U7522 ( .A1(n8530), .A2(n6606), .ZN(n5889) );
  NAND2_X1 U7523 ( .A1(n6932), .A2(n5891), .ZN(n8825) );
  INV_X1 U7524 ( .A(n6932), .ZN(n9961) );
  NAND2_X1 U7525 ( .A1(n9961), .A2(n7427), .ZN(n8636) );
  AND2_X1 U7526 ( .A1(n8825), .A2(n8636), .ZN(n8627) );
  NAND2_X1 U7527 ( .A1(n6900), .A2(n8746), .ZN(n6899) );
  NAND2_X1 U7528 ( .A1(n6932), .A2(n7427), .ZN(n5892) );
  NAND2_X1 U7529 ( .A1(n6899), .A2(n5892), .ZN(n6930) );
  NAND2_X1 U7530 ( .A1(n8536), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5897) );
  NOR2_X1 U7531 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5893) );
  NOR2_X1 U7532 ( .A1(n5905), .A2(n5893), .ZN(n7446) );
  NAND2_X1 U7533 ( .A1(n6154), .A2(n7446), .ZN(n5896) );
  NAND2_X1 U7534 ( .A1(n8537), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7535 ( .A1(n6198), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5894) );
  OR2_X1 U7536 ( .A1(n6610), .A2(n5913), .ZN(n5904) );
  INV_X1 U7537 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U7538 ( .A1(n5898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5899) );
  MUX2_X1 U7539 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5899), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5900) );
  NAND2_X1 U7540 ( .A1(n5900), .A2(n5914), .ZN(n6788) );
  OAI22_X1 U7541 ( .A1(n8530), .A2(n9232), .B1(n5901), .B2(n6788), .ZN(n5902)
         );
  INV_X1 U7542 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7543 ( .A1(n5904), .A2(n5903), .ZN(n6937) );
  NAND2_X1 U7544 ( .A1(n7134), .A2(n6937), .ZN(n8635) );
  INV_X1 U7545 ( .A(n7134), .ZN(n9960) );
  INV_X1 U7546 ( .A(n6937), .ZN(n7449) );
  NAND2_X1 U7547 ( .A1(n9960), .A2(n7449), .ZN(n8637) );
  NAND2_X1 U7548 ( .A1(n8635), .A2(n8637), .ZN(n8745) );
  NOR2_X1 U7549 ( .A1(n5905), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U7550 ( .A1(n5923), .A2(n5906), .ZN(n7691) );
  NAND2_X1 U7551 ( .A1(n6154), .A2(n7691), .ZN(n5912) );
  NAND2_X1 U7552 ( .A1(n8536), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7553 ( .A1(n5907), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7554 ( .A1(n5908), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5909) );
  NAND4_X1 U7555 ( .A1(n5912), .A2(n5911), .A3(n5910), .A4(n5909), .ZN(n9959)
         );
  INV_X1 U7556 ( .A(n9959), .ZN(n6933) );
  NAND2_X1 U7557 ( .A1(n5914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5915) );
  XNOR2_X1 U7558 ( .A(n5915), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U7559 ( .A1(n6049), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6634), .B2(
        n6674), .ZN(n5916) );
  NAND2_X1 U7560 ( .A1(n6933), .A2(n7692), .ZN(n8634) );
  NAND2_X1 U7561 ( .A1(n7341), .A2(n9959), .ZN(n8638) );
  AND2_X1 U7562 ( .A1(n8634), .A2(n8638), .ZN(n8750) );
  INV_X1 U7563 ( .A(n8750), .ZN(n7130) );
  AND2_X1 U7564 ( .A1(n8745), .A2(n7130), .ZN(n5917) );
  NAND2_X1 U7565 ( .A1(n6930), .A2(n5917), .ZN(n7125) );
  NAND2_X1 U7566 ( .A1(n7134), .A2(n7449), .ZN(n7122) );
  OR2_X1 U7567 ( .A1(n8750), .A2(n7122), .ZN(n7124) );
  NAND2_X1 U7568 ( .A1(n6933), .A2(n7341), .ZN(n5918) );
  AND2_X1 U7569 ( .A1(n7124), .A2(n5918), .ZN(n5919) );
  NAND2_X1 U7570 ( .A1(n6617), .A2(n8529), .ZN(n5922) );
  OR2_X1 U7571 ( .A1(n5920), .A2(n5801), .ZN(n5932) );
  XNOR2_X1 U7572 ( .A(n5932), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10028) );
  AOI22_X1 U7573 ( .A1(n6049), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6634), .B2(
        n10028), .ZN(n5921) );
  INV_X1 U7574 ( .A(n5923), .ZN(n5925) );
  INV_X1 U7575 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7576 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  NAND2_X1 U7577 ( .A1(n5936), .A2(n5926), .ZN(n10424) );
  INV_X1 U7578 ( .A(n10424), .ZN(n10453) );
  NAND2_X1 U7579 ( .A1(n6154), .A2(n10453), .ZN(n5930) );
  NAND2_X1 U7580 ( .A1(n8536), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7581 ( .A1(n6198), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7582 ( .A1(n8537), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5927) );
  OR2_X1 U7583 ( .A1(n10449), .A2(n7362), .ZN(n8748) );
  NAND2_X1 U7584 ( .A1(n10449), .A2(n7362), .ZN(n8641) );
  NAND2_X1 U7585 ( .A1(n8748), .A2(n8641), .ZN(n7249) );
  NAND2_X1 U7586 ( .A1(n6623), .A2(n8529), .ZN(n5935) );
  NAND2_X1 U7587 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  NAND2_X1 U7588 ( .A1(n5933), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5944) );
  XNOR2_X1 U7589 ( .A(n5944), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7590 ( .A1(n6049), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6634), .B2(
        n6667), .ZN(n5934) );
  INV_X1 U7591 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U7592 ( .A1(n5936), .A2(n6695), .ZN(n5937) );
  AND2_X1 U7593 ( .A1(n5950), .A2(n5937), .ZN(n10440) );
  NAND2_X1 U7594 ( .A1(n6154), .A2(n10440), .ZN(n5941) );
  NAND2_X1 U7595 ( .A1(n8536), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7596 ( .A1(n8537), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7597 ( .A1(n6198), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7598 ( .A1(n10442), .A2(n7641), .ZN(n7636) );
  AND2_X1 U7599 ( .A1(n7249), .A2(n7376), .ZN(n5943) );
  INV_X1 U7600 ( .A(n7376), .ZN(n5942) );
  INV_X1 U7601 ( .A(n7362), .ZN(n9958) );
  OR2_X1 U7602 ( .A1(n10449), .A2(n9958), .ZN(n7370) );
  INV_X1 U7603 ( .A(n7641), .ZN(n9957) );
  INV_X1 U7604 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U7605 ( .A1(n5944), .A2(n9062), .ZN(n5945) );
  NAND2_X1 U7606 ( .A1(n5945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7607 ( .A(n5946), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U7608 ( .A1(n6049), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6634), .B2(
        n6709), .ZN(n5947) );
  NAND2_X1 U7609 ( .A1(n8536), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5955) );
  INV_X1 U7610 ( .A(n5948), .ZN(n5963) );
  INV_X1 U7611 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7612 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  AND2_X1 U7613 ( .A1(n5963), .A2(n5951), .ZN(n7704) );
  NAND2_X1 U7614 ( .A1(n6154), .A2(n7704), .ZN(n5954) );
  NAND2_X1 U7615 ( .A1(n8537), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7616 ( .A1(n6198), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5952) );
  INV_X1 U7617 ( .A(n7678), .ZN(n9956) );
  NAND2_X1 U7618 ( .A1(n10477), .A2(n9956), .ZN(n5956) );
  NAND2_X1 U7619 ( .A1(n6630), .A2(n8529), .ZN(n5960) );
  OR2_X1 U7620 ( .A1(n5957), .A2(n5801), .ZN(n5958) );
  XNOR2_X1 U7621 ( .A(n5958), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7622 ( .A1(n6049), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6634), .B2(
        n6721), .ZN(n5959) );
  INV_X1 U7623 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7624 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  AND2_X1 U7625 ( .A1(n5974), .A2(n5964), .ZN(n7673) );
  NAND2_X1 U7626 ( .A1(n6154), .A2(n7673), .ZN(n5968) );
  NAND2_X1 U7627 ( .A1(n8536), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7628 ( .A1(n6198), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7629 ( .A1(n8537), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7630 ( .A1(n10486), .A2(n7640), .ZN(n8652) );
  NAND2_X1 U7631 ( .A1(n8658), .A2(n8652), .ZN(n7677) );
  NAND2_X1 U7632 ( .A1(n7672), .A2(n7677), .ZN(n5970) );
  INV_X1 U7633 ( .A(n7640), .ZN(n9955) );
  OR2_X1 U7634 ( .A1(n10486), .A2(n9955), .ZN(n5969) );
  NAND2_X1 U7635 ( .A1(n5970), .A2(n5969), .ZN(n7602) );
  NAND2_X1 U7636 ( .A1(n6638), .A2(n8529), .ZN(n5973) );
  NAND2_X1 U7637 ( .A1(n5971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5982) );
  XNOR2_X1 U7638 ( .A(n5982), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U7639 ( .A1(n6049), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6634), .B2(
        n6764), .ZN(n5972) );
  NAND2_X1 U7640 ( .A1(n6198), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7641 ( .A1(n5974), .A2(n7820), .ZN(n5975) );
  AND2_X1 U7642 ( .A1(n5987), .A2(n5975), .ZN(n7824) );
  NAND2_X1 U7643 ( .A1(n6154), .A2(n7824), .ZN(n5978) );
  NAND2_X1 U7644 ( .A1(n8536), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7645 ( .A1(n8537), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5976) );
  NAND4_X1 U7646 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n9954)
         );
  AND2_X1 U7647 ( .A1(n10494), .A2(n9954), .ZN(n8832) );
  INV_X1 U7648 ( .A(n8832), .ZN(n5980) );
  INV_X1 U7649 ( .A(n10494), .ZN(n7612) );
  INV_X1 U7650 ( .A(n9954), .ZN(n6376) );
  AND2_X1 U7651 ( .A1(n7612), .A2(n6376), .ZN(n8660) );
  INV_X1 U7652 ( .A(n8755), .ZN(n7603) );
  NAND2_X1 U7653 ( .A1(n10494), .A2(n6376), .ZN(n5981) );
  NAND2_X1 U7654 ( .A1(n6732), .A2(n8529), .ZN(n5986) );
  NAND2_X1 U7655 ( .A1(n5982), .A2(n5771), .ZN(n5983) );
  NAND2_X1 U7656 ( .A1(n5983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U7657 ( .A(n5984), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U7658 ( .A1(n6049), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6634), .B2(
        n6817), .ZN(n5985) );
  NAND2_X1 U7659 ( .A1(n5986), .A2(n5985), .ZN(n7916) );
  INV_X1 U7660 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U7661 ( .A1(n5987), .A2(n6768), .ZN(n5988) );
  AND2_X1 U7662 ( .A1(n5989), .A2(n5988), .ZN(n7514) );
  NAND2_X1 U7663 ( .A1(n6154), .A2(n7514), .ZN(n5993) );
  NAND2_X1 U7664 ( .A1(n8536), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7665 ( .A1(n6198), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7666 ( .A1(n8537), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5990) );
  NOR2_X1 U7667 ( .A1(n7916), .A2(n9952), .ZN(n8664) );
  INV_X1 U7668 ( .A(n8664), .ZN(n8655) );
  NAND2_X1 U7669 ( .A1(n7916), .A2(n9952), .ZN(n8663) );
  INV_X1 U7670 ( .A(n7916), .ZN(n10501) );
  NAND2_X1 U7671 ( .A1(n7505), .A2(n4565), .ZN(n7619) );
  OR2_X1 U7672 ( .A1(n7768), .A2(n9950), .ZN(n8666) );
  NAND2_X1 U7673 ( .A1(n7768), .A2(n9950), .ZN(n8838) );
  NAND2_X1 U7674 ( .A1(n8666), .A2(n8838), .ZN(n8758) );
  NOR2_X1 U7675 ( .A1(n7619), .A2(n7620), .ZN(n7618) );
  AOI21_X1 U7676 ( .B1(n10511), .B2(n9950), .A(n7618), .ZN(n10431) );
  NAND2_X1 U7677 ( .A1(n6857), .A2(n8529), .ZN(n5999) );
  NOR2_X1 U7678 ( .A1(n5995), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6008) );
  INV_X1 U7679 ( .A(n6008), .ZN(n5996) );
  NAND2_X1 U7680 ( .A1(n5996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7681 ( .A(n5997), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U7682 ( .A1(n6049), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6634), .B2(
        n7234), .ZN(n5998) );
  NAND2_X1 U7683 ( .A1(n8536), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6006) );
  INV_X1 U7684 ( .A(n6000), .ZN(n6013) );
  NAND2_X1 U7685 ( .A1(n6001), .A2(n7190), .ZN(n6002) );
  AND2_X1 U7686 ( .A1(n6013), .A2(n6002), .ZN(n10429) );
  NAND2_X1 U7687 ( .A1(n6154), .A2(n10429), .ZN(n6005) );
  NAND2_X1 U7688 ( .A1(n8537), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7689 ( .A1(n6198), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6003) );
  OR2_X1 U7690 ( .A1(n10432), .A2(n7868), .ZN(n8682) );
  NAND2_X1 U7691 ( .A1(n10432), .A2(n7868), .ZN(n8837) );
  INV_X1 U7692 ( .A(n7868), .ZN(n9949) );
  NAND2_X1 U7693 ( .A1(n6897), .A2(n8529), .ZN(n6011) );
  NAND2_X1 U7694 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7695 ( .A1(n6009), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  XNOR2_X1 U7696 ( .A(n6020), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7389) );
  AOI22_X1 U7697 ( .A1(n7389), .A2(n6634), .B1(n6049), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7698 ( .A1(n8536), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6018) );
  INV_X1 U7699 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7700 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  AND2_X1 U7701 ( .A1(n6025), .A2(n6014), .ZN(n8041) );
  NAND2_X1 U7702 ( .A1(n6154), .A2(n8041), .ZN(n6017) );
  NAND2_X1 U7703 ( .A1(n8537), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7704 ( .A1(n6198), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6015) );
  INV_X1 U7705 ( .A(n7856), .ZN(n9948) );
  NAND2_X1 U7706 ( .A1(n7042), .A2(n8529), .ZN(n6024) );
  NAND2_X1 U7707 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7708 ( .A1(n6021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7709 ( .A(n6022), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7713) );
  AOI22_X1 U7710 ( .A1(n7713), .A2(n6634), .B1(n6049), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6023) );
  INV_X1 U7711 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U7712 ( .A1(n6025), .A2(n9924), .ZN(n6026) );
  NAND2_X1 U7713 ( .A1(n6039), .A2(n6026), .ZN(n7860) );
  INV_X1 U7714 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6027) );
  OAI22_X1 U7715 ( .A1(n7860), .A2(n6111), .B1(n6152), .B2(n6027), .ZN(n6031)
         );
  INV_X1 U7716 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6029) );
  INV_X1 U7717 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6028) );
  OAI22_X1 U7718 ( .A1(n8540), .A2(n6029), .B1(n6124), .B2(n6028), .ZN(n6030)
         );
  NAND2_X1 U7719 ( .A1(n6032), .A2(n8675), .ZN(n6033) );
  NAND2_X1 U7720 ( .A1(n7213), .A2(n8529), .ZN(n6037) );
  INV_X1 U7721 ( .A(n4511), .ZN(n6034) );
  NAND2_X1 U7722 ( .A1(n6034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6035) );
  XNOR2_X1 U7723 ( .A(n6035), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7808) );
  AOI22_X1 U7724 ( .A1(n6049), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6634), .B2(
        n7808), .ZN(n6036) );
  NAND2_X1 U7725 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  AND2_X1 U7726 ( .A1(n6041), .A2(n6040), .ZN(n9843) );
  NAND2_X1 U7727 ( .A1(n9843), .A2(n6154), .ZN(n6044) );
  AOI22_X1 U7728 ( .A1(n8536), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8537), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7729 ( .A1(n6198), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7730 ( .A1(n9848), .A2(n8153), .ZN(n8688) );
  NAND2_X1 U7731 ( .A1(n9848), .A2(n8153), .ZN(n8689) );
  NAND2_X1 U7732 ( .A1(n8688), .A2(n8689), .ZN(n8763) );
  INV_X1 U7733 ( .A(n8153), .ZN(n9946) );
  NAND2_X1 U7734 ( .A1(n7314), .A2(n8529), .ZN(n6051) );
  OR2_X1 U7735 ( .A1(n6046), .A2(n6160), .ZN(n6047) );
  AND2_X1 U7736 ( .A1(n6048), .A2(n6047), .ZN(n8106) );
  AOI22_X1 U7737 ( .A1(n6049), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6634), .B2(
        n8106), .ZN(n6050) );
  XNOR2_X1 U7738 ( .A(n6052), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U7739 ( .A1(n9901), .A2(n6154), .ZN(n6057) );
  INV_X1 U7740 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U7741 ( .A1(n6198), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7742 ( .A1(n8537), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6053) );
  OAI211_X1 U7743 ( .C1(n10271), .C2(n6152), .A(n6054), .B(n6053), .ZN(n6055)
         );
  INV_X1 U7744 ( .A(n6055), .ZN(n6056) );
  INV_X1 U7745 ( .A(n9815), .ZN(n9944) );
  NAND2_X1 U7746 ( .A1(n10208), .A2(n6059), .ZN(n6060) );
  NAND2_X1 U7747 ( .A1(n10206), .A2(n6060), .ZN(n6061) );
  NAND2_X1 U7748 ( .A1(n7523), .A2(n8529), .ZN(n6063) );
  OR2_X1 U7749 ( .A1(n8530), .A2(n7524), .ZN(n6062) );
  INV_X1 U7750 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7751 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  AND2_X1 U7752 ( .A1(n6077), .A2(n6066), .ZN(n10178) );
  NAND2_X1 U7753 ( .A1(n10178), .A2(n6154), .ZN(n6071) );
  INV_X1 U7754 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U7755 ( .A1(n8536), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7756 ( .A1(n8537), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U7757 ( .C1(n8540), .C2(n9236), .A(n6068), .B(n6067), .ZN(n6069)
         );
  INV_X1 U7758 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7759 ( .A1(n10177), .A2(n5021), .ZN(n6072) );
  NAND2_X1 U7760 ( .A1(n7812), .A2(n8529), .ZN(n6074) );
  OR2_X1 U7761 ( .A1(n8530), .A2(n7813), .ZN(n6073) );
  NAND2_X2 U7762 ( .A1(n6074), .A2(n6073), .ZN(n10159) );
  INV_X1 U7763 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7764 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  NAND2_X1 U7765 ( .A1(n6087), .A2(n6078), .ZN(n10160) );
  OR2_X1 U7766 ( .A1(n10160), .A2(n6111), .ZN(n6083) );
  INV_X1 U7767 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U7768 ( .A1(n6198), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7769 ( .A1(n8537), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6079) );
  OAI211_X1 U7770 ( .C1(n10250), .C2(n6152), .A(n6080), .B(n6079), .ZN(n6081)
         );
  INV_X1 U7771 ( .A(n6081), .ZN(n6082) );
  NAND2_X1 U7772 ( .A1(n6206), .A2(n9827), .ZN(n6084) );
  AOI22_X1 U7773 ( .A1(n10155), .A2(n6084), .B1(n9941), .B2(n10159), .ZN(
        n10139) );
  NAND2_X1 U7774 ( .A1(n7778), .A2(n8529), .ZN(n6086) );
  OR2_X1 U7775 ( .A1(n8530), .A2(n9285), .ZN(n6085) );
  NAND2_X1 U7776 ( .A1(n6086), .A2(n6085), .ZN(n6190) );
  INV_X1 U7777 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U7778 ( .A1(n6087), .A2(n9808), .ZN(n6088) );
  AND2_X1 U7779 ( .A1(n6099), .A2(n6088), .ZN(n10143) );
  INV_X1 U7780 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U7781 ( .A1(n6198), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7782 ( .A1(n8537), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7783 ( .C1(n10245), .C2(n6152), .A(n6090), .B(n6089), .ZN(n6091)
         );
  AOI21_X1 U7784 ( .B1(n10143), .B2(n6154), .A(n6091), .ZN(n9886) );
  INV_X1 U7785 ( .A(n9886), .ZN(n9940) );
  NAND2_X1 U7786 ( .A1(n10142), .A2(n9940), .ZN(n6093) );
  NOR2_X1 U7787 ( .A1(n10142), .A2(n9940), .ZN(n6092) );
  AOI21_X1 U7788 ( .B1(n10139), .B2(n6093), .A(n6092), .ZN(n10123) );
  NAND2_X1 U7789 ( .A1(n6094), .A2(n8529), .ZN(n6096) );
  OR2_X1 U7790 ( .A1(n8530), .A2(n7884), .ZN(n6095) );
  INV_X1 U7791 ( .A(n6099), .ZN(n6097) );
  NAND2_X1 U7792 ( .A1(n6097), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6109) );
  INV_X1 U7793 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7794 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  NAND2_X1 U7795 ( .A1(n6109), .A2(n6100), .ZN(n10125) );
  OR2_X1 U7796 ( .A1(n10125), .A2(n6111), .ZN(n6105) );
  INV_X1 U7797 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U7798 ( .A1(n6198), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7799 ( .A1(n8537), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U7800 ( .C1(n10240), .C2(n6152), .A(n6102), .B(n6101), .ZN(n6103)
         );
  INV_X1 U7801 ( .A(n6103), .ZN(n6104) );
  NAND2_X1 U7802 ( .A1(n4881), .A2(n9834), .ZN(n6106) );
  NAND2_X1 U7803 ( .A1(n7956), .A2(n8529), .ZN(n6108) );
  OR2_X1 U7804 ( .A1(n8530), .A2(n7958), .ZN(n6107) );
  INV_X1 U7805 ( .A(n10304), .ZN(n10113) );
  INV_X1 U7806 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U7807 ( .A1(n6109), .A2(n9836), .ZN(n6110) );
  NAND2_X1 U7808 ( .A1(n6120), .A2(n6110), .ZN(n10109) );
  INV_X1 U7809 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U7810 ( .A1(n8536), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7811 ( .A1(n6198), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7812 ( .C1(n6124), .C2(n10302), .A(n6113), .B(n6112), .ZN(n6114)
         );
  INV_X1 U7813 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7814 ( .A1(n6116), .A2(n6115), .ZN(n9938) );
  NAND2_X1 U7815 ( .A1(n10113), .A2(n9938), .ZN(n6117) );
  NAND2_X1 U7816 ( .A1(n8055), .A2(n8529), .ZN(n6119) );
  OR2_X1 U7817 ( .A1(n8530), .A2(n9258), .ZN(n6118) );
  INV_X1 U7818 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U7819 ( .A1(n6120), .A2(n9913), .ZN(n6121) );
  NAND2_X1 U7820 ( .A1(n10096), .A2(n6154), .ZN(n6127) );
  INV_X1 U7821 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U7822 ( .A1(n8536), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7823 ( .A1(n6198), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6122) );
  OAI211_X1 U7824 ( .C1(n6124), .C2(n10298), .A(n6123), .B(n6122), .ZN(n6125)
         );
  INV_X1 U7825 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7826 ( .A1(n10300), .A2(n9835), .ZN(n6128) );
  NAND2_X1 U7827 ( .A1(n8091), .A2(n8529), .ZN(n6130) );
  OR2_X1 U7828 ( .A1(n8530), .A2(n8141), .ZN(n6129) );
  XNOR2_X1 U7829 ( .A(n6141), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n10081) );
  INV_X1 U7830 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10224) );
  NAND2_X1 U7831 ( .A1(n8537), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7832 ( .A1(n6198), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6131) );
  OAI211_X1 U7833 ( .C1(n6152), .C2(n10224), .A(n6132), .B(n6131), .ZN(n6133)
         );
  AOI21_X1 U7834 ( .B1(n10081), .B2(n6154), .A(n6133), .ZN(n9909) );
  INV_X1 U7835 ( .A(n9909), .ZN(n9936) );
  INV_X1 U7836 ( .A(n8785), .ZN(n6134) );
  NAND2_X1 U7837 ( .A1(n10080), .A2(n9909), .ZN(n6246) );
  NAND2_X1 U7838 ( .A1(n6134), .A2(n6246), .ZN(n10075) );
  NAND2_X1 U7839 ( .A1(n10074), .A2(n6135), .ZN(n6245) );
  NAND2_X1 U7840 ( .A1(n8190), .A2(n8529), .ZN(n6137) );
  OR2_X1 U7841 ( .A1(n8530), .A2(n8892), .ZN(n6136) );
  INV_X1 U7842 ( .A(n6141), .ZN(n6139) );
  AND2_X1 U7843 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6138) );
  NAND2_X1 U7844 ( .A1(n6139), .A2(n6138), .ZN(n10049) );
  INV_X1 U7845 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6568) );
  INV_X1 U7846 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7847 ( .B1(n6141), .B2(n6568), .A(n6140), .ZN(n6142) );
  INV_X1 U7848 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7849 ( .A1(n8537), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7850 ( .A1(n6198), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6143) );
  OAI211_X1 U7851 ( .C1(n6152), .C2(n6554), .A(n6144), .B(n6143), .ZN(n6145)
         );
  AOI21_X1 U7852 ( .B1(n10059), .B2(n6154), .A(n6145), .ZN(n6565) );
  INV_X1 U7853 ( .A(n6565), .ZN(n9935) );
  NAND2_X1 U7854 ( .A1(n6548), .A2(n9935), .ZN(n6147) );
  NOR2_X1 U7855 ( .A1(n6548), .A2(n9935), .ZN(n6146) );
  AOI21_X1 U7856 ( .B1(n6245), .B2(n6147), .A(n6146), .ZN(n6156) );
  NAND2_X1 U7857 ( .A1(n8881), .A2(n8529), .ZN(n6149) );
  OR2_X1 U7858 ( .A1(n8530), .A2(n8882), .ZN(n6148) );
  INV_X1 U7859 ( .A(n10049), .ZN(n6155) );
  INV_X1 U7860 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7861 ( .A1(n8537), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7862 ( .A1(n6198), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6150) );
  OAI211_X1 U7863 ( .C1(n6152), .C2(n6241), .A(n6151), .B(n6150), .ZN(n6153)
         );
  AOI21_X1 U7864 ( .B1(n6155), .B2(n6154), .A(n6153), .ZN(n6248) );
  NAND2_X1 U7865 ( .A1(n10053), .A2(n6248), .ZN(n8802) );
  OR2_X1 U7866 ( .A1(n10053), .A2(n6248), .ZN(n8800) );
  INV_X1 U7867 ( .A(n8732), .ZN(n8777) );
  XNOR2_X1 U7868 ( .A(n6156), .B(n8777), .ZN(n10047) );
  NAND2_X1 U7869 ( .A1(n6162), .A2(n6161), .ZN(n6167) );
  NAND2_X1 U7870 ( .A1(n6164), .A2(n6163), .ZN(n6223) );
  NAND2_X1 U7871 ( .A1(n6167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6168) );
  MUX2_X1 U7872 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6168), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6169) );
  NAND2_X1 U7873 ( .A1(n6169), .A2(n4532), .ZN(n6532) );
  INV_X1 U7874 ( .A(n6265), .ZN(n8876) );
  NAND2_X1 U7875 ( .A1(n4532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7876 ( .A(n6170), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7877 ( .A1(n8876), .A2(n4526), .ZN(n8807) );
  INV_X1 U7878 ( .A(n8807), .ZN(n6636) );
  NAND2_X1 U7879 ( .A1(n6636), .A2(n6266), .ZN(n8873) );
  NAND2_X1 U7880 ( .A1(n6265), .A2(n6166), .ZN(n8737) );
  OR2_X1 U7881 ( .A1(n10477), .A2(n7678), .ZN(n7674) );
  NAND2_X1 U7882 ( .A1(n8658), .A2(n7674), .ZN(n8753) );
  NAND2_X1 U7883 ( .A1(n10477), .A2(n7678), .ZN(n8648) );
  AND2_X1 U7884 ( .A1(n8648), .A2(n7636), .ZN(n8646) );
  OR2_X1 U7885 ( .A1(n8753), .A2(n8646), .ZN(n6171) );
  NAND2_X1 U7886 ( .A1(n6171), .A2(n8652), .ZN(n6180) );
  INV_X1 U7887 ( .A(n8641), .ZN(n6172) );
  NAND2_X1 U7888 ( .A1(n8823), .A2(n8822), .ZN(n6173) );
  INV_X1 U7889 ( .A(n8631), .ZN(n6175) );
  NAND2_X1 U7890 ( .A1(n6175), .A2(n8824), .ZN(n8820) );
  OAI21_X1 U7891 ( .B1(n8820), .B2(n8746), .A(n8825), .ZN(n6931) );
  NAND2_X1 U7892 ( .A1(n6931), .A2(n8637), .ZN(n7129) );
  INV_X1 U7893 ( .A(n8635), .ZN(n6176) );
  NOR2_X1 U7894 ( .A1(n7130), .A2(n6176), .ZN(n6177) );
  NAND2_X1 U7895 ( .A1(n7129), .A2(n6177), .ZN(n7132) );
  AND2_X2 U7896 ( .A1(n7132), .A2(n8638), .ZN(n7377) );
  NAND2_X1 U7897 ( .A1(n8749), .A2(n8748), .ZN(n6178) );
  NOR2_X1 U7898 ( .A1(n8753), .A2(n6178), .ZN(n6179) );
  OR2_X1 U7899 ( .A1(n6180), .A2(n6179), .ZN(n8830) );
  NAND2_X1 U7900 ( .A1(n6181), .A2(n8837), .ZN(n7867) );
  OR2_X1 U7901 ( .A1(n7874), .A2(n7856), .ZN(n8683) );
  AND2_X1 U7902 ( .A1(n7874), .A2(n7856), .ZN(n8685) );
  INV_X1 U7903 ( .A(n8685), .ZN(n8671) );
  NAND2_X1 U7904 ( .A1(n7866), .A2(n8671), .ZN(n7855) );
  XNOR2_X1 U7905 ( .A(n10281), .B(n8675), .ZN(n8762) );
  NAND2_X1 U7906 ( .A1(n6032), .A2(n9947), .ZN(n8687) );
  NAND2_X1 U7907 ( .A1(n10275), .A2(n8205), .ZN(n8701) );
  INV_X1 U7908 ( .A(n8765), .ZN(n6183) );
  INV_X1 U7909 ( .A(n8689), .ZN(n6182) );
  NOR2_X1 U7910 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  OR2_X1 U7911 ( .A1(n8212), .A2(n9815), .ZN(n8705) );
  NAND2_X1 U7912 ( .A1(n8212), .A2(n9815), .ZN(n8702) );
  AND2_X1 U7913 ( .A1(n8705), .A2(n8702), .ZN(n8766) );
  OR2_X1 U7914 ( .A1(n10208), .A2(n6441), .ZN(n8706) );
  AND2_X1 U7915 ( .A1(n10208), .A2(n6441), .ZN(n8707) );
  INV_X1 U7916 ( .A(n8707), .ZN(n8856) );
  NAND2_X1 U7917 ( .A1(n8706), .A2(n8856), .ZN(n10205) );
  AND2_X1 U7918 ( .A1(n10322), .A2(n9943), .ZN(n8700) );
  AND2_X1 U7919 ( .A1(n10197), .A2(n9826), .ZN(n8708) );
  INV_X1 U7920 ( .A(n8708), .ZN(n6187) );
  NAND2_X1 U7921 ( .A1(n6188), .A2(n8712), .ZN(n10167) );
  OR2_X2 U7922 ( .A1(n10167), .A2(n10174), .ZN(n10169) );
  NAND2_X1 U7923 ( .A1(n10177), .A2(n9888), .ZN(n8697) );
  OR2_X1 U7924 ( .A1(n10159), .A2(n9827), .ZN(n8613) );
  NAND2_X1 U7925 ( .A1(n10159), .A2(n9827), .ZN(n8787) );
  NAND2_X1 U7926 ( .A1(n8613), .A2(n8787), .ZN(n8616) );
  NAND2_X1 U7927 ( .A1(n10149), .A2(n10154), .ZN(n6189) );
  NAND2_X1 U7928 ( .A1(n6189), .A2(n8787), .ZN(n10133) );
  NAND2_X1 U7929 ( .A1(n6190), .A2(n9886), .ZN(n10116) );
  NAND2_X1 U7930 ( .A1(n8615), .A2(n10116), .ZN(n10138) );
  INV_X1 U7931 ( .A(n10138), .ZN(n10134) );
  NAND2_X1 U7932 ( .A1(n10124), .A2(n9834), .ZN(n8789) );
  NAND2_X1 U7933 ( .A1(n10102), .A2(n8789), .ZN(n10117) );
  INV_X1 U7934 ( .A(n10116), .ZN(n8790) );
  NOR2_X1 U7935 ( .A1(n10117), .A2(n8790), .ZN(n6191) );
  NAND2_X1 U7936 ( .A1(n10132), .A2(n6191), .ZN(n10119) );
  AND2_X1 U7937 ( .A1(n10304), .A2(n9938), .ZN(n8721) );
  NAND2_X1 U7938 ( .A1(n4785), .A2(n10102), .ZN(n8797) );
  INV_X1 U7939 ( .A(n8797), .ZN(n6192) );
  NAND2_X1 U7940 ( .A1(n10119), .A2(n6192), .ZN(n6193) );
  NAND2_X1 U7941 ( .A1(n10113), .A2(n6500), .ZN(n8792) );
  NAND2_X1 U7942 ( .A1(n6193), .A2(n8792), .ZN(n10088) );
  OR2_X1 U7943 ( .A1(n10095), .A2(n9835), .ZN(n8725) );
  NAND2_X1 U7944 ( .A1(n10095), .A2(n9835), .ZN(n8818) );
  NAND2_X1 U7945 ( .A1(n8725), .A2(n8818), .ZN(n10087) );
  INV_X1 U7946 ( .A(n10087), .ZN(n10092) );
  INV_X1 U7947 ( .A(n10075), .ZN(n10069) );
  NAND2_X1 U7948 ( .A1(n6548), .A2(n6565), .ZN(n6244) );
  AND2_X1 U7949 ( .A1(n6244), .A2(n6246), .ZN(n8735) );
  OR2_X1 U7950 ( .A1(n6548), .A2(n6565), .ZN(n8799) );
  OR2_X1 U7951 ( .A1(n6265), .A2(n8816), .ZN(n6196) );
  NAND2_X1 U7952 ( .A1(n4526), .A2(n8871), .ZN(n6195) );
  NAND2_X1 U7953 ( .A1(n8536), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7954 ( .A1(n6198), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7955 ( .A1(n8537), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6199) );
  AND3_X1 U7956 ( .A1(n6201), .A2(n6200), .A3(n6199), .ZN(n8775) );
  OR2_X1 U7957 ( .A1(n8142), .A2(n6211), .ZN(n6202) );
  NAND2_X1 U7958 ( .A1(n9865), .A2(n6202), .ZN(n8535) );
  OAI22_X1 U7959 ( .A1(n6565), .A2(n9887), .B1(n8775), .B2(n8535), .ZN(n6203)
         );
  AOI21_X1 U7960 ( .B1(n6204), .B2(n10427), .A(n6203), .ZN(n10056) );
  INV_X1 U7961 ( .A(n10053), .ZN(n6593) );
  NAND2_X1 U7962 ( .A1(n6205), .A2(n7492), .ZN(n7491) );
  NAND2_X1 U7963 ( .A1(n6901), .A2(n7427), .ZN(n6936) );
  OAI211_X1 U7964 ( .C1(n6593), .C2(n4550), .A(n10435), .B(n10042), .ZN(n10050) );
  NAND2_X1 U7965 ( .A1(n10056), .A2(n10050), .ZN(n6207) );
  AOI21_X1 U7966 ( .B1(n10047), .B2(n10520), .A(n6207), .ZN(n6597) );
  INV_X1 U7967 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7968 ( .A1(n6209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6210) );
  NOR2_X1 U7969 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6212) );
  NAND2_X1 U7970 ( .A1(n6213), .A2(n6212), .ZN(n6217) );
  NOR2_X1 U7971 ( .A1(n5801), .A2(n5779), .ZN(n6216) );
  MUX2_X1 U7972 ( .A(P1_B_REG_SCAN_IN), .B(n6218), .S(n7885), .Z(n6220) );
  OR2_X1 U7973 ( .A1(n6239), .A2(n7957), .ZN(n10335) );
  OAI21_X1 U7974 ( .B1(n10334), .B2(P1_D_REG_1__SCAN_IN), .A(n10335), .ZN(
        n6521) );
  NOR2_X1 U7975 ( .A1(n8807), .A2(n6266), .ZN(n6535) );
  NOR2_X1 U7976 ( .A1(n7406), .A2(n6528), .ZN(n6236) );
  NOR4_X1 U7977 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6234) );
  NOR4_X1 U7978 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6233) );
  INV_X1 U7979 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10467) );
  INV_X1 U7980 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10466) );
  INV_X1 U7981 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10463) );
  INV_X1 U7982 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U7983 ( .A1(n10467), .A2(n10466), .A3(n10463), .A4(n10465), .ZN(
        n6231) );
  NOR4_X1 U7984 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6229) );
  NOR4_X1 U7985 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7986 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6227) );
  NOR4_X1 U7987 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6226) );
  NAND4_X1 U7988 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6230)
         );
  NOR4_X1 U7989 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6231), .A4(n6230), .ZN(n6232) );
  NAND3_X1 U7990 ( .A1(n6234), .A2(n6233), .A3(n6232), .ZN(n6235) );
  NAND2_X1 U7991 ( .A1(n6238), .A2(n6235), .ZN(n6522) );
  INV_X1 U7992 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7993 ( .A1(n6238), .A2(n6237), .ZN(n6240) );
  INV_X1 U7994 ( .A(n6239), .ZN(n8056) );
  NAND2_X1 U7995 ( .A1(n7885), .A2(n8056), .ZN(n10336) );
  OAI21_X1 U7996 ( .B1(n6597), .B2(n10534), .A(n6243), .ZN(P1_U3551) );
  NAND2_X1 U7997 ( .A1(n8799), .A2(n6244), .ZN(n8774) );
  AOI211_X1 U7998 ( .C1(n6548), .C2(n10077), .A(n10502), .B(n4550), .ZN(n10063) );
  NAND2_X1 U7999 ( .A1(n10067), .A2(n6246), .ZN(n6247) );
  XNOR2_X1 U8000 ( .A(n6247), .B(n8774), .ZN(n6249) );
  INV_X1 U8001 ( .A(n6248), .ZN(n9934) );
  AOI22_X1 U8002 ( .A1(n9936), .A2(n9910), .B1(n9934), .B2(n9865), .ZN(n6543)
         );
  OAI21_X1 U8003 ( .B1(n6249), .B2(n10203), .A(n6543), .ZN(n10057) );
  INV_X1 U8004 ( .A(n7407), .ZN(n6251) );
  INV_X1 U8005 ( .A(n6548), .ZN(n10061) );
  INV_X1 U8006 ( .A(n10517), .ZN(n10282) );
  INV_X1 U8007 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6252) );
  XNOR2_X1 U8008 ( .A(n6255), .B(n8507), .ZN(n6259) );
  MUX2_X1 U8009 ( .A(n6260), .B(n9674), .S(n10649), .Z(n6263) );
  NAND2_X1 U8010 ( .A1(n8601), .A2(n6261), .ZN(n6262) );
  NAND2_X1 U8011 ( .A1(n6263), .A2(n6262), .ZN(P2_U3454) );
  INV_X1 U8012 ( .A(n6264), .ZN(n6266) );
  AND2_X2 U8013 ( .A1(n6267), .A2(n6532), .ZN(n6272) );
  NAND3_X4 U8014 ( .A1(n6268), .A2(n6274), .A3(n7493), .ZN(n6514) );
  NAND2_X1 U8015 ( .A1(n9963), .A2(n6327), .ZN(n6270) );
  NAND2_X1 U8016 ( .A1(n6354), .A2(n8822), .ZN(n6269) );
  INV_X1 U8017 ( .A(n6272), .ZN(n6273) );
  NAND2_X4 U8018 ( .A1(n6276), .A2(n6275), .ZN(n6517) );
  NAND2_X1 U8019 ( .A1(n4521), .A2(n6277), .ZN(n6279) );
  NAND2_X1 U8020 ( .A1(n9963), .A2(n6354), .ZN(n6278) );
  NAND2_X1 U8021 ( .A1(n6279), .A2(n6278), .ZN(n6280) );
  OAI21_X1 U8022 ( .B1(n6282), .B2(n6281), .A(n6295), .ZN(n6803) );
  INV_X1 U8023 ( .A(n6803), .ZN(n6294) );
  NAND2_X1 U8024 ( .A1(n9964), .A2(n6327), .ZN(n6286) );
  INV_X1 U8025 ( .A(n6274), .ZN(n6536) );
  NAND2_X1 U8026 ( .A1(n6536), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U8027 ( .A1(n6286), .A2(n6285), .ZN(n6779) );
  NAND2_X1 U8028 ( .A1(n6296), .A2(n7435), .ZN(n6288) );
  NAND2_X1 U8029 ( .A1(n9964), .A2(n6354), .ZN(n6287) );
  AND2_X1 U8030 ( .A1(n6288), .A2(n6287), .ZN(n6290) );
  NAND2_X1 U8031 ( .A1(n6536), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U8032 ( .A1(n6290), .A2(n6289), .ZN(n6778) );
  NAND2_X1 U8033 ( .A1(n6779), .A2(n6778), .ZN(n6292) );
  NAND2_X1 U8034 ( .A1(n6290), .A2(n4514), .ZN(n6291) );
  NAND2_X1 U8035 ( .A1(n6292), .A2(n6291), .ZN(n6805) );
  NAND2_X1 U8036 ( .A1(n6294), .A2(n6293), .ZN(n6804) );
  INV_X1 U8037 ( .A(n6295), .ZN(n6828) );
  NAND2_X1 U8038 ( .A1(n6804), .A2(n6295), .ZN(n6307) );
  NAND2_X1 U8039 ( .A1(n6296), .A2(n5879), .ZN(n6298) );
  NAND2_X1 U8040 ( .A1(n9962), .A2(n6354), .ZN(n6297) );
  NAND2_X1 U8041 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  INV_X1 U8042 ( .A(n6305), .ZN(n6303) );
  NAND2_X1 U8043 ( .A1(n9962), .A2(n6327), .ZN(n6301) );
  NAND2_X1 U8044 ( .A1(n6354), .A2(n5879), .ZN(n6300) );
  AND2_X1 U8045 ( .A1(n6301), .A2(n6300), .ZN(n6304) );
  INV_X1 U8046 ( .A(n6304), .ZN(n6302) );
  NAND2_X1 U8047 ( .A1(n6303), .A2(n6302), .ZN(n6306) );
  NAND2_X1 U8048 ( .A1(n6305), .A2(n6304), .ZN(n6308) );
  AND2_X1 U8049 ( .A1(n6306), .A2(n6308), .ZN(n6827) );
  NAND2_X1 U8050 ( .A1(n6307), .A2(n6827), .ZN(n6830) );
  NAND2_X1 U8051 ( .A1(n6830), .A2(n6308), .ZN(n6871) );
  NAND2_X1 U8052 ( .A1(n6296), .A2(n5891), .ZN(n6309) );
  OAI21_X1 U8053 ( .B1(n6932), .B2(n4527), .A(n6309), .ZN(n6310) );
  XNOR2_X1 U8054 ( .A(n6310), .B(n4514), .ZN(n6315) );
  OR2_X1 U8055 ( .A1(n6932), .A2(n6514), .ZN(n6312) );
  NAND2_X1 U8056 ( .A1(n6354), .A2(n5891), .ZN(n6311) );
  NAND2_X1 U8057 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  XNOR2_X1 U8058 ( .A(n6315), .B(n6313), .ZN(n6872) );
  INV_X1 U8059 ( .A(n6313), .ZN(n6314) );
  NAND2_X1 U8060 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U8061 ( .A1(n6296), .A2(n6937), .ZN(n6317) );
  OAI21_X1 U8062 ( .B1(n7134), .B2(n4527), .A(n6317), .ZN(n6318) );
  XNOR2_X1 U8063 ( .A(n6318), .B(n6517), .ZN(n6323) );
  OR2_X1 U8064 ( .A1(n7134), .A2(n6514), .ZN(n6320) );
  NAND2_X1 U8065 ( .A1(n6354), .A2(n6937), .ZN(n6319) );
  NAND2_X1 U8066 ( .A1(n6320), .A2(n6319), .ZN(n6322) );
  XNOR2_X1 U8067 ( .A(n6323), .B(n6322), .ZN(n7229) );
  NAND2_X1 U8068 ( .A1(n6323), .A2(n6322), .ZN(n6330) );
  INV_X1 U8069 ( .A(n6296), .ZN(n6498) );
  NAND2_X1 U8070 ( .A1(n9959), .A2(n6354), .ZN(n6324) );
  OAI21_X1 U8071 ( .B1(n7341), .B2(n6498), .A(n6324), .ZN(n6325) );
  XNOR2_X1 U8072 ( .A(n6325), .B(n4514), .ZN(n6331) );
  AND2_X1 U8073 ( .A1(n6330), .A2(n6331), .ZN(n6326) );
  NAND2_X1 U8074 ( .A1(n7227), .A2(n6326), .ZN(n7342) );
  OR2_X1 U8075 ( .A1(n7341), .A2(n4527), .ZN(n6329) );
  NAND2_X1 U8076 ( .A1(n9959), .A2(n6327), .ZN(n6328) );
  NAND2_X1 U8077 ( .A1(n6329), .A2(n6328), .ZN(n7345) );
  NAND2_X1 U8078 ( .A1(n7342), .A2(n7345), .ZN(n6334) );
  NAND2_X1 U8079 ( .A1(n7227), .A2(n6330), .ZN(n6333) );
  INV_X1 U8080 ( .A(n6331), .ZN(n6332) );
  NAND2_X1 U8081 ( .A1(n6333), .A2(n6332), .ZN(n7343) );
  NAND2_X1 U8082 ( .A1(n10449), .A2(n6479), .ZN(n6336) );
  OR2_X1 U8083 ( .A1(n7362), .A2(n4527), .ZN(n6335) );
  NAND2_X1 U8084 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  XNOR2_X1 U8085 ( .A(n6337), .B(n4514), .ZN(n6340) );
  NAND2_X1 U8086 ( .A1(n10449), .A2(n6354), .ZN(n6339) );
  OR2_X1 U8087 ( .A1(n7362), .A2(n6514), .ZN(n6338) );
  AND2_X1 U8088 ( .A1(n6339), .A2(n6338), .ZN(n6341) );
  NAND2_X1 U8089 ( .A1(n6340), .A2(n6341), .ZN(n6346) );
  INV_X1 U8090 ( .A(n6340), .ZN(n6343) );
  INV_X1 U8091 ( .A(n6341), .ZN(n6342) );
  NAND2_X1 U8092 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  NAND2_X1 U8093 ( .A1(n6346), .A2(n6344), .ZN(n10414) );
  INV_X1 U8094 ( .A(n10414), .ZN(n6345) );
  NAND2_X1 U8095 ( .A1(n10442), .A2(n6479), .ZN(n6348) );
  OR2_X1 U8096 ( .A1(n7641), .A2(n4527), .ZN(n6347) );
  NAND2_X1 U8097 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  XNOR2_X1 U8098 ( .A(n6349), .B(n4514), .ZN(n6352) );
  NOR2_X1 U8099 ( .A1(n7641), .A2(n6514), .ZN(n6350) );
  AOI21_X1 U8100 ( .B1(n10442), .B2(n6354), .A(n6350), .ZN(n6351) );
  NAND2_X1 U8101 ( .A1(n6352), .A2(n6351), .ZN(n7358) );
  NAND2_X1 U8102 ( .A1(n7360), .A2(n7358), .ZN(n6353) );
  OR2_X1 U8103 ( .A1(n6352), .A2(n6351), .ZN(n7359) );
  NAND2_X1 U8104 ( .A1(n10486), .A2(n6296), .ZN(n6356) );
  OR2_X1 U8105 ( .A1(n7640), .A2(n4527), .ZN(n6355) );
  NAND2_X1 U8106 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  XNOR2_X1 U8107 ( .A(n6357), .B(n4514), .ZN(n7788) );
  NAND2_X1 U8108 ( .A1(n10486), .A2(n6354), .ZN(n6359) );
  OR2_X1 U8109 ( .A1(n7640), .A2(n6514), .ZN(n6358) );
  NAND2_X1 U8110 ( .A1(n6359), .A2(n6358), .ZN(n6366) );
  INV_X1 U8111 ( .A(n6366), .ZN(n7787) );
  NAND2_X1 U8112 ( .A1(n10477), .A2(n6354), .ZN(n6361) );
  OR2_X1 U8113 ( .A1(n7678), .A2(n6514), .ZN(n6360) );
  NAND2_X1 U8114 ( .A1(n6361), .A2(n6360), .ZN(n6365) );
  INV_X1 U8115 ( .A(n6365), .ZN(n7703) );
  NAND2_X1 U8116 ( .A1(n10477), .A2(n6296), .ZN(n6363) );
  OR2_X1 U8117 ( .A1(n7678), .A2(n4527), .ZN(n6362) );
  NAND2_X1 U8118 ( .A1(n6363), .A2(n6362), .ZN(n6364) );
  XNOR2_X1 U8119 ( .A(n6364), .B(n6517), .ZN(n7786) );
  INV_X1 U8120 ( .A(n7786), .ZN(n7701) );
  OAI22_X1 U8121 ( .A1(n7788), .A2(n7787), .B1(n7703), .B2(n7701), .ZN(n6370)
         );
  OAI21_X1 U8122 ( .B1(n7786), .B2(n6365), .A(n6366), .ZN(n6368) );
  NOR2_X1 U8123 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  AOI22_X1 U8124 ( .A1(n7788), .A2(n6368), .B1(n6367), .B2(n7701), .ZN(n6369)
         );
  NAND2_X1 U8125 ( .A1(n7916), .A2(n6479), .ZN(n6372) );
  OR2_X1 U8126 ( .A1(n9952), .A2(n4527), .ZN(n6371) );
  NAND2_X1 U8127 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  XNOR2_X1 U8128 ( .A(n6373), .B(n6517), .ZN(n6381) );
  NAND2_X1 U8129 ( .A1(n7916), .A2(n6354), .ZN(n6375) );
  OR2_X1 U8130 ( .A1(n9952), .A2(n6514), .ZN(n6374) );
  NAND2_X1 U8131 ( .A1(n6375), .A2(n6374), .ZN(n7908) );
  OAI22_X1 U8132 ( .A1(n10494), .A2(n6498), .B1(n6376), .B2(n4527), .ZN(n6377)
         );
  XNOR2_X1 U8133 ( .A(n6377), .B(n6517), .ZN(n6382) );
  OR2_X1 U8134 ( .A1(n10494), .A2(n4527), .ZN(n6379) );
  NAND2_X1 U8135 ( .A1(n9954), .A2(n6327), .ZN(n6378) );
  NAND2_X1 U8136 ( .A1(n6379), .A2(n6378), .ZN(n7818) );
  AOI22_X1 U8137 ( .A1(n6381), .A2(n7908), .B1(n6382), .B2(n7818), .ZN(n6380)
         );
  OAI21_X1 U8138 ( .B1(n6382), .B2(n7818), .A(n7908), .ZN(n6384) );
  INV_X1 U8139 ( .A(n6381), .ZN(n7909) );
  INV_X1 U8140 ( .A(n6382), .ZN(n7907) );
  NOR2_X1 U8141 ( .A1(n7908), .A2(n7818), .ZN(n6383) );
  AOI22_X1 U8142 ( .A1(n6384), .A2(n7909), .B1(n7907), .B2(n6383), .ZN(n6385)
         );
  NAND2_X1 U8143 ( .A1(n7768), .A2(n6479), .ZN(n6387) );
  OR2_X1 U8144 ( .A1(n9950), .A2(n4527), .ZN(n6386) );
  NAND2_X1 U8145 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  XNOR2_X1 U8146 ( .A(n6388), .B(n6517), .ZN(n6390) );
  NOR2_X1 U8147 ( .A1(n9950), .A2(n6514), .ZN(n6389) );
  AOI21_X1 U8148 ( .B1(n7768), .B2(n6354), .A(n6389), .ZN(n6391) );
  XNOR2_X1 U8149 ( .A(n6390), .B(n6391), .ZN(n7761) );
  INV_X1 U8150 ( .A(n6390), .ZN(n6392) );
  NAND2_X1 U8151 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  NAND2_X1 U8152 ( .A1(n10432), .A2(n6479), .ZN(n6395) );
  OR2_X1 U8153 ( .A1(n7868), .A2(n4527), .ZN(n6394) );
  NAND2_X1 U8154 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  XNOR2_X1 U8155 ( .A(n6396), .B(n6517), .ZN(n6398) );
  NOR2_X1 U8156 ( .A1(n7868), .A2(n6514), .ZN(n6397) );
  AOI21_X1 U8157 ( .B1(n10432), .B2(n6354), .A(n6397), .ZN(n6399) );
  XNOR2_X1 U8158 ( .A(n6398), .B(n6399), .ZN(n7836) );
  NAND2_X1 U8159 ( .A1(n7835), .A2(n7836), .ZN(n6402) );
  INV_X1 U8160 ( .A(n6398), .ZN(n6400) );
  NAND2_X1 U8161 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  NAND2_X1 U8162 ( .A1(n6402), .A2(n6401), .ZN(n6407) );
  NAND2_X1 U8163 ( .A1(n7874), .A2(n6479), .ZN(n6404) );
  OR2_X1 U8164 ( .A1(n7856), .A2(n4527), .ZN(n6403) );
  NAND2_X1 U8165 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  XNOR2_X1 U8166 ( .A(n6405), .B(n6517), .ZN(n6408) );
  XNOR2_X1 U8167 ( .A(n6407), .B(n6408), .ZN(n8037) );
  NOR2_X1 U8168 ( .A1(n7856), .A2(n6514), .ZN(n6406) );
  AOI21_X1 U8169 ( .B1(n7874), .B2(n6354), .A(n6406), .ZN(n8039) );
  NAND2_X1 U8170 ( .A1(n8037), .A2(n8039), .ZN(n8038) );
  INV_X1 U8171 ( .A(n6408), .ZN(n6409) );
  NAND2_X1 U8172 ( .A1(n6407), .A2(n6409), .ZN(n6410) );
  NAND2_X1 U8173 ( .A1(n10281), .A2(n6479), .ZN(n6412) );
  NAND2_X1 U8174 ( .A1(n9947), .A2(n6354), .ZN(n6411) );
  NAND2_X1 U8175 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  XNOR2_X1 U8176 ( .A(n6413), .B(n6517), .ZN(n6415) );
  AND2_X1 U8177 ( .A1(n9947), .A2(n6327), .ZN(n6414) );
  AOI21_X1 U8178 ( .B1(n10281), .B2(n6354), .A(n6414), .ZN(n9921) );
  INV_X1 U8179 ( .A(n6415), .ZN(n6416) );
  NAND2_X1 U8180 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  NAND2_X1 U8181 ( .A1(n9848), .A2(n6479), .ZN(n6420) );
  OR2_X1 U8182 ( .A1(n8153), .A2(n4527), .ZN(n6419) );
  NAND2_X1 U8183 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  XNOR2_X1 U8184 ( .A(n6421), .B(n6517), .ZN(n6423) );
  NOR2_X1 U8185 ( .A1(n8153), .A2(n6514), .ZN(n6422) );
  AOI21_X1 U8186 ( .B1(n9848), .B2(n6354), .A(n6422), .ZN(n6424) );
  XNOR2_X1 U8187 ( .A(n6423), .B(n6424), .ZN(n9842) );
  INV_X1 U8188 ( .A(n6423), .ZN(n6425) );
  NAND2_X1 U8189 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  NAND2_X1 U8190 ( .A1(n10275), .A2(n6479), .ZN(n6428) );
  NAND2_X1 U8191 ( .A1(n9945), .A2(n6354), .ZN(n6427) );
  NAND2_X1 U8192 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  XNOR2_X1 U8193 ( .A(n6429), .B(n6517), .ZN(n6431) );
  NOR2_X1 U8194 ( .A1(n8205), .A2(n6514), .ZN(n6430) );
  AOI21_X1 U8195 ( .B1(n10275), .B2(n6354), .A(n6430), .ZN(n6432) );
  XNOR2_X1 U8196 ( .A(n6431), .B(n6432), .ZN(n9852) );
  INV_X1 U8197 ( .A(n6431), .ZN(n6433) );
  NAND2_X1 U8198 ( .A1(n8212), .A2(n6479), .ZN(n6435) );
  OR2_X1 U8199 ( .A1(n9815), .A2(n4527), .ZN(n6434) );
  NAND2_X1 U8200 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  XNOR2_X1 U8201 ( .A(n6436), .B(n6517), .ZN(n6448) );
  XNOR2_X1 U8202 ( .A(n6450), .B(n6448), .ZN(n9812) );
  NOR2_X1 U8203 ( .A1(n9815), .A2(n6514), .ZN(n6437) );
  AOI21_X1 U8204 ( .B1(n8212), .B2(n6354), .A(n6437), .ZN(n9896) );
  NAND2_X1 U8205 ( .A1(n10208), .A2(n6479), .ZN(n6439) );
  NAND2_X1 U8206 ( .A1(n6059), .A2(n6354), .ZN(n6438) );
  NAND2_X1 U8207 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  XNOR2_X1 U8208 ( .A(n6440), .B(n6517), .ZN(n6445) );
  INV_X1 U8209 ( .A(n6445), .ZN(n6443) );
  NOR2_X1 U8210 ( .A1(n6441), .A2(n6514), .ZN(n6442) );
  AOI21_X1 U8211 ( .B1(n10208), .B2(n6354), .A(n6442), .ZN(n6444) );
  NAND2_X1 U8212 ( .A1(n6443), .A2(n6444), .ZN(n6451) );
  INV_X1 U8213 ( .A(n6451), .ZN(n6446) );
  XNOR2_X1 U8214 ( .A(n6445), .B(n6444), .ZN(n9814) );
  OR2_X1 U8215 ( .A1(n6446), .A2(n9814), .ZN(n6453) );
  AND2_X1 U8216 ( .A1(n9896), .A2(n6453), .ZN(n6447) );
  NAND2_X1 U8217 ( .A1(n9812), .A2(n6447), .ZN(n6455) );
  INV_X1 U8218 ( .A(n6448), .ZN(n6449) );
  NAND2_X1 U8219 ( .A1(n6450), .A2(n6449), .ZN(n9813) );
  NAND2_X1 U8220 ( .A1(n9813), .A2(n6451), .ZN(n6452) );
  NAND2_X1 U8221 ( .A1(n10197), .A2(n6479), .ZN(n6457) );
  NAND2_X1 U8222 ( .A1(n9943), .A2(n6354), .ZN(n6456) );
  NAND2_X1 U8223 ( .A1(n6457), .A2(n6456), .ZN(n6458) );
  XNOR2_X1 U8224 ( .A(n6458), .B(n4514), .ZN(n9872) );
  NOR2_X1 U8225 ( .A1(n9826), .A2(n6514), .ZN(n6459) );
  AOI21_X1 U8226 ( .B1(n10197), .B2(n6354), .A(n6459), .ZN(n9871) );
  NAND2_X1 U8227 ( .A1(n10177), .A2(n6479), .ZN(n6461) );
  OR2_X1 U8228 ( .A1(n9888), .A2(n4527), .ZN(n6460) );
  NAND2_X1 U8229 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  XNOR2_X1 U8230 ( .A(n6462), .B(n4514), .ZN(n6469) );
  NOR2_X1 U8231 ( .A1(n9888), .A2(n6514), .ZN(n6463) );
  AOI21_X1 U8232 ( .B1(n10177), .B2(n6354), .A(n6463), .ZN(n6468) );
  XNOR2_X1 U8233 ( .A(n6469), .B(n6468), .ZN(n9825) );
  INV_X1 U8234 ( .A(n9825), .ZN(n6466) );
  INV_X1 U8235 ( .A(n9872), .ZN(n6465) );
  INV_X1 U8236 ( .A(n9871), .ZN(n6464) );
  NAND2_X1 U8237 ( .A1(n6465), .A2(n6464), .ZN(n9823) );
  AND2_X1 U8238 ( .A1(n6466), .A2(n9823), .ZN(n6467) );
  NAND2_X1 U8239 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  NAND2_X1 U8240 ( .A1(n6471), .A2(n6470), .ZN(n6478) );
  NAND2_X1 U8241 ( .A1(n10159), .A2(n6479), .ZN(n6473) );
  NAND2_X1 U8242 ( .A1(n9941), .A2(n6354), .ZN(n6472) );
  NAND2_X1 U8243 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  XNOR2_X1 U8244 ( .A(n6474), .B(n4514), .ZN(n6477) );
  NAND2_X1 U8245 ( .A1(n10159), .A2(n6354), .ZN(n6476) );
  NAND2_X1 U8246 ( .A1(n9941), .A2(n6327), .ZN(n6475) );
  NAND2_X1 U8247 ( .A1(n6476), .A2(n6475), .ZN(n9883) );
  NAND2_X1 U8248 ( .A1(n10142), .A2(n6479), .ZN(n6481) );
  OR2_X1 U8249 ( .A1(n9886), .A2(n4527), .ZN(n6480) );
  NAND2_X1 U8250 ( .A1(n6481), .A2(n6480), .ZN(n6482) );
  XNOR2_X1 U8251 ( .A(n6482), .B(n4514), .ZN(n6485) );
  NOR2_X1 U8252 ( .A1(n9886), .A2(n6514), .ZN(n6483) );
  AOI21_X1 U8253 ( .B1(n10142), .B2(n6354), .A(n6483), .ZN(n6484) );
  NAND2_X1 U8254 ( .A1(n6485), .A2(n6484), .ZN(n9861) );
  OR2_X1 U8255 ( .A1(n6485), .A2(n6484), .ZN(n6486) );
  AND2_X1 U8256 ( .A1(n9861), .A2(n6486), .ZN(n9804) );
  NAND2_X1 U8257 ( .A1(n10124), .A2(n6479), .ZN(n6488) );
  NAND2_X1 U8258 ( .A1(n9939), .A2(n6354), .ZN(n6487) );
  NAND2_X1 U8259 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  XNOR2_X1 U8260 ( .A(n6489), .B(n4514), .ZN(n6491) );
  NOR2_X1 U8261 ( .A1(n9834), .A2(n6514), .ZN(n6490) );
  AOI21_X1 U8262 ( .B1(n10124), .B2(n6354), .A(n6490), .ZN(n6492) );
  NAND2_X1 U8263 ( .A1(n6491), .A2(n6492), .ZN(n6496) );
  INV_X1 U8264 ( .A(n6491), .ZN(n6494) );
  INV_X1 U8265 ( .A(n6492), .ZN(n6493) );
  NAND2_X1 U8266 ( .A1(n6494), .A2(n6493), .ZN(n6495) );
  NAND2_X1 U8267 ( .A1(n6496), .A2(n6495), .ZN(n9860) );
  INV_X1 U8268 ( .A(n6496), .ZN(n6497) );
  OAI22_X1 U8269 ( .A1(n10304), .A2(n6498), .B1(n6500), .B2(n4527), .ZN(n6499)
         );
  XNOR2_X1 U8270 ( .A(n6499), .B(n6517), .ZN(n6502) );
  OAI22_X1 U8271 ( .A1(n10304), .A2(n4527), .B1(n6500), .B2(n6514), .ZN(n6501)
         );
  XNOR2_X1 U8272 ( .A(n6502), .B(n6501), .ZN(n9833) );
  NOR2_X1 U8273 ( .A1(n6502), .A2(n6501), .ZN(n9905) );
  NAND2_X1 U8274 ( .A1(n10095), .A2(n6479), .ZN(n6504) );
  NAND2_X1 U8275 ( .A1(n9937), .A2(n6354), .ZN(n6503) );
  NAND2_X1 U8276 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  XNOR2_X1 U8277 ( .A(n6505), .B(n4514), .ZN(n6507) );
  NOR2_X1 U8278 ( .A1(n9835), .A2(n6514), .ZN(n6506) );
  AOI21_X1 U8279 ( .B1(n10095), .B2(n6354), .A(n6506), .ZN(n6508) );
  XNOR2_X1 U8280 ( .A(n6507), .B(n6508), .ZN(n9904) );
  INV_X1 U8281 ( .A(n6507), .ZN(n6510) );
  INV_X1 U8282 ( .A(n6508), .ZN(n6509) );
  AOI22_X1 U8283 ( .A1(n10080), .A2(n6479), .B1(n6354), .B2(n9936), .ZN(n6511)
         );
  XNOR2_X1 U8284 ( .A(n6511), .B(n6517), .ZN(n6513) );
  AOI22_X1 U8285 ( .A1(n10080), .A2(n6354), .B1(n6327), .B2(n9936), .ZN(n6512)
         );
  NAND2_X1 U8286 ( .A1(n6513), .A2(n6512), .ZN(n6544) );
  OAI21_X1 U8287 ( .B1(n6513), .B2(n6512), .A(n6544), .ZN(n6560) );
  NAND2_X1 U8288 ( .A1(n6548), .A2(n6354), .ZN(n6516) );
  OR2_X1 U8289 ( .A1(n6565), .A2(n6514), .ZN(n6515) );
  NAND2_X1 U8290 ( .A1(n6516), .A2(n6515), .ZN(n6518) );
  XNOR2_X1 U8291 ( .A(n6518), .B(n6517), .ZN(n6520) );
  AOI22_X1 U8292 ( .A1(n6548), .A2(n6479), .B1(n6354), .B2(n9935), .ZN(n6519)
         );
  XNOR2_X1 U8293 ( .A(n6520), .B(n6519), .ZN(n6527) );
  INV_X1 U8294 ( .A(n6527), .ZN(n6545) );
  INV_X1 U8295 ( .A(n6521), .ZN(n6523) );
  INV_X1 U8296 ( .A(n7409), .ZN(n6525) );
  INV_X1 U8297 ( .A(n8875), .ZN(n10333) );
  NAND2_X1 U8298 ( .A1(n7407), .A2(n10333), .ZN(n6524) );
  AND2_X1 U8299 ( .A1(n10517), .A2(n8807), .ZN(n6526) );
  AND2_X1 U8300 ( .A1(n6527), .A2(n9922), .ZN(n6551) );
  NOR2_X1 U8301 ( .A1(n7436), .A2(n6532), .ZN(n7411) );
  NAND2_X1 U8302 ( .A1(n6531), .A2(n7411), .ZN(n6530) );
  INV_X1 U8303 ( .A(n6528), .ZN(n6529) );
  NAND2_X1 U8304 ( .A1(n7409), .A2(n7407), .ZN(n6534) );
  OR2_X1 U8305 ( .A1(n6532), .A2(P1_U3086), .ZN(n7403) );
  NAND2_X1 U8306 ( .A1(n10282), .A2(n7403), .ZN(n6533) );
  NAND2_X1 U8307 ( .A1(n6534), .A2(n6533), .ZN(n6800) );
  NOR2_X1 U8308 ( .A1(n6536), .A2(n6535), .ZN(n6537) );
  NAND2_X1 U8309 ( .A1(n6800), .A2(n6537), .ZN(n6540) );
  INV_X1 U8310 ( .A(n6635), .ZN(n6538) );
  NAND2_X1 U8311 ( .A1(n6538), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8879) );
  INV_X1 U8312 ( .A(n8879), .ZN(n6539) );
  AOI21_X2 U8313 ( .B1(n6540), .B2(P1_STATE_REG_SCAN_IN), .A(n6539), .ZN(
        n10423) );
  INV_X1 U8314 ( .A(n10423), .ZN(n9927) );
  AOI22_X1 U8315 ( .A1(n10059), .A2(n9927), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6542) );
  OAI21_X1 U8316 ( .B1(n6543), .B2(n10413), .A(n6542), .ZN(n6547) );
  NOR3_X1 U8317 ( .A1(n6545), .A2(n10416), .A3(n6544), .ZN(n6546) );
  AOI211_X1 U8318 ( .C1(n6548), .C2(n10421), .A(n6547), .B(n6546), .ZN(n6549)
         );
  AOI21_X1 U8319 ( .B1(n6563), .B2(n6551), .A(n6550), .ZN(n6552) );
  NAND2_X1 U8320 ( .A1(n6553), .A2(n6552), .ZN(P1_U3220) );
  NOR2_X1 U8321 ( .A1(n10537), .A2(n6554), .ZN(n6556) );
  INV_X1 U8322 ( .A(n6559), .ZN(n6562) );
  INV_X1 U8323 ( .A(n6560), .ZN(n6561) );
  AOI21_X1 U8324 ( .B1(n5064), .B2(n6562), .A(n6561), .ZN(n6564) );
  OAI21_X1 U8325 ( .B1(n6564), .B2(n6563), .A(n9922), .ZN(n6574) );
  OR2_X1 U8326 ( .A1(n6565), .A2(n9908), .ZN(n6567) );
  NAND2_X1 U8327 ( .A1(n9937), .A2(n9910), .ZN(n6566) );
  NAND2_X1 U8328 ( .A1(n6567), .A2(n6566), .ZN(n10071) );
  INV_X1 U8329 ( .A(n10081), .ZN(n6569) );
  OAI22_X1 U8330 ( .A1(n6569), .A2(n10423), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6568), .ZN(n6570) );
  AOI21_X1 U8331 ( .B1(n10071), .B2(n9916), .A(n6570), .ZN(n6571) );
  INV_X1 U8332 ( .A(n6572), .ZN(n6573) );
  NAND2_X1 U8333 ( .A1(n6574), .A2(n6573), .ZN(P1_U3214) );
  INV_X1 U8334 ( .A(n6575), .ZN(n6576) );
  NOR2_X1 U8335 ( .A1(n8453), .A2(n6576), .ZN(n6948) );
  NOR2_X1 U8336 ( .A1(n6577), .A2(n6948), .ZN(n6578) );
  NAND2_X1 U8337 ( .A1(n6579), .A2(n8516), .ZN(n6580) );
  AND2_X1 U8338 ( .A1(n6580), .A2(n8453), .ZN(n6581) );
  NAND2_X1 U8339 ( .A1(n6640), .A2(n6581), .ZN(n6838) );
  NOR2_X1 U8340 ( .A1(n9737), .A2(n8513), .ZN(n6841) );
  INV_X1 U8341 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8342 ( .A1(n6583), .A2(n6582), .ZN(n6836) );
  OAI21_X1 U8343 ( .B1(n6838), .B2(n6841), .A(n6836), .ZN(n6585) );
  NAND2_X1 U8344 ( .A1(n6586), .A2(n9744), .ZN(n6591) );
  NAND2_X1 U8345 ( .A1(n9743), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6587) );
  INV_X1 U8346 ( .A(n6589), .ZN(n6590) );
  NAND2_X1 U8347 ( .A1(n6591), .A2(n6590), .ZN(P2_U3488) );
  INV_X1 U8348 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6592) );
  OAI21_X1 U8349 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(P1_U3519) );
  INV_X1 U8350 ( .A(n6598), .ZN(n6599) );
  INV_X1 U8351 ( .A(n7020), .ZN(n6600) );
  NAND2_X1 U8352 ( .A1(n7057), .A2(n8453), .ZN(n6601) );
  NAND2_X1 U8353 ( .A1(n6601), .A2(n7055), .ZN(n7067) );
  NAND2_X1 U8354 ( .A1(n7067), .A2(n6602), .ZN(n6603) );
  NAND2_X1 U8355 ( .A1(n6603), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U8356 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8357 ( .A(n6740), .B(n6604), .S(P1_U3086), .Z(n6605) );
  INV_X1 U8358 ( .A(n6605), .ZN(P1_U3355) );
  NAND2_X1 U8359 ( .A1(n4518), .A2(P1_U3086), .ZN(n8891) );
  NOR2_X1 U8360 ( .A1(n4518), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10343) );
  INV_X2 U8361 ( .A(n10343), .ZN(n8546) );
  OAI222_X1 U8362 ( .A1(n8891), .A2(n4826), .B1(n8546), .B2(n6622), .C1(
        P1_U3086), .C2(n9969), .ZN(P1_U3354) );
  INV_X1 U8363 ( .A(n8891), .ZN(n6618) );
  INV_X1 U8364 ( .A(n6618), .ZN(n10338) );
  OAI222_X1 U8365 ( .A1(n10338), .A2(n9232), .B1(n8546), .B2(n6610), .C1(
        P1_U3086), .C2(n6788), .ZN(P1_U3351) );
  OAI222_X1 U8366 ( .A1(n10338), .A2(n6606), .B1(n8546), .B2(n6612), .C1(
        P1_U3086), .C2(n9996), .ZN(P1_U3352) );
  INV_X1 U8367 ( .A(n9983), .ZN(n6607) );
  OAI222_X1 U8368 ( .A1(n10338), .A2(n6608), .B1(n8546), .B2(n6613), .C1(
        P1_U3086), .C2(n6607), .ZN(P1_U3353) );
  INV_X1 U8369 ( .A(n7165), .ZN(n7304) );
  NAND2_X1 U8370 ( .A1(n4518), .A2(P2_U3151), .ZN(n9801) );
  NOR2_X1 U8371 ( .A1(n4518), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9795) );
  INV_X2 U8372 ( .A(n9795), .ZN(n9798) );
  OAI222_X1 U8373 ( .A1(n7304), .A2(P2_U3151), .B1(n9801), .B2(n6610), .C1(
        n6609), .C2(n9798), .ZN(P2_U3291) );
  INV_X1 U8374 ( .A(n7051), .ZN(n7145) );
  OAI222_X1 U8375 ( .A1(n7145), .A2(P2_U3151), .B1(n9801), .B2(n6612), .C1(
        n6611), .C2(n9798), .ZN(P2_U3292) );
  INV_X1 U8376 ( .A(n10570), .ZN(n7071) );
  OAI222_X1 U8377 ( .A1(n9798), .A2(n6614), .B1(n9801), .B2(n6613), .C1(n7071), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  INV_X1 U8378 ( .A(n6674), .ZN(n10006) );
  OAI222_X1 U8379 ( .A1(n10338), .A2(n6615), .B1(n8546), .B2(n6616), .C1(
        P1_U3086), .C2(n10006), .ZN(P1_U3350) );
  OAI222_X1 U8380 ( .A1(n7279), .A2(P2_U3151), .B1(n9801), .B2(n6616), .C1(
        n9234), .C2(n9798), .ZN(P2_U3290) );
  INV_X1 U8381 ( .A(n6617), .ZN(n6620) );
  AOI22_X1 U8382 ( .A1(n10028), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n6618), .ZN(n6619) );
  OAI21_X1 U8383 ( .B1(n6620), .B2(n8546), .A(n6619), .ZN(P1_U3349) );
  INV_X1 U8384 ( .A(n7172), .ZN(n7537) );
  INV_X1 U8385 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9214) );
  OAI222_X1 U8386 ( .A1(n7537), .A2(P2_U3151), .B1(n9801), .B2(n6620), .C1(
        n9214), .C2(n9798), .ZN(P2_U3289) );
  INV_X1 U8387 ( .A(n9801), .ZN(n7775) );
  INV_X1 U8388 ( .A(n7775), .ZN(n8274) );
  INV_X1 U8389 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6621) );
  OAI222_X1 U8390 ( .A1(P2_U3151), .A2(n4751), .B1(n8274), .B2(n6622), .C1(
        n6621), .C2(n9798), .ZN(P2_U3294) );
  INV_X1 U8391 ( .A(n6623), .ZN(n6625) );
  AOI22_X1 U8392 ( .A1(n10585), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9795), .ZN(n6624) );
  OAI21_X1 U8393 ( .B1(n6625), .B2(n9801), .A(n6624), .ZN(P2_U3288) );
  INV_X1 U8394 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6626) );
  INV_X1 U8395 ( .A(n6667), .ZN(n6699) );
  OAI222_X1 U8396 ( .A1(n10338), .A2(n6626), .B1(n8546), .B2(n6625), .C1(
        P1_U3086), .C2(n6699), .ZN(P1_U3348) );
  INV_X1 U8397 ( .A(n6627), .ZN(n6629) );
  INV_X1 U8398 ( .A(n6709), .ZN(n6686) );
  OAI222_X1 U8399 ( .A1(n10338), .A2(n6628), .B1(n8546), .B2(n6629), .C1(
        P1_U3086), .C2(n6686), .ZN(P1_U3347) );
  INV_X1 U8400 ( .A(n7751), .ZN(n7741) );
  OAI222_X1 U8401 ( .A1(n7741), .A2(P2_U3151), .B1(n9801), .B2(n6629), .C1(
        n9206), .C2(n9798), .ZN(P2_U3287) );
  INV_X1 U8402 ( .A(n6630), .ZN(n6633) );
  INV_X1 U8403 ( .A(n6721), .ZN(n6707) );
  OAI222_X1 U8404 ( .A1(n8546), .A2(n6633), .B1(n6707), .B2(P1_U3086), .C1(
        n6631), .C2(n10338), .ZN(P1_U3346) );
  INV_X1 U8405 ( .A(n7985), .ZN(n7977) );
  OAI222_X1 U8406 ( .A1(P2_U3151), .A2(n7977), .B1(n8274), .B2(n6633), .C1(
        n6632), .C2(n9798), .ZN(P2_U3286) );
  NAND2_X1 U8407 ( .A1(n8875), .A2(n8879), .ZN(n6662) );
  INV_X1 U8408 ( .A(n6662), .ZN(n6637) );
  AOI21_X1 U8409 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6661) );
  NOR2_X2 U8410 ( .A1(n6637), .A2(n6661), .ZN(n10021) );
  NOR2_X1 U8411 ( .A1(n10021), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8412 ( .A(n6638), .ZN(n6643) );
  INV_X1 U8413 ( .A(n6764), .ZN(n6771) );
  OAI222_X1 U8414 ( .A1(n8546), .A2(n6643), .B1(n6771), .B2(P1_U3086), .C1(
        n6639), .C2(n10338), .ZN(P1_U3345) );
  INV_X1 U8415 ( .A(n6640), .ZN(n6641) );
  NAND2_X1 U8416 ( .A1(n6641), .A2(n6952), .ZN(n6642) );
  OAI21_X1 U8417 ( .B1(n6952), .B2(n5716), .A(n6642), .ZN(P2_U3377) );
  OAI222_X1 U8418 ( .A1(P2_U3151), .A2(n7988), .B1(n8274), .B2(n6643), .C1(
        n8970), .C2(n9798), .ZN(P2_U3285) );
  NAND2_X1 U8419 ( .A1(n9500), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n6644) );
  OAI21_X1 U8420 ( .B1(n9500), .B2(n8563), .A(n6644), .ZN(P2_U3507) );
  NAND2_X1 U8421 ( .A1(n6952), .A2(n6645), .ZN(n6750) );
  INV_X1 U8422 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6647) );
  INV_X1 U8423 ( .A(n6975), .ZN(n6646) );
  AOI22_X1 U8424 ( .A1(n6750), .A2(n6647), .B1(n7020), .B2(n6646), .ZN(
        P2_U3376) );
  INV_X1 U8425 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6648) );
  XNOR2_X1 U8426 ( .A(n9983), .B(n6648), .ZN(n9986) );
  XNOR2_X1 U8427 ( .A(n9969), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U8428 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6781) );
  INV_X1 U8429 ( .A(n6781), .ZN(n9975) );
  NAND2_X1 U8430 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  INV_X1 U8431 ( .A(n9969), .ZN(n9968) );
  NAND2_X1 U8432 ( .A1(n9968), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8433 ( .A1(n9974), .A2(n6649), .ZN(n9985) );
  NAND2_X1 U8434 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U8435 ( .A1(n9983), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U8436 ( .A1(n9984), .A2(n6650), .ZN(n9994) );
  XNOR2_X1 U8437 ( .A(n9996), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U8438 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  INV_X1 U8439 ( .A(n9996), .ZN(n6651) );
  NAND2_X1 U8440 ( .A1(n6651), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8441 ( .A1(n9993), .A2(n6652), .ZN(n6786) );
  XNOR2_X1 U8442 ( .A(n6788), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8443 ( .A1(n6786), .A2(n6785), .ZN(n6654) );
  INV_X1 U8444 ( .A(n6788), .ZN(n6796) );
  NAND2_X1 U8445 ( .A1(n6796), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8446 ( .A1(n6654), .A2(n6653), .ZN(n10011) );
  INV_X1 U8447 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6655) );
  MUX2_X1 U8448 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6655), .S(n6674), .Z(n10012)
         );
  NAND2_X1 U8449 ( .A1(n10011), .A2(n10012), .ZN(n10010) );
  NAND2_X1 U8450 ( .A1(n6674), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8451 ( .A1(n10010), .A2(n6656), .ZN(n10026) );
  OR2_X1 U8452 ( .A1(n10028), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U8453 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n10028), .ZN(n6657) );
  AND2_X1 U8454 ( .A1(n6658), .A2(n6657), .ZN(n10027) );
  AND2_X1 U8455 ( .A1(n10026), .A2(n10027), .ZN(n10023) );
  AOI21_X1 U8456 ( .B1(n10028), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10023), .ZN(
        n6691) );
  INV_X1 U8457 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U8458 ( .A1(n6667), .A2(n6659), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6699), .ZN(n6690) );
  NOR2_X1 U8459 ( .A1(n6691), .A2(n6690), .ZN(n6689) );
  AOI21_X1 U8460 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6667), .A(n6689), .ZN(
        n6664) );
  NAND2_X1 U8461 ( .A1(n6709), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U8462 ( .B1(n6709), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6660), .ZN(
        n6663) );
  NOR2_X1 U8463 ( .A1(n6664), .A2(n6663), .ZN(n6708) );
  NAND2_X1 U8464 ( .A1(n6662), .A2(n6661), .ZN(n6739) );
  INV_X1 U8465 ( .A(n8142), .ZN(n6780) );
  NAND2_X1 U8466 ( .A1(n6665), .A2(n6780), .ZN(n8874) );
  AOI211_X1 U8467 ( .C1(n6664), .C2(n6663), .A(n6708), .B(n7948), .ZN(n6688)
         );
  AND2_X1 U8468 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6666) );
  AOI21_X1 U8469 ( .B1(n10021), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6666), .ZN(
        n6685) );
  INV_X1 U8470 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6679) );
  MUX2_X1 U8471 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6679), .S(n6667), .Z(n6693)
         );
  XOR2_X1 U8472 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9983), .Z(n9980) );
  INV_X1 U8473 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10524) );
  NAND2_X1 U8474 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9970) );
  AOI21_X1 U8475 ( .B1(n9969), .B2(n10524), .A(n9970), .ZN(n6668) );
  OR2_X1 U8476 ( .A1(n9969), .A2(n10524), .ZN(n6669) );
  NAND2_X1 U8477 ( .A1(n6668), .A2(n6669), .ZN(n9973) );
  NAND2_X1 U8478 ( .A1(n9973), .A2(n6669), .ZN(n9981) );
  AOI22_X1 U8479 ( .A1(n9980), .A2(n9981), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n9983), .ZN(n9997) );
  INV_X1 U8480 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6670) );
  MUX2_X1 U8481 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6670), .S(n9996), .Z(n6671)
         );
  NOR2_X1 U8482 ( .A1(n9997), .A2(n6671), .ZN(n9998) );
  NOR2_X1 U8483 ( .A1(n9996), .A2(n6670), .ZN(n6787) );
  INV_X1 U8484 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8485 ( .A(n6672), .B(P1_REG1_REG_4__SCAN_IN), .S(n6788), .Z(n6673)
         );
  OAI21_X1 U8486 ( .B1(n9998), .B2(n6787), .A(n6673), .ZN(n10015) );
  NAND2_X1 U8487 ( .A1(n6796), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10014) );
  INV_X1 U8488 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6675) );
  MUX2_X1 U8489 ( .A(n6675), .B(P1_REG1_REG_5__SCAN_IN), .S(n6674), .Z(n10013)
         );
  AOI21_X1 U8490 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10035) );
  NOR2_X1 U8491 ( .A1(n10006), .A2(n6675), .ZN(n10029) );
  INV_X1 U8492 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U8493 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6676), .S(n10028), .Z(n6677)
         );
  OAI21_X1 U8494 ( .B1(n10035), .B2(n10029), .A(n6677), .ZN(n10032) );
  NAND2_X1 U8495 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n10028), .ZN(n6678) );
  NAND2_X1 U8496 ( .A1(n10032), .A2(n6678), .ZN(n6694) );
  NAND2_X1 U8497 ( .A1(n6693), .A2(n6694), .ZN(n6692) );
  OAI21_X1 U8498 ( .B1(n6699), .B2(n6679), .A(n6692), .ZN(n6683) );
  INV_X1 U8499 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U8500 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6680), .S(n6709), .Z(n6682)
         );
  INV_X1 U8501 ( .A(n6739), .ZN(n6681) );
  NAND2_X1 U8502 ( .A1(n6682), .A2(n6683), .ZN(n6702) );
  OAI211_X1 U8503 ( .C1(n6683), .C2(n6682), .A(n10033), .B(n6702), .ZN(n6684)
         );
  OAI211_X1 U8504 ( .C1(n10007), .C2(n6686), .A(n6685), .B(n6684), .ZN(n6687)
         );
  OR2_X1 U8505 ( .A1(n6688), .A2(n6687), .ZN(P1_U3251) );
  AOI211_X1 U8506 ( .C1(n6691), .C2(n6690), .A(n6689), .B(n7948), .ZN(n6701)
         );
  OAI211_X1 U8507 ( .C1(n6694), .C2(n6693), .A(n6692), .B(n10033), .ZN(n6698)
         );
  NOR2_X1 U8508 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6695), .ZN(n6696) );
  AOI21_X1 U8509 ( .B1(n10021), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6696), .ZN(
        n6697) );
  OAI211_X1 U8510 ( .C1(n10007), .C2(n6699), .A(n6698), .B(n6697), .ZN(n6700)
         );
  OR2_X1 U8511 ( .A1(n6701), .A2(n6700), .ZN(P1_U3250) );
  INV_X1 U8512 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U8513 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6707), .B1(n6721), .B2(
        n10527), .ZN(n6705) );
  NAND2_X1 U8514 ( .A1(n6709), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6703) );
  NAND2_X1 U8515 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  NOR2_X1 U8516 ( .A1(n6705), .A2(n6704), .ZN(n6723) );
  AOI21_X1 U8517 ( .B1(n6705), .B2(n6704), .A(n6723), .ZN(n6717) );
  INV_X1 U8518 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U8519 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6721), .B1(n6707), .B2(
        n6706), .ZN(n6711) );
  AOI21_X1 U8520 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6709), .A(n6708), .ZN(
        n6710) );
  NAND2_X1 U8521 ( .A1(n6711), .A2(n6710), .ZN(n6718) );
  OAI21_X1 U8522 ( .B1(n6711), .B2(n6710), .A(n6718), .ZN(n6712) );
  NAND2_X1 U8523 ( .A1(n6712), .A2(n10025), .ZN(n6716) );
  INV_X1 U8524 ( .A(n10007), .ZN(n10022) );
  INV_X1 U8525 ( .A(n10021), .ZN(n9966) );
  INV_X1 U8526 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8527 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7794) );
  OAI21_X1 U8528 ( .B1(n9966), .B2(n6713), .A(n7794), .ZN(n6714) );
  AOI21_X1 U8529 ( .B1(n6721), .B2(n10022), .A(n6714), .ZN(n6715) );
  OAI211_X1 U8530 ( .C1(n6717), .C2(n8109), .A(n6716), .B(n6715), .ZN(P1_U3252) );
  INV_X1 U8531 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8951) );
  AOI22_X1 U8532 ( .A1(n6764), .A2(n8951), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6771), .ZN(n6720) );
  OAI21_X1 U8533 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6721), .A(n6718), .ZN(
        n6719) );
  NOR2_X1 U8534 ( .A1(n6720), .A2(n6719), .ZN(n6763) );
  AOI211_X1 U8535 ( .C1(n6720), .C2(n6719), .A(n6763), .B(n7948), .ZN(n6731)
         );
  NOR2_X1 U8536 ( .A1(n6721), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6722) );
  NOR2_X1 U8537 ( .A1(n6723), .A2(n6722), .ZN(n6726) );
  INV_X1 U8538 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6724) );
  MUX2_X1 U8539 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6724), .S(n6764), .Z(n6725)
         );
  NAND2_X1 U8540 ( .A1(n6725), .A2(n6726), .ZN(n6770) );
  OAI211_X1 U8541 ( .C1(n6726), .C2(n6725), .A(n6770), .B(n10033), .ZN(n6729)
         );
  AND2_X1 U8542 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6727) );
  AOI21_X1 U8543 ( .B1(n10021), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6727), .ZN(
        n6728) );
  OAI211_X1 U8544 ( .C1(n10007), .C2(n6771), .A(n6729), .B(n6728), .ZN(n6730)
         );
  OR2_X1 U8545 ( .A1(n6731), .A2(n6730), .ZN(P1_U3253) );
  INV_X1 U8546 ( .A(n6732), .ZN(n6734) );
  AOI22_X1 U8547 ( .A1(n8177), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9795), .ZN(n6733) );
  OAI21_X1 U8548 ( .B1(n6734), .B2(n9801), .A(n6733), .ZN(P2_U3284) );
  INV_X1 U8549 ( .A(n6817), .ZN(n6812) );
  OAI222_X1 U8550 ( .A1(n10338), .A2(n6735), .B1(n8546), .B2(n6734), .C1(
        P1_U3086), .C2(n6812), .ZN(P1_U3344) );
  INV_X1 U8551 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6736) );
  AOI21_X1 U8552 ( .B1(n6780), .B2(n6736), .A(n8893), .ZN(n6782) );
  OAI21_X1 U8553 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n6780), .A(n6782), .ZN(
        n6737) );
  MUX2_X1 U8554 ( .A(n6782), .B(n6737), .S(n6740), .Z(n6738) );
  INV_X1 U8555 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7440) );
  OAI22_X1 U8556 ( .A1(n6739), .A2(n6738), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7440), .ZN(n6742) );
  NOR3_X1 U8557 ( .A1(n8109), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6740), .ZN(
        n6741) );
  AOI211_X1 U8558 ( .C1(n10021), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n6742), .B(
        n6741), .ZN(n6743) );
  INV_X1 U8559 ( .A(n6743), .ZN(P1_U3243) );
  INV_X1 U8560 ( .A(n6744), .ZN(n6762) );
  INV_X1 U8561 ( .A(n7192), .ZN(n6822) );
  OAI222_X1 U8562 ( .A1(n8546), .A2(n6762), .B1(n6822), .B2(P1_U3086), .C1(
        n6745), .C2(n10338), .ZN(P1_U3343) );
  INV_X1 U8563 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6749) );
  INV_X1 U8564 ( .A(n7486), .ZN(n6746) );
  NAND2_X1 U8565 ( .A1(n9964), .A2(n7492), .ZN(n8821) );
  AND2_X1 U8566 ( .A1(n6746), .A2(n8821), .ZN(n8743) );
  INV_X1 U8567 ( .A(n8743), .ZN(n7437) );
  OAI21_X1 U8568 ( .B1(n10520), .B2(n10427), .A(n7437), .ZN(n6747) );
  NAND2_X1 U8569 ( .A1(n9963), .A2(n9865), .ZN(n7438) );
  OAI211_X1 U8570 ( .C1(n7436), .C2(n7492), .A(n6747), .B(n7438), .ZN(n10286)
         );
  NAND2_X1 U8571 ( .A1(n10286), .A2(n10523), .ZN(n6748) );
  OAI21_X1 U8572 ( .B1(n10523), .B2(n6749), .A(n6748), .ZN(P1_U3453) );
  INV_X1 U8573 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U8574 ( .A1(n6915), .A2(n6751), .ZN(P2_U3248) );
  INV_X1 U8575 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6752) );
  NOR2_X1 U8576 ( .A1(n6915), .A2(n6752), .ZN(P2_U3250) );
  INV_X1 U8577 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6753) );
  NOR2_X1 U8578 ( .A1(n6915), .A2(n6753), .ZN(P2_U3254) );
  INV_X1 U8579 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n8971) );
  NOR2_X1 U8580 ( .A1(n6915), .A2(n8971), .ZN(P2_U3252) );
  INV_X1 U8581 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6754) );
  NOR2_X1 U8582 ( .A1(n6915), .A2(n6754), .ZN(P2_U3255) );
  INV_X1 U8583 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9204) );
  NOR2_X1 U8584 ( .A1(n6915), .A2(n9204), .ZN(P2_U3253) );
  INV_X1 U8585 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6755) );
  NOR2_X1 U8586 ( .A1(n6915), .A2(n6755), .ZN(P2_U3249) );
  INV_X1 U8587 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6756) );
  NOR2_X1 U8588 ( .A1(n6915), .A2(n6756), .ZN(P2_U3247) );
  INV_X1 U8589 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6757) );
  NOR2_X1 U8590 ( .A1(n6915), .A2(n6757), .ZN(P2_U3257) );
  INV_X1 U8591 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6758) );
  NOR2_X1 U8592 ( .A1(n6915), .A2(n6758), .ZN(P2_U3246) );
  INV_X1 U8593 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6759) );
  NOR2_X1 U8594 ( .A1(n6915), .A2(n6759), .ZN(P2_U3256) );
  INV_X1 U8595 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U8596 ( .A1(n6915), .A2(n6760), .ZN(P2_U3251) );
  INV_X1 U8597 ( .A(n8174), .ZN(n9405) );
  OAI222_X1 U8598 ( .A1(P2_U3151), .A2(n9405), .B1(n8274), .B2(n6762), .C1(
        n6761), .C2(n9798), .ZN(P2_U3283) );
  AOI21_X1 U8599 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6764), .A(n6763), .ZN(
        n6767) );
  NAND2_X1 U8600 ( .A1(n6817), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6765) );
  OAI21_X1 U8601 ( .B1(n6817), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6765), .ZN(
        n6766) );
  NOR2_X1 U8602 ( .A1(n6767), .A2(n6766), .ZN(n6816) );
  AOI211_X1 U8603 ( .C1(n6767), .C2(n6766), .A(n6816), .B(n7948), .ZN(n6777)
         );
  NOR2_X1 U8604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6768), .ZN(n6769) );
  AOI21_X1 U8605 ( .B1(n10021), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6769), .ZN(
        n6775) );
  OAI21_X1 U8606 ( .B1(n6771), .B2(n6724), .A(n6770), .ZN(n6773) );
  MUX2_X1 U8607 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10530), .S(n6817), .Z(n6772) );
  NAND2_X1 U8608 ( .A1(n6772), .A2(n6773), .ZN(n6811) );
  OAI211_X1 U8609 ( .C1(n6773), .C2(n6772), .A(n10033), .B(n6811), .ZN(n6774)
         );
  OAI211_X1 U8610 ( .C1(n10007), .C2(n6812), .A(n6775), .B(n6774), .ZN(n6776)
         );
  OR2_X1 U8611 ( .A1(n6777), .A2(n6776), .ZN(P1_U3254) );
  XOR2_X1 U8612 ( .A(n6779), .B(n6778), .Z(n6798) );
  NOR3_X1 U8613 ( .A1(n6798), .A2(n6780), .A3(n8893), .ZN(n6784) );
  OAI22_X1 U8614 ( .A1(n6782), .A2(P1_IR_REG_0__SCAN_IN), .B1(n6781), .B2(
        n8874), .ZN(n6783) );
  OR3_X1 U8615 ( .A1(n6784), .A2(n9942), .A3(n6783), .ZN(n9990) );
  XNOR2_X1 U8616 ( .A(n6786), .B(n6785), .ZN(n6793) );
  INV_X1 U8617 ( .A(n6787), .ZN(n6790) );
  MUX2_X1 U8618 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6672), .S(n6788), .Z(n6789)
         );
  NAND2_X1 U8619 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  OAI211_X1 U8620 ( .C1(n9998), .C2(n6791), .A(n10033), .B(n10015), .ZN(n6792)
         );
  OAI21_X1 U8621 ( .B1(n6793), .B2(n7948), .A(n6792), .ZN(n6795) );
  INV_X1 U8622 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U8623 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7225) );
  OAI21_X1 U8624 ( .B1(n9966), .B2(n10357), .A(n7225), .ZN(n6794) );
  AOI211_X1 U8625 ( .C1(n6796), .C2(n10022), .A(n6795), .B(n6794), .ZN(n6797)
         );
  NAND2_X1 U8626 ( .A1(n9990), .A2(n6797), .ZN(P1_U3247) );
  AOI22_X1 U8627 ( .A1(n10421), .A2(n7435), .B1(n9922), .B2(n6798), .ZN(n6802)
         );
  INV_X1 U8628 ( .A(n7406), .ZN(n6799) );
  NAND2_X1 U8629 ( .A1(n6800), .A2(n6799), .ZN(n6833) );
  NAND2_X1 U8630 ( .A1(n6833), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6801) );
  OAI211_X1 U8631 ( .C1(n10413), .C2(n7438), .A(n6802), .B(n6801), .ZN(
        P1_U3232) );
  INV_X1 U8632 ( .A(n6804), .ZN(n6829) );
  AOI21_X1 U8633 ( .B1(n6805), .B2(n6803), .A(n6829), .ZN(n6810) );
  NAND2_X1 U8634 ( .A1(n9964), .A2(n9910), .ZN(n6807) );
  NAND2_X1 U8635 ( .A1(n9962), .A2(n9865), .ZN(n6806) );
  NAND2_X1 U8636 ( .A1(n6807), .A2(n6806), .ZN(n7487) );
  AOI22_X1 U8637 ( .A1(n9916), .A2(n7487), .B1(n6833), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U8638 ( .A1(n10421), .A2(n8822), .ZN(n6808) );
  OAI211_X1 U8639 ( .C1(n6810), .C2(n10416), .A(n6809), .B(n6808), .ZN(
        P1_U3222) );
  INV_X1 U8640 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10530) );
  OAI21_X1 U8641 ( .B1(n10530), .B2(n6812), .A(n6811), .ZN(n6814) );
  INV_X1 U8642 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U8643 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6822), .B1(n7192), .B2(
        n10532), .ZN(n6813) );
  NOR2_X1 U8644 ( .A1(n6814), .A2(n6813), .ZN(n7187) );
  AOI21_X1 U8645 ( .B1(n6814), .B2(n6813), .A(n7187), .ZN(n6826) );
  NOR2_X1 U8646 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7192), .ZN(n6815) );
  AOI21_X1 U8647 ( .B1(n7192), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6815), .ZN(
        n6819) );
  AOI21_X1 U8648 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6817), .A(n6816), .ZN(
        n6818) );
  NAND2_X1 U8649 ( .A1(n6819), .A2(n6818), .ZN(n7191) );
  OAI21_X1 U8650 ( .B1(n6819), .B2(n6818), .A(n7191), .ZN(n6820) );
  NAND2_X1 U8651 ( .A1(n6820), .A2(n10025), .ZN(n6825) );
  NOR2_X1 U8652 ( .A1(n6821), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7763) );
  NOR2_X1 U8653 ( .A1(n10007), .A2(n6822), .ZN(n6823) );
  AOI211_X1 U8654 ( .C1(n10021), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7763), .B(
        n6823), .ZN(n6824) );
  OAI211_X1 U8655 ( .C1(n6826), .C2(n8109), .A(n6825), .B(n6824), .ZN(P1_U3255) );
  NOR3_X1 U8656 ( .A1(n6829), .A2(n6828), .A3(n6827), .ZN(n6832) );
  INV_X1 U8657 ( .A(n6830), .ZN(n6831) );
  OAI21_X1 U8658 ( .B1(n6832), .B2(n6831), .A(n9922), .ZN(n6835) );
  OAI22_X1 U8659 ( .A1(n8823), .A2(n9887), .B1(n6932), .B2(n9908), .ZN(n6853)
         );
  AOI22_X1 U8660 ( .A1(n9916), .A2(n6853), .B1(n6833), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6834) );
  OAI211_X1 U8661 ( .C1(n7417), .C2(n9931), .A(n6835), .B(n6834), .ZN(P1_U3237) );
  INV_X1 U8662 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6847) );
  AND2_X1 U8663 ( .A1(n6837), .A2(n6836), .ZN(n6839) );
  NAND3_X1 U8664 ( .A1(n6840), .A2(n6839), .A3(n6838), .ZN(n6844) );
  AND2_X1 U8665 ( .A1(n5679), .A2(n7044), .ZN(n8282) );
  NOR2_X1 U8666 ( .A1(n4638), .A2(n8282), .ZN(n8480) );
  INV_X1 U8667 ( .A(n6842), .ZN(n6959) );
  NOR3_X1 U8668 ( .A1(n8480), .A2(n6959), .A3(n9739), .ZN(n6843) );
  NOR2_X1 U8669 ( .A1(n7099), .A2(n9646), .ZN(n6910) );
  OAI21_X1 U8670 ( .B1(n6843), .B2(n6910), .A(n10629), .ZN(n6846) );
  NOR2_X2 U8671 ( .A1(n6844), .A2(n10622), .ZN(n9651) );
  AOI22_X1 U8672 ( .A1(n9651), .A2(n6976), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10628), .ZN(n6845) );
  OAI211_X1 U8673 ( .C1(n6847), .C2(n10629), .A(n6846), .B(n6845), .ZN(
        P2_U3233) );
  OAI21_X1 U8674 ( .B1(n6849), .B2(n6852), .A(n6848), .ZN(n7419) );
  NAND2_X1 U8675 ( .A1(n7491), .A2(n5879), .ZN(n6850) );
  NAND2_X1 U8676 ( .A1(n6850), .A2(n10435), .ZN(n6851) );
  NOR2_X1 U8677 ( .A1(n6901), .A2(n6851), .ZN(n7414) );
  XNOR2_X1 U8678 ( .A(n8624), .B(n6852), .ZN(n6855) );
  INV_X1 U8679 ( .A(n6853), .ZN(n6854) );
  OAI21_X1 U8680 ( .B1(n6855), .B2(n10203), .A(n6854), .ZN(n7410) );
  AOI211_X1 U8681 ( .C1(n10520), .C2(n7419), .A(n7414), .B(n7410), .ZN(n6883)
         );
  AOI22_X1 U8682 ( .A1(n8889), .A2(n5879), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n10534), .ZN(n6856) );
  OAI21_X1 U8683 ( .B1(n6883), .B2(n10534), .A(n6856), .ZN(P1_U3524) );
  INV_X1 U8684 ( .A(n6857), .ZN(n6859) );
  INV_X1 U8685 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6858) );
  OAI222_X1 U8686 ( .A1(n9410), .A2(P2_U3151), .B1(n8274), .B2(n6859), .C1(
        n6858), .C2(n9798), .ZN(P2_U3282) );
  INV_X1 U8687 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6860) );
  INV_X1 U8688 ( .A(n7234), .ZN(n7199) );
  OAI222_X1 U8689 ( .A1(n10338), .A2(n6860), .B1(n8546), .B2(n6859), .C1(
        P1_U3086), .C2(n7199), .ZN(P1_U3342) );
  INV_X1 U8690 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10553) );
  XNOR2_X1 U8691 ( .A(n6861), .B(n8289), .ZN(n7200) );
  NOR2_X1 U8692 ( .A1(n6862), .A2(n9716), .ZN(n6868) );
  NAND2_X1 U8693 ( .A1(n6976), .A2(n9730), .ZN(n6864) );
  OAI21_X1 U8694 ( .B1(n6861), .B2(n6864), .A(n9644), .ZN(n6865) );
  NAND2_X1 U8695 ( .A1(n6865), .A2(n5679), .ZN(n6867) );
  NAND2_X1 U8696 ( .A1(n9387), .A2(n6257), .ZN(n6866) );
  OAI211_X1 U8697 ( .C1(n6863), .C2(n9642), .A(n6867), .B(n6866), .ZN(n7201)
         );
  AOI211_X1 U8698 ( .C1(n9711), .C2(n7200), .A(n6868), .B(n7201), .ZN(n10633)
         );
  OR2_X1 U8699 ( .A1(n10633), .A2(n9743), .ZN(n6869) );
  OAI21_X1 U8700 ( .B1(n9744), .B2(n10553), .A(n6869), .ZN(P2_U3460) );
  OAI21_X1 U8701 ( .B1(n6872), .B2(n6871), .A(n6870), .ZN(n6878) );
  OR2_X1 U8702 ( .A1(n7134), .A2(n9908), .ZN(n6874) );
  NAND2_X1 U8703 ( .A1(n9962), .A2(n9910), .ZN(n6873) );
  NAND2_X1 U8704 ( .A1(n6874), .A2(n6873), .ZN(n6903) );
  AOI22_X1 U8705 ( .A1(n9916), .A2(n6903), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n6875) );
  OAI21_X1 U8706 ( .B1(n7427), .B2(n9931), .A(n6875), .ZN(n6877) );
  NOR2_X1 U8707 ( .A1(n10423), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6876) );
  AOI211_X1 U8708 ( .C1(n9922), .C2(n6878), .A(n6877), .B(n6876), .ZN(n6879)
         );
  INV_X1 U8709 ( .A(n6879), .ZN(P1_U3218) );
  INV_X1 U8710 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6880) );
  OAI22_X1 U8711 ( .A1(n10329), .A2(n7417), .B1(n10523), .B2(n6880), .ZN(n6881) );
  INV_X1 U8712 ( .A(n6881), .ZN(n6882) );
  OAI21_X1 U8713 ( .B1(n6883), .B2(n6596), .A(n6882), .ZN(P1_U3459) );
  INV_X1 U8714 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9076) );
  NAND3_X1 U8715 ( .A1(n6885), .A2(n8292), .A3(n6887), .ZN(n6886) );
  NAND2_X1 U8716 ( .A1(n6884), .A2(n6886), .ZN(n7112) );
  NOR2_X1 U8717 ( .A1(n7108), .A2(n9716), .ZN(n6895) );
  NAND2_X1 U8718 ( .A1(n6888), .A2(n6887), .ZN(n7013) );
  NAND3_X1 U8719 ( .A1(n6889), .A2(n8478), .A3(n6890), .ZN(n6891) );
  NAND2_X1 U8720 ( .A1(n7013), .A2(n6891), .ZN(n6892) );
  NAND2_X1 U8721 ( .A1(n6892), .A2(n9730), .ZN(n6894) );
  INV_X1 U8722 ( .A(n9644), .ZN(n9724) );
  AOI22_X1 U8723 ( .A1(n9724), .A2(n9387), .B1(n5305), .B2(n6257), .ZN(n6893)
         );
  NAND2_X1 U8724 ( .A1(n6894), .A2(n6893), .ZN(n7109) );
  AOI211_X1 U8725 ( .C1(n9711), .C2(n7112), .A(n6895), .B(n7109), .ZN(n10637)
         );
  OR2_X1 U8726 ( .A1(n10637), .A2(n9743), .ZN(n6896) );
  OAI21_X1 U8727 ( .B1(n9744), .B2(n9076), .A(n6896), .ZN(P2_U3462) );
  INV_X1 U8728 ( .A(n6897), .ZN(n6898) );
  OAI222_X1 U8729 ( .A1(n9433), .A2(P2_U3151), .B1(n8274), .B2(n6898), .C1(
        n9278), .C2(n9798), .ZN(P2_U3281) );
  INV_X1 U8730 ( .A(n7389), .ZN(n7397) );
  OAI222_X1 U8731 ( .A1(n10338), .A2(n9269), .B1(n8546), .B2(n6898), .C1(
        P1_U3086), .C2(n7397), .ZN(P1_U3341) );
  OAI21_X1 U8732 ( .B1(n6900), .B2(n8746), .A(n6899), .ZN(n7429) );
  INV_X1 U8733 ( .A(n6901), .ZN(n6902) );
  AOI211_X1 U8734 ( .C1(n5891), .C2(n6902), .A(n10502), .B(n4893), .ZN(n7424)
         );
  XNOR2_X1 U8735 ( .A(n8820), .B(n8627), .ZN(n6905) );
  INV_X1 U8736 ( .A(n6903), .ZN(n6904) );
  OAI21_X1 U8737 ( .B1(n6905), .B2(n10203), .A(n6904), .ZN(n7422) );
  AOI211_X1 U8738 ( .C1(n10520), .C2(n7429), .A(n7424), .B(n7422), .ZN(n6908)
         );
  AOI22_X1 U8739 ( .A1(n8889), .A2(n5891), .B1(n10534), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6906) );
  OAI21_X1 U8740 ( .B1(n6908), .B2(n10534), .A(n6906), .ZN(P1_U3525) );
  INV_X1 U8741 ( .A(n10329), .ZN(n8098) );
  AOI22_X1 U8742 ( .A1(n8098), .A2(n5891), .B1(P1_REG0_REG_3__SCAN_IN), .B2(
        n6596), .ZN(n6907) );
  OAI21_X1 U8743 ( .B1(n6908), .B2(n6596), .A(n6907), .ZN(P1_U3462) );
  INV_X1 U8744 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6914) );
  INV_X1 U8745 ( .A(n8480), .ZN(n6909) );
  OAI21_X1 U8746 ( .B1(n9711), .B2(n9730), .A(n6909), .ZN(n6912) );
  INV_X1 U8747 ( .A(n6910), .ZN(n6911) );
  OAI211_X1 U8748 ( .C1(n9716), .C2(n7044), .A(n6912), .B(n6911), .ZN(n9745)
         );
  NAND2_X1 U8749 ( .A1(n10649), .A2(n9745), .ZN(n6913) );
  OAI21_X1 U8750 ( .B1(n10649), .B2(n6914), .A(n6913), .ZN(P2_U3390) );
  INV_X1 U8751 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9241) );
  NOR2_X1 U8752 ( .A1(n6915), .A2(n9241), .ZN(P2_U3259) );
  INV_X1 U8753 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9270) );
  NOR2_X1 U8754 ( .A1(n6915), .A2(n9270), .ZN(P2_U3258) );
  INV_X1 U8755 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6916) );
  NOR2_X1 U8756 ( .A1(n6915), .A2(n6916), .ZN(P2_U3263) );
  INV_X1 U8757 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6917) );
  NOR2_X1 U8758 ( .A1(n6915), .A2(n6917), .ZN(P2_U3262) );
  INV_X1 U8759 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U8760 ( .A1(n6915), .A2(n6918), .ZN(P2_U3261) );
  INV_X1 U8761 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6919) );
  NOR2_X1 U8762 ( .A1(n6915), .A2(n6919), .ZN(P2_U3260) );
  INV_X1 U8763 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U8764 ( .A1(n6915), .A2(n6920), .ZN(P2_U3245) );
  INV_X1 U8765 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8766 ( .A1(n6915), .A2(n6921), .ZN(P2_U3244) );
  INV_X1 U8767 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6922) );
  NOR2_X1 U8768 ( .A1(n6915), .A2(n6922), .ZN(P2_U3238) );
  INV_X1 U8769 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U8770 ( .A1(n6915), .A2(n6923), .ZN(P2_U3243) );
  INV_X1 U8771 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8772 ( .A1(n6915), .A2(n6924), .ZN(P2_U3242) );
  INV_X1 U8773 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U8774 ( .A1(n6915), .A2(n6925), .ZN(P2_U3241) );
  INV_X1 U8775 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U8776 ( .A1(n6915), .A2(n6926), .ZN(P2_U3240) );
  INV_X1 U8777 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U8778 ( .A1(n6915), .A2(n6927), .ZN(P2_U3239) );
  INV_X1 U8779 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9259) );
  NOR2_X1 U8780 ( .A1(n6915), .A2(n9259), .ZN(P2_U3236) );
  INV_X1 U8781 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6928) );
  NOR2_X1 U8782 ( .A1(n6915), .A2(n6928), .ZN(P2_U3237) );
  INV_X1 U8783 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9191) );
  NOR2_X1 U8784 ( .A1(n6915), .A2(n9191), .ZN(P2_U3234) );
  INV_X1 U8785 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6929) );
  NOR2_X1 U8786 ( .A1(n6915), .A2(n6929), .ZN(P2_U3235) );
  INV_X1 U8787 ( .A(n10520), .ZN(n10284) );
  NAND2_X1 U8788 ( .A1(n6930), .A2(n8745), .ZN(n7123) );
  OAI21_X1 U8789 ( .B1(n6930), .B2(n8745), .A(n7123), .ZN(n7451) );
  INV_X1 U8790 ( .A(n7451), .ZN(n6939) );
  XOR2_X1 U8791 ( .A(n6931), .B(n8745), .Z(n6934) );
  OAI22_X1 U8792 ( .A1(n6933), .A2(n9908), .B1(n6932), .B2(n9887), .ZN(n7223)
         );
  AOI21_X1 U8793 ( .B1(n6934), .B2(n10427), .A(n7223), .ZN(n7453) );
  INV_X1 U8794 ( .A(n5127), .ZN(n6935) );
  AOI21_X1 U8795 ( .B1(n6937), .B2(n6936), .A(n6935), .ZN(n7444) );
  AOI22_X1 U8796 ( .A1(n7444), .A2(n10435), .B1(n10282), .B2(n6937), .ZN(n6938) );
  OAI211_X1 U8797 ( .C1(n10284), .C2(n6939), .A(n7453), .B(n6938), .ZN(n6941)
         );
  NAND2_X1 U8798 ( .A1(n6941), .A2(n10537), .ZN(n6940) );
  OAI21_X1 U8799 ( .B1(n10537), .B2(n6672), .A(n6940), .ZN(P1_U3526) );
  INV_X1 U8800 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8801 ( .A1(n6941), .A2(n10523), .ZN(n6942) );
  OAI21_X1 U8802 ( .B1(n10523), .B2(n6943), .A(n6942), .ZN(P1_U3465) );
  INV_X1 U8803 ( .A(n6944), .ZN(n6945) );
  OR2_X1 U8804 ( .A1(n6946), .A2(n6945), .ZN(n6951) );
  INV_X1 U8805 ( .A(n6947), .ZN(n6987) );
  NAND2_X1 U8806 ( .A1(n6953), .A2(n6987), .ZN(n6950) );
  INV_X1 U8807 ( .A(n6948), .ZN(n6949) );
  NAND4_X1 U8808 ( .A1(n6951), .A2(n7057), .A3(n6950), .A4(n6949), .ZN(n6956)
         );
  NAND2_X1 U8809 ( .A1(n6952), .A2(n6959), .ZN(n8522) );
  INV_X1 U8810 ( .A(n8522), .ZN(n6954) );
  AND2_X1 U8811 ( .A1(n6954), .A2(n6953), .ZN(n6955) );
  AOI21_X1 U8812 ( .B1(n6956), .B2(P2_STATE_REG_SCAN_IN), .A(n6955), .ZN(n7021) );
  OR2_X1 U8813 ( .A1(n7055), .A2(P2_U3151), .ZN(n8526) );
  INV_X1 U8814 ( .A(n9355), .ZN(n7335) );
  OR2_X1 U8815 ( .A1(n6986), .A2(n10622), .ZN(n6957) );
  NOR2_X1 U8816 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6958), .ZN(n7079) );
  AND2_X1 U8817 ( .A1(n6988), .A2(n6959), .ZN(n6960) );
  INV_X1 U8818 ( .A(n9387), .ZN(n7026) );
  INV_X1 U8819 ( .A(n6960), .ZN(n6962) );
  OAI22_X1 U8820 ( .A1(n9358), .A2(n5304), .B1(n7026), .B2(n9327), .ZN(n6963)
         );
  AOI211_X1 U8821 ( .C1(n6964), .C2(n9360), .A(n7079), .B(n6963), .ZN(n6996)
         );
  NOR2_X1 U8822 ( .A1(n8070), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6966) );
  INV_X1 U8823 ( .A(n6968), .ZN(n6970) );
  AOI21_X1 U8824 ( .B1(n6971), .B2(n6970), .A(n6969), .ZN(n6972) );
  NAND2_X1 U8825 ( .A1(n7023), .A2(n7024), .ZN(n7022) );
  INV_X1 U8826 ( .A(n6982), .ZN(n6983) );
  NAND2_X1 U8827 ( .A1(n7022), .A2(n6983), .ZN(n7101) );
  XNOR2_X1 U8828 ( .A(n4513), .B(n10623), .ZN(n6984) );
  XNOR2_X1 U8829 ( .A(n6984), .B(n9387), .ZN(n7102) );
  NAND2_X1 U8830 ( .A1(n7101), .A2(n7102), .ZN(n6992) );
  NAND2_X1 U8831 ( .A1(n7026), .A2(n6984), .ZN(n6991) );
  AND2_X1 U8832 ( .A1(n6992), .A2(n6991), .ZN(n6994) );
  OR2_X1 U8833 ( .A1(n6986), .A2(n6985), .ZN(n6990) );
  NAND2_X1 U8834 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  INV_X1 U8835 ( .A(n9363), .ZN(n9342) );
  OAI211_X1 U8836 ( .C1(n6994), .C2(n6993), .A(n9342), .B(n6999), .ZN(n6995)
         );
  OAI211_X1 U8837 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7335), .A(n6996), .B(
        n6995), .ZN(P2_U3158) );
  INV_X1 U8838 ( .A(n9726), .ZN(n7017) );
  OR2_X1 U8839 ( .A1(n6997), .A2(n7017), .ZN(n6998) );
  XNOR2_X1 U8840 ( .A(n4513), .B(n7116), .ZN(n7000) );
  NAND2_X1 U8841 ( .A1(n5304), .A2(n7000), .ZN(n7317) );
  OAI21_X1 U8842 ( .B1(n5304), .B2(n7000), .A(n7317), .ZN(n7001) );
  AOI21_X1 U8843 ( .B1(n7002), .B2(n7001), .A(n7319), .ZN(n7007) );
  INV_X1 U8844 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7003) );
  NOR2_X1 U8845 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7003), .ZN(n7296) );
  OAI22_X1 U8846 ( .A1(n9358), .A2(n7321), .B1(n7017), .B2(n9327), .ZN(n7004)
         );
  AOI211_X1 U8847 ( .C1(n5303), .C2(n9360), .A(n7296), .B(n7004), .ZN(n7006)
         );
  NAND2_X1 U8848 ( .A1(n9355), .A2(n7114), .ZN(n7005) );
  OAI211_X1 U8849 ( .C1(n7007), .C2(n9363), .A(n7006), .B(n7005), .ZN(P2_U3170) );
  INV_X1 U8850 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7153) );
  NAND3_X1 U8851 ( .A1(n6884), .A2(n8483), .A3(n8309), .ZN(n7008) );
  NAND2_X1 U8852 ( .A1(n7009), .A2(n7008), .ZN(n7120) );
  NOR2_X1 U8853 ( .A1(n7116), .A2(n9716), .ZN(n7018) );
  AND2_X1 U8854 ( .A1(n7011), .A2(n7010), .ZN(n7015) );
  NAND3_X1 U8855 ( .A1(n7013), .A2(n8299), .A3(n7012), .ZN(n7014) );
  AND2_X1 U8856 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  OAI222_X1 U8857 ( .A1(n9644), .A2(n7017), .B1(n9646), .B2(n7321), .C1(n9642), 
        .C2(n7016), .ZN(n7117) );
  AOI211_X1 U8858 ( .C1(n9711), .C2(n7120), .A(n7018), .B(n7117), .ZN(n10639)
         );
  OR2_X1 U8859 ( .A1(n10639), .A2(n9743), .ZN(n7019) );
  OAI21_X1 U8860 ( .B1(n9744), .B2(n7153), .A(n7019), .ZN(P2_U3463) );
  AND2_X1 U8861 ( .A1(n7021), .A2(n7020), .ZN(n7107) );
  INV_X1 U8862 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7030) );
  OAI21_X1 U8863 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7028) );
  AOI22_X1 U8864 ( .A1(n9354), .A2(n5679), .B1(n6978), .B2(n9360), .ZN(n7025)
         );
  OAI21_X1 U8865 ( .B1(n7026), .B2(n9358), .A(n7025), .ZN(n7027) );
  AOI21_X1 U8866 ( .B1(n9342), .B2(n7028), .A(n7027), .ZN(n7029) );
  OAI21_X1 U8867 ( .B1(n7107), .B2(n7030), .A(n7029), .ZN(P2_U3162) );
  AND2_X1 U8868 ( .A1(n5698), .A2(n8513), .ZN(n10621) );
  NAND2_X1 U8869 ( .A1(n10629), .A2(n10621), .ZN(n7221) );
  INV_X1 U8870 ( .A(n7031), .ZN(n9734) );
  NAND2_X1 U8871 ( .A1(n10629), .A2(n9734), .ZN(n7032) );
  NAND2_X1 U8872 ( .A1(n7088), .A2(n8303), .ZN(n7033) );
  INV_X1 U8873 ( .A(n8482), .ZN(n7034) );
  XNOR2_X1 U8874 ( .A(n7033), .B(n7034), .ZN(n7183) );
  INV_X1 U8875 ( .A(n7183), .ZN(n7041) );
  INV_X1 U8876 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7171) );
  AOI21_X1 U8877 ( .B1(n7035), .B2(n7034), .A(n9642), .ZN(n7038) );
  OAI22_X1 U8878 ( .A1(n7463), .A2(n9646), .B1(n7321), .B2(n9644), .ZN(n7037)
         );
  AOI21_X1 U8879 ( .B1(n7038), .B2(n7036), .A(n7037), .ZN(n7181) );
  MUX2_X1 U8880 ( .A(n7171), .B(n7181), .S(n10629), .Z(n7040) );
  AOI22_X1 U8881 ( .A1(n9651), .A2(n9345), .B1(n10628), .B2(n9347), .ZN(n7039)
         );
  OAI211_X1 U8882 ( .C1(n8900), .C2(n7041), .A(n7040), .B(n7039), .ZN(P2_U3227) );
  INV_X1 U8883 ( .A(n7042), .ZN(n7098) );
  OAI222_X1 U8884 ( .A1(n8546), .A2(n7098), .B1(n7723), .B2(P1_U3086), .C1(
        n7043), .C2(n10338), .ZN(P1_U3340) );
  INV_X1 U8885 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7208) );
  INV_X1 U8886 ( .A(n9360), .ZN(n8930) );
  OAI22_X1 U8887 ( .A1(n8930), .A2(n7044), .B1(n9363), .B2(n8480), .ZN(n7045)
         );
  AOI21_X1 U8888 ( .B1(n9346), .B2(n9725), .A(n7045), .ZN(n7046) );
  OAI21_X1 U8889 ( .B1(n7107), .B2(n7208), .A(n7046), .ZN(P2_U3172) );
  NOR2_X1 U8890 ( .A1(n9521), .A2(P2_U3151), .ZN(n8092) );
  NAND2_X1 U8891 ( .A1(n7067), .A2(n8092), .ZN(n7048) );
  MUX2_X1 U8892 ( .A(n7048), .B(n9500), .S(n7047), .Z(n10598) );
  MUX2_X1 U8893 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5669), .Z(n7050) );
  AOI21_X1 U8894 ( .B1(n7049), .B2(n4751), .A(n10542), .ZN(n10562) );
  XOR2_X1 U8895 ( .A(n10570), .B(n7050), .Z(n10563) );
  NOR2_X1 U8896 ( .A1(n10562), .A2(n10563), .ZN(n10560) );
  MUX2_X1 U8897 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9521), .Z(n7146) );
  XNOR2_X1 U8898 ( .A(n7146), .B(n7051), .ZN(n7052) );
  OAI21_X1 U8899 ( .B1(n7053), .B2(n7052), .A(n7144), .ZN(n7054) );
  NAND2_X1 U8900 ( .A1(n7054), .A2(n10612), .ZN(n7085) );
  INV_X1 U8901 ( .A(n7055), .ZN(n7056) );
  NOR2_X1 U8902 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  INV_X1 U8903 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7059) );
  MUX2_X1 U8904 ( .A(n7059), .B(P2_REG1_REG_2__SCAN_IN), .S(n10570), .Z(n10573) );
  NAND2_X1 U8905 ( .A1(n4642), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7060) );
  NAND2_X1 U8906 ( .A1(n10549), .A2(n7060), .ZN(n7062) );
  NAND2_X1 U8907 ( .A1(n7061), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U8908 ( .A1(n7062), .A2(n7063), .ZN(n10552) );
  OR2_X1 U8909 ( .A1(n10552), .A2(n10553), .ZN(n10550) );
  NAND2_X1 U8910 ( .A1(n10550), .A2(n7063), .ZN(n10572) );
  NAND2_X1 U8911 ( .A1(n7071), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U8912 ( .A1(n7065), .A2(n9076), .ZN(n7066) );
  AND2_X1 U8913 ( .A1(n7287), .A2(n7066), .ZN(n7082) );
  NOR2_X1 U8914 ( .A1(n5668), .A2(P2_U3151), .ZN(n8191) );
  AND2_X1 U8915 ( .A1(n7067), .A2(n8191), .ZN(n7206) );
  INV_X1 U8916 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U8917 ( .A1(n4642), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U8918 ( .A1(n10549), .A2(n7068), .ZN(n7069) );
  NAND2_X1 U8919 ( .A1(n7061), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7070) );
  NAND2_X1 U8920 ( .A1(n7069), .A2(n7070), .ZN(n10540) );
  INV_X1 U8921 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10541) );
  OR2_X1 U8922 ( .A1(n10540), .A2(n10541), .ZN(n10538) );
  NAND2_X1 U8923 ( .A1(n10538), .A2(n7070), .ZN(n10558) );
  NAND2_X1 U8924 ( .A1(n7071), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7072) );
  OAI21_X1 U8925 ( .B1(n7073), .B2(n7145), .A(n7291), .ZN(n7076) );
  INV_X1 U8926 ( .A(n7076), .ZN(n7074) );
  INV_X1 U8927 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8928 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  NAND2_X1 U8929 ( .A1(n7292), .A2(n7077), .ZN(n7078) );
  NAND2_X1 U8930 ( .A1(n10566), .A2(n7078), .ZN(n7081) );
  INV_X1 U8931 ( .A(n7079), .ZN(n7080) );
  OAI211_X1 U8932 ( .C1(n7082), .C2(n10606), .A(n7081), .B(n7080), .ZN(n7083)
         );
  AOI21_X1 U8933 ( .B1(n7301), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7083), .ZN(
        n7084) );
  OAI211_X1 U8934 ( .C1(n10598), .C2(n7145), .A(n7085), .B(n7084), .ZN(
        P2_U3185) );
  OR2_X1 U8935 ( .A1(n7086), .A2(n7089), .ZN(n7087) );
  OAI22_X1 U8936 ( .A1(n7222), .A2(n9737), .B1(n7320), .B2(n9716), .ZN(n7095)
         );
  XNOR2_X1 U8937 ( .A(n7090), .B(n7089), .ZN(n7094) );
  INV_X1 U8938 ( .A(n7222), .ZN(n7091) );
  NAND2_X1 U8939 ( .A1(n7091), .A2(n9734), .ZN(n7093) );
  AOI22_X1 U8940 ( .A1(n9724), .A2(n5305), .B1(n9385), .B2(n6257), .ZN(n7092)
         );
  OAI211_X1 U8941 ( .C1(n9642), .C2(n7094), .A(n7093), .B(n7092), .ZN(n7217)
         );
  NOR2_X1 U8942 ( .A1(n7095), .A2(n7217), .ZN(n10641) );
  INV_X1 U8943 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7268) );
  OR2_X1 U8944 ( .A1(n9744), .A2(n7268), .ZN(n7096) );
  OAI21_X1 U8945 ( .B1(n10641), .B2(n9743), .A(n7096), .ZN(P2_U3464) );
  INV_X1 U8946 ( .A(n9456), .ZN(n9446) );
  OAI222_X1 U8947 ( .A1(P2_U3151), .A2(n9446), .B1(n8274), .B2(n7098), .C1(
        n7097), .C2(n9798), .ZN(P2_U3280) );
  INV_X1 U8948 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7106) );
  OAI22_X1 U8949 ( .A1(n8930), .A2(n10623), .B1(n9327), .B2(n7099), .ZN(n7100)
         );
  AOI21_X1 U8950 ( .B1(n9346), .B2(n9726), .A(n7100), .ZN(n7105) );
  OAI21_X1 U8951 ( .B1(n7102), .B2(n7101), .A(n6992), .ZN(n7103) );
  NAND2_X1 U8952 ( .A1(n7103), .A2(n9342), .ZN(n7104) );
  OAI211_X1 U8953 ( .C1(n7107), .C2(n7106), .A(n7105), .B(n7104), .ZN(P2_U3177) );
  OAI22_X1 U8954 ( .A1(n9637), .A2(n7108), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8222), .ZN(n7111) );
  MUX2_X1 U8955 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7109), .S(n10629), .Z(n7110)
         );
  AOI211_X1 U8956 ( .C1(n9657), .C2(n7112), .A(n7111), .B(n7110), .ZN(n7113)
         );
  INV_X1 U8957 ( .A(n7113), .ZN(P2_U3230) );
  INV_X1 U8958 ( .A(n7114), .ZN(n7115) );
  OAI22_X1 U8959 ( .A1(n9637), .A2(n7116), .B1(n7115), .B2(n8222), .ZN(n7119)
         );
  MUX2_X1 U8960 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7117), .S(n10629), .Z(n7118)
         );
  AOI211_X1 U8961 ( .C1(n9657), .C2(n7120), .A(n7119), .B(n7118), .ZN(n7121)
         );
  INV_X1 U8962 ( .A(n7121), .ZN(P2_U3229) );
  NAND2_X1 U8963 ( .A1(n7123), .A2(n7122), .ZN(n7127) );
  AND2_X1 U8964 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  OAI21_X1 U8965 ( .B1(n7127), .B2(n7130), .A(n7126), .ZN(n7698) );
  INV_X1 U8966 ( .A(n7248), .ZN(n7128) );
  NAND2_X1 U8967 ( .A1(n7129), .A2(n8635), .ZN(n7131) );
  NAND2_X1 U8968 ( .A1(n7131), .A2(n7130), .ZN(n7133) );
  NAND3_X1 U8969 ( .A1(n7133), .A2(n7132), .A3(n10427), .ZN(n7138) );
  OR2_X1 U8970 ( .A1(n7362), .A2(n9908), .ZN(n7136) );
  OR2_X1 U8971 ( .A1(n7134), .A2(n9887), .ZN(n7135) );
  NAND2_X1 U8972 ( .A1(n7136), .A2(n7135), .ZN(n7339) );
  INV_X1 U8973 ( .A(n7339), .ZN(n7137) );
  NAND2_X1 U8974 ( .A1(n7138), .A2(n7137), .ZN(n7695) );
  AOI211_X1 U8975 ( .C1(n10520), .C2(n7698), .A(n7690), .B(n7695), .ZN(n7143)
         );
  INV_X1 U8976 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7139) );
  OAI22_X1 U8977 ( .A1(n10329), .A2(n7341), .B1(n10523), .B2(n7139), .ZN(n7140) );
  INV_X1 U8978 ( .A(n7140), .ZN(n7141) );
  OAI21_X1 U8979 ( .B1(n7143), .B2(n6596), .A(n7141), .ZN(P1_U3468) );
  AOI22_X1 U8980 ( .A1(n8889), .A2(n7692), .B1(n10534), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7142) );
  OAI21_X1 U8981 ( .B1(n7143), .B2(n10534), .A(n7142), .ZN(P1_U3527) );
  MUX2_X1 U8982 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9521), .Z(n7149) );
  MUX2_X1 U8983 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9521), .Z(n7147) );
  XOR2_X1 U8984 ( .A(n7165), .B(n7147), .Z(n7282) );
  AOI21_X1 U8985 ( .B1(n7147), .B2(n7304), .A(n7280), .ZN(n7264) );
  XOR2_X1 U8986 ( .A(n7148), .B(n7149), .Z(n7265) );
  NOR2_X1 U8987 ( .A1(n7264), .A2(n7265), .ZN(n7263) );
  MUX2_X1 U8988 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9521), .Z(n7538) );
  XNOR2_X1 U8989 ( .A(n7538), .B(n7172), .ZN(n7150) );
  OAI21_X1 U8990 ( .B1(n7151), .B2(n7150), .A(n7539), .ZN(n7152) );
  NAND2_X1 U8991 ( .A1(n7152), .A2(n10612), .ZN(n7180) );
  MUX2_X1 U8992 ( .A(n7153), .B(P2_REG1_REG_4__SCAN_IN), .S(n7165), .Z(n7284)
         );
  NAND2_X1 U8993 ( .A1(n7154), .A2(n7284), .ZN(n7289) );
  OR2_X1 U8994 ( .A1(n7165), .A2(n7153), .ZN(n7155) );
  NAND2_X1 U8995 ( .A1(n4583), .A2(n7157), .ZN(n7269) );
  INV_X1 U8996 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7158) );
  OR2_X1 U8997 ( .A1(n7172), .A2(n7158), .ZN(n7548) );
  NAND2_X1 U8998 ( .A1(n7172), .A2(n7158), .ZN(n7159) );
  NAND2_X1 U8999 ( .A1(n7548), .A2(n7159), .ZN(n7160) );
  AOI21_X1 U9000 ( .B1(n4615), .B2(n7160), .A(n7550), .ZN(n7163) );
  INV_X1 U9001 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7161) );
  NOR2_X1 U9002 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7161), .ZN(n9344) );
  INV_X1 U9003 ( .A(n9344), .ZN(n7162) );
  OAI21_X1 U9004 ( .B1(n10606), .B2(n7163), .A(n7162), .ZN(n7178) );
  INV_X1 U9005 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7164) );
  MUX2_X1 U9006 ( .A(n7164), .B(P2_REG2_REG_4__SCAN_IN), .S(n7165), .Z(n7290)
         );
  OR2_X1 U9007 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  INV_X1 U9008 ( .A(n7170), .ZN(n7169) );
  OR2_X1 U9009 ( .A1(n7167), .A2(n7279), .ZN(n7168) );
  NAND2_X1 U9010 ( .A1(n7169), .A2(n7168), .ZN(n7271) );
  INV_X1 U9011 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7270) );
  NOR2_X1 U9012 ( .A1(n7271), .A2(n7270), .ZN(n7273) );
  NOR2_X1 U9013 ( .A1(n7170), .A2(n7273), .ZN(n7175) );
  OR2_X1 U9014 ( .A1(n7172), .A2(n7171), .ZN(n7525) );
  NAND2_X1 U9015 ( .A1(n7172), .A2(n7171), .ZN(n7173) );
  NAND2_X1 U9016 ( .A1(n7525), .A2(n7173), .ZN(n7174) );
  AOI21_X1 U9017 ( .B1(n7175), .B2(n7174), .A(n7527), .ZN(n7176) );
  NOR2_X1 U9018 ( .A1(n10615), .A2(n7176), .ZN(n7177) );
  AOI211_X1 U9019 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n7301), .A(n7178), .B(
        n7177), .ZN(n7179) );
  OAI211_X1 U9020 ( .C1(n10598), .C2(n7537), .A(n7180), .B(n7179), .ZN(
        P2_U3188) );
  OAI21_X1 U9021 ( .B1(n7316), .B2(n9716), .A(n7181), .ZN(n7182) );
  AOI21_X1 U9022 ( .B1(n7183), .B2(n9711), .A(n7182), .ZN(n10643) );
  OR2_X1 U9023 ( .A1(n9744), .A2(n7158), .ZN(n7184) );
  OAI21_X1 U9024 ( .B1(n10643), .B2(n9743), .A(n7184), .ZN(P2_U3465) );
  NOR2_X1 U9025 ( .A1(n7192), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7186) );
  INV_X1 U9026 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10535) );
  MUX2_X1 U9027 ( .A(n10535), .B(P1_REG1_REG_13__SCAN_IN), .S(n7234), .Z(n7185) );
  NOR3_X1 U9028 ( .A1(n7187), .A2(n7186), .A3(n7185), .ZN(n7233) );
  INV_X1 U9029 ( .A(n7233), .ZN(n7189) );
  OAI21_X1 U9030 ( .B1(n7187), .B2(n7186), .A(n7185), .ZN(n7188) );
  NAND3_X1 U9031 ( .A1(n7189), .A2(n10033), .A3(n7188), .ZN(n7198) );
  NOR2_X1 U9032 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7190), .ZN(n7196) );
  NAND2_X1 U9033 ( .A1(n7234), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7237) );
  OAI21_X1 U9034 ( .B1(n7234), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7237), .ZN(
        n7194) );
  OAI21_X1 U9035 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7192), .A(n7191), .ZN(
        n7193) );
  NOR2_X1 U9036 ( .A1(n7193), .A2(n7194), .ZN(n7239) );
  AOI211_X1 U9037 ( .C1(n7194), .C2(n7193), .A(n7239), .B(n7948), .ZN(n7195)
         );
  AOI211_X1 U9038 ( .C1(n10021), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7196), .B(
        n7195), .ZN(n7197) );
  OAI211_X1 U9039 ( .C1(n10007), .C2(n7199), .A(n7198), .B(n7197), .ZN(
        P1_U3256) );
  INV_X1 U9040 ( .A(n7200), .ZN(n7205) );
  INV_X1 U9041 ( .A(n7201), .ZN(n7202) );
  MUX2_X1 U9042 ( .A(n7202), .B(n10541), .S(n10632), .Z(n7204) );
  AOI22_X1 U9043 ( .A1(n9651), .A2(n6978), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10628), .ZN(n7203) );
  OAI211_X1 U9044 ( .C1(n8900), .C2(n7205), .A(n7204), .B(n7203), .ZN(P2_U3232) );
  NOR2_X1 U9045 ( .A1(n10612), .A2(n7206), .ZN(n7210) );
  AOI21_X1 U9046 ( .B1(n4642), .B2(n7207), .A(n10543), .ZN(n7209) );
  OAI22_X1 U9047 ( .A1(n7210), .A2(n7209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7208), .ZN(n7211) );
  AOI21_X1 U9048 ( .B1(n7301), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7211), .ZN(
        n7212) );
  OAI21_X1 U9049 ( .B1(n4642), .B2(n10598), .A(n7212), .ZN(P2_U3182) );
  INV_X1 U9050 ( .A(n7213), .ZN(n7216) );
  INV_X1 U9051 ( .A(n7808), .ZN(n7717) );
  OAI222_X1 U9052 ( .A1(n8891), .A2(n7214), .B1(n8546), .B2(n7216), .C1(
        P1_U3086), .C2(n7717), .ZN(P1_U3339) );
  OAI222_X1 U9053 ( .A1(n9475), .A2(P2_U3151), .B1(n8274), .B2(n7216), .C1(
        n7215), .C2(n9798), .ZN(P2_U3279) );
  MUX2_X1 U9054 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7217), .S(n10629), .Z(n7218)
         );
  INV_X1 U9055 ( .A(n7218), .ZN(n7220) );
  INV_X1 U9056 ( .A(n7320), .ZN(n9308) );
  AOI22_X1 U9057 ( .A1(n9651), .A2(n9308), .B1(n10628), .B2(n9309), .ZN(n7219)
         );
  OAI211_X1 U9058 ( .C1(n7222), .C2(n7221), .A(n7220), .B(n7219), .ZN(P2_U3228) );
  NAND2_X1 U9059 ( .A1(n9916), .A2(n7223), .ZN(n7224) );
  OAI211_X1 U9060 ( .C1(n9931), .C2(n7449), .A(n7225), .B(n7224), .ZN(n7231)
         );
  INV_X1 U9061 ( .A(n7227), .ZN(n7228) );
  AOI211_X1 U9062 ( .C1(n7229), .C2(n7226), .A(n10416), .B(n7228), .ZN(n7230)
         );
  AOI211_X1 U9063 ( .C1(n7446), .C2(n9927), .A(n7231), .B(n7230), .ZN(n7232)
         );
  INV_X1 U9064 ( .A(n7232), .ZN(P1_U3230) );
  AOI21_X1 U9065 ( .B1(n7234), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7233), .ZN(
        n7392) );
  XNOR2_X1 U9066 ( .A(n7397), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7394) );
  XNOR2_X1 U9067 ( .A(n7392), .B(n7394), .ZN(n7245) );
  AND2_X1 U9068 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7235) );
  AOI21_X1 U9069 ( .B1(n10021), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7235), .ZN(
        n7236) );
  OAI21_X1 U9070 ( .B1(n7397), .B2(n10007), .A(n7236), .ZN(n7244) );
  INV_X1 U9071 ( .A(n7237), .ZN(n7238) );
  NOR2_X1 U9072 ( .A1(n7239), .A2(n7238), .ZN(n7242) );
  NAND2_X1 U9073 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n7389), .ZN(n7240) );
  OAI21_X1 U9074 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7389), .A(n7240), .ZN(
        n7241) );
  NOR2_X1 U9075 ( .A1(n7242), .A2(n7241), .ZN(n7388) );
  AOI211_X1 U9076 ( .C1(n7242), .C2(n7241), .A(n7388), .B(n7948), .ZN(n7243)
         );
  AOI211_X1 U9077 ( .C1(n10033), .C2(n7245), .A(n7244), .B(n7243), .ZN(n7246)
         );
  INV_X1 U9078 ( .A(n7246), .ZN(P1_U3257) );
  NAND2_X1 U9079 ( .A1(n7247), .A2(n7249), .ZN(n7371) );
  OAI21_X1 U9080 ( .B1(n7247), .B2(n7249), .A(n7371), .ZN(n10459) );
  AOI211_X1 U9081 ( .C1(n10449), .C2(n7248), .A(n10502), .B(n7373), .ZN(n10451) );
  XOR2_X1 U9082 ( .A(n7377), .B(n7249), .Z(n7251) );
  AOI22_X1 U9083 ( .A1(n9957), .A2(n9865), .B1(n9910), .B2(n9959), .ZN(n10412)
         );
  INV_X1 U9084 ( .A(n10412), .ZN(n7250) );
  AOI21_X1 U9085 ( .B1(n7251), .B2(n10427), .A(n7250), .ZN(n10461) );
  INV_X1 U9086 ( .A(n10461), .ZN(n7252) );
  AOI211_X1 U9087 ( .C1(n10520), .C2(n10459), .A(n10451), .B(n7252), .ZN(n7257) );
  INV_X1 U9088 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7253) );
  NOR2_X1 U9089 ( .A1(n10523), .A2(n7253), .ZN(n7254) );
  AOI21_X1 U9090 ( .B1(n8098), .B2(n10449), .A(n7254), .ZN(n7255) );
  OAI21_X1 U9091 ( .B1(n7257), .B2(n6596), .A(n7255), .ZN(P1_U3471) );
  AOI22_X1 U9092 ( .A1(n8889), .A2(n10449), .B1(n10534), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7256) );
  OAI21_X1 U9093 ( .B1(n7257), .B2(n10534), .A(n7256), .ZN(P1_U3528) );
  INV_X1 U9094 ( .A(n9507), .ZN(n9494) );
  INV_X1 U9095 ( .A(n7258), .ZN(n7260) );
  OAI222_X1 U9096 ( .A1(P2_U3151), .A2(n9494), .B1(n8274), .B2(n7260), .C1(
        n7259), .C2(n9798), .ZN(P2_U3278) );
  INV_X1 U9097 ( .A(n7937), .ZN(n7732) );
  OAI222_X1 U9098 ( .A1(n8891), .A2(n7261), .B1(n7732), .B2(P1_U3086), .C1(
        n8546), .C2(n7260), .ZN(P1_U3338) );
  NAND2_X1 U9099 ( .A1(n9500), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7262) );
  OAI21_X1 U9100 ( .B1(n9500), .B2(n8449), .A(n7262), .ZN(P2_U3521) );
  INV_X1 U9101 ( .A(n10612), .ZN(n10561) );
  AOI211_X1 U9102 ( .C1(n7265), .C2(n7264), .A(n10561), .B(n7263), .ZN(n7266)
         );
  INV_X1 U9103 ( .A(n7266), .ZN(n7278) );
  AOI21_X1 U9104 ( .B1(n7269), .B2(n7268), .A(n7267), .ZN(n7275) );
  AND2_X1 U9105 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  OAI21_X1 U9106 ( .B1(n7273), .B2(n7272), .A(n10566), .ZN(n7274) );
  NAND2_X1 U9107 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9306) );
  OAI211_X1 U9108 ( .C1(n7275), .C2(n10606), .A(n7274), .B(n9306), .ZN(n7276)
         );
  AOI21_X1 U9109 ( .B1(n7301), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7276), .ZN(
        n7277) );
  OAI211_X1 U9110 ( .C1(n10598), .C2(n7279), .A(n7278), .B(n7277), .ZN(
        P2_U3187) );
  AOI211_X1 U9111 ( .C1(n7282), .C2(n7281), .A(n10561), .B(n7280), .ZN(n7283)
         );
  INV_X1 U9112 ( .A(n7283), .ZN(n7303) );
  INV_X1 U9113 ( .A(n7284), .ZN(n7286) );
  NAND3_X1 U9114 ( .A1(n7287), .A2(n7286), .A3(n7285), .ZN(n7288) );
  AND2_X1 U9115 ( .A1(n7289), .A2(n7288), .ZN(n7299) );
  NAND3_X1 U9116 ( .A1(n7292), .A2(n4925), .A3(n7291), .ZN(n7293) );
  NAND2_X1 U9117 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  NAND2_X1 U9118 ( .A1(n10566), .A2(n7295), .ZN(n7298) );
  INV_X1 U9119 ( .A(n7296), .ZN(n7297) );
  OAI211_X1 U9120 ( .C1(n7299), .C2(n10606), .A(n7298), .B(n7297), .ZN(n7300)
         );
  AOI21_X1 U9121 ( .B1(n7301), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7300), .ZN(
        n7302) );
  OAI211_X1 U9122 ( .C1(n10598), .C2(n7304), .A(n7303), .B(n7302), .ZN(
        P2_U3186) );
  XNOR2_X1 U9123 ( .A(n7306), .B(n7305), .ZN(n7350) );
  INV_X1 U9124 ( .A(n9385), .ZN(n7330) );
  INV_X1 U9125 ( .A(n7307), .ZN(n7308) );
  AOI21_X1 U9126 ( .B1(n8487), .B2(n7309), .A(n7308), .ZN(n7310) );
  OAI222_X1 U9127 ( .A1(n9646), .A2(n7468), .B1(n9644), .B2(n7330), .C1(n9642), 
        .C2(n7310), .ZN(n7351) );
  AOI21_X1 U9128 ( .B1(n9711), .B2(n7350), .A(n7351), .ZN(n7313) );
  INV_X1 U9129 ( .A(n9715), .ZN(n9670) );
  INV_X1 U9130 ( .A(n7331), .ZN(n7354) );
  AOI22_X1 U9131 ( .A1(n9670), .A2(n7354), .B1(n9743), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7311) );
  OAI21_X1 U9132 ( .B1(n7313), .B2(n9743), .A(n7311), .ZN(P2_U3466) );
  AOI22_X1 U9133 ( .A1(n6261), .A2(n7354), .B1(n10652), .B2(
        P2_REG0_REG_7__SCAN_IN), .ZN(n7312) );
  OAI21_X1 U9134 ( .B1(n7313), .B2(n10652), .A(n7312), .ZN(P2_U3411) );
  INV_X1 U9135 ( .A(n7314), .ZN(n7337) );
  INV_X1 U9136 ( .A(n9514), .ZN(n9525) );
  OAI222_X1 U9137 ( .A1(n9798), .A2(n7315), .B1(n8274), .B2(n7337), .C1(
        P2_U3151), .C2(n9525), .ZN(P2_U3277) );
  INV_X1 U9138 ( .A(n7353), .ZN(n7336) );
  XNOR2_X1 U9139 ( .A(n7316), .B(n8600), .ZN(n7324) );
  INV_X1 U9140 ( .A(n7324), .ZN(n7325) );
  INV_X1 U9141 ( .A(n7317), .ZN(n7318) );
  XNOR2_X1 U9142 ( .A(n8600), .B(n7320), .ZN(n7322) );
  XNOR2_X1 U9143 ( .A(n7321), .B(n7322), .ZN(n9303) );
  NOR2_X1 U9144 ( .A1(n9304), .A2(n9303), .ZN(n9340) );
  INV_X1 U9145 ( .A(n7322), .ZN(n7323) );
  NOR2_X1 U9146 ( .A1(n7323), .A2(n9386), .ZN(n9339) );
  XOR2_X1 U9147 ( .A(n9385), .B(n7324), .Z(n9338) );
  NOR3_X1 U9148 ( .A1(n9340), .A2(n9339), .A3(n9338), .ZN(n9337) );
  AOI21_X1 U9149 ( .B1(n9385), .B2(n7325), .A(n9337), .ZN(n7328) );
  XNOR2_X1 U9150 ( .A(n7331), .B(n8244), .ZN(n7326) );
  NOR2_X1 U9151 ( .A1(n7326), .A2(n9384), .ZN(n7454) );
  AOI21_X1 U9152 ( .B1(n9384), .B2(n7326), .A(n7454), .ZN(n7327) );
  NAND2_X1 U9153 ( .A1(n7328), .A2(n7327), .ZN(n7456) );
  OAI21_X1 U9154 ( .B1(n7328), .B2(n7327), .A(n7456), .ZN(n7329) );
  NAND2_X1 U9155 ( .A1(n7329), .A2(n9342), .ZN(n7334) );
  AND2_X1 U9156 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10584) );
  OAI22_X1 U9157 ( .A1(n8930), .A2(n7331), .B1(n9327), .B2(n7330), .ZN(n7332)
         );
  AOI211_X1 U9158 ( .C1(n9346), .C2(n9383), .A(n10584), .B(n7332), .ZN(n7333)
         );
  OAI211_X1 U9159 ( .C1(n7336), .C2(n7335), .A(n7334), .B(n7333), .ZN(P2_U3153) );
  INV_X1 U9160 ( .A(n8106), .ZN(n7955) );
  OAI222_X1 U9161 ( .A1(n8891), .A2(n7338), .B1(n7955), .B2(P1_U3086), .C1(
        n8546), .C2(n7337), .ZN(P1_U3337) );
  AOI22_X1 U9162 ( .A1(n9916), .A2(n7339), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7340) );
  OAI21_X1 U9163 ( .B1(n7341), .B2(n9931), .A(n7340), .ZN(n7348) );
  NAND2_X1 U9164 ( .A1(n7343), .A2(n7342), .ZN(n7344) );
  XOR2_X1 U9165 ( .A(n7345), .B(n7344), .Z(n7346) );
  NOR2_X1 U9166 ( .A1(n7346), .A2(n10416), .ZN(n7347) );
  AOI211_X1 U9167 ( .C1(n7691), .C2(n9927), .A(n7348), .B(n7347), .ZN(n7349)
         );
  INV_X1 U9168 ( .A(n7349), .ZN(P1_U3227) );
  INV_X1 U9169 ( .A(n7350), .ZN(n7357) );
  INV_X1 U9170 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7535) );
  INV_X1 U9171 ( .A(n7351), .ZN(n7352) );
  MUX2_X1 U9172 ( .A(n7535), .B(n7352), .S(n10629), .Z(n7356) );
  AOI22_X1 U9173 ( .A1(n9651), .A2(n7354), .B1(n10628), .B2(n7353), .ZN(n7355)
         );
  OAI211_X1 U9174 ( .C1(n8900), .C2(n7357), .A(n7356), .B(n7355), .ZN(P2_U3226) );
  NAND2_X1 U9175 ( .A1(n7359), .A2(n7358), .ZN(n7361) );
  XOR2_X1 U9176 ( .A(n7361), .B(n7360), .Z(n7369) );
  INV_X1 U9177 ( .A(n10440), .ZN(n7366) );
  OR2_X1 U9178 ( .A1(n7678), .A2(n9908), .ZN(n7364) );
  OR2_X1 U9179 ( .A1(n7362), .A2(n9887), .ZN(n7363) );
  NAND2_X1 U9180 ( .A1(n7364), .A2(n7363), .ZN(n7382) );
  AOI22_X1 U9181 ( .A1(n9916), .A2(n7382), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7365) );
  OAI21_X1 U9182 ( .B1(n10423), .B2(n7366), .A(n7365), .ZN(n7367) );
  AOI21_X1 U9183 ( .B1(n10442), .B2(n10421), .A(n7367), .ZN(n7368) );
  OAI21_X1 U9184 ( .B1(n7369), .B2(n10416), .A(n7368), .ZN(P1_U3213) );
  INV_X1 U9185 ( .A(n10499), .ZN(n10481) );
  NAND2_X1 U9186 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  OAI21_X1 U9187 ( .B1(n7372), .B2(n7376), .A(n4612), .ZN(n10445) );
  INV_X1 U9188 ( .A(n7373), .ZN(n7375) );
  INV_X1 U9189 ( .A(n7647), .ZN(n7374) );
  AOI211_X1 U9190 ( .C1(n10442), .C2(n7375), .A(n10502), .B(n7374), .ZN(n10443) );
  NAND2_X1 U9191 ( .A1(n7377), .A2(n8748), .ZN(n7378) );
  NAND2_X1 U9192 ( .A1(n7378), .A2(n8641), .ZN(n7379) );
  NAND2_X1 U9193 ( .A1(n7379), .A2(n5942), .ZN(n7675) );
  OAI21_X1 U9194 ( .B1(n5942), .B2(n7379), .A(n7675), .ZN(n7383) );
  INV_X1 U9195 ( .A(n10445), .ZN(n7380) );
  NOR2_X1 U9196 ( .A1(n7380), .A2(n7871), .ZN(n7381) );
  AOI211_X1 U9197 ( .C1(n10427), .C2(n7383), .A(n7382), .B(n7381), .ZN(n10448)
         );
  INV_X1 U9198 ( .A(n10448), .ZN(n7384) );
  AOI211_X1 U9199 ( .C1(n10481), .C2(n10445), .A(n10443), .B(n7384), .ZN(n7387) );
  AOI22_X1 U9200 ( .A1(n8098), .A2(n10442), .B1(n6596), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n7385) );
  OAI21_X1 U9201 ( .B1(n7387), .B2(n6596), .A(n7385), .ZN(P1_U3474) );
  AOI22_X1 U9202 ( .A1(n8889), .A2(n10442), .B1(n10534), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7386) );
  OAI21_X1 U9203 ( .B1(n7387), .B2(n10534), .A(n7386), .ZN(P1_U3529) );
  AOI21_X1 U9204 ( .B1(n7389), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7388), .ZN(
        n7724) );
  XNOR2_X1 U9205 ( .A(n7724), .B(n7723), .ZN(n7390) );
  NOR2_X1 U9206 ( .A1(n6029), .A2(n7390), .ZN(n7725) );
  AOI211_X1 U9207 ( .C1(n6029), .C2(n7390), .A(n7725), .B(n7948), .ZN(n7402)
         );
  NOR2_X1 U9208 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9924), .ZN(n7391) );
  AOI21_X1 U9209 ( .B1(n10021), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7391), .ZN(
        n7400) );
  INV_X1 U9210 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7396) );
  INV_X1 U9211 ( .A(n7392), .ZN(n7393) );
  NAND2_X1 U9212 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  OAI21_X1 U9213 ( .B1(n7397), .B2(n7396), .A(n7395), .ZN(n7712) );
  XNOR2_X1 U9214 ( .A(n7723), .B(n7712), .ZN(n7398) );
  NAND2_X1 U9215 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7398), .ZN(n7714) );
  OAI211_X1 U9216 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7398), .A(n10033), .B(
        n7714), .ZN(n7399) );
  OAI211_X1 U9217 ( .C1(n10007), .C2(n7723), .A(n7400), .B(n7399), .ZN(n7401)
         );
  OR2_X1 U9218 ( .A1(n7402), .A2(n7401), .ZN(P1_U3258) );
  NAND2_X1 U9219 ( .A1(n8271), .A2(n10343), .ZN(n7404) );
  OAI211_X1 U9220 ( .C1(n7405), .C2(n10338), .A(n7404), .B(n7403), .ZN(
        P1_U3335) );
  NOR2_X1 U9221 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  NAND2_X1 U9222 ( .A1(n7409), .A2(n7408), .ZN(n7413) );
  INV_X1 U9223 ( .A(n7410), .ZN(n7421) );
  AOI21_X2 U9224 ( .B1(n7493), .B2(n7871), .A(n10215), .ZN(n10458) );
  INV_X1 U9225 ( .A(n7411), .ZN(n7412) );
  AOI22_X1 U9226 ( .A1(n10450), .A2(n7414), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n10452), .ZN(n7416) );
  NAND2_X1 U9227 ( .A1(n10215), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7415) );
  OAI211_X1 U9228 ( .C1(n7417), .C2(n10456), .A(n7416), .B(n7415), .ZN(n7418)
         );
  AOI21_X1 U9229 ( .B1(n10458), .B2(n7419), .A(n7418), .ZN(n7420) );
  OAI21_X1 U9230 ( .B1(n10462), .B2(n7421), .A(n7420), .ZN(P1_U3291) );
  INV_X1 U9231 ( .A(n7422), .ZN(n7431) );
  AOI22_X1 U9232 ( .A1(n7424), .A2(n10450), .B1(n10452), .B2(n7423), .ZN(n7426) );
  NAND2_X1 U9233 ( .A1(n10215), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7425) );
  OAI211_X1 U9234 ( .C1(n7427), .C2(n10456), .A(n7426), .B(n7425), .ZN(n7428)
         );
  AOI21_X1 U9235 ( .B1(n10458), .B2(n7429), .A(n7428), .ZN(n7430) );
  OAI21_X1 U9236 ( .B1(n10462), .B2(n7431), .A(n7430), .ZN(P1_U3290) );
  INV_X1 U9237 ( .A(n7432), .ZN(n7434) );
  OAI222_X1 U9238 ( .A1(n8891), .A2(n7433), .B1(n8546), .B2(n7434), .C1(
        P1_U3086), .C2(n8816), .ZN(P1_U3336) );
  OAI222_X1 U9239 ( .A1(P2_U3151), .A2(n5694), .B1(n8274), .B2(n7434), .C1(
        n9197), .C2(n9798), .ZN(P2_U3276) );
  NAND2_X1 U9240 ( .A1(n10450), .A2(n10435), .ZN(n7517) );
  INV_X1 U9241 ( .A(n7517), .ZN(n7445) );
  OAI21_X1 U9242 ( .B1(n7445), .B2(n10441), .A(n7435), .ZN(n7443) );
  NAND3_X1 U9243 ( .A1(n7437), .A2(n8873), .A3(n7436), .ZN(n7439) );
  OAI211_X1 U9244 ( .C1(n10190), .C2(n7440), .A(n7439), .B(n7438), .ZN(n7441)
         );
  NAND2_X1 U9245 ( .A1(n8066), .A2(n7441), .ZN(n7442) );
  OAI211_X1 U9246 ( .C1(n6736), .C2(n8066), .A(n7443), .B(n7442), .ZN(P1_U3293) );
  NAND2_X1 U9247 ( .A1(n7445), .A2(n7444), .ZN(n7448) );
  AOI22_X1 U9248 ( .A1(n10462), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7446), .B2(
        n10452), .ZN(n7447) );
  OAI211_X1 U9249 ( .C1(n7449), .C2(n10456), .A(n7448), .B(n7447), .ZN(n7450)
         );
  AOI21_X1 U9250 ( .B1(n10458), .B2(n7451), .A(n7450), .ZN(n7452) );
  OAI21_X1 U9251 ( .B1(n7453), .B2(n10462), .A(n7452), .ZN(P1_U3289) );
  XNOR2_X1 U9252 ( .A(n8266), .B(n8600), .ZN(n7467) );
  XNOR2_X1 U9253 ( .A(n7467), .B(n7468), .ZN(n7458) );
  INV_X1 U9254 ( .A(n7454), .ZN(n7455) );
  NAND2_X1 U9255 ( .A1(n7456), .A2(n7455), .ZN(n7457) );
  OAI21_X1 U9256 ( .B1(n7458), .B2(n7457), .A(n7473), .ZN(n7459) );
  NAND2_X1 U9257 ( .A1(n7459), .A2(n9342), .ZN(n7466) );
  NAND2_X1 U9258 ( .A1(n9355), .A2(n8265), .ZN(n7462) );
  NOR2_X1 U9259 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7460), .ZN(n7533) );
  AOI21_X1 U9260 ( .B1(n9346), .B2(n4672), .A(n7533), .ZN(n7461) );
  OAI211_X1 U9261 ( .C1(n7463), .C2(n9327), .A(n7462), .B(n7461), .ZN(n7464)
         );
  AOI21_X1 U9262 ( .B1(n8266), .B2(n9360), .A(n7464), .ZN(n7465) );
  NAND2_X1 U9263 ( .A1(n7466), .A2(n7465), .ZN(P2_U3161) );
  XNOR2_X1 U9264 ( .A(n7579), .B(n8600), .ZN(n7842) );
  XNOR2_X1 U9265 ( .A(n7842), .B(n7843), .ZN(n7471) );
  INV_X1 U9266 ( .A(n7467), .ZN(n7469) );
  NAND2_X1 U9267 ( .A1(n7469), .A2(n7468), .ZN(n7472) );
  NAND2_X1 U9268 ( .A1(n7845), .A2(n9342), .ZN(n7479) );
  AOI21_X1 U9269 ( .B1(n7473), .B2(n7472), .A(n7471), .ZN(n7478) );
  AND2_X1 U9270 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7747) );
  AOI21_X1 U9271 ( .B1(n9354), .B2(n9383), .A(n7747), .ZN(n7475) );
  NAND2_X1 U9272 ( .A1(n9355), .A2(n7578), .ZN(n7474) );
  OAI211_X1 U9273 ( .C1(n9358), .C2(n7892), .A(n7475), .B(n7474), .ZN(n7476)
         );
  AOI21_X1 U9274 ( .B1(n7579), .B2(n9360), .A(n7476), .ZN(n7477) );
  OAI21_X1 U9275 ( .B1(n7479), .B2(n7478), .A(n7477), .ZN(P2_U3171) );
  INV_X1 U9276 ( .A(n7481), .ZN(n7482) );
  NAND2_X1 U9277 ( .A1(n8741), .A2(n7482), .ZN(n7483) );
  AND2_X1 U9278 ( .A1(n7484), .A2(n7483), .ZN(n7494) );
  INV_X1 U9279 ( .A(n7494), .ZN(n10473) );
  INV_X1 U9280 ( .A(n7871), .ZN(n7635) );
  NAND2_X1 U9281 ( .A1(n10473), .A2(n7635), .ZN(n7490) );
  OAI21_X1 U9282 ( .B1(n7486), .B2(n8741), .A(n7485), .ZN(n7488) );
  AOI21_X1 U9283 ( .B1(n7488), .B2(n10427), .A(n7487), .ZN(n7489) );
  AND2_X1 U9284 ( .A1(n7490), .A2(n7489), .ZN(n10474) );
  OAI211_X1 U9285 ( .C1(n6205), .C2(n7492), .A(n10435), .B(n7491), .ZN(n10471)
         );
  INV_X1 U9286 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9965) );
  OAI22_X1 U9287 ( .A1(n10194), .A2(n10471), .B1(n9965), .B2(n10190), .ZN(
        n7496) );
  NOR2_X1 U9288 ( .A1(n10215), .A2(n7493), .ZN(n10444) );
  INV_X1 U9289 ( .A(n10444), .ZN(n7522) );
  OAI22_X1 U9290 ( .A1(n7522), .A2(n7494), .B1(n6205), .B2(n10456), .ZN(n7495)
         );
  AOI211_X1 U9291 ( .C1(P1_REG2_REG_1__SCAN_IN), .C2(n10215), .A(n7496), .B(
        n7495), .ZN(n7497) );
  OAI21_X1 U9292 ( .B1(n10215), .B2(n10474), .A(n7497), .ZN(P1_U3292) );
  INV_X1 U9293 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7504) );
  XNOR2_X1 U9294 ( .A(n7498), .B(n8485), .ZN(n8268) );
  NOR2_X1 U9295 ( .A1(n8268), .A2(n9718), .ZN(n7502) );
  OR2_X1 U9296 ( .A1(n7584), .A2(n8485), .ZN(n7567) );
  NAND2_X1 U9297 ( .A1(n7584), .A2(n8485), .ZN(n7499) );
  NAND3_X1 U9298 ( .A1(n7567), .A2(n9730), .A3(n7499), .ZN(n7501) );
  AOI22_X1 U9299 ( .A1(n4672), .A2(n6257), .B1(n9724), .B2(n9384), .ZN(n7500)
         );
  NAND2_X1 U9300 ( .A1(n7501), .A2(n7500), .ZN(n8264) );
  AOI211_X1 U9301 ( .C1(n9739), .C2(n8266), .A(n7502), .B(n8264), .ZN(n10645)
         );
  OR2_X1 U9302 ( .A1(n10645), .A2(n9743), .ZN(n7503) );
  OAI21_X1 U9303 ( .B1(n9744), .B2(n7504), .A(n7503), .ZN(P2_U3467) );
  NAND2_X1 U9304 ( .A1(n7506), .A2(n8756), .ZN(n7507) );
  NAND2_X1 U9305 ( .A1(n7505), .A2(n7507), .ZN(n10500) );
  OR2_X1 U9306 ( .A1(n10500), .A2(n7871), .ZN(n7513) );
  NAND3_X1 U9307 ( .A1(n7604), .A2(n8653), .A3(n5994), .ZN(n7508) );
  NAND2_X1 U9308 ( .A1(n7621), .A2(n7508), .ZN(n7511) );
  OR2_X1 U9309 ( .A1(n9950), .A2(n9908), .ZN(n7510) );
  NAND2_X1 U9310 ( .A1(n9954), .A2(n9910), .ZN(n7509) );
  NAND2_X1 U9311 ( .A1(n7510), .A2(n7509), .ZN(n7912) );
  AOI21_X1 U9312 ( .B1(n7511), .B2(n10427), .A(n7912), .ZN(n7512) );
  NAND2_X1 U9313 ( .A1(n7513), .A2(n7512), .ZN(n10506) );
  NAND2_X1 U9314 ( .A1(n10506), .A2(n8066), .ZN(n7521) );
  INV_X1 U9315 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7515) );
  INV_X1 U9316 ( .A(n7514), .ZN(n7914) );
  OAI22_X1 U9317 ( .A1(n8066), .A2(n7515), .B1(n7914), .B2(n10190), .ZN(n7519)
         );
  OR2_X1 U9318 ( .A1(n7610), .A2(n10501), .ZN(n7516) );
  NAND2_X1 U9319 ( .A1(n7627), .A2(n7516), .ZN(n10503) );
  NOR2_X1 U9320 ( .A1(n10503), .A2(n7517), .ZN(n7518) );
  AOI211_X1 U9321 ( .C1(n10441), .C2(n7916), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI211_X1 U9322 ( .C1(n10500), .C2(n7522), .A(n7521), .B(n7520), .ZN(
        P1_U3282) );
  INV_X1 U9323 ( .A(n7523), .ZN(n7563) );
  OAI222_X1 U9324 ( .A1(n8546), .A2(n7563), .B1(n8742), .B2(P1_U3086), .C1(
        n7524), .C2(n10338), .ZN(P1_U3334) );
  INV_X1 U9325 ( .A(n7525), .ZN(n7526) );
  NOR2_X2 U9326 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  NOR2_X1 U9327 ( .A1(n10585), .A2(n7528), .ZN(n7529) );
  INV_X1 U9328 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7750) );
  MUX2_X1 U9329 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7750), .S(n7751), .Z(n7531)
         );
  INV_X1 U9330 ( .A(n7753), .ZN(n7530) );
  AOI21_X1 U9331 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7561) );
  INV_X1 U9332 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7547) );
  INV_X1 U9333 ( .A(n7533), .ZN(n7546) );
  INV_X1 U9334 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7534) );
  MUX2_X1 U9335 ( .A(n7535), .B(n7534), .S(n9521), .Z(n7536) );
  NAND2_X1 U9336 ( .A1(n7536), .A2(n10585), .ZN(n7541) );
  XOR2_X1 U9337 ( .A(n10585), .B(n7536), .Z(n10592) );
  OR2_X1 U9338 ( .A1(n7538), .A2(n7537), .ZN(n7540) );
  NAND2_X1 U9339 ( .A1(n7541), .A2(n10590), .ZN(n7543) );
  MUX2_X1 U9340 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9521), .Z(n7742) );
  XNOR2_X1 U9341 ( .A(n7742), .B(n7751), .ZN(n7542) );
  NAND2_X1 U9342 ( .A1(n7542), .A2(n7543), .ZN(n7743) );
  OAI21_X1 U9343 ( .B1(n7543), .B2(n7542), .A(n7743), .ZN(n7544) );
  NAND2_X1 U9344 ( .A1(n10612), .A2(n7544), .ZN(n7545) );
  OAI211_X1 U9345 ( .C1(n10597), .C2(n7547), .A(n7546), .B(n7545), .ZN(n7559)
         );
  INV_X1 U9346 ( .A(n7548), .ZN(n7549) );
  NOR2_X1 U9347 ( .A1(n7534), .A2(n10579), .ZN(n10578) );
  NOR2_X1 U9348 ( .A1(n10585), .A2(n7551), .ZN(n7552) );
  MUX2_X1 U9349 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7504), .S(n7751), .Z(n7555)
         );
  NAND2_X1 U9350 ( .A1(n7556), .A2(n7555), .ZN(n7557) );
  AOI21_X1 U9351 ( .B1(n7738), .B2(n7557), .A(n10606), .ZN(n7558) );
  AOI211_X1 U9352 ( .C1(n10586), .C2(n7751), .A(n7559), .B(n7558), .ZN(n7560)
         );
  OAI21_X1 U9353 ( .B1(n7561), .B2(n10615), .A(n7560), .ZN(P2_U3190) );
  OAI222_X1 U9354 ( .A1(n6970), .A2(P2_U3151), .B1(n8274), .B2(n7563), .C1(
        n7562), .C2(n9798), .ZN(P2_U3274) );
  XNOR2_X1 U9355 ( .A(n7564), .B(n8486), .ZN(n7582) );
  AND2_X1 U9356 ( .A1(n7567), .A2(n7565), .ZN(n7570) );
  NAND2_X1 U9357 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  OAI21_X1 U9358 ( .B1(n7570), .B2(n7569), .A(n7568), .ZN(n7571) );
  AOI222_X1 U9359 ( .A1(n9730), .A2(n7571), .B1(n9382), .B2(n6257), .C1(n9383), 
        .C2(n9724), .ZN(n7576) );
  OAI21_X1 U9360 ( .B1(n9718), .B2(n7582), .A(n7576), .ZN(n7572) );
  INV_X1 U9361 ( .A(n7572), .ZN(n7575) );
  AOI22_X1 U9362 ( .A1(n6261), .A2(n7579), .B1(n10652), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7573) );
  OAI21_X1 U9363 ( .B1(n7575), .B2(n10652), .A(n7573), .ZN(P2_U3417) );
  AOI22_X1 U9364 ( .A1(n9670), .A2(n7579), .B1(n9743), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U9365 ( .B1(n7575), .B2(n9743), .A(n7574), .ZN(P2_U3468) );
  INV_X1 U9366 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7577) );
  MUX2_X1 U9367 ( .A(n7577), .B(n7576), .S(n10629), .Z(n7581) );
  AOI22_X1 U9368 ( .A1(n9651), .A2(n7579), .B1(n10628), .B2(n7578), .ZN(n7580)
         );
  OAI211_X1 U9369 ( .C1(n8900), .C2(n7582), .A(n7581), .B(n7580), .ZN(P2_U3224) );
  OR2_X1 U9370 ( .A1(n7584), .A2(n7583), .ZN(n7586) );
  AND2_X1 U9371 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  XOR2_X1 U9372 ( .A(n8490), .B(n7587), .Z(n7588) );
  OAI222_X1 U9373 ( .A1(n9646), .A2(n8011), .B1(n9644), .B2(n7843), .C1(n9642), 
        .C2(n7588), .ZN(n7662) );
  INV_X1 U9374 ( .A(n7662), .ZN(n7593) );
  XNOR2_X1 U9375 ( .A(n7589), .B(n8490), .ZN(n7663) );
  INV_X1 U9376 ( .A(n7851), .ZN(n7665) );
  AOI22_X1 U9377 ( .A1(n10632), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10628), 
        .B2(n7847), .ZN(n7590) );
  OAI21_X1 U9378 ( .B1(n7665), .B2(n9637), .A(n7590), .ZN(n7591) );
  AOI21_X1 U9379 ( .B1(n7663), .B2(n9657), .A(n7591), .ZN(n7592) );
  OAI21_X1 U9380 ( .B1(n7593), .B2(n10632), .A(n7592), .ZN(P2_U3223) );
  XNOR2_X1 U9381 ( .A(n7594), .B(n8477), .ZN(n7595) );
  OAI222_X1 U9382 ( .A1(n9646), .A2(n8074), .B1(n9644), .B2(n7892), .C1(n9642), 
        .C2(n7595), .ZN(n7781) );
  INV_X1 U9383 ( .A(n7781), .ZN(n7601) );
  OAI21_X1 U9384 ( .B1(n7597), .B2(n8477), .A(n7596), .ZN(n7783) );
  AOI22_X1 U9385 ( .A1(n10632), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10628), 
        .B2(n8071), .ZN(n7598) );
  OAI21_X1 U9386 ( .B1(n7780), .B2(n9637), .A(n7598), .ZN(n7599) );
  AOI21_X1 U9387 ( .B1(n7783), .B2(n9657), .A(n7599), .ZN(n7600) );
  OAI21_X1 U9388 ( .B1(n7601), .B2(n10632), .A(n7600), .ZN(P2_U3222) );
  XNOR2_X1 U9389 ( .A(n7602), .B(n7603), .ZN(n10497) );
  INV_X1 U9390 ( .A(n10497), .ZN(n7617) );
  OAI21_X1 U9391 ( .B1(n8755), .B2(n7605), .A(n7604), .ZN(n7606) );
  NAND2_X1 U9392 ( .A1(n7606), .A2(n10427), .ZN(n7609) );
  OR2_X1 U9393 ( .A1(n7640), .A2(n9887), .ZN(n7608) );
  OR2_X1 U9394 ( .A1(n9952), .A2(n9908), .ZN(n7607) );
  AND2_X1 U9395 ( .A1(n7608), .A2(n7607), .ZN(n7821) );
  NAND2_X1 U9396 ( .A1(n7609), .A2(n7821), .ZN(n10496) );
  INV_X1 U9397 ( .A(n7610), .ZN(n7611) );
  OAI211_X1 U9398 ( .C1(n10494), .C2(n7681), .A(n7611), .B(n10435), .ZN(n10493) );
  AOI22_X1 U9399 ( .A1(n10462), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7824), .B2(
        n10452), .ZN(n7614) );
  NAND2_X1 U9400 ( .A1(n7612), .A2(n10441), .ZN(n7613) );
  OAI211_X1 U9401 ( .C1(n10493), .C2(n10194), .A(n7614), .B(n7613), .ZN(n7615)
         );
  AOI21_X1 U9402 ( .B1(n10496), .B2(n8066), .A(n7615), .ZN(n7616) );
  OAI21_X1 U9403 ( .B1(n7617), .B2(n8158), .A(n7616), .ZN(P1_U3283) );
  AOI21_X1 U9404 ( .B1(n7620), .B2(n7619), .A(n7618), .ZN(n10508) );
  NAND3_X1 U9405 ( .A1(n7621), .A2(n8663), .A3(n8758), .ZN(n7622) );
  NAND2_X1 U9406 ( .A1(n7623), .A2(n7622), .ZN(n7626) );
  OR2_X1 U9407 ( .A1(n9952), .A2(n9887), .ZN(n7625) );
  OR2_X1 U9408 ( .A1(n7868), .A2(n9908), .ZN(n7624) );
  NAND2_X1 U9409 ( .A1(n7625), .A2(n7624), .ZN(n7764) );
  AOI21_X1 U9410 ( .B1(n7626), .B2(n10427), .A(n7764), .ZN(n10510) );
  INV_X1 U9411 ( .A(n10510), .ZN(n7632) );
  INV_X1 U9412 ( .A(n7627), .ZN(n7628) );
  OAI211_X1 U9413 ( .C1(n7628), .C2(n10511), .A(n10435), .B(n10433), .ZN(
        n10509) );
  AOI22_X1 U9414 ( .A1(n10462), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7762), .B2(
        n10452), .ZN(n7630) );
  NAND2_X1 U9415 ( .A1(n7768), .A2(n10441), .ZN(n7629) );
  OAI211_X1 U9416 ( .C1(n10509), .C2(n10194), .A(n7630), .B(n7629), .ZN(n7631)
         );
  AOI21_X1 U9417 ( .B1(n7632), .B2(n8066), .A(n7631), .ZN(n7633) );
  OAI21_X1 U9418 ( .B1(n10508), .B2(n8158), .A(n7633), .ZN(P1_U3281) );
  XNOR2_X1 U9419 ( .A(n10477), .B(n7678), .ZN(n7637) );
  XNOR2_X1 U9420 ( .A(n7634), .B(n7637), .ZN(n10482) );
  NAND2_X1 U9421 ( .A1(n10482), .A2(n7635), .ZN(n7646) );
  NAND2_X1 U9422 ( .A1(n7675), .A2(n7636), .ZN(n7639) );
  INV_X1 U9423 ( .A(n7637), .ZN(n7638) );
  XNOR2_X1 U9424 ( .A(n7639), .B(n7638), .ZN(n7644) );
  OR2_X1 U9425 ( .A1(n7640), .A2(n9908), .ZN(n7643) );
  OR2_X1 U9426 ( .A1(n7641), .A2(n9887), .ZN(n7642) );
  NAND2_X1 U9427 ( .A1(n7643), .A2(n7642), .ZN(n7705) );
  AOI21_X1 U9428 ( .B1(n7644), .B2(n10427), .A(n7705), .ZN(n7645) );
  AND2_X1 U9429 ( .A1(n7646), .A2(n7645), .ZN(n10484) );
  AOI21_X1 U9430 ( .B1(n7647), .B2(n10477), .A(n10502), .ZN(n7648) );
  NAND2_X1 U9431 ( .A1(n7648), .A2(n5118), .ZN(n10478) );
  AOI22_X1 U9432 ( .A1(n10462), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7704), .B2(
        n10452), .ZN(n7650) );
  NAND2_X1 U9433 ( .A1(n10441), .A2(n10477), .ZN(n7649) );
  OAI211_X1 U9434 ( .C1(n10478), .C2(n10194), .A(n7650), .B(n7649), .ZN(n7651)
         );
  AOI21_X1 U9435 ( .B1(n10482), .B2(n10444), .A(n7651), .ZN(n7652) );
  OAI21_X1 U9436 ( .B1(n10484), .B2(n10462), .A(n7652), .ZN(P1_U3285) );
  INV_X1 U9437 ( .A(n7596), .ZN(n7653) );
  OAI21_X1 U9438 ( .B1(n7653), .B2(n8340), .A(n8492), .ZN(n7655) );
  NAND2_X1 U9439 ( .A1(n7655), .A2(n7654), .ZN(n7771) );
  XNOR2_X1 U9440 ( .A(n7656), .B(n8492), .ZN(n7657) );
  OAI222_X1 U9441 ( .A1(n9646), .A2(n8022), .B1(n9644), .B2(n8011), .C1(n7657), 
        .C2(n9642), .ZN(n7772) );
  NAND2_X1 U9442 ( .A1(n7772), .A2(n10629), .ZN(n7661) );
  INV_X1 U9443 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8169) );
  INV_X1 U9444 ( .A(n8019), .ZN(n7658) );
  OAI22_X1 U9445 ( .A1(n10629), .A2(n8169), .B1(n7658), .B2(n8222), .ZN(n7659)
         );
  AOI21_X1 U9446 ( .B1(n8024), .B2(n9651), .A(n7659), .ZN(n7660) );
  OAI211_X1 U9447 ( .C1(n8900), .C2(n7771), .A(n7661), .B(n7660), .ZN(P2_U3221) );
  AOI21_X1 U9448 ( .B1(n9711), .B2(n7663), .A(n7662), .ZN(n7671) );
  INV_X1 U9449 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7664) );
  OAI22_X1 U9450 ( .A1(n7665), .A2(n9789), .B1(n10649), .B2(n7664), .ZN(n7666)
         );
  INV_X1 U9451 ( .A(n7666), .ZN(n7667) );
  OAI21_X1 U9452 ( .B1(n7671), .B2(n10652), .A(n7667), .ZN(P2_U3420) );
  INV_X1 U9453 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7668) );
  NOR2_X1 U9454 ( .A1(n9744), .A2(n7668), .ZN(n7669) );
  AOI21_X1 U9455 ( .B1(n9670), .B2(n7851), .A(n7669), .ZN(n7670) );
  OAI21_X1 U9456 ( .B1(n7671), .B2(n9743), .A(n7670), .ZN(P2_U3469) );
  XNOR2_X1 U9457 ( .A(n7672), .B(n7677), .ZN(n10491) );
  INV_X1 U9458 ( .A(n10491), .ZN(n7689) );
  INV_X1 U9459 ( .A(n7673), .ZN(n7795) );
  INV_X1 U9460 ( .A(n7674), .ZN(n8645) );
  AOI21_X1 U9461 ( .B1(n7675), .B2(n8646), .A(n8645), .ZN(n7676) );
  XOR2_X1 U9462 ( .A(n7677), .B(n7676), .Z(n7679) );
  NOR2_X1 U9463 ( .A1(n7678), .A2(n9887), .ZN(n7791) );
  AOI21_X1 U9464 ( .B1(n7679), .B2(n10427), .A(n7791), .ZN(n10488) );
  OAI21_X1 U9465 ( .B1(n7795), .B2(n10190), .A(n10488), .ZN(n7687) );
  NAND2_X1 U9466 ( .A1(n5118), .A2(n10486), .ZN(n7680) );
  NAND2_X1 U9467 ( .A1(n7680), .A2(n10435), .ZN(n7682) );
  OR2_X1 U9468 ( .A1(n7682), .A2(n7681), .ZN(n7684) );
  AND2_X1 U9469 ( .A1(n9954), .A2(n9865), .ZN(n7792) );
  INV_X1 U9470 ( .A(n7792), .ZN(n7683) );
  AND2_X1 U9471 ( .A1(n7684), .A2(n7683), .ZN(n10487) );
  AOI22_X1 U9472 ( .A1(n10441), .A2(n10486), .B1(P1_REG2_REG_9__SCAN_IN), .B2(
        n10462), .ZN(n7685) );
  OAI21_X1 U9473 ( .B1(n10487), .B2(n10194), .A(n7685), .ZN(n7686) );
  AOI21_X1 U9474 ( .B1(n7687), .B2(n8066), .A(n7686), .ZN(n7688) );
  OAI21_X1 U9475 ( .B1(n7689), .B2(n8158), .A(n7688), .ZN(P1_U3284) );
  INV_X1 U9476 ( .A(n7690), .ZN(n7694) );
  AOI22_X1 U9477 ( .A1(n10441), .A2(n7692), .B1(n10452), .B2(n7691), .ZN(n7693) );
  OAI21_X1 U9478 ( .B1(n7694), .B2(n10194), .A(n7693), .ZN(n7697) );
  MUX2_X1 U9479 ( .A(n7695), .B(P1_REG2_REG_5__SCAN_IN), .S(n10215), .Z(n7696)
         );
  AOI211_X1 U9480 ( .C1(n10458), .C2(n7698), .A(n7697), .B(n7696), .ZN(n7699)
         );
  INV_X1 U9481 ( .A(n7699), .ZN(P1_U3288) );
  XNOR2_X1 U9482 ( .A(n7700), .B(n7701), .ZN(n7702) );
  NAND2_X1 U9483 ( .A1(n7702), .A2(n7703), .ZN(n7785) );
  OAI21_X1 U9484 ( .B1(n7703), .B2(n7702), .A(n7785), .ZN(n7710) );
  INV_X1 U9485 ( .A(n7704), .ZN(n7708) );
  AOI22_X1 U9486 ( .A1(n9916), .A2(n7705), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7707) );
  NAND2_X1 U9487 ( .A1(n10421), .A2(n10477), .ZN(n7706) );
  OAI211_X1 U9488 ( .C1(n10423), .C2(n7708), .A(n7707), .B(n7706), .ZN(n7709)
         );
  AOI21_X1 U9489 ( .B1(n7710), .B2(n9922), .A(n7709), .ZN(n7711) );
  INV_X1 U9490 ( .A(n7711), .ZN(P1_U3221) );
  NAND2_X1 U9491 ( .A1(n7713), .A2(n7712), .ZN(n7715) );
  NAND2_X1 U9492 ( .A1(n7715), .A2(n7714), .ZN(n7801) );
  INV_X1 U9493 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U9494 ( .A1(n7717), .A2(n7716), .ZN(n7718) );
  OAI21_X1 U9495 ( .B1(n7717), .B2(n7716), .A(n7718), .ZN(n7800) );
  NOR2_X1 U9496 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  INV_X1 U9497 ( .A(n7718), .ZN(n7719) );
  NOR2_X1 U9498 ( .A1(n7799), .A2(n7719), .ZN(n7721) );
  XNOR2_X1 U9499 ( .A(n7937), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7720) );
  NOR2_X1 U9500 ( .A1(n7721), .A2(n7720), .ZN(n7940) );
  AOI21_X1 U9501 ( .B1(n7721), .B2(n7720), .A(n7940), .ZN(n7736) );
  OR2_X1 U9502 ( .A1(n7937), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U9503 ( .A1(n7937), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7722) );
  AND2_X1 U9504 ( .A1(n7943), .A2(n7722), .ZN(n7730) );
  NOR2_X1 U9505 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  NOR2_X1 U9506 ( .A1(n7726), .A2(n7725), .ZN(n7805) );
  NAND2_X1 U9507 ( .A1(n7808), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7728) );
  OR2_X1 U9508 ( .A1(n7808), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U9509 ( .A1(n7728), .A2(n7727), .ZN(n7804) );
  OR2_X1 U9510 ( .A1(n7805), .A2(n7804), .ZN(n7802) );
  NAND2_X1 U9511 ( .A1(n7729), .A2(n7730), .ZN(n7944) );
  OAI21_X1 U9512 ( .B1(n7730), .B2(n7729), .A(n7944), .ZN(n7731) );
  NAND2_X1 U9513 ( .A1(n7731), .A2(n10025), .ZN(n7735) );
  NOR2_X1 U9514 ( .A1(n9272), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9853) );
  NOR2_X1 U9515 ( .A1(n10007), .A2(n7732), .ZN(n7733) );
  AOI211_X1 U9516 ( .C1(n10021), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9853), .B(
        n7733), .ZN(n7734) );
  OAI211_X1 U9517 ( .C1(n7736), .C2(n8109), .A(n7735), .B(n7734), .ZN(P1_U3260) );
  OR2_X1 U9518 ( .A1(n7751), .A2(n7504), .ZN(n7737) );
  INV_X1 U9519 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7739) );
  AOI21_X1 U9520 ( .B1(n7740), .B2(n7739), .A(n7986), .ZN(n7759) );
  INV_X1 U9521 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10372) );
  MUX2_X1 U9522 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9521), .Z(n7978) );
  XNOR2_X1 U9523 ( .A(n7978), .B(n7985), .ZN(n7746) );
  OR2_X1 U9524 ( .A1(n7742), .A2(n7741), .ZN(n7744) );
  OAI21_X1 U9525 ( .B1(n7746), .B2(n7745), .A(n7976), .ZN(n7748) );
  AOI21_X1 U9526 ( .B1(n10612), .B2(n7748), .A(n7747), .ZN(n7749) );
  OAI21_X1 U9527 ( .B1(n10597), .B2(n10372), .A(n7749), .ZN(n7757) );
  OR2_X1 U9528 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  AOI21_X1 U9529 ( .B1(n7577), .B2(n7754), .A(n7969), .ZN(n7755) );
  NOR2_X1 U9530 ( .A1(n7755), .A2(n10615), .ZN(n7756) );
  AOI211_X1 U9531 ( .C1(n10586), .C2(n7985), .A(n7757), .B(n7756), .ZN(n7758)
         );
  OAI21_X1 U9532 ( .B1(n7759), .B2(n10606), .A(n7758), .ZN(P2_U3191) );
  XOR2_X1 U9533 ( .A(n7760), .B(n7761), .Z(n7770) );
  INV_X1 U9534 ( .A(n7762), .ZN(n7766) );
  AOI21_X1 U9535 ( .B1(n9916), .B2(n7764), .A(n7763), .ZN(n7765) );
  OAI21_X1 U9536 ( .B1(n10423), .B2(n7766), .A(n7765), .ZN(n7767) );
  AOI21_X1 U9537 ( .B1(n7768), .B2(n10421), .A(n7767), .ZN(n7769) );
  OAI21_X1 U9538 ( .B1(n7770), .B2(n10416), .A(n7769), .ZN(P1_U3224) );
  NOR2_X1 U9539 ( .A1(n7771), .A2(n9718), .ZN(n7773) );
  AOI211_X1 U9540 ( .C1(n9739), .C2(n8024), .A(n7773), .B(n7772), .ZN(n10650)
         );
  NAND2_X1 U9541 ( .A1(n9743), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7774) );
  OAI21_X1 U9542 ( .B1(n10650), .B2(n9743), .A(n7774), .ZN(P2_U3471) );
  NAND2_X1 U9543 ( .A1(n7778), .A2(n7775), .ZN(n7776) );
  OAI211_X1 U9544 ( .C1(n7777), .C2(n9798), .A(n7776), .B(n8526), .ZN(P2_U3272) );
  NAND2_X1 U9545 ( .A1(n7778), .A2(n10343), .ZN(n7779) );
  OAI211_X1 U9546 ( .C1(n9285), .C2(n10338), .A(n7779), .B(n8879), .ZN(
        P1_U3332) );
  INV_X1 U9547 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8119) );
  NOR2_X1 U9548 ( .A1(n7780), .A2(n9716), .ZN(n7782) );
  AOI211_X1 U9549 ( .C1(n9711), .C2(n7783), .A(n7782), .B(n7781), .ZN(n10647)
         );
  OR2_X1 U9550 ( .A1(n10647), .A2(n9743), .ZN(n7784) );
  OAI21_X1 U9551 ( .B1(n9744), .B2(n8119), .A(n7784), .ZN(P2_U3470) );
  OAI21_X1 U9552 ( .B1(n7786), .B2(n7700), .A(n7785), .ZN(n7790) );
  XNOR2_X1 U9553 ( .A(n7788), .B(n7787), .ZN(n7789) );
  XNOR2_X1 U9554 ( .A(n7790), .B(n7789), .ZN(n7798) );
  OAI21_X1 U9555 ( .B1(n7792), .B2(n7791), .A(n9916), .ZN(n7793) );
  OAI211_X1 U9556 ( .C1(n10423), .C2(n7795), .A(n7794), .B(n7793), .ZN(n7796)
         );
  AOI21_X1 U9557 ( .B1(n10486), .B2(n10421), .A(n7796), .ZN(n7797) );
  OAI21_X1 U9558 ( .B1(n7798), .B2(n10416), .A(n7797), .ZN(P1_U3231) );
  AOI21_X1 U9559 ( .B1(n7801), .B2(n7800), .A(n7799), .ZN(n7811) );
  AND2_X1 U9560 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7807) );
  INV_X1 U9561 ( .A(n7802), .ZN(n7803) );
  AOI211_X1 U9562 ( .C1(n7805), .C2(n7804), .A(n7803), .B(n7948), .ZN(n7806)
         );
  AOI211_X1 U9563 ( .C1(n10021), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n7807), .B(
        n7806), .ZN(n7810) );
  NAND2_X1 U9564 ( .A1(n10022), .A2(n7808), .ZN(n7809) );
  OAI211_X1 U9565 ( .C1(n7811), .C2(n8109), .A(n7810), .B(n7809), .ZN(P1_U3259) );
  INV_X1 U9566 ( .A(n7812), .ZN(n7815) );
  OAI222_X1 U9567 ( .A1(n8891), .A2(n7813), .B1(n8546), .B2(n7815), .C1(
        P1_U3086), .C2(n6265), .ZN(P1_U3333) );
  OAI222_X1 U9568 ( .A1(P2_U3151), .A2(n7816), .B1(n9801), .B2(n7815), .C1(
        n7814), .C2(n9798), .ZN(P2_U3273) );
  XNOR2_X1 U9569 ( .A(n7817), .B(n7907), .ZN(n7819) );
  NOR2_X1 U9570 ( .A1(n7819), .A2(n7818), .ZN(n7906) );
  AOI21_X1 U9571 ( .B1(n7819), .B2(n7818), .A(n7906), .ZN(n7826) );
  OAI22_X1 U9572 ( .A1(n10413), .A2(n7821), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7820), .ZN(n7823) );
  NOR2_X1 U9573 ( .A1(n10494), .A2(n9931), .ZN(n7822) );
  AOI211_X1 U9574 ( .C1(n7824), .C2(n9927), .A(n7823), .B(n7822), .ZN(n7825)
         );
  OAI21_X1 U9575 ( .B1(n7826), .B2(n10416), .A(n7825), .ZN(P1_U3217) );
  NAND2_X1 U9576 ( .A1(n4827), .A2(n8348), .ZN(n8493) );
  XNOR2_X1 U9577 ( .A(n7827), .B(n8493), .ZN(n7880) );
  XOR2_X1 U9578 ( .A(n7828), .B(n8493), .Z(n7829) );
  OAI222_X1 U9579 ( .A1(n9646), .A2(n8236), .B1(n9644), .B2(n8074), .C1(n9642), 
        .C2(n7829), .ZN(n7881) );
  INV_X1 U9580 ( .A(n8349), .ZN(n7831) );
  INV_X1 U9581 ( .A(n7900), .ZN(n7830) );
  OAI22_X1 U9582 ( .A1(n7831), .A2(n10622), .B1(n7830), .B2(n8222), .ZN(n7832)
         );
  OAI21_X1 U9583 ( .B1(n7881), .B2(n7832), .A(n10629), .ZN(n7834) );
  NAND2_X1 U9584 ( .A1(n10632), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7833) );
  OAI211_X1 U9585 ( .C1(n8900), .C2(n7880), .A(n7834), .B(n7833), .ZN(P2_U3220) );
  XOR2_X1 U9586 ( .A(n7835), .B(n7836), .Z(n7841) );
  INV_X1 U9587 ( .A(n10429), .ZN(n7838) );
  OAI22_X1 U9588 ( .A1(n7856), .A2(n9908), .B1(n9950), .B2(n9887), .ZN(n10426)
         );
  AOI22_X1 U9589 ( .A1(n9916), .A2(n10426), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n7837) );
  OAI21_X1 U9590 ( .B1(n10423), .B2(n7838), .A(n7837), .ZN(n7839) );
  AOI21_X1 U9591 ( .B1(n10432), .B2(n10421), .A(n7839), .ZN(n7840) );
  OAI21_X1 U9592 ( .B1(n7841), .B2(n10416), .A(n7840), .ZN(P1_U3234) );
  XNOR2_X1 U9593 ( .A(n7851), .B(n8600), .ZN(n7891) );
  XNOR2_X1 U9594 ( .A(n8010), .B(n9382), .ZN(n7846) );
  NOR2_X1 U9595 ( .A1(n7846), .A2(n7891), .ZN(n8076) );
  AOI21_X1 U9596 ( .B1(n7891), .B2(n7846), .A(n8076), .ZN(n7853) );
  INV_X1 U9597 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8962) );
  NOR2_X1 U9598 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8962), .ZN(n7980) );
  AOI21_X1 U9599 ( .B1(n9354), .B2(n4672), .A(n7980), .ZN(n7849) );
  NAND2_X1 U9600 ( .A1(n9355), .A2(n7847), .ZN(n7848) );
  OAI211_X1 U9601 ( .C1(n9358), .C2(n8011), .A(n7849), .B(n7848), .ZN(n7850)
         );
  AOI21_X1 U9602 ( .B1(n7851), .B2(n9360), .A(n7850), .ZN(n7852) );
  OAI21_X1 U9603 ( .B1(n7853), .B2(n9363), .A(n7852), .ZN(P2_U3157) );
  XNOR2_X1 U9604 ( .A(n7854), .B(n8762), .ZN(n10285) );
  XNOR2_X1 U9605 ( .A(n7855), .B(n8762), .ZN(n7858) );
  NOR2_X1 U9606 ( .A1(n7856), .A2(n9887), .ZN(n7857) );
  AOI21_X1 U9607 ( .B1(n9946), .B2(n9865), .A(n7857), .ZN(n9925) );
  OAI21_X1 U9608 ( .B1(n7858), .B2(n10203), .A(n9925), .ZN(n10279) );
  INV_X1 U9609 ( .A(n5126), .ZN(n7859) );
  AOI211_X1 U9610 ( .C1(n10281), .C2(n7873), .A(n10502), .B(n7859), .ZN(n10280) );
  NAND2_X1 U9611 ( .A1(n10280), .A2(n10450), .ZN(n7862) );
  INV_X1 U9612 ( .A(n7860), .ZN(n9928) );
  AOI22_X1 U9613 ( .A1(n10462), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9928), .B2(
        n10452), .ZN(n7861) );
  OAI211_X1 U9614 ( .C1(n6032), .C2(n10456), .A(n7862), .B(n7861), .ZN(n7863)
         );
  AOI21_X1 U9615 ( .B1(n10279), .B2(n8066), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9616 ( .B1(n10285), .B2(n8158), .A(n7864), .ZN(P1_U3278) );
  XNOR2_X1 U9617 ( .A(n7865), .B(n8760), .ZN(n7872) );
  OAI21_X1 U9618 ( .B1(n8760), .B2(n7867), .A(n7866), .ZN(n7869) );
  OAI22_X1 U9619 ( .A1(n8675), .A2(n9908), .B1(n7868), .B2(n9887), .ZN(n8040)
         );
  AOI21_X1 U9620 ( .B1(n7869), .B2(n10427), .A(n8040), .ZN(n7870) );
  OAI21_X1 U9621 ( .B1(n7872), .B2(n7871), .A(n7870), .ZN(n7961) );
  INV_X1 U9622 ( .A(n7961), .ZN(n7879) );
  INV_X1 U9623 ( .A(n7872), .ZN(n7963) );
  OAI211_X1 U9624 ( .C1(n8044), .C2(n10434), .A(n7873), .B(n10435), .ZN(n7960)
         );
  AOI22_X1 U9625 ( .A1(n10462), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8041), .B2(
        n10452), .ZN(n7876) );
  NAND2_X1 U9626 ( .A1(n7874), .A2(n10441), .ZN(n7875) );
  OAI211_X1 U9627 ( .C1(n7960), .C2(n10194), .A(n7876), .B(n7875), .ZN(n7877)
         );
  AOI21_X1 U9628 ( .B1(n7963), .B2(n10444), .A(n7877), .ZN(n7878) );
  OAI21_X1 U9629 ( .B1(n7879), .B2(n10462), .A(n7878), .ZN(P1_U3279) );
  NOR2_X1 U9630 ( .A1(n7880), .A2(n9718), .ZN(n7882) );
  AOI211_X1 U9631 ( .C1(n9739), .C2(n8349), .A(n7882), .B(n7881), .ZN(n10408)
         );
  NAND2_X1 U9632 ( .A1(n9743), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7883) );
  OAI21_X1 U9633 ( .B1(n10408), .B2(n9743), .A(n7883), .ZN(P2_U3472) );
  INV_X1 U9634 ( .A(n6094), .ZN(n7887) );
  OAI222_X1 U9635 ( .A1(n8546), .A2(n7887), .B1(P1_U3086), .B2(n7885), .C1(
        n7884), .C2(n10338), .ZN(P1_U3331) );
  OAI222_X1 U9636 ( .A1(n5735), .A2(P2_U3151), .B1(n9801), .B2(n7887), .C1(
        n7886), .C2(n9798), .ZN(P2_U3271) );
  XNOR2_X1 U9637 ( .A(n8082), .B(n8244), .ZN(n8012) );
  NOR2_X1 U9638 ( .A1(n8012), .A2(n8011), .ZN(n8013) );
  INV_X1 U9639 ( .A(n8013), .ZN(n7889) );
  NAND2_X1 U9640 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  INV_X1 U9641 ( .A(n7891), .ZN(n7893) );
  AND2_X1 U9642 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  INV_X1 U9643 ( .A(n7894), .ZN(n7896) );
  XNOR2_X1 U9644 ( .A(n8024), .B(n8244), .ZN(n7897) );
  NAND2_X1 U9645 ( .A1(n7897), .A2(n8074), .ZN(n8014) );
  OAI21_X1 U9646 ( .B1(n7894), .B2(n8011), .A(n8012), .ZN(n7895) );
  OAI211_X1 U9647 ( .C1(n9381), .C2(n7896), .A(n8014), .B(n7895), .ZN(n7899)
         );
  INV_X1 U9648 ( .A(n7897), .ZN(n7898) );
  NAND2_X1 U9649 ( .A1(n7898), .A2(n9380), .ZN(n8015) );
  XNOR2_X1 U9650 ( .A(n8349), .B(n8600), .ZN(n8027) );
  XNOR2_X1 U9651 ( .A(n8027), .B(n9379), .ZN(n8028) );
  XOR2_X1 U9652 ( .A(n8029), .B(n8028), .Z(n7905) );
  AOI22_X1 U9653 ( .A1(n9346), .A2(n9378), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n7902) );
  NAND2_X1 U9654 ( .A1(n9355), .A2(n7900), .ZN(n7901) );
  OAI211_X1 U9655 ( .C1(n8074), .C2(n9327), .A(n7902), .B(n7901), .ZN(n7903)
         );
  AOI21_X1 U9656 ( .B1(n8349), .B2(n9360), .A(n7903), .ZN(n7904) );
  OAI21_X1 U9657 ( .B1(n7905), .B2(n9363), .A(n7904), .ZN(P2_U3174) );
  AOI21_X1 U9658 ( .B1(n7907), .B2(n7817), .A(n7906), .ZN(n7911) );
  XNOR2_X1 U9659 ( .A(n7909), .B(n7908), .ZN(n7910) );
  XNOR2_X1 U9660 ( .A(n7911), .B(n7910), .ZN(n7918) );
  AOI22_X1 U9661 ( .A1(n9916), .A2(n7912), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7913) );
  OAI21_X1 U9662 ( .B1(n10423), .B2(n7914), .A(n7913), .ZN(n7915) );
  AOI21_X1 U9663 ( .B1(n7916), .B2(n10421), .A(n7915), .ZN(n7917) );
  OAI21_X1 U9664 ( .B1(n7918), .B2(n10416), .A(n7917), .ZN(P1_U3236) );
  XNOR2_X1 U9665 ( .A(n9717), .B(n8240), .ZN(n8497) );
  XNOR2_X1 U9666 ( .A(n7919), .B(n8497), .ZN(n9719) );
  INV_X1 U9667 ( .A(n8497), .ZN(n8355) );
  XNOR2_X1 U9668 ( .A(n7920), .B(n8355), .ZN(n7921) );
  NAND2_X1 U9669 ( .A1(n7921), .A2(n9730), .ZN(n7924) );
  OAI22_X1 U9670 ( .A1(n8563), .A2(n9646), .B1(n8236), .B2(n9644), .ZN(n7922)
         );
  INV_X1 U9671 ( .A(n7922), .ZN(n7923) );
  NAND2_X1 U9672 ( .A1(n7924), .A2(n7923), .ZN(n9721) );
  NAND2_X1 U9673 ( .A1(n9721), .A2(n10629), .ZN(n7929) );
  INV_X1 U9674 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9424) );
  INV_X1 U9675 ( .A(n8565), .ZN(n7925) );
  OAI22_X1 U9676 ( .A1(n10629), .A2(n9424), .B1(n7925), .B2(n8222), .ZN(n7926)
         );
  AOI21_X1 U9677 ( .B1(n7927), .B2(n9651), .A(n7926), .ZN(n7928) );
  OAI211_X1 U9678 ( .C1(n8900), .C2(n9719), .A(n7929), .B(n7928), .ZN(P2_U3218) );
  INV_X1 U9679 ( .A(n8034), .ZN(n8007) );
  NOR2_X1 U9680 ( .A1(n8007), .A2(n10622), .ZN(n7933) );
  OAI211_X1 U9681 ( .C1(n4606), .C2(n4671), .A(n9730), .B(n7930), .ZN(n7932)
         );
  NAND2_X1 U9682 ( .A1(n8240), .A2(n6257), .ZN(n7931) );
  OAI211_X1 U9683 ( .C1(n8022), .C2(n9644), .A(n7932), .B(n7931), .ZN(n8000)
         );
  AOI211_X1 U9684 ( .C1(n10628), .C2(n8030), .A(n7933), .B(n8000), .ZN(n7936)
         );
  XNOR2_X1 U9685 ( .A(n7934), .B(n8495), .ZN(n8001) );
  AOI22_X1 U9686 ( .A1(n8001), .A2(n9657), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10632), .ZN(n7935) );
  OAI21_X1 U9687 ( .B1(n7936), .B2(n10632), .A(n7935), .ZN(P2_U3219) );
  NOR2_X1 U9688 ( .A1(n7937), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7939) );
  XNOR2_X1 U9689 ( .A(n8106), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n7938) );
  NOR3_X1 U9690 ( .A1(n7940), .A2(n7939), .A3(n7938), .ZN(n8105) );
  INV_X1 U9691 ( .A(n8105), .ZN(n7942) );
  OAI21_X1 U9692 ( .B1(n7940), .B2(n7939), .A(n7938), .ZN(n7941) );
  NAND3_X1 U9693 ( .A1(n7942), .A2(n10033), .A3(n7941), .ZN(n7954) );
  AND2_X1 U9694 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9695 ( .A1(n7944), .A2(n7943), .ZN(n7950) );
  NAND2_X1 U9696 ( .A1(n7955), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7947) );
  INV_X1 U9697 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U9698 ( .A1(n8106), .A2(n7945), .ZN(n7946) );
  AND2_X1 U9699 ( .A1(n7947), .A2(n7946), .ZN(n7949) );
  NOR2_X1 U9700 ( .A1(n7950), .A2(n7949), .ZN(n8102) );
  AOI211_X1 U9701 ( .C1(n7950), .C2(n7949), .A(n8102), .B(n7948), .ZN(n7951)
         );
  AOI211_X1 U9702 ( .C1(n10021), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n7952), .B(
        n7951), .ZN(n7953) );
  OAI211_X1 U9703 ( .C1(n10007), .C2(n7955), .A(n7954), .B(n7953), .ZN(
        P1_U3261) );
  INV_X1 U9704 ( .A(n7956), .ZN(n8008) );
  INV_X1 U9705 ( .A(n7957), .ZN(n7959) );
  OAI222_X1 U9706 ( .A1(n8546), .A2(n8008), .B1(P1_U3086), .B2(n7959), .C1(
        n7958), .C2(n10338), .ZN(P1_U3330) );
  OAI21_X1 U9707 ( .B1(n8044), .B2(n10517), .A(n7960), .ZN(n7962) );
  AOI211_X1 U9708 ( .C1(n10481), .C2(n7963), .A(n7962), .B(n7961), .ZN(n7966)
         );
  NAND2_X1 U9709 ( .A1(n10534), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7964) );
  OAI21_X1 U9710 ( .B1(n7966), .B2(n10534), .A(n7964), .ZN(P1_U3536) );
  NAND2_X1 U9711 ( .A1(n6596), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7965) );
  OAI21_X1 U9712 ( .B1(n7966), .B2(n6596), .A(n7965), .ZN(P1_U3495) );
  NOR2_X1 U9713 ( .A1(n7985), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U9714 ( .A1(n7988), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8131) );
  INV_X1 U9715 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U9716 ( .A1(n7997), .A2(n7971), .ZN(n7972) );
  NAND2_X1 U9717 ( .A1(n8131), .A2(n7972), .ZN(n7974) );
  INV_X1 U9718 ( .A(n8132), .ZN(n7973) );
  AOI21_X1 U9719 ( .B1(n7975), .B2(n7974), .A(n7973), .ZN(n7999) );
  INV_X1 U9720 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10375) );
  MUX2_X1 U9721 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9521), .Z(n8121) );
  NAND2_X1 U9722 ( .A1(n7979), .A2(n7997), .ZN(n8124) );
  OAI21_X1 U9723 ( .B1(n7997), .B2(n7979), .A(n8124), .ZN(n7981) );
  AOI21_X1 U9724 ( .B1(n10612), .B2(n7981), .A(n7980), .ZN(n7982) );
  OAI21_X1 U9725 ( .B1(n10597), .B2(n10375), .A(n7982), .ZN(n7996) );
  INV_X1 U9726 ( .A(n7983), .ZN(n7984) );
  NOR2_X1 U9727 ( .A1(n7985), .A2(n7984), .ZN(n7987) );
  NAND2_X1 U9728 ( .A1(n7988), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U9729 ( .A1(n7997), .A2(n7668), .ZN(n7989) );
  NAND2_X1 U9730 ( .A1(n8117), .A2(n7989), .ZN(n7992) );
  NAND2_X1 U9731 ( .A1(n7993), .A2(n7992), .ZN(n7994) );
  AOI21_X1 U9732 ( .B1(n8118), .B2(n7994), .A(n10606), .ZN(n7995) );
  AOI211_X1 U9733 ( .C1(n10586), .C2(n7997), .A(n7996), .B(n7995), .ZN(n7998)
         );
  OAI21_X1 U9734 ( .B1(n7999), .B2(n10615), .A(n7998), .ZN(P2_U3192) );
  INV_X1 U9735 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8002) );
  AOI21_X1 U9736 ( .B1(n8001), .B2(n9711), .A(n8000), .ZN(n8004) );
  MUX2_X1 U9737 ( .A(n8002), .B(n8004), .S(n9744), .Z(n8003) );
  OAI21_X1 U9738 ( .B1(n8007), .B2(n9715), .A(n8003), .ZN(P2_U3473) );
  INV_X1 U9739 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8005) );
  MUX2_X1 U9740 ( .A(n8005), .B(n8004), .S(n10649), .Z(n8006) );
  OAI21_X1 U9741 ( .B1(n8007), .B2(n9789), .A(n8006), .ZN(P2_U3432) );
  OAI222_X1 U9742 ( .A1(n8009), .A2(P2_U3151), .B1(n8274), .B2(n8008), .C1(
        n8964), .C2(n9798), .ZN(P2_U3270) );
  NOR2_X1 U9743 ( .A1(n8010), .A2(n9382), .ZN(n8075) );
  XNOR2_X1 U9744 ( .A(n8012), .B(n8011), .ZN(n8079) );
  NOR3_X1 U9745 ( .A1(n8076), .A2(n8075), .A3(n8079), .ZN(n8077) );
  NOR2_X1 U9746 ( .A1(n8077), .A2(n8013), .ZN(n8017) );
  NAND2_X1 U9747 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  XNOR2_X1 U9748 ( .A(n8017), .B(n8016), .ZN(n8026) );
  INV_X1 U9749 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8018) );
  NOR2_X1 U9750 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8018), .ZN(n8182) );
  AOI21_X1 U9751 ( .B1(n9354), .B2(n9381), .A(n8182), .ZN(n8021) );
  NAND2_X1 U9752 ( .A1(n9355), .A2(n8019), .ZN(n8020) );
  OAI211_X1 U9753 ( .C1(n9358), .C2(n8022), .A(n8021), .B(n8020), .ZN(n8023)
         );
  AOI21_X1 U9754 ( .B1(n8024), .B2(n9360), .A(n8023), .ZN(n8025) );
  OAI21_X1 U9755 ( .B1(n8026), .B2(n9363), .A(n8025), .ZN(P2_U3164) );
  XNOR2_X1 U9756 ( .A(n8034), .B(n8600), .ZN(n8234) );
  XNOR2_X1 U9757 ( .A(n8234), .B(n8236), .ZN(n8237) );
  XOR2_X1 U9758 ( .A(n8238), .B(n8237), .Z(n8036) );
  AOI22_X1 U9759 ( .A1(n9354), .A2(n9379), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8032) );
  NAND2_X1 U9760 ( .A1(n9355), .A2(n8030), .ZN(n8031) );
  OAI211_X1 U9761 ( .C1(n8554), .C2(n9358), .A(n8032), .B(n8031), .ZN(n8033)
         );
  AOI21_X1 U9762 ( .B1(n8034), .B2(n9360), .A(n8033), .ZN(n8035) );
  OAI21_X1 U9763 ( .B1(n8036), .B2(n9363), .A(n8035), .ZN(P2_U3155) );
  OAI21_X1 U9764 ( .B1(n8039), .B2(n8037), .A(n8038), .ZN(n8046) );
  AOI22_X1 U9765 ( .A1(n9916), .A2(n8040), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8043) );
  NAND2_X1 U9766 ( .A1(n9927), .A2(n8041), .ZN(n8042) );
  OAI211_X1 U9767 ( .C1(n8044), .C2(n9931), .A(n8043), .B(n8042), .ZN(n8045)
         );
  AOI21_X1 U9768 ( .B1(n8046), .B2(n9922), .A(n8045), .ZN(n8047) );
  INV_X1 U9769 ( .A(n8047), .ZN(P1_U3215) );
  XNOR2_X1 U9770 ( .A(n8048), .B(n8496), .ZN(n8049) );
  OAI222_X1 U9771 ( .A1(n9644), .A2(n8554), .B1(n9646), .B2(n8259), .C1(n8049), 
        .C2(n9642), .ZN(n8193) );
  INV_X1 U9772 ( .A(n8193), .ZN(n8054) );
  XOR2_X1 U9773 ( .A(n8050), .B(n8496), .Z(n8194) );
  AOI22_X1 U9774 ( .A1(n10632), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10628), 
        .B2(n8551), .ZN(n8051) );
  OAI21_X1 U9775 ( .B1(n8200), .B2(n9637), .A(n8051), .ZN(n8052) );
  AOI21_X1 U9776 ( .B1(n8194), .B2(n9657), .A(n8052), .ZN(n8053) );
  OAI21_X1 U9777 ( .B1(n8054), .B2(n10632), .A(n8053), .ZN(P2_U3217) );
  INV_X1 U9778 ( .A(n8055), .ZN(n8069) );
  OAI222_X1 U9779 ( .A1(n8546), .A2(n8069), .B1(P1_U3086), .B2(n8056), .C1(
        n9258), .C2(n8891), .ZN(P1_U3329) );
  XOR2_X1 U9780 ( .A(n8057), .B(n8763), .Z(n8096) );
  INV_X1 U9781 ( .A(n8096), .ZN(n8068) );
  INV_X1 U9782 ( .A(n8151), .ZN(n8058) );
  AOI21_X1 U9783 ( .B1(n8763), .B2(n8059), .A(n8058), .ZN(n8061) );
  OAI22_X1 U9784 ( .A1(n8205), .A2(n9908), .B1(n8675), .B2(n9887), .ZN(n9844)
         );
  INV_X1 U9785 ( .A(n9844), .ZN(n8060) );
  OAI21_X1 U9786 ( .B1(n8061), .B2(n10203), .A(n8060), .ZN(n8094) );
  INV_X1 U9787 ( .A(n9848), .ZN(n8064) );
  AOI211_X1 U9788 ( .C1(n9848), .C2(n5126), .A(n10502), .B(n8145), .ZN(n8095)
         );
  NAND2_X1 U9789 ( .A1(n8095), .A2(n10450), .ZN(n8063) );
  AOI22_X1 U9790 ( .A1(n10462), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9843), .B2(
        n10452), .ZN(n8062) );
  OAI211_X1 U9791 ( .C1(n8064), .C2(n10456), .A(n8063), .B(n8062), .ZN(n8065)
         );
  AOI21_X1 U9792 ( .B1(n8094), .B2(n8066), .A(n8065), .ZN(n8067) );
  OAI21_X1 U9793 ( .B1(n8068), .B2(n8158), .A(n8067), .ZN(P1_U3277) );
  OAI222_X1 U9794 ( .A1(n8070), .A2(P2_U3151), .B1(n9801), .B2(n8069), .C1(
        n9061), .C2(n9798), .ZN(P2_U3269) );
  AND2_X1 U9795 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8128) );
  AOI21_X1 U9796 ( .B1(n9354), .B2(n9382), .A(n8128), .ZN(n8073) );
  NAND2_X1 U9797 ( .A1(n9355), .A2(n8071), .ZN(n8072) );
  OAI211_X1 U9798 ( .C1(n9358), .C2(n8074), .A(n8073), .B(n8072), .ZN(n8081)
         );
  OR2_X1 U9799 ( .A1(n8076), .A2(n8075), .ZN(n8078) );
  AOI211_X1 U9800 ( .C1(n8079), .C2(n8078), .A(n9363), .B(n8077), .ZN(n8080)
         );
  AOI211_X1 U9801 ( .C1(n8082), .C2(n9360), .A(n8081), .B(n8080), .ZN(n8083)
         );
  INV_X1 U9802 ( .A(n8083), .ZN(P2_U3176) );
  XNOR2_X1 U9803 ( .A(n8084), .B(n8498), .ZN(n8085) );
  OAI222_X1 U9804 ( .A1(n9644), .A2(n8563), .B1(n9646), .B2(n9645), .C1(n8085), 
        .C2(n9642), .ZN(n8228) );
  INV_X1 U9805 ( .A(n8228), .ZN(n8090) );
  XNOR2_X1 U9806 ( .A(n8086), .B(n8498), .ZN(n8229) );
  INV_X1 U9807 ( .A(n8250), .ZN(n8233) );
  AOI22_X1 U9808 ( .A1(n10632), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n10628), 
        .B2(n8246), .ZN(n8087) );
  OAI21_X1 U9809 ( .B1(n8233), .B2(n9637), .A(n8087), .ZN(n8088) );
  AOI21_X1 U9810 ( .B1(n8229), .B2(n9657), .A(n8088), .ZN(n8089) );
  OAI21_X1 U9811 ( .B1(n8090), .B2(n10632), .A(n8089), .ZN(P2_U3216) );
  INV_X1 U9812 ( .A(n8091), .ZN(n8143) );
  AOI21_X1 U9813 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9795), .A(n8092), .ZN(
        n8093) );
  OAI21_X1 U9814 ( .B1(n8143), .B2(n9801), .A(n8093), .ZN(P2_U3268) );
  AOI211_X1 U9815 ( .C1(n8096), .C2(n10520), .A(n8095), .B(n8094), .ZN(n8100)
         );
  AOI22_X1 U9816 ( .A1(n9848), .A2(n8889), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n10534), .ZN(n8097) );
  OAI21_X1 U9817 ( .B1(n8100), .B2(n10534), .A(n8097), .ZN(P1_U3538) );
  AOI22_X1 U9818 ( .A1(n9848), .A2(n8098), .B1(P1_REG0_REG_16__SCAN_IN), .B2(
        n6596), .ZN(n8099) );
  OAI21_X1 U9819 ( .B1(n8100), .B2(n6596), .A(n8099), .ZN(P1_U3501) );
  INV_X1 U9820 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8116) );
  AND2_X1 U9821 ( .A1(n8106), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8101) );
  OR2_X1 U9822 ( .A1(n8102), .A2(n8101), .ZN(n8104) );
  INV_X1 U9823 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8103) );
  XNOR2_X1 U9824 ( .A(n8104), .B(n8103), .ZN(n8108) );
  AOI21_X1 U9825 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8106), .A(n8105), .ZN(
        n8107) );
  XNOR2_X1 U9826 ( .A(n8107), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8110) );
  AOI22_X1 U9827 ( .A1(n8108), .A2(n10025), .B1(n10033), .B2(n8110), .ZN(n8114) );
  INV_X1 U9828 ( .A(n8108), .ZN(n8112) );
  OAI21_X1 U9829 ( .B1(n8110), .B2(n8109), .A(n10007), .ZN(n8111) );
  AOI21_X1 U9830 ( .B1(n8112), .B2(n10025), .A(n8111), .ZN(n8113) );
  MUX2_X1 U9831 ( .A(n8114), .B(n8113), .S(n6166), .Z(n8115) );
  NAND2_X1 U9832 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9817) );
  OAI211_X1 U9833 ( .C1(n8116), .C2(n9966), .A(n8115), .B(n9817), .ZN(P1_U3262) );
  AOI21_X1 U9834 ( .B1(n8120), .B2(n8119), .A(n8161), .ZN(n8140) );
  INV_X1 U9835 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10380) );
  MUX2_X1 U9836 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9521), .Z(n8175) );
  XNOR2_X1 U9837 ( .A(n8175), .B(n8177), .ZN(n8127) );
  INV_X1 U9838 ( .A(n8121), .ZN(n8123) );
  NAND2_X1 U9839 ( .A1(n8123), .A2(n8122), .ZN(n8125) );
  NAND2_X1 U9840 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  NAND2_X1 U9841 ( .A1(n8127), .A2(n8126), .ZN(n8178) );
  OAI21_X1 U9842 ( .B1(n8127), .B2(n8126), .A(n8178), .ZN(n8129) );
  AOI21_X1 U9843 ( .B1(n10612), .B2(n8129), .A(n8128), .ZN(n8130) );
  OAI21_X1 U9844 ( .B1(n10597), .B2(n10380), .A(n8130), .ZN(n8138) );
  INV_X1 U9845 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8135) );
  INV_X1 U9846 ( .A(n8177), .ZN(n8133) );
  AOI21_X1 U9847 ( .B1(n8135), .B2(n8134), .A(n8167), .ZN(n8136) );
  NOR2_X1 U9848 ( .A1(n8136), .A2(n10615), .ZN(n8137) );
  AOI211_X1 U9849 ( .C1(n10586), .C2(n8177), .A(n8138), .B(n8137), .ZN(n8139)
         );
  OAI21_X1 U9850 ( .B1(n8140), .B2(n10606), .A(n8139), .ZN(P2_U3193) );
  OAI222_X1 U9851 ( .A1(n8546), .A2(n8143), .B1(P1_U3086), .B2(n8142), .C1(
        n8141), .C2(n10338), .ZN(P1_U3328) );
  XNOR2_X1 U9852 ( .A(n8144), .B(n8765), .ZN(n10278) );
  INV_X1 U9853 ( .A(n8145), .ZN(n8147) );
  INV_X1 U9854 ( .A(n8211), .ZN(n8146) );
  AOI211_X1 U9855 ( .C1(n10275), .C2(n8147), .A(n10502), .B(n8146), .ZN(n10274) );
  INV_X1 U9856 ( .A(n9856), .ZN(n8148) );
  AOI22_X1 U9857 ( .A1(n10215), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8148), .B2(
        n10452), .ZN(n8149) );
  OAI21_X1 U9858 ( .B1(n8150), .B2(n10456), .A(n8149), .ZN(n8156) );
  NAND2_X1 U9859 ( .A1(n8151), .A2(n8689), .ZN(n8152) );
  XNOR2_X1 U9860 ( .A(n8152), .B(n8765), .ZN(n8154) );
  OAI22_X1 U9861 ( .A1(n9815), .A2(n9908), .B1(n8153), .B2(n9887), .ZN(n9854)
         );
  AOI21_X1 U9862 ( .B1(n8154), .B2(n10427), .A(n9854), .ZN(n10277) );
  NOR2_X1 U9863 ( .A1(n10277), .A2(n10215), .ZN(n8155) );
  AOI211_X1 U9864 ( .C1(n10274), .C2(n10450), .A(n8156), .B(n8155), .ZN(n8157)
         );
  OAI21_X1 U9865 ( .B1(n10278), .B2(n8158), .A(n8157), .ZN(P1_U3276) );
  INV_X1 U9866 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8162) );
  MUX2_X1 U9867 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8162), .S(n8174), .Z(n8164)
         );
  INV_X1 U9868 ( .A(n9389), .ZN(n8163) );
  AOI21_X1 U9869 ( .B1(n4611), .B2(n8164), .A(n8163), .ZN(n8189) );
  NOR2_X1 U9870 ( .A1(n8177), .A2(n8166), .ZN(n8168) );
  INV_X1 U9871 ( .A(n8171), .ZN(n8173) );
  MUX2_X1 U9872 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8169), .S(n8174), .Z(n8170)
         );
  INV_X1 U9873 ( .A(n8170), .ZN(n8172) );
  OAI21_X1 U9874 ( .B1(n8173), .B2(n8172), .A(n9407), .ZN(n8187) );
  INV_X1 U9875 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U9876 ( .A1(n10586), .A2(n8174), .ZN(n8185) );
  MUX2_X1 U9877 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9521), .Z(n9395) );
  XNOR2_X1 U9878 ( .A(n8174), .B(n9395), .ZN(n8181) );
  INV_X1 U9879 ( .A(n8175), .ZN(n8176) );
  NAND2_X1 U9880 ( .A1(n8177), .A2(n8176), .ZN(n8179) );
  NAND2_X1 U9881 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND2_X1 U9882 ( .A1(n8181), .A2(n8180), .ZN(n9396) );
  OAI21_X1 U9883 ( .B1(n8181), .B2(n8180), .A(n9396), .ZN(n8183) );
  AOI21_X1 U9884 ( .B1(n10612), .B2(n8183), .A(n8182), .ZN(n8184) );
  OAI211_X1 U9885 ( .C1(n10382), .C2(n10597), .A(n8185), .B(n8184), .ZN(n8186)
         );
  AOI21_X1 U9886 ( .B1(n8187), .B2(n10566), .A(n8186), .ZN(n8188) );
  OAI21_X1 U9887 ( .B1(n8189), .B2(n10606), .A(n8188), .ZN(P2_U3194) );
  INV_X1 U9888 ( .A(n8190), .ZN(n8894) );
  AOI21_X1 U9889 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9795), .A(n8191), .ZN(
        n8192) );
  OAI21_X1 U9890 ( .B1(n8894), .B2(n8274), .A(n8192), .ZN(P2_U3267) );
  INV_X1 U9891 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8195) );
  AOI21_X1 U9892 ( .B1(n9711), .B2(n8194), .A(n8193), .ZN(n8197) );
  MUX2_X1 U9893 ( .A(n8195), .B(n8197), .S(n9744), .Z(n8196) );
  OAI21_X1 U9894 ( .B1(n8200), .B2(n9715), .A(n8196), .ZN(P2_U3475) );
  INV_X1 U9895 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8198) );
  MUX2_X1 U9896 ( .A(n8198), .B(n8197), .S(n10649), .Z(n8199) );
  OAI21_X1 U9897 ( .B1(n8200), .B2(n9789), .A(n8199), .ZN(P2_U3438) );
  NAND2_X1 U9898 ( .A1(n8201), .A2(n8208), .ZN(n8202) );
  NAND2_X1 U9899 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  NAND2_X1 U9900 ( .A1(n8204), .A2(n10427), .ZN(n8207) );
  NOR2_X1 U9901 ( .A1(n8205), .A2(n9887), .ZN(n8206) );
  AOI21_X1 U9902 ( .B1(n6059), .B2(n9865), .A(n8206), .ZN(n9899) );
  NAND2_X1 U9903 ( .A1(n8207), .A2(n9899), .ZN(n10268) );
  INV_X1 U9904 ( .A(n10268), .ZN(n8217) );
  XNOR2_X1 U9905 ( .A(n8209), .B(n8208), .ZN(n10270) );
  NAND2_X1 U9906 ( .A1(n10270), .A2(n10458), .ZN(n8216) );
  INV_X1 U9907 ( .A(n10207), .ZN(n8210) );
  AOI211_X1 U9908 ( .C1(n8212), .C2(n8211), .A(n10502), .B(n8210), .ZN(n10269)
         );
  AOI22_X1 U9909 ( .A1(n10462), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9901), .B2(
        n10452), .ZN(n8213) );
  OAI21_X1 U9910 ( .B1(n10330), .B2(n10456), .A(n8213), .ZN(n8214) );
  AOI21_X1 U9911 ( .B1(n10269), .B2(n10450), .A(n8214), .ZN(n8215) );
  OAI211_X1 U9912 ( .C1(n10215), .C2(n8217), .A(n8216), .B(n8215), .ZN(
        P1_U3275) );
  NAND2_X1 U9913 ( .A1(n8218), .A2(n8500), .ZN(n8219) );
  INV_X1 U9914 ( .A(n9712), .ZN(n8227) );
  XOR2_X1 U9915 ( .A(n4559), .B(n8500), .Z(n8221) );
  OAI222_X1 U9916 ( .A1(n9644), .A2(n8259), .B1(n9646), .B2(n9630), .C1(n8221), 
        .C2(n9642), .ZN(n9710) );
  NAND2_X1 U9917 ( .A1(n9710), .A2(n10629), .ZN(n8226) );
  INV_X1 U9918 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9496) );
  INV_X1 U9919 ( .A(n8256), .ZN(n8223) );
  OAI22_X1 U9920 ( .A1(n10629), .A2(n9496), .B1(n8223), .B2(n8222), .ZN(n8224)
         );
  AOI21_X1 U9921 ( .B1(n8261), .B2(n9651), .A(n8224), .ZN(n8225) );
  OAI211_X1 U9922 ( .C1(n8900), .C2(n8227), .A(n8226), .B(n8225), .ZN(P2_U3215) );
  INV_X1 U9923 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9476) );
  AOI21_X1 U9924 ( .B1(n9711), .B2(n8229), .A(n8228), .ZN(n8231) );
  MUX2_X1 U9925 ( .A(n9476), .B(n8231), .S(n9744), .Z(n8230) );
  OAI21_X1 U9926 ( .B1(n8233), .B2(n9715), .A(n8230), .ZN(P2_U3476) );
  INV_X1 U9927 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8961) );
  MUX2_X1 U9928 ( .A(n8961), .B(n8231), .S(n10649), .Z(n8232) );
  OAI21_X1 U9929 ( .B1(n8233), .B2(n9789), .A(n8232), .ZN(P2_U3441) );
  INV_X1 U9930 ( .A(n8234), .ZN(n8235) );
  XNOR2_X1 U9931 ( .A(n9717), .B(n8600), .ZN(n8239) );
  XNOR2_X1 U9932 ( .A(n8239), .B(n8240), .ZN(n8560) );
  INV_X1 U9933 ( .A(n8239), .ZN(n8241) );
  XNOR2_X1 U9934 ( .A(n8556), .B(n8600), .ZN(n8549) );
  INV_X1 U9935 ( .A(n8549), .ZN(n8243) );
  XNOR2_X1 U9936 ( .A(n8250), .B(n8244), .ZN(n8253) );
  XNOR2_X1 U9937 ( .A(n8253), .B(n9377), .ZN(n8245) );
  XNOR2_X1 U9938 ( .A(n8255), .B(n8245), .ZN(n8252) );
  NAND2_X1 U9939 ( .A1(n9355), .A2(n8246), .ZN(n8248) );
  AND2_X1 U9940 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9481) );
  AOI21_X1 U9941 ( .B1(n9346), .B2(n9376), .A(n9481), .ZN(n8247) );
  OAI211_X1 U9942 ( .C1(n8563), .C2(n9327), .A(n8248), .B(n8247), .ZN(n8249)
         );
  AOI21_X1 U9943 ( .B1(n8250), .B2(n9360), .A(n8249), .ZN(n8251) );
  OAI21_X1 U9944 ( .B1(n8252), .B2(n9363), .A(n8251), .ZN(P2_U3168) );
  XNOR2_X1 U9945 ( .A(n9790), .B(n8600), .ZN(n8568) );
  XNOR2_X1 U9946 ( .A(n8568), .B(n9376), .ZN(n8571) );
  INV_X1 U9947 ( .A(n8253), .ZN(n8254) );
  XOR2_X1 U9948 ( .A(n8571), .B(n8572), .Z(n8263) );
  AOI22_X1 U9949 ( .A1(n9346), .A2(n9375), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8258) );
  NAND2_X1 U9950 ( .A1(n9355), .A2(n8256), .ZN(n8257) );
  OAI211_X1 U9951 ( .C1(n8259), .C2(n9327), .A(n8258), .B(n8257), .ZN(n8260)
         );
  AOI21_X1 U9952 ( .B1(n8261), .B2(n9360), .A(n8260), .ZN(n8262) );
  OAI21_X1 U9953 ( .B1(n8263), .B2(n9363), .A(n8262), .ZN(P2_U3178) );
  MUX2_X1 U9954 ( .A(n8264), .B(P2_REG2_REG_8__SCAN_IN), .S(n10632), .Z(n8270)
         );
  AOI22_X1 U9955 ( .A1(n9651), .A2(n8266), .B1(n10628), .B2(n8265), .ZN(n8267)
         );
  OAI21_X1 U9956 ( .B1(n8268), .B2(n8900), .A(n8267), .ZN(n8269) );
  OR2_X1 U9957 ( .A1(n8270), .A2(n8269), .ZN(P2_U3225) );
  INV_X1 U9958 ( .A(n8271), .ZN(n8273) );
  OAI222_X1 U9959 ( .A1(n6967), .A2(P2_U3151), .B1(n8274), .B2(n8273), .C1(
        n8272), .C2(n9798), .ZN(P2_U3275) );
  MUX2_X1 U9960 ( .A(n8912), .B(n9548), .S(n8453), .Z(n8451) );
  AND2_X1 U9961 ( .A1(n8381), .A2(n8371), .ZN(n8369) );
  NAND2_X1 U9962 ( .A1(n5689), .A2(n8453), .ZN(n8277) );
  OAI211_X1 U9963 ( .C1(n8278), .C2(n8453), .A(n8277), .B(n8276), .ZN(n8279)
         );
  INV_X1 U9964 ( .A(n8279), .ZN(n8366) );
  MUX2_X1 U9965 ( .A(n8285), .B(n8280), .S(n8453), .Z(n8291) );
  INV_X1 U9966 ( .A(n8282), .ZN(n8283) );
  NAND2_X1 U9967 ( .A1(n8283), .A2(n8523), .ZN(n8287) );
  NAND2_X1 U9968 ( .A1(n8283), .A2(n8513), .ZN(n8284) );
  NAND3_X1 U9969 ( .A1(n8285), .A2(n8284), .A3(n8453), .ZN(n8286) );
  OAI21_X1 U9970 ( .B1(n6861), .B2(n8287), .A(n8286), .ZN(n8288) );
  OAI21_X1 U9971 ( .B1(n8513), .B2(n8289), .A(n8288), .ZN(n8290) );
  NAND3_X1 U9972 ( .A1(n8291), .A2(n8281), .A3(n8290), .ZN(n8298) );
  NAND2_X1 U9973 ( .A1(n8309), .A2(n8292), .ZN(n8295) );
  NAND2_X1 U9974 ( .A1(n8301), .A2(n8293), .ZN(n8294) );
  MUX2_X1 U9975 ( .A(n8295), .B(n8294), .S(n8448), .Z(n8296) );
  INV_X1 U9976 ( .A(n8296), .ZN(n8297) );
  NAND2_X1 U9977 ( .A1(n8298), .A2(n8297), .ZN(n8300) );
  NAND2_X1 U9978 ( .A1(n8300), .A2(n8299), .ZN(n8312) );
  INV_X1 U9979 ( .A(n8301), .ZN(n8304) );
  OAI211_X1 U9980 ( .C1(n8312), .C2(n8304), .A(n8303), .B(n8302), .ZN(n8308)
         );
  AND2_X1 U9981 ( .A1(n8313), .A2(n8310), .ZN(n8307) );
  INV_X1 U9982 ( .A(n8305), .ZN(n8306) );
  AOI21_X1 U9983 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8317) );
  OAI211_X1 U9984 ( .C1(n8312), .C2(n4636), .A(n8311), .B(n8310), .ZN(n8315)
         );
  AOI21_X1 U9985 ( .B1(n8315), .B2(n8314), .A(n4648), .ZN(n8316) );
  MUX2_X1 U9986 ( .A(n8317), .B(n8316), .S(n8448), .Z(n8318) );
  NAND3_X1 U9987 ( .A1(n8318), .A2(n8487), .A3(n8329), .ZN(n8333) );
  NAND2_X1 U9988 ( .A1(n8320), .A2(n8319), .ZN(n8323) );
  NAND2_X1 U9989 ( .A1(n8338), .A2(n8321), .ZN(n8322) );
  AOI21_X1 U9990 ( .B1(n8329), .B2(n8323), .A(n8322), .ZN(n8331) );
  NAND2_X1 U9991 ( .A1(n8325), .A2(n8324), .ZN(n8328) );
  NAND2_X1 U9992 ( .A1(n8334), .A2(n8326), .ZN(n8327) );
  AOI21_X1 U9993 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(n8330) );
  MUX2_X1 U9994 ( .A(n8331), .B(n8330), .S(n8448), .Z(n8332) );
  NAND2_X1 U9995 ( .A1(n8333), .A2(n8332), .ZN(n8342) );
  NAND2_X1 U9996 ( .A1(n8342), .A2(n8334), .ZN(n8335) );
  NAND2_X1 U9997 ( .A1(n8335), .A2(n8339), .ZN(n8337) );
  NAND2_X1 U9998 ( .A1(n8337), .A2(n8336), .ZN(n8344) );
  AND2_X1 U9999 ( .A1(n8339), .A2(n8338), .ZN(n8341) );
  AOI21_X1 U10000 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8343) );
  MUX2_X1 U10001 ( .A(n8346), .B(n8345), .S(n8448), .Z(n8347) );
  MUX2_X1 U10002 ( .A(n9379), .B(n8349), .S(n8448), .Z(n8350) );
  MUX2_X1 U10003 ( .A(n8353), .B(n8352), .S(n8453), .Z(n8354) );
  NAND3_X1 U10004 ( .A1(n8356), .A2(n8355), .A3(n8354), .ZN(n8361) );
  INV_X1 U10005 ( .A(n8357), .ZN(n8359) );
  MUX2_X1 U10006 ( .A(n8359), .B(n8358), .S(n8453), .Z(n8360) );
  INV_X1 U10007 ( .A(n8498), .ZN(n8365) );
  MUX2_X1 U10008 ( .A(n8363), .B(n8362), .S(n8453), .Z(n8364) );
  NAND2_X1 U10009 ( .A1(n9645), .A2(n8453), .ZN(n8367) );
  OAI21_X1 U10010 ( .B1(n9790), .B2(n8367), .A(n8379), .ZN(n8368) );
  NAND2_X1 U10011 ( .A1(n8369), .A2(n8368), .ZN(n8374) );
  AOI21_X1 U10012 ( .B1(n8371), .B2(n8370), .A(n8453), .ZN(n8372) );
  INV_X1 U10013 ( .A(n8372), .ZN(n8373) );
  INV_X1 U10014 ( .A(n8380), .ZN(n8378) );
  INV_X1 U10015 ( .A(n8375), .ZN(n8377) );
  INV_X1 U10016 ( .A(n8384), .ZN(n8376) );
  AOI21_X1 U10017 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8387) );
  INV_X1 U10018 ( .A(n8382), .ZN(n8383) );
  AOI21_X1 U10019 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8386) );
  NAND2_X1 U10020 ( .A1(n9586), .A2(n8388), .ZN(n8391) );
  NAND2_X1 U10021 ( .A1(n8475), .A2(n8389), .ZN(n8390) );
  MUX2_X1 U10022 ( .A(n8391), .B(n8390), .S(n8448), .Z(n8392) );
  INV_X1 U10023 ( .A(n8392), .ZN(n8393) );
  NAND2_X1 U10024 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  INV_X1 U10025 ( .A(n8396), .ZN(n8399) );
  NAND3_X1 U10026 ( .A1(n8398), .A2(n9575), .A3(n8397), .ZN(n8400) );
  NAND2_X1 U10027 ( .A1(n8400), .A2(n8399), .ZN(n8408) );
  AOI21_X1 U10028 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(n8406) );
  INV_X1 U10029 ( .A(n9575), .ZN(n8405) );
  OAI21_X1 U10030 ( .B1(n8406), .B2(n8405), .A(n8404), .ZN(n8407) );
  MUX2_X1 U10031 ( .A(n8408), .B(n8407), .S(n8448), .Z(n8414) );
  INV_X1 U10032 ( .A(n8409), .ZN(n8411) );
  INV_X1 U10033 ( .A(n9563), .ZN(n8505) );
  MUX2_X1 U10034 ( .A(n8411), .B(n8410), .S(n8448), .Z(n8412) );
  OR2_X1 U10035 ( .A1(n8507), .A2(n8412), .ZN(n8413) );
  AOI21_X1 U10036 ( .B1(n8414), .B2(n8505), .A(n8413), .ZN(n8418) );
  INV_X1 U10037 ( .A(n8415), .ZN(n8417) );
  MUX2_X1 U10038 ( .A(n9367), .B(n8601), .S(n8453), .Z(n8416) );
  INV_X1 U10039 ( .A(SI_29_), .ZN(n8419) );
  INV_X1 U10040 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8547) );
  INV_X1 U10041 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10042 ( .A(n8547), .B(n8895), .S(n4518), .Z(n8426) );
  INV_X1 U10043 ( .A(SI_30_), .ZN(n8425) );
  NAND2_X1 U10044 ( .A1(n8426), .A2(n8425), .ZN(n8432) );
  INV_X1 U10045 ( .A(n8426), .ZN(n8427) );
  NAND2_X1 U10046 ( .A1(n8427), .A2(SI_30_), .ZN(n8428) );
  NAND2_X1 U10047 ( .A1(n8432), .A2(n8428), .ZN(n8433) );
  NAND2_X1 U10048 ( .A1(n8544), .A2(n8438), .ZN(n8430) );
  OR2_X1 U10049 ( .A1(n5333), .A2(n8895), .ZN(n8429) );
  NAND2_X1 U10050 ( .A1(n8430), .A2(n8429), .ZN(n9750) );
  NAND2_X1 U10051 ( .A1(n9750), .A2(n8449), .ZN(n8510) );
  NAND2_X1 U10052 ( .A1(n8510), .A2(n8431), .ZN(n8466) );
  AOI21_X1 U10053 ( .B1(n8461), .B2(n8912), .A(n8466), .ZN(n8458) );
  INV_X1 U10054 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10339) );
  INV_X1 U10055 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8439) );
  MUX2_X1 U10056 ( .A(n10339), .B(n8439), .S(n4518), .Z(n8435) );
  XNOR2_X1 U10057 ( .A(n8435), .B(SI_31_), .ZN(n8436) );
  NAND2_X1 U10058 ( .A1(n10344), .A2(n8438), .ZN(n8441) );
  OR2_X1 U10059 ( .A1(n5333), .A2(n8439), .ZN(n8440) );
  NAND2_X1 U10060 ( .A1(n4519), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10061 ( .A1(n4525), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10062 ( .A1(n4520), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8443) );
  NAND4_X1 U10063 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n9540)
         );
  INV_X1 U10064 ( .A(n9540), .ZN(n8447) );
  NAND2_X1 U10065 ( .A1(n8510), .A2(n8448), .ZN(n8450) );
  OR2_X1 U10066 ( .A1(n9750), .A2(n8449), .ZN(n8509) );
  NAND2_X1 U10067 ( .A1(n8450), .A2(n8509), .ZN(n8462) );
  NOR2_X1 U10068 ( .A1(n4546), .A2(n8462), .ZN(n8455) );
  INV_X1 U10069 ( .A(n8455), .ZN(n8457) );
  NAND2_X1 U10070 ( .A1(n9662), .A2(n9540), .ZN(n8470) );
  INV_X1 U10071 ( .A(n8470), .ZN(n8473) );
  NOR3_X1 U10072 ( .A1(n4546), .A2(n8456), .A3(n8453), .ZN(n8454) );
  INV_X1 U10073 ( .A(n8467), .ZN(n8460) );
  INV_X1 U10074 ( .A(n8509), .ZN(n8459) );
  NAND2_X1 U10075 ( .A1(n8470), .A2(n8462), .ZN(n8463) );
  AOI21_X1 U10076 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8471) );
  INV_X1 U10077 ( .A(n9750), .ZN(n9665) );
  NOR2_X1 U10078 ( .A1(n8509), .A2(n9662), .ZN(n8472) );
  NOR2_X1 U10079 ( .A1(n4546), .A2(n8473), .ZN(n8512) );
  INV_X1 U10080 ( .A(n8474), .ZN(n8604) );
  NAND2_X1 U10081 ( .A1(n8475), .A2(n9586), .ZN(n9595) );
  INV_X1 U10082 ( .A(n9619), .ZN(n9613) );
  INV_X1 U10083 ( .A(n9632), .ZN(n8502) );
  INV_X1 U10084 ( .A(n8477), .ZN(n8491) );
  INV_X1 U10085 ( .A(n6861), .ZN(n8479) );
  NAND4_X1 U10086 ( .A1(n8281), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n8484)
         );
  NOR4_X1 U10087 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n8488)
         );
  NAND4_X1 U10088 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n8489)
         );
  NOR4_X1 U10089 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n8494)
         );
  NAND4_X1 U10090 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(n8499)
         );
  NOR4_X1 U10091 ( .A1(n8500), .A2(n8499), .A3(n8498), .A4(n8497), .ZN(n8501)
         );
  NAND4_X1 U10092 ( .A1(n9613), .A2(n8502), .A3(n9654), .A4(n8501), .ZN(n8503)
         );
  NOR4_X1 U10093 ( .A1(n9589), .A2(n9595), .A3(n9605), .A4(n8503), .ZN(n8504)
         );
  NAND3_X1 U10094 ( .A1(n8505), .A2(n9575), .A3(n8504), .ZN(n8506) );
  NOR4_X1 U10095 ( .A1(n8508), .A2(n8507), .A3(n8604), .A4(n8506), .ZN(n8511)
         );
  NAND4_X1 U10096 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n8514)
         );
  NAND2_X1 U10097 ( .A1(n8517), .A2(n8516), .ZN(n8518) );
  NAND2_X1 U10098 ( .A1(n8519), .A2(n8518), .ZN(n8520) );
  XNOR2_X1 U10099 ( .A(n8520), .B(n5694), .ZN(n8527) );
  NOR3_X1 U10100 ( .A1(n8522), .A2(n8521), .A3(n5668), .ZN(n8525) );
  OAI21_X1 U10101 ( .B1(n8526), .B2(n8523), .A(P2_B_REG_SCAN_IN), .ZN(n8524)
         );
  OAI22_X1 U10102 ( .A1(n8527), .A2(n8526), .B1(n8525), .B2(n8524), .ZN(
        P2_U3296) );
  NOR2_X1 U10103 ( .A1(n8530), .A2(n10339), .ZN(n8528) );
  NAND2_X1 U10104 ( .A1(n8544), .A2(n8529), .ZN(n8532) );
  OR2_X1 U10105 ( .A1(n8530), .A2(n8547), .ZN(n8531) );
  NAND2_X1 U10106 ( .A1(n8533), .A2(n4741), .ZN(n10040) );
  XNOR2_X1 U10107 ( .A(n10289), .B(n10040), .ZN(n8534) );
  INV_X1 U10108 ( .A(n8535), .ZN(n8541) );
  INV_X1 U10109 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U10110 ( .A1(n8536), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10111 ( .A1(n8537), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8538) );
  OAI211_X1 U10112 ( .C1(n8540), .C2(n9194), .A(n8539), .B(n8538), .ZN(n9932)
         );
  NAND2_X1 U10113 ( .A1(n8541), .A2(n9932), .ZN(n10216) );
  NOR2_X1 U10114 ( .A1(n10215), .A2(n10216), .ZN(n10044) );
  NOR2_X1 U10115 ( .A1(n10289), .A2(n10456), .ZN(n8542) );
  AOI211_X1 U10116 ( .C1(n10215), .C2(P1_REG2_REG_31__SCAN_IN), .A(n10044), 
        .B(n8542), .ZN(n8543) );
  OAI21_X1 U10117 ( .B1(n8884), .B2(n10194), .A(n8543), .ZN(P1_U3263) );
  INV_X1 U10118 ( .A(n8544), .ZN(n8896) );
  OAI222_X1 U10119 ( .A1(n10338), .A2(n8547), .B1(n8546), .B2(n8896), .C1(
        P1_U3086), .C2(n8545), .ZN(P1_U3325) );
  XNOR2_X1 U10120 ( .A(n8549), .B(n8563), .ZN(n8550) );
  XNOR2_X1 U10121 ( .A(n8548), .B(n8550), .ZN(n8558) );
  NAND2_X1 U10122 ( .A1(n9355), .A2(n8551), .ZN(n8553) );
  NOR2_X1 U10123 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9192), .ZN(n9452) );
  AOI21_X1 U10124 ( .B1(n9346), .B2(n9377), .A(n9452), .ZN(n8552) );
  OAI211_X1 U10125 ( .C1(n8554), .C2(n9327), .A(n8553), .B(n8552), .ZN(n8555)
         );
  AOI21_X1 U10126 ( .B1(n8556), .B2(n9360), .A(n8555), .ZN(n8557) );
  OAI21_X1 U10127 ( .B1(n8558), .B2(n9363), .A(n8557), .ZN(P2_U3166) );
  OAI211_X1 U10128 ( .C1(n8561), .C2(n8560), .A(n8559), .B(n9342), .ZN(n8567)
         );
  AND2_X1 U10129 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9430) );
  AOI21_X1 U10130 ( .B1(n9354), .B2(n9378), .A(n9430), .ZN(n8562) );
  OAI21_X1 U10131 ( .B1(n9358), .B2(n8563), .A(n8562), .ZN(n8564) );
  AOI21_X1 U10132 ( .B1(n8565), .B2(n9355), .A(n8564), .ZN(n8566) );
  OAI211_X1 U10133 ( .C1(n9717), .C2(n8930), .A(n8567), .B(n8566), .ZN(
        P2_U3181) );
  INV_X1 U10134 ( .A(n8568), .ZN(n8569) );
  NOR2_X1 U10135 ( .A1(n8569), .A2(n9376), .ZN(n8570) );
  AOI21_X1 U10136 ( .B1(n8572), .B2(n8571), .A(n8570), .ZN(n8925) );
  XNOR2_X1 U10137 ( .A(n9652), .B(n8600), .ZN(n8573) );
  XNOR2_X1 U10138 ( .A(n8573), .B(n9630), .ZN(n8924) );
  NAND2_X1 U10139 ( .A1(n8925), .A2(n8924), .ZN(n8923) );
  NAND2_X1 U10140 ( .A1(n8573), .A2(n9375), .ZN(n8574) );
  NAND2_X1 U10141 ( .A1(n8923), .A2(n8574), .ZN(n9323) );
  INV_X1 U10142 ( .A(n9323), .ZN(n8576) );
  XNOR2_X1 U10143 ( .A(n9634), .B(n8600), .ZN(n8577) );
  XNOR2_X1 U10144 ( .A(n8577), .B(n9374), .ZN(n9324) );
  INV_X1 U10145 ( .A(n8577), .ZN(n8578) );
  NAND2_X1 U10146 ( .A1(n8578), .A2(n9647), .ZN(n8579) );
  XNOR2_X1 U10147 ( .A(n8936), .B(n8600), .ZN(n8580) );
  XNOR2_X1 U10148 ( .A(n8580), .B(n9631), .ZN(n8931) );
  INV_X1 U10149 ( .A(n8580), .ZN(n8581) );
  XNOR2_X1 U10150 ( .A(n9607), .B(n8600), .ZN(n8583) );
  XNOR2_X1 U10151 ( .A(n8582), .B(n8583), .ZN(n9331) );
  NAND2_X1 U10152 ( .A1(n9331), .A2(n9616), .ZN(n8586) );
  INV_X1 U10153 ( .A(n8583), .ZN(n8584) );
  NAND2_X1 U10154 ( .A1(n8582), .A2(n8584), .ZN(n8585) );
  NAND2_X1 U10155 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  XNOR2_X1 U10156 ( .A(n8920), .B(n4513), .ZN(n8588) );
  XNOR2_X1 U10157 ( .A(n8587), .B(n8588), .ZN(n8916) );
  NAND2_X1 U10158 ( .A1(n8916), .A2(n9604), .ZN(n8591) );
  INV_X1 U10159 ( .A(n8587), .ZN(n8589) );
  NAND2_X1 U10160 ( .A1(n8591), .A2(n8590), .ZN(n9314) );
  XNOR2_X1 U10161 ( .A(n9580), .B(n8600), .ZN(n8592) );
  XNOR2_X1 U10162 ( .A(n8592), .B(n9594), .ZN(n9315) );
  INV_X1 U10163 ( .A(n8592), .ZN(n8593) );
  NAND2_X1 U10164 ( .A1(n8593), .A2(n9594), .ZN(n8594) );
  XNOR2_X1 U10165 ( .A(n9572), .B(n4513), .ZN(n8595) );
  XNOR2_X1 U10166 ( .A(n8595), .B(n9583), .ZN(n8940) );
  NOR2_X1 U10167 ( .A1(n8595), .A2(n9369), .ZN(n8596) );
  XNOR2_X1 U10168 ( .A(n9361), .B(n8600), .ZN(n8597) );
  INV_X1 U10169 ( .A(n8597), .ZN(n8598) );
  NAND2_X1 U10170 ( .A1(n8598), .A2(n9571), .ZN(n8599) );
  XNOR2_X1 U10171 ( .A(n8601), .B(n4513), .ZN(n8602) );
  NAND2_X1 U10172 ( .A1(n8602), .A2(n9367), .ZN(n8603) );
  OAI21_X1 U10173 ( .B1(n8602), .B2(n9367), .A(n8603), .ZN(n8908) );
  NAND2_X1 U10174 ( .A1(n8909), .A2(n8603), .ZN(n8606) );
  XNOR2_X1 U10175 ( .A(n8604), .B(n4513), .ZN(n8605) );
  XNOR2_X1 U10176 ( .A(n8606), .B(n8605), .ZN(n8612) );
  INV_X1 U10177 ( .A(n8607), .ZN(n9365) );
  AOI22_X1 U10178 ( .A1(n9346), .A2(n9365), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8609) );
  NAND2_X1 U10179 ( .A1(n9355), .A2(n9546), .ZN(n8608) );
  OAI211_X1 U10180 ( .C1(n9562), .C2(n9327), .A(n8609), .B(n8608), .ZN(n8610)
         );
  AOI21_X1 U10181 ( .B1(n9671), .B2(n9360), .A(n8610), .ZN(n8611) );
  OAI21_X1 U10182 ( .B1(n8612), .B2(n9363), .A(n8611), .ZN(P2_U3160) );
  INV_X1 U10183 ( .A(n8775), .ZN(n9933) );
  OAI21_X1 U10184 ( .B1(n10289), .B2(n9933), .A(n9932), .ZN(n8740) );
  NAND2_X1 U10185 ( .A1(n8615), .A2(n8613), .ZN(n8796) );
  OR2_X1 U10186 ( .A1(n10177), .A2(n9888), .ZN(n8713) );
  NAND2_X1 U10187 ( .A1(n8713), .A2(n8708), .ZN(n8614) );
  NAND2_X1 U10188 ( .A1(n8614), .A2(n8697), .ZN(n8786) );
  OAI21_X1 U10189 ( .B1(n8616), .B2(n8786), .A(n8629), .ZN(n8619) );
  MUX2_X1 U10190 ( .A(n10116), .B(n8615), .S(n8737), .Z(n8618) );
  AND2_X1 U10191 ( .A1(n8787), .A2(n8737), .ZN(n8621) );
  NAND3_X1 U10192 ( .A1(n10116), .A2(n8621), .A3(n8616), .ZN(n8617) );
  OAI211_X1 U10193 ( .C1(n8796), .C2(n8619), .A(n8618), .B(n8617), .ZN(n8620)
         );
  INV_X1 U10194 ( .A(n8620), .ZN(n8720) );
  INV_X1 U10195 ( .A(n8621), .ZN(n8622) );
  OAI22_X1 U10196 ( .A1(n8796), .A2(n8737), .B1(n8790), .B2(n8622), .ZN(n8718)
         );
  AOI21_X1 U10197 ( .B1(n8624), .B2(n8824), .A(n8623), .ZN(n8630) );
  INV_X1 U10198 ( .A(n8824), .ZN(n8625) );
  NAND2_X1 U10199 ( .A1(n8637), .A2(n8636), .ZN(n8639) );
  INV_X1 U10200 ( .A(n8749), .ZN(n8644) );
  NOR2_X1 U10201 ( .A1(n8645), .A2(n8644), .ZN(n8647) );
  MUX2_X1 U10202 ( .A(n8647), .B(n8646), .S(n8737), .Z(n8651) );
  NAND2_X1 U10203 ( .A1(n8652), .A2(n8648), .ZN(n8649) );
  MUX2_X1 U10204 ( .A(n8649), .B(n8753), .S(n8737), .Z(n8650) );
  NAND2_X1 U10205 ( .A1(n8663), .A2(n8653), .ZN(n8835) );
  NOR2_X1 U10206 ( .A1(n8654), .A2(n8835), .ZN(n8656) );
  NAND2_X1 U10207 ( .A1(n8666), .A2(n8655), .ZN(n8839) );
  OAI21_X1 U10208 ( .B1(n8656), .B2(n8839), .A(n8838), .ZN(n8657) );
  NAND2_X1 U10209 ( .A1(n8657), .A2(n8737), .ZN(n8670) );
  INV_X1 U10210 ( .A(n8658), .ZN(n8659) );
  OAI211_X1 U10211 ( .C1(n8665), .C2(n8664), .A(n8838), .B(n8663), .ZN(n8667)
         );
  NAND2_X1 U10212 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  INV_X1 U10213 ( .A(n8684), .ZN(n8673) );
  INV_X1 U10214 ( .A(n8682), .ZN(n8672) );
  OAI211_X1 U10215 ( .C1(n8673), .C2(n8672), .A(n8837), .B(n8671), .ZN(n8674)
         );
  NAND3_X1 U10216 ( .A1(n8674), .A2(n8683), .A3(n8687), .ZN(n8678) );
  NAND2_X1 U10217 ( .A1(n10281), .A2(n8675), .ZN(n8676) );
  NAND2_X1 U10218 ( .A1(n8689), .A2(n8676), .ZN(n8686) );
  INV_X1 U10219 ( .A(n8686), .ZN(n8677) );
  INV_X1 U10220 ( .A(n8688), .ZN(n8679) );
  NOR2_X1 U10221 ( .A1(n8679), .A2(n8629), .ZN(n8680) );
  NAND2_X1 U10222 ( .A1(n8681), .A2(n8680), .ZN(n8694) );
  NAND2_X1 U10223 ( .A1(n8683), .A2(n8682), .ZN(n8841) );
  AOI21_X1 U10224 ( .B1(n8684), .B2(n8837), .A(n8841), .ZN(n8691) );
  OR2_X1 U10225 ( .A1(n8686), .A2(n8685), .ZN(n8819) );
  NAND2_X1 U10226 ( .A1(n8688), .A2(n8687), .ZN(n8690) );
  NAND2_X1 U10227 ( .A1(n8690), .A2(n8689), .ZN(n8844) );
  OAI21_X1 U10228 ( .B1(n8691), .B2(n8819), .A(n8844), .ZN(n8692) );
  NAND2_X1 U10229 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  INV_X1 U10230 ( .A(n8705), .ZN(n8696) );
  NOR2_X1 U10231 ( .A1(n8696), .A2(n8703), .ZN(n8845) );
  AOI211_X1 U10232 ( .C1(n8704), .C2(n8845), .A(n8707), .B(n4993), .ZN(n8698)
         );
  NAND2_X1 U10233 ( .A1(n8697), .A2(n8737), .ZN(n8714) );
  OAI21_X1 U10234 ( .B1(n8698), .B2(n10174), .A(n8714), .ZN(n8711) );
  INV_X1 U10235 ( .A(n8706), .ZN(n8699) );
  OAI21_X1 U10236 ( .B1(n8700), .B2(n8699), .A(n8629), .ZN(n8710) );
  AND2_X1 U10237 ( .A1(n8702), .A2(n8701), .ZN(n8850) );
  AND2_X1 U10238 ( .A1(n8706), .A2(n8705), .ZN(n8851) );
  INV_X1 U10239 ( .A(n10102), .ZN(n8719) );
  NAND2_X1 U10240 ( .A1(n8818), .A2(n8792), .ZN(n8723) );
  NAND2_X1 U10241 ( .A1(n8722), .A2(n8737), .ZN(n8729) );
  AOI21_X1 U10242 ( .B1(n8724), .B2(n4785), .A(n8723), .ZN(n8726) );
  INV_X1 U10243 ( .A(n8725), .ZN(n8784) );
  NOR2_X1 U10244 ( .A1(n8726), .A2(n8784), .ZN(n8727) );
  NAND2_X1 U10245 ( .A1(n8727), .A2(n8629), .ZN(n8728) );
  NAND2_X1 U10246 ( .A1(n8729), .A2(n8728), .ZN(n8734) );
  INV_X1 U10247 ( .A(n8734), .ZN(n8730) );
  OAI21_X1 U10248 ( .B1(n8730), .B2(n8785), .A(n8735), .ZN(n8731) );
  AOI21_X1 U10249 ( .B1(n8731), .B2(n8799), .A(n8737), .ZN(n8733) );
  NOR2_X1 U10250 ( .A1(n8734), .A2(n8785), .ZN(n8736) );
  INV_X1 U10251 ( .A(n8735), .ZN(n8794) );
  OAI211_X1 U10252 ( .C1(n8736), .C2(n8794), .A(n8737), .B(n8799), .ZN(n8739)
         );
  INV_X1 U10253 ( .A(n8800), .ZN(n8738) );
  INV_X1 U10254 ( .A(n9932), .ZN(n8804) );
  AND2_X1 U10255 ( .A1(n4940), .A2(n8804), .ZN(n8808) );
  OAI21_X1 U10256 ( .B1(n8780), .B2(n6265), .A(n4526), .ZN(n8779) );
  OR2_X1 U10257 ( .A1(n10043), .A2(n8775), .ZN(n8863) );
  NAND2_X1 U10258 ( .A1(n4785), .A2(n8792), .ZN(n10106) );
  NAND4_X1 U10259 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n8747)
         );
  NOR3_X1 U10260 ( .A1(n8747), .A2(n8746), .A3(n8745), .ZN(n8751) );
  NAND4_X1 U10261 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n8752)
         );
  NOR2_X1 U10262 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  NAND4_X1 U10263 ( .A1(n8756), .A2(n8834), .A3(n8755), .A4(n8754), .ZN(n8757)
         );
  NOR2_X1 U10264 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NAND3_X1 U10265 ( .A1(n8760), .A2(n10430), .A3(n8759), .ZN(n8761) );
  NOR3_X1 U10266 ( .A1(n8763), .A2(n8762), .A3(n8761), .ZN(n8764) );
  NAND3_X1 U10267 ( .A1(n8766), .A2(n8765), .A3(n8764), .ZN(n8767) );
  NOR2_X1 U10268 ( .A1(n10205), .A2(n8767), .ZN(n8769) );
  INV_X1 U10269 ( .A(n10174), .ZN(n8768) );
  NAND4_X1 U10270 ( .A1(n10154), .A2(n10189), .A3(n8769), .A4(n8768), .ZN(
        n8770) );
  NOR2_X1 U10271 ( .A1(n10138), .A2(n8770), .ZN(n8771) );
  NAND2_X1 U10272 ( .A1(n4796), .A2(n8771), .ZN(n8772) );
  OR4_X1 U10273 ( .A1(n10075), .A2(n10087), .A3(n10106), .A4(n8772), .ZN(n8773) );
  NOR2_X1 U10274 ( .A1(n8774), .A2(n8773), .ZN(n8776) );
  NAND2_X1 U10275 ( .A1(n10043), .A2(n8775), .ZN(n8803) );
  AND4_X1 U10276 ( .A1(n8777), .A2(n8863), .A3(n8776), .A4(n8803), .ZN(n8778)
         );
  NAND3_X1 U10277 ( .A1(n8866), .A2(n8778), .A3(n4936), .ZN(n8809) );
  NAND2_X1 U10278 ( .A1(n8779), .A2(n8809), .ZN(n8817) );
  OAI211_X1 U10279 ( .C1(n8866), .C2(n8816), .A(n4526), .B(n6265), .ZN(n8781)
         );
  INV_X1 U10280 ( .A(n8781), .ZN(n8782) );
  NAND2_X1 U10281 ( .A1(n8783), .A2(n8782), .ZN(n8815) );
  NOR2_X1 U10282 ( .A1(n8785), .A2(n8784), .ZN(n8857) );
  INV_X1 U10283 ( .A(n8786), .ZN(n8788) );
  AOI21_X1 U10284 ( .B1(n8788), .B2(n8787), .A(n8796), .ZN(n8791) );
  NOR3_X1 U10285 ( .A1(n8791), .A2(n4790), .A3(n8790), .ZN(n8793) );
  OAI21_X1 U10286 ( .B1(n8793), .B2(n8797), .A(n8792), .ZN(n8795) );
  AOI21_X1 U10287 ( .B1(n8857), .B2(n8795), .A(n8794), .ZN(n8862) );
  OR3_X1 U10288 ( .A1(n8797), .A2(n5123), .A3(n8796), .ZN(n8854) );
  OAI21_X1 U10289 ( .B1(n8854), .B2(n10185), .A(n8818), .ZN(n8798) );
  NAND2_X1 U10290 ( .A1(n8857), .A2(n8798), .ZN(n8801) );
  NAND2_X1 U10291 ( .A1(n8800), .A2(n8799), .ZN(n8860) );
  AOI21_X1 U10292 ( .B1(n8862), .B2(n8801), .A(n8860), .ZN(n8805) );
  NAND2_X1 U10293 ( .A1(n8803), .A2(n8802), .ZN(n8864) );
  OAI22_X1 U10294 ( .A1(n8805), .A2(n8864), .B1(n8804), .B2(n8863), .ZN(n8806)
         );
  OAI211_X1 U10295 ( .C1(n4741), .C2(n9932), .A(n8806), .B(n8866), .ZN(n8812)
         );
  NOR2_X1 U10296 ( .A1(n8808), .A2(n8807), .ZN(n8811) );
  INV_X1 U10297 ( .A(n8809), .ZN(n8810) );
  AOI21_X1 U10298 ( .B1(n8812), .B2(n8811), .A(n8810), .ZN(n8813) );
  OAI211_X1 U10299 ( .C1(n8817), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8872)
         );
  NOR2_X1 U10300 ( .A1(n8816), .A2(n8871), .ZN(n8869) );
  INV_X1 U10301 ( .A(n8818), .ZN(n8859) );
  INV_X1 U10302 ( .A(n8819), .ZN(n8849) );
  INV_X1 U10303 ( .A(n8820), .ZN(n8829) );
  OAI211_X1 U10304 ( .C1(n8823), .C2(n8822), .A(n4526), .B(n8821), .ZN(n8827)
         );
  OAI211_X1 U10305 ( .C1(n8827), .C2(n8625), .A(n8826), .B(n8825), .ZN(n8828)
         );
  OAI21_X1 U10306 ( .B1(n8829), .B2(n8828), .A(n4609), .ZN(n8833) );
  INV_X1 U10307 ( .A(n8830), .ZN(n8831) );
  NOR2_X1 U10308 ( .A1(n8836), .A2(n8835), .ZN(n8840) );
  OAI211_X1 U10309 ( .C1(n8840), .C2(n8839), .A(n8838), .B(n8837), .ZN(n8843)
         );
  INV_X1 U10310 ( .A(n8841), .ZN(n8842) );
  NAND2_X1 U10311 ( .A1(n8843), .A2(n8842), .ZN(n8848) );
  INV_X1 U10312 ( .A(n8844), .ZN(n8847) );
  INV_X1 U10313 ( .A(n8845), .ZN(n8846) );
  AOI211_X1 U10314 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8853)
         );
  INV_X1 U10315 ( .A(n8850), .ZN(n8852) );
  OAI21_X1 U10316 ( .B1(n8853), .B2(n8852), .A(n8851), .ZN(n8855) );
  AOI21_X1 U10317 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8858) );
  OAI21_X1 U10318 ( .B1(n8859), .B2(n8858), .A(n8857), .ZN(n8861) );
  AOI21_X1 U10319 ( .B1(n8862), .B2(n8861), .A(n8860), .ZN(n8865) );
  OAI211_X1 U10320 ( .C1(n8865), .C2(n8864), .A(n4936), .B(n8863), .ZN(n8867)
         );
  NAND2_X1 U10321 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  MUX2_X1 U10322 ( .A(n8869), .B(n6266), .S(n8868), .Z(n8870) );
  AOI21_X1 U10323 ( .B1(n8872), .B2(n8871), .A(n8870), .ZN(n8880) );
  NOR3_X1 U10324 ( .A1(n8875), .A2(n8874), .A3(n8873), .ZN(n8878) );
  OAI21_X1 U10325 ( .B1(n8879), .B2(n8876), .A(P1_B_REG_SCAN_IN), .ZN(n8877)
         );
  OAI22_X1 U10326 ( .A1(n8880), .A2(n8879), .B1(n8878), .B2(n8877), .ZN(
        P1_U3242) );
  INV_X1 U10327 ( .A(n8881), .ZN(n9800) );
  OAI222_X1 U10328 ( .A1(n8546), .A2(n9800), .B1(n8883), .B2(P1_U3086), .C1(
        n8882), .C2(n8891), .ZN(P1_U3326) );
  INV_X1 U10329 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8885) );
  OR2_X1 U10330 ( .A1(n10537), .A2(n8885), .ZN(n8886) );
  AOI21_X1 U10331 ( .B1(n8889), .B2(n4940), .A(n8888), .ZN(n8890) );
  INV_X1 U10332 ( .A(n8890), .ZN(P1_U3553) );
  OAI222_X1 U10333 ( .A1(n8546), .A2(n8894), .B1(n8893), .B2(P1_U3086), .C1(
        n8892), .C2(n8891), .ZN(P1_U3327) );
  OAI222_X1 U10334 ( .A1(n8897), .A2(P2_U3151), .B1(n9801), .B2(n8896), .C1(
        n8895), .C2(n9798), .ZN(P2_U3265) );
  INV_X1 U10335 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U10336 ( .A1(n10628), .A2(n8898), .ZN(n9541) );
  OAI21_X1 U10337 ( .B1(n10629), .B2(n8899), .A(n9541), .ZN(n8903) );
  NOR2_X1 U10338 ( .A1(n8901), .A2(n8900), .ZN(n8902) );
  AOI211_X1 U10339 ( .C1(n9651), .C2(n8904), .A(n8903), .B(n8902), .ZN(n8905)
         );
  OAI21_X1 U10340 ( .B1(n8906), .B2(n10632), .A(n8905), .ZN(P2_U3204) );
  AOI21_X1 U10341 ( .B1(n8907), .B2(n8908), .A(n9363), .ZN(n8910) );
  NAND2_X1 U10342 ( .A1(n8910), .A2(n8909), .ZN(n8915) );
  AOI22_X1 U10343 ( .A1(n9368), .A2(n9354), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8911) );
  OAI21_X1 U10344 ( .B1(n8912), .B2(n9358), .A(n8911), .ZN(n8913) );
  AOI21_X1 U10345 ( .B1(n9554), .B2(n9355), .A(n8913), .ZN(n8914) );
  OAI211_X1 U10346 ( .C1(n9677), .C2(n8930), .A(n8915), .B(n8914), .ZN(
        P2_U3154) );
  XNOR2_X1 U10347 ( .A(n8916), .B(n9371), .ZN(n8922) );
  AOI22_X1 U10348 ( .A1(n9354), .A2(n9372), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8918) );
  NAND2_X1 U10349 ( .A1(n9355), .A2(n9597), .ZN(n8917) );
  OAI211_X1 U10350 ( .C1(n9594), .C2(n9358), .A(n8918), .B(n8917), .ZN(n8919)
         );
  AOI21_X1 U10351 ( .B1(n8920), .B2(n9360), .A(n8919), .ZN(n8921) );
  OAI21_X1 U10352 ( .B1(n8922), .B2(n9363), .A(n8921), .ZN(P2_U3156) );
  INV_X1 U10353 ( .A(n9652), .ZN(n9785) );
  OAI211_X1 U10354 ( .C1(n8925), .C2(n8924), .A(n8923), .B(n9342), .ZN(n8929)
         );
  NAND2_X1 U10355 ( .A1(n9346), .A2(n9374), .ZN(n8926) );
  NAND2_X1 U10356 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9530) );
  OAI211_X1 U10357 ( .C1(n9645), .C2(n9327), .A(n8926), .B(n9530), .ZN(n8927)
         );
  AOI21_X1 U10358 ( .B1(n9650), .B2(n9355), .A(n8927), .ZN(n8928) );
  OAI211_X1 U10359 ( .C1(n9785), .C2(n8930), .A(n8929), .B(n8928), .ZN(
        P2_U3159) );
  XOR2_X1 U10360 ( .A(n8932), .B(n8931), .Z(n8938) );
  AOI22_X1 U10361 ( .A1(n9354), .A2(n9374), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8934) );
  NAND2_X1 U10362 ( .A1(n9355), .A2(n9621), .ZN(n8933) );
  OAI211_X1 U10363 ( .C1(n9616), .C2(n9358), .A(n8934), .B(n8933), .ZN(n8935)
         );
  AOI21_X1 U10364 ( .B1(n8936), .B2(n9360), .A(n8935), .ZN(n8937) );
  OAI21_X1 U10365 ( .B1(n8938), .B2(n9363), .A(n8937), .ZN(P2_U3163) );
  XOR2_X1 U10366 ( .A(n8940), .B(n8939), .Z(n8945) );
  AOI22_X1 U10367 ( .A1(n9368), .A2(n9346), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8942) );
  NAND2_X1 U10368 ( .A1(n9574), .A2(n9355), .ZN(n8941) );
  OAI211_X1 U10369 ( .C1(n9594), .C2(n9327), .A(n8942), .B(n8941), .ZN(n8943)
         );
  AOI21_X1 U10370 ( .B1(n9572), .B2(n9360), .A(n8943), .ZN(n8944) );
  OAI21_X1 U10371 ( .B1(n8945), .B2(n9363), .A(n8944), .ZN(n9302) );
  OAI22_X1 U10372 ( .A1(n9285), .A2(keyinput142), .B1(n8947), .B2(keyinput249), 
        .ZN(n8946) );
  AOI221_X1 U10373 ( .B1(n9285), .B2(keyinput142), .C1(keyinput249), .C2(n8947), .A(n8946), .ZN(n8956) );
  OAI22_X1 U10374 ( .A1(n9232), .A2(keyinput168), .B1(n10532), .B2(keyinput133), .ZN(n8948) );
  AOI221_X1 U10375 ( .B1(n9232), .B2(keyinput168), .C1(keyinput133), .C2(
        n10532), .A(n8948), .ZN(n8955) );
  INV_X1 U10376 ( .A(SI_5_), .ZN(n9277) );
  OAI22_X1 U10377 ( .A1(n9277), .A2(keyinput215), .B1(n9272), .B2(keyinput224), 
        .ZN(n8949) );
  AOI221_X1 U10378 ( .B1(n9277), .B2(keyinput215), .C1(keyinput224), .C2(n9272), .A(n8949), .ZN(n8954) );
  OAI22_X1 U10379 ( .A1(n8952), .A2(keyinput245), .B1(n8951), .B2(keyinput159), 
        .ZN(n8950) );
  AOI221_X1 U10380 ( .B1(n8952), .B2(keyinput245), .C1(keyinput159), .C2(n8951), .A(n8950), .ZN(n8953) );
  NAND4_X1 U10381 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n8984)
         );
  OAI22_X1 U10382 ( .A1(n9234), .A2(keyinput248), .B1(n10381), .B2(keyinput193), .ZN(n8957) );
  AOI221_X1 U10383 ( .B1(n9234), .B2(keyinput248), .C1(keyinput193), .C2(
        n10381), .A(n8957), .ZN(n8968) );
  OAI22_X1 U10384 ( .A1(n8959), .A2(keyinput200), .B1(n10631), .B2(keyinput243), .ZN(n8958) );
  AOI221_X1 U10385 ( .B1(n8959), .B2(keyinput200), .C1(keyinput243), .C2(
        n10631), .A(n8958), .ZN(n8967) );
  OAI22_X1 U10386 ( .A1(n8962), .A2(keyinput239), .B1(n8961), .B2(keyinput241), 
        .ZN(n8960) );
  AOI221_X1 U10387 ( .B1(n8962), .B2(keyinput239), .C1(keyinput241), .C2(n8961), .A(n8960), .ZN(n8966) );
  OAI22_X1 U10388 ( .A1(n8964), .A2(keyinput175), .B1(n9236), .B2(keyinput228), 
        .ZN(n8963) );
  AOI221_X1 U10389 ( .B1(n8964), .B2(keyinput175), .C1(keyinput228), .C2(n9236), .A(n8963), .ZN(n8965) );
  NAND4_X1 U10390 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n8983)
         );
  AOI22_X1 U10391 ( .A1(n6724), .A2(keyinput219), .B1(n8970), .B2(keyinput216), 
        .ZN(n8969) );
  OAI221_X1 U10392 ( .B1(n6724), .B2(keyinput219), .C1(n8970), .C2(keyinput216), .A(n8969), .ZN(n8982) );
  XOR2_X1 U10393 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput184), .Z(n8975) );
  XNOR2_X1 U10394 ( .A(n8971), .B(keyinput130), .ZN(n8974) );
  XOR2_X1 U10395 ( .A(SI_0_), .B(keyinput194), .Z(n8973) );
  INV_X1 U10396 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9434) );
  XNOR2_X1 U10397 ( .A(n9434), .B(keyinput254), .ZN(n8972) );
  NOR4_X1 U10398 ( .A1(n8975), .A2(n8974), .A3(n8973), .A4(n8972), .ZN(n8980)
         );
  INV_X1 U10399 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8978) );
  INV_X1 U10400 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8977) );
  OAI22_X1 U10401 ( .A1(n8978), .A2(keyinput234), .B1(n8977), .B2(keyinput145), 
        .ZN(n8976) );
  AOI221_X1 U10402 ( .B1(n8978), .B2(keyinput234), .C1(keyinput145), .C2(n8977), .A(n8976), .ZN(n8979) );
  NAND2_X1 U10403 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NOR4_X1 U10404 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n9117)
         );
  OAI22_X1 U10405 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(keyinput212), .B1(
        P1_REG2_REG_4__SCAN_IN), .B2(keyinput141), .ZN(n8985) );
  AOI221_X1 U10406 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput212), .C1(
        keyinput141), .C2(P1_REG2_REG_4__SCAN_IN), .A(n8985), .ZN(n8992) );
  OAI22_X1 U10407 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput162), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput163), .ZN(n8986) );
  AOI221_X1 U10408 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput162), .C1(
        keyinput163), .C2(P1_REG0_REG_7__SCAN_IN), .A(n8986), .ZN(n8991) );
  OAI22_X1 U10409 ( .A1(P2_D_REG_5__SCAN_IN), .A2(keyinput185), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput231), .ZN(n8987) );
  AOI221_X1 U10410 ( .B1(P2_D_REG_5__SCAN_IN), .B2(keyinput185), .C1(
        keyinput231), .C2(P1_D_REG_12__SCAN_IN), .A(n8987), .ZN(n8990) );
  OAI22_X1 U10411 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(keyinput220), .B1(
        keyinput181), .B2(P1_REG3_REG_1__SCAN_IN), .ZN(n8988) );
  AOI221_X1 U10412 ( .B1(P1_DATAO_REG_3__SCAN_IN), .B2(keyinput220), .C1(
        P1_REG3_REG_1__SCAN_IN), .C2(keyinput181), .A(n8988), .ZN(n8989) );
  NAND4_X1 U10413 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(n8989), .ZN(n9020)
         );
  OAI22_X1 U10414 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput154), .B1(
        keyinput152), .B2(P2_REG0_REG_18__SCAN_IN), .ZN(n8993) );
  AOI221_X1 U10415 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput154), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput152), .A(n8993), .ZN(n9000) );
  OAI22_X1 U10416 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(keyinput251), .B1(
        keyinput196), .B2(P1_REG1_REG_20__SCAN_IN), .ZN(n8994) );
  AOI221_X1 U10417 ( .B1(P2_IR_REG_26__SCAN_IN), .B2(keyinput251), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput196), .A(n8994), .ZN(n8999) );
  OAI22_X1 U10418 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput213), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput137), .ZN(n8995) );
  AOI221_X1 U10419 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput213), .C1(
        keyinput137), .C2(P1_D_REG_20__SCAN_IN), .A(n8995), .ZN(n8998) );
  OAI22_X1 U10420 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput191), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput235), .ZN(n8996) );
  AOI221_X1 U10421 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput191), .C1(
        keyinput235), .C2(P1_IR_REG_24__SCAN_IN), .A(n8996), .ZN(n8997) );
  NAND4_X1 U10422 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n9019)
         );
  OAI22_X1 U10423 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput236), .B1(
        P1_REG0_REG_20__SCAN_IN), .B2(keyinput203), .ZN(n9001) );
  AOI221_X1 U10424 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput236), .C1(
        keyinput203), .C2(P1_REG0_REG_20__SCAN_IN), .A(n9001), .ZN(n9008) );
  OAI22_X1 U10425 ( .A1(P2_REG0_REG_28__SCAN_IN), .A2(keyinput138), .B1(
        keyinput208), .B2(P1_REG0_REG_14__SCAN_IN), .ZN(n9002) );
  AOI221_X1 U10426 ( .B1(P2_REG0_REG_28__SCAN_IN), .B2(keyinput138), .C1(
        P1_REG0_REG_14__SCAN_IN), .C2(keyinput208), .A(n9002), .ZN(n9007) );
  OAI22_X1 U10427 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput244), .B1(
        keyinput204), .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9003) );
  AOI221_X1 U10428 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput244), .C1(
        P1_DATAO_REG_6__SCAN_IN), .C2(keyinput204), .A(n9003), .ZN(n9006) );
  OAI22_X1 U10429 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput164), .B1(
        P1_ADDR_REG_2__SCAN_IN), .B2(keyinput136), .ZN(n9004) );
  AOI221_X1 U10430 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput164), .C1(
        keyinput136), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9004), .ZN(n9005) );
  NAND4_X1 U10431 ( .A1(n9008), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n9018)
         );
  OAI22_X1 U10432 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(keyinput169), .B1(
        keyinput144), .B2(P2_REG2_REG_1__SCAN_IN), .ZN(n9009) );
  AOI221_X1 U10433 ( .B1(P2_REG0_REG_19__SCAN_IN), .B2(keyinput169), .C1(
        P2_REG2_REG_1__SCAN_IN), .C2(keyinput144), .A(n9009), .ZN(n9016) );
  OAI22_X1 U10434 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput214), .B1(
        keyinput188), .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9010) );
  AOI221_X1 U10435 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput214), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput188), .A(n9010), .ZN(n9015) );
  OAI22_X1 U10436 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(keyinput173), .B1(
        keyinput176), .B2(P1_REG1_REG_1__SCAN_IN), .ZN(n9011) );
  AOI221_X1 U10437 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(keyinput173), .C1(
        P1_REG1_REG_1__SCAN_IN), .C2(keyinput176), .A(n9011), .ZN(n9014) );
  OAI22_X1 U10438 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(keyinput172), .B1(
        keyinput178), .B2(P2_REG2_REG_13__SCAN_IN), .ZN(n9012) );
  AOI221_X1 U10439 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(keyinput172), .C1(
        P2_REG2_REG_13__SCAN_IN), .C2(keyinput178), .A(n9012), .ZN(n9013) );
  NAND4_X1 U10440 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n9017)
         );
  NOR4_X1 U10441 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n9116)
         );
  OAI22_X1 U10442 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput146), .B1(
        keyinput198), .B2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9021) );
  AOI221_X1 U10443 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput146), .C1(
        P1_ADDR_REG_5__SCAN_IN), .C2(keyinput198), .A(n9021), .ZN(n9028) );
  OAI22_X1 U10444 ( .A1(P2_REG1_REG_28__SCAN_IN), .A2(keyinput139), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput207), .ZN(n9022) );
  AOI221_X1 U10445 ( .B1(P2_REG1_REG_28__SCAN_IN), .B2(keyinput139), .C1(
        keyinput207), .C2(P1_REG0_REG_26__SCAN_IN), .A(n9022), .ZN(n9027) );
  OAI22_X1 U10446 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput158), .B1(
        keyinput153), .B2(SI_4_), .ZN(n9023) );
  AOI221_X1 U10447 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput158), .C1(
        SI_4_), .C2(keyinput153), .A(n9023), .ZN(n9026) );
  OAI22_X1 U10448 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(keyinput179), .B1(
        P2_D_REG_7__SCAN_IN), .B2(keyinput238), .ZN(n9024) );
  AOI221_X1 U10449 ( .B1(P2_IR_REG_21__SCAN_IN), .B2(keyinput179), .C1(
        keyinput238), .C2(P2_D_REG_7__SCAN_IN), .A(n9024), .ZN(n9025) );
  NAND4_X1 U10450 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n9056)
         );
  OAI22_X1 U10451 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput183), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(keyinput217), .ZN(n9029) );
  AOI221_X1 U10452 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput183), .C1(
        keyinput217), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9029), .ZN(n9036) );
  OAI22_X1 U10453 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput186), .B1(keyinput250), 
        .B2(P2_D_REG_12__SCAN_IN), .ZN(n9030) );
  AOI221_X1 U10454 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput186), .C1(
        P2_D_REG_12__SCAN_IN), .C2(keyinput250), .A(n9030), .ZN(n9035) );
  OAI22_X1 U10455 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput143), .B1(
        keyinput199), .B2(P1_IR_REG_12__SCAN_IN), .ZN(n9031) );
  AOI221_X1 U10456 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput143), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput199), .A(n9031), .ZN(n9034) );
  OAI22_X1 U10457 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput160), .B1(
        keyinput135), .B2(P1_D_REG_8__SCAN_IN), .ZN(n9032) );
  AOI221_X1 U10458 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput160), .C1(
        P1_D_REG_8__SCAN_IN), .C2(keyinput135), .A(n9032), .ZN(n9033) );
  NAND4_X1 U10459 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n9055)
         );
  OAI22_X1 U10460 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(keyinput166), .B1(
        keyinput177), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n9037) );
  AOI221_X1 U10461 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(keyinput166), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput177), .A(n9037), .ZN(n9044) );
  OAI22_X1 U10462 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(keyinput157), .B1(
        keyinput170), .B2(P1_REG1_REG_23__SCAN_IN), .ZN(n9038) );
  AOI221_X1 U10463 ( .B1(P2_REG1_REG_19__SCAN_IN), .B2(keyinput157), .C1(
        P1_REG1_REG_23__SCAN_IN), .C2(keyinput170), .A(n9038), .ZN(n9043) );
  OAI22_X1 U10464 ( .A1(P2_D_REG_31__SCAN_IN), .A2(keyinput171), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput165), .ZN(n9039) );
  AOI221_X1 U10465 ( .B1(P2_D_REG_31__SCAN_IN), .B2(keyinput171), .C1(
        keyinput165), .C2(P2_DATAO_REG_26__SCAN_IN), .A(n9039), .ZN(n9042) );
  OAI22_X1 U10466 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput197), .B1(
        P2_ADDR_REG_7__SCAN_IN), .B2(keyinput180), .ZN(n9040) );
  AOI221_X1 U10467 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput197), .C1(
        keyinput180), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n9040), .ZN(n9041) );
  NAND4_X1 U10468 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n9054)
         );
  OAI22_X1 U10469 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput149), .B1(
        keyinput190), .B2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9045) );
  AOI221_X1 U10470 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput149), .C1(
        P1_ADDR_REG_4__SCAN_IN), .C2(keyinput190), .A(n9045), .ZN(n9052) );
  OAI22_X1 U10471 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(keyinput232), .B1(
        P2_REG0_REG_22__SCAN_IN), .B2(keyinput252), .ZN(n9046) );
  AOI221_X1 U10472 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(keyinput232), .C1(
        keyinput252), .C2(P2_REG0_REG_22__SCAN_IN), .A(n9046), .ZN(n9051) );
  OAI22_X1 U10473 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput209), .B1(
        keyinput156), .B2(P1_REG2_REG_30__SCAN_IN), .ZN(n9047) );
  AOI221_X1 U10474 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput209), .C1(
        P1_REG2_REG_30__SCAN_IN), .C2(keyinput156), .A(n9047), .ZN(n9050) );
  OAI22_X1 U10475 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(keyinput218), .B1(
        keyinput131), .B2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9048) );
  AOI221_X1 U10476 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(keyinput218), .C1(
        P1_ADDR_REG_14__SCAN_IN), .C2(keyinput131), .A(n9048), .ZN(n9049) );
  NAND4_X1 U10477 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(n9053)
         );
  NOR4_X1 U10478 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n9115)
         );
  INV_X1 U10479 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9198) );
  AOI22_X1 U10480 ( .A1(n9198), .A2(keyinput223), .B1(keyinput229), .B2(n7577), 
        .ZN(n9057) );
  OAI221_X1 U10481 ( .B1(n9198), .B2(keyinput223), .C1(n7577), .C2(keyinput229), .A(n9057), .ZN(n9067) );
  AOI22_X1 U10482 ( .A1(n9059), .A2(keyinput255), .B1(n9192), .B2(keyinput247), 
        .ZN(n9058) );
  OAI221_X1 U10483 ( .B1(n9059), .B2(keyinput255), .C1(n9192), .C2(keyinput247), .A(n9058), .ZN(n9066) );
  AOI22_X1 U10484 ( .A1(n9062), .A2(keyinput237), .B1(n9061), .B2(keyinput129), 
        .ZN(n9060) );
  OAI221_X1 U10485 ( .B1(n9062), .B2(keyinput237), .C1(n9061), .C2(keyinput129), .A(n9060), .ZN(n9065) );
  INV_X1 U10486 ( .A(SI_10_), .ZN(n9275) );
  AOI22_X1 U10487 ( .A1(n9275), .A2(keyinput195), .B1(n9259), .B2(keyinput201), 
        .ZN(n9063) );
  OAI221_X1 U10488 ( .B1(n9275), .B2(keyinput195), .C1(n9259), .C2(keyinput201), .A(n9063), .ZN(n9064) );
  NOR4_X1 U10489 ( .A1(n9067), .A2(n9066), .A3(n9065), .A4(n9064), .ZN(n9113)
         );
  XNOR2_X1 U10490 ( .A(n10467), .B(keyinput233), .ZN(n9069) );
  INV_X1 U10491 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10391) );
  XNOR2_X1 U10492 ( .A(n10391), .B(keyinput132), .ZN(n9068) );
  NOR2_X1 U10493 ( .A1(n9069), .A2(n9068), .ZN(n9112) );
  AOI22_X1 U10494 ( .A1(P1_U3086), .A2(keyinput240), .B1(n5854), .B2(
        keyinput167), .ZN(n9070) );
  OAI221_X1 U10495 ( .B1(P1_U3086), .B2(keyinput240), .C1(n5854), .C2(
        keyinput167), .A(n9070), .ZN(n9074) );
  AOI22_X1 U10496 ( .A1(n7534), .A2(keyinput227), .B1(keyinput210), .B2(n10266), .ZN(n9071) );
  OAI221_X1 U10497 ( .B1(n7534), .B2(keyinput227), .C1(n10266), .C2(
        keyinput210), .A(n9071), .ZN(n9073) );
  INV_X1 U10498 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10464) );
  XNOR2_X1 U10499 ( .A(n10464), .B(keyinput206), .ZN(n9072) );
  NOR3_X1 U10500 ( .A1(n9074), .A2(n9073), .A3(n9072), .ZN(n9111) );
  AOI22_X1 U10501 ( .A1(n9076), .A2(keyinput221), .B1(keyinput226), .B2(n7423), 
        .ZN(n9075) );
  OAI221_X1 U10502 ( .B1(n9076), .B2(keyinput221), .C1(n7423), .C2(keyinput226), .A(n9075), .ZN(n9081) );
  AOI22_X1 U10503 ( .A1(n5771), .A2(keyinput192), .B1(n9206), .B2(keyinput187), 
        .ZN(n9077) );
  OAI221_X1 U10504 ( .B1(n5771), .B2(keyinput192), .C1(n9206), .C2(keyinput187), .A(n9077), .ZN(n9080) );
  AOI22_X1 U10505 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(keyinput148), .B1(
        P1_REG2_REG_31__SCAN_IN), .B2(keyinput211), .ZN(n9078) );
  OAI221_X1 U10506 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(keyinput148), .C1(
        P1_REG2_REG_31__SCAN_IN), .C2(keyinput211), .A(n9078), .ZN(n9079) );
  NOR3_X1 U10507 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9109) );
  AOI22_X1 U10508 ( .A1(n9241), .A2(keyinput189), .B1(keyinput155), .B2(n10302), .ZN(n9082) );
  OAI221_X1 U10509 ( .B1(n9241), .B2(keyinput189), .C1(n10302), .C2(
        keyinput155), .A(n9082), .ZN(n9088) );
  XNOR2_X1 U10510 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput222), .ZN(n9086) );
  XNOR2_X1 U10511 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput151), .ZN(n9085) );
  XNOR2_X1 U10512 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput128), .ZN(n9084) );
  XNOR2_X1 U10513 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput253), .ZN(n9083) );
  NAND4_X1 U10514 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9087)
         );
  NOR2_X1 U10515 ( .A1(n9088), .A2(n9087), .ZN(n9097) );
  INV_X1 U10516 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9090) );
  AOI22_X1 U10517 ( .A1(n9090), .A2(keyinput134), .B1(n9278), .B2(keyinput182), 
        .ZN(n9089) );
  OAI221_X1 U10518 ( .B1(n9090), .B2(keyinput134), .C1(n9278), .C2(keyinput182), .A(n9089), .ZN(n9095) );
  XNOR2_X1 U10519 ( .A(P1_REG0_REG_15__SCAN_IN), .B(keyinput230), .ZN(n9093)
         );
  XNOR2_X1 U10520 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput246), .ZN(n9092) );
  XNOR2_X1 U10521 ( .A(keyinput242), .B(P1_REG0_REG_3__SCAN_IN), .ZN(n9091) );
  NAND3_X1 U10522 ( .A1(n9093), .A2(n9092), .A3(n9091), .ZN(n9094) );
  NOR2_X1 U10523 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  AND2_X1 U10524 ( .A1(n9097), .A2(n9096), .ZN(n9108) );
  INV_X1 U10525 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10394) );
  INV_X1 U10526 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U10527 ( .A1(n10394), .A2(keyinput174), .B1(keyinput202), .B2(
        n10348), .ZN(n9098) );
  OAI221_X1 U10528 ( .B1(n10394), .B2(keyinput174), .C1(n10348), .C2(
        keyinput202), .A(n9098), .ZN(n9101) );
  INV_X1 U10529 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U10530 ( .A1(n10372), .A2(keyinput140), .B1(keyinput205), .B2(
        n10386), .ZN(n9099) );
  OAI221_X1 U10531 ( .B1(n10372), .B2(keyinput140), .C1(n10386), .C2(
        keyinput205), .A(n9099), .ZN(n9100) );
  NOR2_X1 U10532 ( .A1(n9101), .A2(n9100), .ZN(n9107) );
  INV_X1 U10533 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10640) );
  INV_X1 U10534 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U10535 ( .A1(n10640), .A2(keyinput147), .B1(keyinput225), .B2(
        n10400), .ZN(n9102) );
  OAI221_X1 U10536 ( .B1(n10640), .B2(keyinput147), .C1(n10400), .C2(
        keyinput225), .A(n9102), .ZN(n9105) );
  AOI22_X1 U10537 ( .A1(n9262), .A2(keyinput161), .B1(keyinput150), .B2(n10463), .ZN(n9103) );
  OAI221_X1 U10538 ( .B1(n9262), .B2(keyinput161), .C1(n10463), .C2(
        keyinput150), .A(n9103), .ZN(n9104) );
  NOR2_X1 U10539 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  AND4_X1 U10540 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n9110)
         );
  AND4_X1 U10541 ( .A1(n9113), .A2(n9112), .A3(n9111), .A4(n9110), .ZN(n9114)
         );
  NAND4_X1 U10542 ( .A1(n9117), .A2(n9116), .A3(n9115), .A4(n9114), .ZN(n9300)
         );
  OAI22_X1 U10543 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput50), .B1(
        keyinput6), .B2(P2_REG0_REG_7__SCAN_IN), .ZN(n9118) );
  AOI221_X1 U10544 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput50), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput6), .A(n9118), .ZN(n9125) );
  OAI22_X1 U10545 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(keyinput26), .B1(
        keyinput55), .B2(P2_REG1_REG_6__SCAN_IN), .ZN(n9119) );
  AOI221_X1 U10546 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(keyinput26), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput55), .A(n9119), .ZN(n9124) );
  OAI22_X1 U10547 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput1), .B1(
        keyinput108), .B2(P2_REG2_REG_23__SCAN_IN), .ZN(n9120) );
  AOI221_X1 U10548 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput1), .C1(
        P2_REG2_REG_23__SCAN_IN), .C2(keyinput108), .A(n9120), .ZN(n9123) );
  OAI22_X1 U10549 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput86), .B1(
        keyinput27), .B2(P1_REG0_REG_25__SCAN_IN), .ZN(n9121) );
  AOI221_X1 U10550 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput86), .C1(
        P1_REG0_REG_25__SCAN_IN), .C2(keyinput27), .A(n9121), .ZN(n9122) );
  NAND4_X1 U10551 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n9122), .ZN(n9153)
         );
  OAI22_X1 U10552 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(keyinput13), .B1(
        keyinput74), .B2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9126) );
  AOI221_X1 U10553 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(keyinput13), .C1(
        P1_ADDR_REG_3__SCAN_IN), .C2(keyinput74), .A(n9126), .ZN(n9133) );
  OAI22_X1 U10554 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(keyinput38), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(keyinput77), .ZN(n9127) );
  AOI221_X1 U10555 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(keyinput38), .C1(
        keyinput77), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9127), .ZN(n9132) );
  OAI22_X1 U10556 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(keyinput125), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput10), .ZN(n9128) );
  AOI221_X1 U10557 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(keyinput125), .C1(
        keyinput10), .C2(P2_REG0_REG_28__SCAN_IN), .A(n9128), .ZN(n9131) );
  OAI22_X1 U10558 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(keyinput84), .B1(
        keyinput64), .B2(P1_IR_REG_10__SCAN_IN), .ZN(n9129) );
  AOI221_X1 U10559 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput84), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput64), .A(n9129), .ZN(n9130) );
  NAND4_X1 U10560 ( .A1(n9133), .A2(n9132), .A3(n9131), .A4(n9130), .ZN(n9152)
         );
  OAI22_X1 U10561 ( .A1(SI_27_), .A2(keyinput127), .B1(keyinput41), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n9134) );
  AOI221_X1 U10562 ( .B1(SI_27_), .B2(keyinput127), .C1(
        P2_REG0_REG_19__SCAN_IN), .C2(keyinput41), .A(n9134), .ZN(n9141) );
  OAI22_X1 U10563 ( .A1(P1_D_REG_13__SCAN_IN), .A2(keyinput105), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput69), .ZN(n9135) );
  AOI221_X1 U10564 ( .B1(P1_D_REG_13__SCAN_IN), .B2(keyinput105), .C1(
        keyinput69), .C2(P1_IR_REG_27__SCAN_IN), .A(n9135), .ZN(n9140) );
  OAI22_X1 U10565 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput112), .B1(
        keyinput21), .B2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9136) );
  AOI221_X1 U10566 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput112), .C1(
        P1_DATAO_REG_31__SCAN_IN), .C2(keyinput21), .A(n9136), .ZN(n9139) );
  OAI22_X1 U10567 ( .A1(P2_REG0_REG_18__SCAN_IN), .A2(keyinput24), .B1(
        P1_D_REG_14__SCAN_IN), .B2(keyinput18), .ZN(n9137) );
  AOI221_X1 U10568 ( .B1(P2_REG0_REG_18__SCAN_IN), .B2(keyinput24), .C1(
        keyinput18), .C2(P1_D_REG_14__SCAN_IN), .A(n9137), .ZN(n9138) );
  NAND4_X1 U10569 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n9151)
         );
  OAI22_X1 U10570 ( .A1(P2_D_REG_5__SCAN_IN), .A2(keyinput57), .B1(keyinput45), 
        .B2(P1_REG3_REG_2__SCAN_IN), .ZN(n9142) );
  AOI221_X1 U10571 ( .B1(P2_D_REG_5__SCAN_IN), .B2(keyinput57), .C1(
        P1_REG3_REG_2__SCAN_IN), .C2(keyinput45), .A(n9142), .ZN(n9149) );
  OAI22_X1 U10572 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(keyinput47), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(keyinput3), .ZN(n9143) );
  AOI221_X1 U10573 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput47), .C1(
        keyinput3), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9143), .ZN(n9148) );
  OAI22_X1 U10574 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput113), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(keyinput4), .ZN(n9144) );
  AOI221_X1 U10575 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput113), .C1(
        keyinput4), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n9144), .ZN(n9147) );
  OAI22_X1 U10576 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput124), .B1(
        keyinput117), .B2(P1_REG3_REG_20__SCAN_IN), .ZN(n9145) );
  AOI221_X1 U10577 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput124), .C1(
        P1_REG3_REG_20__SCAN_IN), .C2(keyinput117), .A(n9145), .ZN(n9146) );
  NAND4_X1 U10578 ( .A1(n9149), .A2(n9148), .A3(n9147), .A4(n9146), .ZN(n9150)
         );
  NOR4_X1 U10579 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(n9299)
         );
  OAI22_X1 U10580 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput5), .B1(
        keyinput48), .B2(P1_REG1_REG_1__SCAN_IN), .ZN(n9154) );
  AOI221_X1 U10581 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput5), .C1(
        P1_REG1_REG_1__SCAN_IN), .C2(keyinput48), .A(n9154), .ZN(n9161) );
  OAI22_X1 U10582 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput2), .B1(keyinput44), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n9155) );
  AOI221_X1 U10583 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput2), .C1(
        P2_REG2_REG_16__SCAN_IN), .C2(keyinput44), .A(n9155), .ZN(n9160) );
  OAI22_X1 U10584 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput115), .B1(
        keyinput53), .B2(P1_REG3_REG_1__SCAN_IN), .ZN(n9156) );
  AOI221_X1 U10585 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput115), .C1(
        P1_REG3_REG_1__SCAN_IN), .C2(keyinput53), .A(n9156), .ZN(n9159) );
  OAI22_X1 U10586 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput22), .B1(
        P1_ADDR_REG_2__SCAN_IN), .B2(keyinput8), .ZN(n9157) );
  AOI221_X1 U10587 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput22), .C1(keyinput8), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9157), .ZN(n9158) );
  NAND4_X1 U10588 ( .A1(n9161), .A2(n9160), .A3(n9159), .A4(n9158), .ZN(n9189)
         );
  OAI22_X1 U10589 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput85), .B1(
        keyinput81), .B2(P1_REG0_REG_11__SCAN_IN), .ZN(n9162) );
  AOI221_X1 U10590 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput85), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput81), .A(n9162), .ZN(n9169) );
  OAI22_X1 U10591 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(keyinput91), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(keyinput46), .ZN(n9163) );
  AOI221_X1 U10592 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(keyinput91), .C1(
        keyinput46), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n9163), .ZN(n9168) );
  OAI22_X1 U10593 ( .A1(SI_0_), .A2(keyinput66), .B1(keyinput107), .B2(
        P1_IR_REG_24__SCAN_IN), .ZN(n9164) );
  AOI221_X1 U10594 ( .B1(SI_0_), .B2(keyinput66), .C1(P1_IR_REG_24__SCAN_IN), 
        .C2(keyinput107), .A(n9164), .ZN(n9167) );
  OAI22_X1 U10595 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput89), .B1(
        P2_ADDR_REG_18__SCAN_IN), .B2(keyinput20), .ZN(n9165) );
  AOI221_X1 U10596 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput89), .C1(
        keyinput20), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n9165), .ZN(n9166) );
  NAND4_X1 U10597 ( .A1(n9169), .A2(n9168), .A3(n9167), .A4(n9166), .ZN(n9188)
         );
  OAI22_X1 U10598 ( .A1(SI_22_), .A2(keyinput72), .B1(P1_DATAO_REG_10__SCAN_IN), .B2(keyinput88), .ZN(n9170) );
  AOI221_X1 U10599 ( .B1(SI_22_), .B2(keyinput72), .C1(keyinput88), .C2(
        P1_DATAO_REG_10__SCAN_IN), .A(n9170), .ZN(n9177) );
  OAI22_X1 U10600 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(keyinput29), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(keyinput65), .ZN(n9171) );
  AOI221_X1 U10601 ( .B1(P2_REG1_REG_19__SCAN_IN), .B2(keyinput29), .C1(
        keyinput65), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9171), .ZN(n9176) );
  OAI22_X1 U10602 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput98), .B1(
        keyinput49), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n9172) );
  AOI221_X1 U10603 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput98), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput49), .A(n9172), .ZN(n9175) );
  OAI22_X1 U10604 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput15), .B1(
        keyinput104), .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9173) );
  AOI221_X1 U10605 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput15), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput104), .A(n9173), .ZN(n9174) );
  NAND4_X1 U10606 ( .A1(n9177), .A2(n9176), .A3(n9175), .A4(n9174), .ZN(n9187)
         );
  OAI22_X1 U10607 ( .A1(SI_20_), .A2(keyinput121), .B1(P1_REG2_REG_10__SCAN_IN), .B2(keyinput31), .ZN(n9178) );
  AOI221_X1 U10608 ( .B1(SI_20_), .B2(keyinput121), .C1(keyinput31), .C2(
        P1_REG2_REG_10__SCAN_IN), .A(n9178), .ZN(n9185) );
  OAI22_X1 U10609 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput58), .B1(
        P1_REG0_REG_14__SCAN_IN), .B2(keyinput80), .ZN(n9179) );
  AOI221_X1 U10610 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput58), .C1(keyinput80), 
        .C2(P1_REG0_REG_14__SCAN_IN), .A(n9179), .ZN(n9184) );
  OAI22_X1 U10611 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput0), .B1(keyinput9), 
        .B2(P1_D_REG_20__SCAN_IN), .ZN(n9180) );
  AOI221_X1 U10612 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput0), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput9), .A(n9180), .ZN(n9183) );
  OAI22_X1 U10613 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(keyinput17), .B1(
        keyinput93), .B2(P2_REG1_REG_3__SCAN_IN), .ZN(n9181) );
  AOI221_X1 U10614 ( .B1(P2_REG0_REG_29__SCAN_IN), .B2(keyinput17), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput93), .A(n9181), .ZN(n9182) );
  NAND4_X1 U10615 ( .A1(n9185), .A2(n9184), .A3(n9183), .A4(n9182), .ZN(n9186)
         );
  NOR4_X1 U10616 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n9298)
         );
  AOI22_X1 U10617 ( .A1(n9192), .A2(keyinput119), .B1(keyinput43), .B2(n9191), 
        .ZN(n9190) );
  OAI221_X1 U10618 ( .B1(n9192), .B2(keyinput119), .C1(n9191), .C2(keyinput43), 
        .A(n9190), .ZN(n9201) );
  AOI22_X1 U10619 ( .A1(n9195), .A2(keyinput25), .B1(keyinput83), .B2(n9194), 
        .ZN(n9193) );
  OAI221_X1 U10620 ( .B1(n9195), .B2(keyinput25), .C1(n9194), .C2(keyinput83), 
        .A(n9193), .ZN(n9200) );
  AOI22_X1 U10621 ( .A1(n9198), .A2(keyinput95), .B1(n9197), .B2(keyinput30), 
        .ZN(n9196) );
  OAI221_X1 U10622 ( .B1(n9198), .B2(keyinput95), .C1(n9197), .C2(keyinput30), 
        .A(n9196), .ZN(n9199) );
  NOR3_X1 U10623 ( .A1(n9201), .A2(n9200), .A3(n9199), .ZN(n9222) );
  INV_X1 U10624 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10596) );
  INV_X1 U10625 ( .A(keyinput52), .ZN(n9202) );
  XNOR2_X1 U10626 ( .A(n10596), .B(n9202), .ZN(n9221) );
  AOI22_X1 U10627 ( .A1(n10298), .A2(keyinput79), .B1(n9204), .B2(keyinput122), 
        .ZN(n9203) );
  OAI221_X1 U10628 ( .B1(n10298), .B2(keyinput79), .C1(n9204), .C2(keyinput122), .A(n9203), .ZN(n9211) );
  AOI22_X1 U10629 ( .A1(n10320), .A2(keyinput75), .B1(n9206), .B2(keyinput59), 
        .ZN(n9205) );
  OAI221_X1 U10630 ( .B1(n10320), .B2(keyinput75), .C1(n9206), .C2(keyinput59), 
        .A(n9205), .ZN(n9210) );
  XNOR2_X1 U10631 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput92), .ZN(n9208) );
  XNOR2_X1 U10632 ( .A(P2_REG0_REG_27__SCAN_IN), .B(keyinput32), .ZN(n9207) );
  NAND2_X1 U10633 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  NOR3_X1 U10634 ( .A1(n9211), .A2(n9210), .A3(n9209), .ZN(n9220) );
  INV_X1 U10635 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9213) );
  AOI22_X1 U10636 ( .A1(n9214), .A2(keyinput76), .B1(keyinput28), .B2(n9213), 
        .ZN(n9212) );
  OAI221_X1 U10637 ( .B1(n9214), .B2(keyinput76), .C1(n9213), .C2(keyinput28), 
        .A(n9212), .ZN(n9218) );
  INV_X1 U10638 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9216) );
  AOI22_X1 U10639 ( .A1(n9216), .A2(keyinput114), .B1(n8162), .B2(keyinput36), 
        .ZN(n9215) );
  OAI221_X1 U10640 ( .B1(n9216), .B2(keyinput114), .C1(n8162), .C2(keyinput36), 
        .A(n9215), .ZN(n9217) );
  NOR2_X1 U10641 ( .A1(n9218), .A2(n9217), .ZN(n9219) );
  AND4_X1 U10642 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(n9256)
         );
  AOI22_X1 U10643 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput68), .ZN(n9223) );
  OAI221_X1 U10644 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput97), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput68), .A(n9223), .ZN(n9230) );
  AOI22_X1 U10645 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput102), .B1(
        P1_REG3_REG_21__SCAN_IN), .B2(keyinput90), .ZN(n9224) );
  OAI221_X1 U10646 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput102), .C1(
        P1_REG3_REG_21__SCAN_IN), .C2(keyinput90), .A(n9224), .ZN(n9229) );
  AOI22_X1 U10647 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(keyinput101), .B1(
        P2_REG1_REG_15__SCAN_IN), .B2(keyinput126), .ZN(n9225) );
  OAI221_X1 U10648 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(keyinput101), .C1(
        P2_REG1_REG_15__SCAN_IN), .C2(keyinput126), .A(n9225), .ZN(n9228) );
  AOI22_X1 U10649 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(keyinput42), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput109), .ZN(n9226) );
  OAI221_X1 U10650 ( .B1(P1_REG1_REG_23__SCAN_IN), .B2(keyinput42), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput109), .A(n9226), .ZN(n9227) );
  NOR4_X1 U10651 ( .A1(n9230), .A2(n9229), .A3(n9228), .A4(n9227), .ZN(n9255)
         );
  AOI22_X1 U10652 ( .A1(n9232), .A2(keyinput40), .B1(keyinput39), .B2(n5854), 
        .ZN(n9231) );
  OAI221_X1 U10653 ( .B1(n9232), .B2(keyinput40), .C1(n5854), .C2(keyinput39), 
        .A(n9231), .ZN(n9240) );
  INV_X1 U10654 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U10655 ( .A1(n10468), .A2(keyinput103), .B1(n9234), .B2(keyinput120), .ZN(n9233) );
  OAI221_X1 U10656 ( .B1(n10468), .B2(keyinput103), .C1(n9234), .C2(
        keyinput120), .A(n9233), .ZN(n9239) );
  INV_X1 U10657 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9237) );
  AOI22_X1 U10658 ( .A1(n9237), .A2(keyinput35), .B1(n9236), .B2(keyinput100), 
        .ZN(n9235) );
  OAI221_X1 U10659 ( .B1(n9237), .B2(keyinput35), .C1(n9236), .C2(keyinput100), 
        .A(n9235), .ZN(n9238) );
  NOR3_X1 U10660 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(n9254) );
  XNOR2_X1 U10661 ( .A(n9241), .B(keyinput61), .ZN(n9252) );
  XNOR2_X1 U10662 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput11), .ZN(n9245) );
  XNOR2_X1 U10663 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput94), .ZN(n9244) );
  XNOR2_X1 U10664 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput56), .ZN(n9243) );
  XNOR2_X1 U10665 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput111), .ZN(n9242)
         );
  NAND4_X1 U10666 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(n9251)
         );
  XNOR2_X1 U10667 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput118), .ZN(n9249) );
  XNOR2_X1 U10668 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput123), .ZN(n9248) );
  XNOR2_X1 U10669 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput23), .ZN(n9247) );
  XNOR2_X1 U10670 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput71), .ZN(n9246) );
  NAND4_X1 U10671 ( .A1(n9249), .A2(n9248), .A3(n9247), .A4(n9246), .ZN(n9250)
         );
  NOR3_X1 U10672 ( .A1(n9252), .A2(n9251), .A3(n9250), .ZN(n9253) );
  AND4_X1 U10673 ( .A1(n9256), .A2(n9255), .A3(n9254), .A4(n9253), .ZN(n9296)
         );
  AOI22_X1 U10674 ( .A1(n9259), .A2(keyinput73), .B1(keyinput37), .B2(n9258), 
        .ZN(n9257) );
  OAI221_X1 U10675 ( .B1(n9259), .B2(keyinput73), .C1(n9258), .C2(keyinput37), 
        .A(n9257), .ZN(n9267) );
  AOI22_X1 U10676 ( .A1(n5256), .A2(keyinput116), .B1(keyinput16), .B2(n10541), 
        .ZN(n9260) );
  OAI221_X1 U10677 ( .B1(n5256), .B2(keyinput116), .C1(n10541), .C2(keyinput16), .A(n9260), .ZN(n9266) );
  AOI22_X1 U10678 ( .A1(n10640), .A2(keyinput19), .B1(n9262), .B2(keyinput33), 
        .ZN(n9261) );
  OAI221_X1 U10679 ( .B1(n10640), .B2(keyinput19), .C1(n9262), .C2(keyinput33), 
        .A(n9261), .ZN(n9265) );
  INV_X1 U10680 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U10681 ( .A1(n10361), .A2(keyinput70), .B1(n10266), .B2(keyinput82), 
        .ZN(n9263) );
  OAI221_X1 U10682 ( .B1(n10361), .B2(keyinput70), .C1(n10266), .C2(keyinput82), .A(n9263), .ZN(n9264) );
  NOR4_X1 U10683 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n9295)
         );
  AOI22_X1 U10684 ( .A1(n9270), .A2(keyinput110), .B1(keyinput60), .B2(n9269), 
        .ZN(n9268) );
  OAI221_X1 U10685 ( .B1(n9270), .B2(keyinput110), .C1(n9269), .C2(keyinput60), 
        .A(n9268), .ZN(n9282) );
  INV_X1 U10686 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9273) );
  AOI22_X1 U10687 ( .A1(n9273), .A2(keyinput63), .B1(keyinput96), .B2(n9272), 
        .ZN(n9271) );
  OAI221_X1 U10688 ( .B1(n9273), .B2(keyinput63), .C1(n9272), .C2(keyinput96), 
        .A(n9271), .ZN(n9281) );
  AOI22_X1 U10689 ( .A1(n10372), .A2(keyinput12), .B1(n9275), .B2(keyinput67), 
        .ZN(n9274) );
  OAI221_X1 U10690 ( .B1(n10372), .B2(keyinput12), .C1(n9275), .C2(keyinput67), 
        .A(n9274), .ZN(n9280) );
  AOI22_X1 U10691 ( .A1(n9278), .A2(keyinput54), .B1(keyinput87), .B2(n9277), 
        .ZN(n9276) );
  OAI221_X1 U10692 ( .B1(n9278), .B2(keyinput54), .C1(n9277), .C2(keyinput87), 
        .A(n9276), .ZN(n9279) );
  NOR4_X1 U10693 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(n9294)
         );
  AOI22_X1 U10694 ( .A1(P1_D_REG_24__SCAN_IN), .A2(keyinput78), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput106), .ZN(n9283) );
  OAI221_X1 U10695 ( .B1(P1_D_REG_24__SCAN_IN), .B2(keyinput78), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput106), .A(n9283), .ZN(n9292) );
  AOI22_X1 U10696 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput7), .B1(n9285), .B2(
        keyinput14), .ZN(n9284) );
  OAI221_X1 U10697 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput7), .C1(n9285), 
        .C2(keyinput14), .A(n9284), .ZN(n9291) );
  AOI22_X1 U10698 ( .A1(n10357), .A2(keyinput62), .B1(n5774), .B2(keyinput34), 
        .ZN(n9286) );
  OAI221_X1 U10699 ( .B1(n10357), .B2(keyinput62), .C1(n5774), .C2(keyinput34), 
        .A(n9286), .ZN(n9290) );
  INV_X1 U10700 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9288) );
  AOI22_X1 U10701 ( .A1(n7534), .A2(keyinput99), .B1(n9288), .B2(keyinput51), 
        .ZN(n9287) );
  OAI221_X1 U10702 ( .B1(n7534), .B2(keyinput99), .C1(n9288), .C2(keyinput51), 
        .A(n9287), .ZN(n9289) );
  NOR4_X1 U10703 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n9293)
         );
  AND4_X1 U10704 ( .A1(n9296), .A2(n9295), .A3(n9294), .A4(n9293), .ZN(n9297)
         );
  NAND4_X1 U10705 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9301)
         );
  XNOR2_X1 U10706 ( .A(n9302), .B(n9301), .ZN(P2_U3165) );
  AOI21_X1 U10707 ( .B1(n9304), .B2(n9303), .A(n9340), .ZN(n9305) );
  OR2_X1 U10708 ( .A1(n9305), .A2(n9363), .ZN(n9313) );
  INV_X1 U10709 ( .A(n9306), .ZN(n9307) );
  AOI21_X1 U10710 ( .B1(n9360), .B2(n9308), .A(n9307), .ZN(n9312) );
  AOI22_X1 U10711 ( .A1(n9354), .A2(n5305), .B1(n9346), .B2(n9385), .ZN(n9311)
         );
  NAND2_X1 U10712 ( .A1(n9355), .A2(n9309), .ZN(n9310) );
  NAND4_X1 U10713 ( .A1(n9313), .A2(n9312), .A3(n9311), .A4(n9310), .ZN(
        P2_U3167) );
  XOR2_X1 U10714 ( .A(n9315), .B(n9314), .Z(n9320) );
  AOI22_X1 U10715 ( .A1(n9369), .A2(n9346), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n9317) );
  NAND2_X1 U10716 ( .A1(n9355), .A2(n9585), .ZN(n9316) );
  OAI211_X1 U10717 ( .C1(n9604), .C2(n9327), .A(n9317), .B(n9316), .ZN(n9318)
         );
  AOI21_X1 U10718 ( .B1(n9580), .B2(n9360), .A(n9318), .ZN(n9319) );
  OAI21_X1 U10719 ( .B1(n9320), .B2(n9363), .A(n9319), .ZN(P2_U3169) );
  INV_X1 U10720 ( .A(n9321), .ZN(n9322) );
  AOI21_X1 U10721 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9330) );
  INV_X1 U10722 ( .A(n9631), .ZN(n9373) );
  AOI22_X1 U10723 ( .A1(n9346), .A2(n9373), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n9326) );
  NAND2_X1 U10724 ( .A1(n9355), .A2(n9635), .ZN(n9325) );
  OAI211_X1 U10725 ( .C1(n9630), .C2(n9327), .A(n9326), .B(n9325), .ZN(n9328)
         );
  AOI21_X1 U10726 ( .B1(n9634), .B2(n9360), .A(n9328), .ZN(n9329) );
  OAI21_X1 U10727 ( .B1(n9330), .B2(n9363), .A(n9329), .ZN(P2_U3173) );
  XNOR2_X1 U10728 ( .A(n9331), .B(n9372), .ZN(n9336) );
  AOI22_X1 U10729 ( .A1(n9354), .A2(n9373), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9333) );
  NAND2_X1 U10730 ( .A1(n9355), .A2(n9608), .ZN(n9332) );
  OAI211_X1 U10731 ( .C1(n9604), .C2(n9358), .A(n9333), .B(n9332), .ZN(n9334)
         );
  AOI21_X1 U10732 ( .B1(n9607), .B2(n9360), .A(n9334), .ZN(n9335) );
  OAI21_X1 U10733 ( .B1(n9336), .B2(n9363), .A(n9335), .ZN(P2_U3175) );
  INV_X1 U10734 ( .A(n9337), .ZN(n9343) );
  OAI21_X1 U10735 ( .B1(n9340), .B2(n9339), .A(n9338), .ZN(n9341) );
  NAND3_X1 U10736 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n9351) );
  AOI21_X1 U10737 ( .B1(n9360), .B2(n9345), .A(n9344), .ZN(n9350) );
  AOI22_X1 U10738 ( .A1(n9354), .A2(n9386), .B1(n9346), .B2(n9384), .ZN(n9349)
         );
  NAND2_X1 U10739 ( .A1(n9355), .A2(n9347), .ZN(n9348) );
  NAND4_X1 U10740 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(
        P2_U3179) );
  XOR2_X1 U10741 ( .A(n9353), .B(n9352), .Z(n9364) );
  AOI22_X1 U10742 ( .A1(n9369), .A2(n9354), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9357) );
  NAND2_X1 U10743 ( .A1(n9565), .A2(n9355), .ZN(n9356) );
  OAI211_X1 U10744 ( .C1(n9562), .C2(n9358), .A(n9357), .B(n9356), .ZN(n9359)
         );
  AOI21_X1 U10745 ( .B1(n9361), .B2(n9360), .A(n9359), .ZN(n9362) );
  OAI21_X1 U10746 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(P2_U3180) );
  MUX2_X1 U10747 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9540), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10748 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9365), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10749 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9366), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10750 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9367), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10751 ( .A(n9368), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9500), .Z(
        P2_U3517) );
  MUX2_X1 U10752 ( .A(n9369), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9500), .Z(
        P2_U3516) );
  MUX2_X1 U10753 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9370), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10754 ( .A(n9371), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9500), .Z(
        P2_U3514) );
  MUX2_X1 U10755 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9372), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10756 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9373), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10757 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9374), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10758 ( .A(n9375), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9500), .Z(
        P2_U3510) );
  MUX2_X1 U10759 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9376), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10760 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9377), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10761 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8240), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10762 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9378), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10763 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9379), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10764 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9380), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10765 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9381), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10766 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9382), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10767 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n4672), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10768 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9383), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10769 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9384), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10770 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9385), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10771 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9386), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10772 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n5305), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10773 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9726), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10774 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9387), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10775 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9725), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10776 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n5679), .S(P2_U3893), .Z(
        P2_U3491) );
  NAND2_X1 U10777 ( .A1(n9405), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9388) );
  NOR2_X1 U10778 ( .A1(n9409), .A2(n9390), .ZN(n9391) );
  INV_X1 U10779 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10605) );
  NOR2_X1 U10780 ( .A1(n10605), .A2(n10604), .ZN(n10603) );
  XNOR2_X1 U10781 ( .A(n9433), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9392) );
  NOR2_X1 U10782 ( .A1(n9393), .A2(n9392), .ZN(n9432) );
  AOI21_X1 U10783 ( .B1(n9393), .B2(n9392), .A(n9432), .ZN(n9421) );
  MUX2_X1 U10784 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9521), .Z(n9425) );
  XNOR2_X1 U10785 ( .A(n9419), .B(n9425), .ZN(n9400) );
  MUX2_X1 U10786 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9521), .Z(n9394) );
  OR2_X1 U10787 ( .A1(n9394), .A2(n9410), .ZN(n9398) );
  XNOR2_X1 U10788 ( .A(n9409), .B(n9394), .ZN(n10610) );
  OR2_X1 U10789 ( .A1(n9395), .A2(n9405), .ZN(n9397) );
  NAND2_X1 U10790 ( .A1(n9397), .A2(n9396), .ZN(n10609) );
  NAND2_X1 U10791 ( .A1(n10610), .A2(n10609), .ZN(n10608) );
  NAND2_X1 U10792 ( .A1(n9398), .A2(n10608), .ZN(n9399) );
  NAND2_X1 U10793 ( .A1(n9400), .A2(n9399), .ZN(n9426) );
  OAI21_X1 U10794 ( .B1(n9400), .B2(n9399), .A(n9426), .ZN(n9403) );
  AND2_X1 U10795 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9402) );
  AOI21_X1 U10796 ( .B1(n10612), .B2(n9403), .A(n9402), .ZN(n9404) );
  OAI21_X1 U10797 ( .B1(n10597), .B2(n10391), .A(n9404), .ZN(n9418) );
  NAND2_X1 U10798 ( .A1(n9405), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9406) );
  NOR2_X1 U10799 ( .A1(n9409), .A2(n9408), .ZN(n9412) );
  INV_X1 U10800 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10602) );
  NOR2_X1 U10801 ( .A1(n10602), .A2(n10601), .ZN(n10600) );
  INV_X1 U10802 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9413) );
  AOI22_X1 U10803 ( .A1(n9419), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9413), .B2(
        n9433), .ZN(n9414) );
  NOR2_X1 U10804 ( .A1(n9415), .A2(n9414), .ZN(n9422) );
  AOI21_X1 U10805 ( .B1(n9415), .B2(n9414), .A(n9422), .ZN(n9416) );
  NOR2_X1 U10806 ( .A1(n9416), .A2(n10615), .ZN(n9417) );
  AOI211_X1 U10807 ( .C1(n10586), .C2(n9419), .A(n9418), .B(n9417), .ZN(n9420)
         );
  OAI21_X1 U10808 ( .B1(n9421), .B2(n10606), .A(n9420), .ZN(P2_U3196) );
  AOI21_X1 U10809 ( .B1(n9424), .B2(n9423), .A(n9457), .ZN(n9441) );
  MUX2_X1 U10810 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9521), .Z(n9447) );
  XNOR2_X1 U10811 ( .A(n9456), .B(n9447), .ZN(n9429) );
  OR2_X1 U10812 ( .A1(n9425), .A2(n9433), .ZN(n9427) );
  NAND2_X1 U10813 ( .A1(n9427), .A2(n9426), .ZN(n9428) );
  NAND2_X1 U10814 ( .A1(n9429), .A2(n9428), .ZN(n9448) );
  OAI21_X1 U10815 ( .B1(n9429), .B2(n9428), .A(n9448), .ZN(n9439) );
  INV_X1 U10816 ( .A(n9430), .ZN(n9431) );
  OAI21_X1 U10817 ( .B1(n10597), .B2(n10394), .A(n9431), .ZN(n9438) );
  AOI21_X1 U10818 ( .B1(n9435), .B2(n9434), .A(n9443), .ZN(n9436) );
  OAI22_X1 U10819 ( .A1(n10598), .A2(n9446), .B1(n9436), .B2(n10606), .ZN(
        n9437) );
  AOI211_X1 U10820 ( .C1(n10612), .C2(n9439), .A(n9438), .B(n9437), .ZN(n9440)
         );
  OAI21_X1 U10821 ( .B1(n9441), .B2(n10615), .A(n9440), .ZN(P2_U3197) );
  NOR2_X1 U10822 ( .A1(n9456), .A2(n9442), .ZN(n9444) );
  XNOR2_X1 U10823 ( .A(n9475), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9445) );
  AOI21_X1 U10824 ( .B1(n4605), .B2(n9445), .A(n9474), .ZN(n9465) );
  INV_X1 U10825 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10396) );
  MUX2_X1 U10826 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9521), .Z(n9469) );
  XNOR2_X1 U10827 ( .A(n9469), .B(n9463), .ZN(n9451) );
  OR2_X1 U10828 ( .A1(n9447), .A2(n9446), .ZN(n9449) );
  NAND2_X1 U10829 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  NAND2_X1 U10830 ( .A1(n9451), .A2(n9450), .ZN(n9470) );
  OAI21_X1 U10831 ( .B1(n9451), .B2(n9450), .A(n9470), .ZN(n9453) );
  AOI21_X1 U10832 ( .B1(n10612), .B2(n9453), .A(n9452), .ZN(n9454) );
  OAI21_X1 U10833 ( .B1(n10597), .B2(n10396), .A(n9454), .ZN(n9462) );
  NOR2_X1 U10834 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  AOI22_X1 U10835 ( .A1(n9463), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n4909), .B2(
        n9475), .ZN(n9459) );
  AOI21_X1 U10836 ( .B1(n4597), .B2(n9459), .A(n9466), .ZN(n9460) );
  NOR2_X1 U10837 ( .A1(n9460), .A2(n10615), .ZN(n9461) );
  AOI211_X1 U10838 ( .C1(n10586), .C2(n9463), .A(n9462), .B(n9461), .ZN(n9464)
         );
  OAI21_X1 U10839 ( .B1(n9465), .B2(n10606), .A(n9464), .ZN(P2_U3198) );
  INV_X1 U10840 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9468) );
  AOI21_X1 U10841 ( .B1(n9468), .B2(n9467), .A(n9509), .ZN(n9487) );
  MUX2_X1 U10842 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9521), .Z(n9495) );
  XNOR2_X1 U10843 ( .A(n9495), .B(n9507), .ZN(n9473) );
  OR2_X1 U10844 ( .A1(n9469), .A2(n9475), .ZN(n9471) );
  NAND2_X1 U10845 ( .A1(n9471), .A2(n9470), .ZN(n9472) );
  NAND2_X1 U10846 ( .A1(n9473), .A2(n9472), .ZN(n9493) );
  OAI21_X1 U10847 ( .B1(n9473), .B2(n9472), .A(n9493), .ZN(n9482) );
  NOR2_X1 U10848 ( .A1(n9476), .A2(n9477), .ZN(n9489) );
  INV_X1 U10849 ( .A(n9489), .ZN(n9479) );
  AOI21_X1 U10850 ( .B1(n9479), .B2(n9478), .A(n10606), .ZN(n9480) );
  AOI21_X1 U10851 ( .B1(n10586), .B2(n9507), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10852 ( .B1(n9487), .B2(n10615), .A(n9486), .ZN(P2_U3199) );
  NOR2_X1 U10853 ( .A1(n9507), .A2(n9488), .ZN(n9490) );
  NAND2_X1 U10854 ( .A1(n9525), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9516) );
  OAI21_X1 U10855 ( .B1(n9525), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9516), .ZN(
        n9491) );
  AOI21_X1 U10856 ( .B1(n9492), .B2(n9491), .A(n9518), .ZN(n9515) );
  OAI21_X1 U10857 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9498) );
  INV_X1 U10858 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9713) );
  MUX2_X1 U10859 ( .A(n9496), .B(n9713), .S(n9521), .Z(n9497) );
  NOR2_X1 U10860 ( .A1(n9498), .A2(n9497), .ZN(n9526) );
  INV_X1 U10861 ( .A(n9526), .ZN(n9499) );
  NAND2_X1 U10862 ( .A1(n9498), .A2(n9497), .ZN(n9524) );
  NAND2_X1 U10863 ( .A1(n9499), .A2(n9524), .ZN(n9501) );
  OAI21_X1 U10864 ( .B1(n9500), .B2(n9501), .A(n10598), .ZN(n9513) );
  INV_X1 U10865 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10404) );
  INV_X1 U10866 ( .A(n9501), .ZN(n9502) );
  NOR2_X1 U10867 ( .A1(n9502), .A2(n9514), .ZN(n9505) );
  INV_X1 U10868 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9503) );
  NOR2_X1 U10869 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9503), .ZN(n9504) );
  NOR2_X1 U10870 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  NAND2_X1 U10871 ( .A1(n9525), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9519) );
  OAI21_X1 U10872 ( .B1(n9525), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9519), .ZN(
        n9510) );
  AOI21_X1 U10873 ( .B1(n4575), .B2(n9511), .A(n10615), .ZN(n9512) );
  XNOR2_X1 U10874 ( .A(n5694), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9522) );
  INV_X1 U10875 ( .A(n9516), .ZN(n9517) );
  XNOR2_X1 U10876 ( .A(n5694), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n9523) );
  NOR2_X1 U10877 ( .A1(n10598), .A2(n5694), .ZN(n9534) );
  INV_X1 U10878 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n9532) );
  MUX2_X1 U10879 ( .A(n9523), .B(n9522), .S(n9521), .Z(n9528) );
  OAI21_X1 U10880 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  XOR2_X1 U10881 ( .A(n9528), .B(n9527), .Z(n9529) );
  NAND2_X1 U10882 ( .A1(n9529), .A2(n10612), .ZN(n9531) );
  OAI211_X1 U10883 ( .C1(n10597), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9533)
         );
  AOI211_X2 U10884 ( .C1(n9535), .C2(n10566), .A(n9534), .B(n9533), .ZN(n9536)
         );
  INV_X1 U10885 ( .A(n9538), .ZN(n9539) );
  NAND2_X1 U10886 ( .A1(n9540), .A2(n9539), .ZN(n9747) );
  OAI21_X1 U10887 ( .B1(n10632), .B2(n9747), .A(n9541), .ZN(n9543) );
  AOI21_X1 U10888 ( .B1(n10632), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9543), .ZN(
        n9542) );
  OAI21_X1 U10889 ( .B1(n9662), .B2(n9637), .A(n9542), .ZN(P2_U3202) );
  AOI21_X1 U10890 ( .B1(n10632), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9543), .ZN(
        n9544) );
  OAI21_X1 U10891 ( .B1(n9665), .B2(n9637), .A(n9544), .ZN(P2_U3203) );
  INV_X1 U10892 ( .A(n9545), .ZN(n9552) );
  AOI22_X1 U10893 ( .A1(n10632), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n10628), 
        .B2(n9546), .ZN(n9547) );
  OAI21_X1 U10894 ( .B1(n9548), .B2(n9637), .A(n9547), .ZN(n9549) );
  AOI21_X1 U10895 ( .B1(n9550), .B2(n9657), .A(n9549), .ZN(n9551) );
  OAI21_X1 U10896 ( .B1(n9552), .B2(n10632), .A(n9551), .ZN(P2_U3205) );
  INV_X1 U10897 ( .A(n9553), .ZN(n9559) );
  AOI22_X1 U10898 ( .A1(n9554), .A2(n10628), .B1(n10632), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9555) );
  OAI21_X1 U10899 ( .B1(n9677), .B2(n9637), .A(n9555), .ZN(n9556) );
  AOI21_X1 U10900 ( .B1(n9557), .B2(n9657), .A(n9556), .ZN(n9558) );
  OAI21_X1 U10901 ( .B1(n9559), .B2(n10632), .A(n9558), .ZN(P2_U3206) );
  XNOR2_X1 U10902 ( .A(n9560), .B(n9563), .ZN(n9561) );
  OAI222_X1 U10903 ( .A1(n9644), .A2(n9583), .B1(n9646), .B2(n9562), .C1(n9642), .C2(n9561), .ZN(n9678) );
  INV_X1 U10904 ( .A(n9678), .ZN(n9569) );
  XNOR2_X1 U10905 ( .A(n9564), .B(n9563), .ZN(n9679) );
  AOI22_X1 U10906 ( .A1(n9565), .A2(n10628), .B1(n10632), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9566) );
  OAI21_X1 U10907 ( .B1(n9757), .B2(n9637), .A(n9566), .ZN(n9567) );
  AOI21_X1 U10908 ( .B1(n9679), .B2(n9657), .A(n9567), .ZN(n9568) );
  OAI21_X1 U10909 ( .B1(n9569), .B2(n10632), .A(n9568), .ZN(P2_U3207) );
  INV_X1 U10910 ( .A(n10622), .ZN(n9573) );
  OAI222_X1 U10911 ( .A1(n9644), .A2(n9594), .B1(n9646), .B2(n9571), .C1(n9570), .C2(n9642), .ZN(n9682) );
  AOI21_X1 U10912 ( .B1(n9573), .B2(n9572), .A(n9682), .ZN(n9579) );
  AOI22_X1 U10913 ( .A1(n9574), .A2(n10628), .B1(n10632), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U10914 ( .A(n9576), .B(n9575), .ZN(n9683) );
  NAND2_X1 U10915 ( .A1(n9683), .A2(n9657), .ZN(n9577) );
  OAI211_X1 U10916 ( .C1(n9579), .C2(n10632), .A(n9578), .B(n9577), .ZN(
        P2_U3208) );
  INV_X1 U10917 ( .A(n9580), .ZN(n9765) );
  NOR2_X1 U10918 ( .A1(n9765), .A2(n10622), .ZN(n9584) );
  XNOR2_X1 U10919 ( .A(n9581), .B(n9589), .ZN(n9582) );
  OAI222_X1 U10920 ( .A1(n9646), .A2(n9583), .B1(n9644), .B2(n9604), .C1(n9582), .C2(n9642), .ZN(n9686) );
  AOI211_X1 U10921 ( .C1(n10628), .C2(n9585), .A(n9584), .B(n9686), .ZN(n9591)
         );
  NAND2_X1 U10922 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  XOR2_X1 U10923 ( .A(n9589), .B(n9588), .Z(n9687) );
  AOI22_X1 U10924 ( .A1(n9687), .A2(n9657), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10632), .ZN(n9590) );
  OAI21_X1 U10925 ( .B1(n9591), .B2(n10632), .A(n9590), .ZN(P2_U3209) );
  XOR2_X1 U10926 ( .A(n9595), .B(n9592), .Z(n9593) );
  OAI222_X1 U10927 ( .A1(n9646), .A2(n9594), .B1(n9644), .B2(n9616), .C1(n9642), .C2(n9593), .ZN(n9690) );
  INV_X1 U10928 ( .A(n9690), .ZN(n9601) );
  XOR2_X1 U10929 ( .A(n9596), .B(n9595), .Z(n9691) );
  AOI22_X1 U10930 ( .A1(n10632), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n10628), 
        .B2(n9597), .ZN(n9598) );
  OAI21_X1 U10931 ( .B1(n9769), .B2(n9637), .A(n9598), .ZN(n9599) );
  AOI21_X1 U10932 ( .B1(n9691), .B2(n9657), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10933 ( .B1(n9601), .B2(n10632), .A(n9600), .ZN(P2_U3210) );
  XNOR2_X1 U10934 ( .A(n9602), .B(n9605), .ZN(n9603) );
  OAI222_X1 U10935 ( .A1(n9646), .A2(n9604), .B1(n9644), .B2(n9631), .C1(n9642), .C2(n9603), .ZN(n9694) );
  INV_X1 U10936 ( .A(n9694), .ZN(n9612) );
  XNOR2_X1 U10937 ( .A(n9606), .B(n9605), .ZN(n9695) );
  INV_X1 U10938 ( .A(n9607), .ZN(n9773) );
  AOI22_X1 U10939 ( .A1(n10632), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n10628), 
        .B2(n9608), .ZN(n9609) );
  OAI21_X1 U10940 ( .B1(n9773), .B2(n9637), .A(n9609), .ZN(n9610) );
  AOI21_X1 U10941 ( .B1(n9695), .B2(n9657), .A(n9610), .ZN(n9611) );
  OAI21_X1 U10942 ( .B1(n9612), .B2(n10632), .A(n9611), .ZN(P2_U3211) );
  XNOR2_X1 U10943 ( .A(n9614), .B(n9613), .ZN(n9615) );
  OAI222_X1 U10944 ( .A1(n9646), .A2(n9616), .B1(n9644), .B2(n9647), .C1(n9642), .C2(n9615), .ZN(n9698) );
  INV_X1 U10945 ( .A(n9698), .ZN(n9625) );
  NOR2_X1 U10946 ( .A1(n9618), .A2(n4702), .ZN(n9620) );
  XNOR2_X1 U10947 ( .A(n9620), .B(n9619), .ZN(n9699) );
  AOI22_X1 U10948 ( .A1(n10632), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n10628), 
        .B2(n9621), .ZN(n9622) );
  OAI21_X1 U10949 ( .B1(n9777), .B2(n9637), .A(n9622), .ZN(n9623) );
  AOI21_X1 U10950 ( .B1(n9699), .B2(n9657), .A(n9623), .ZN(n9624) );
  OAI21_X1 U10951 ( .B1(n9625), .B2(n10632), .A(n9624), .ZN(P2_U3212) );
  OAI21_X1 U10952 ( .B1(n9627), .B2(n9632), .A(n9626), .ZN(n9628) );
  INV_X1 U10953 ( .A(n9628), .ZN(n9629) );
  OAI222_X1 U10954 ( .A1(n9646), .A2(n9631), .B1(n9644), .B2(n9630), .C1(n9642), .C2(n9629), .ZN(n9702) );
  INV_X1 U10955 ( .A(n9702), .ZN(n9640) );
  XNOR2_X1 U10956 ( .A(n9633), .B(n9632), .ZN(n9703) );
  INV_X1 U10957 ( .A(n9634), .ZN(n9781) );
  AOI22_X1 U10958 ( .A1(n10632), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n10628), 
        .B2(n9635), .ZN(n9636) );
  OAI21_X1 U10959 ( .B1(n9781), .B2(n9637), .A(n9636), .ZN(n9638) );
  AOI21_X1 U10960 ( .B1(n9703), .B2(n9657), .A(n9638), .ZN(n9639) );
  OAI21_X1 U10961 ( .B1(n9640), .B2(n10632), .A(n9639), .ZN(P2_U3213) );
  AOI211_X1 U10962 ( .C1(n9654), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9649)
         );
  OAI22_X1 U10963 ( .A1(n9647), .A2(n9646), .B1(n9645), .B2(n9644), .ZN(n9648)
         );
  OR2_X1 U10964 ( .A1(n9649), .A2(n9648), .ZN(n9706) );
  AOI21_X1 U10965 ( .B1(n10628), .B2(n9650), .A(n9706), .ZN(n9660) );
  AOI22_X1 U10966 ( .A1(n9652), .A2(n9651), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10632), .ZN(n9659) );
  OAI21_X1 U10967 ( .B1(n9655), .B2(n9654), .A(n9653), .ZN(n9656) );
  INV_X1 U10968 ( .A(n9656), .ZN(n9707) );
  NAND2_X1 U10969 ( .A1(n9707), .A2(n9657), .ZN(n9658) );
  OAI211_X1 U10970 ( .C1(n9660), .C2(n10632), .A(n9659), .B(n9658), .ZN(
        P2_U3214) );
  NOR2_X1 U10971 ( .A1(n9743), .A2(n9747), .ZN(n9663) );
  AOI21_X1 U10972 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n9743), .A(n9663), .ZN(
        n9661) );
  OAI21_X1 U10973 ( .B1(n9662), .B2(n9715), .A(n9661), .ZN(P2_U3490) );
  AOI21_X1 U10974 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n9743), .A(n9663), .ZN(
        n9664) );
  OAI21_X1 U10975 ( .B1(n9665), .B2(n9715), .A(n9664), .ZN(P2_U3489) );
  NAND2_X1 U10976 ( .A1(n9666), .A2(n9744), .ZN(n9669) );
  INV_X1 U10977 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U10978 ( .A1(n9743), .A2(n9667), .ZN(n9668) );
  NAND2_X1 U10979 ( .A1(n9669), .A2(n9668), .ZN(n9673) );
  NAND2_X1 U10980 ( .A1(n9671), .A2(n9670), .ZN(n9672) );
  NAND2_X1 U10981 ( .A1(n9673), .A2(n9672), .ZN(P2_U3487) );
  INV_X1 U10982 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9675) );
  MUX2_X1 U10983 ( .A(n9675), .B(n9674), .S(n9744), .Z(n9676) );
  OAI21_X1 U10984 ( .B1(n9677), .B2(n9715), .A(n9676), .ZN(P2_U3486) );
  INV_X1 U10985 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9680) );
  AOI21_X1 U10986 ( .B1(n9711), .B2(n9679), .A(n9678), .ZN(n9754) );
  MUX2_X1 U10987 ( .A(n9680), .B(n9754), .S(n9744), .Z(n9681) );
  OAI21_X1 U10988 ( .B1(n9757), .B2(n9715), .A(n9681), .ZN(P2_U3485) );
  INV_X1 U10989 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9684) );
  AOI21_X1 U10990 ( .B1(n9711), .B2(n9683), .A(n9682), .ZN(n9758) );
  MUX2_X1 U10991 ( .A(n9684), .B(n9758), .S(n9744), .Z(n9685) );
  OAI21_X1 U10992 ( .B1(n9761), .B2(n9715), .A(n9685), .ZN(P2_U3484) );
  INV_X1 U10993 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9688) );
  AOI21_X1 U10994 ( .B1(n9687), .B2(n9711), .A(n9686), .ZN(n9762) );
  MUX2_X1 U10995 ( .A(n9688), .B(n9762), .S(n9744), .Z(n9689) );
  OAI21_X1 U10996 ( .B1(n9765), .B2(n9715), .A(n9689), .ZN(P2_U3483) );
  INV_X1 U10997 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9692) );
  AOI21_X1 U10998 ( .B1(n9711), .B2(n9691), .A(n9690), .ZN(n9766) );
  MUX2_X1 U10999 ( .A(n9692), .B(n9766), .S(n9744), .Z(n9693) );
  OAI21_X1 U11000 ( .B1(n9769), .B2(n9715), .A(n9693), .ZN(P2_U3482) );
  INV_X1 U11001 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9696) );
  AOI21_X1 U11002 ( .B1(n9711), .B2(n9695), .A(n9694), .ZN(n9770) );
  MUX2_X1 U11003 ( .A(n9696), .B(n9770), .S(n9744), .Z(n9697) );
  OAI21_X1 U11004 ( .B1(n9773), .B2(n9715), .A(n9697), .ZN(P2_U3481) );
  INV_X1 U11005 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9700) );
  AOI21_X1 U11006 ( .B1(n9699), .B2(n9711), .A(n9698), .ZN(n9774) );
  MUX2_X1 U11007 ( .A(n9700), .B(n9774), .S(n9744), .Z(n9701) );
  OAI21_X1 U11008 ( .B1(n9777), .B2(n9715), .A(n9701), .ZN(P2_U3480) );
  INV_X1 U11009 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9704) );
  AOI21_X1 U11010 ( .B1(n9711), .B2(n9703), .A(n9702), .ZN(n9778) );
  MUX2_X1 U11011 ( .A(n9704), .B(n9778), .S(n9744), .Z(n9705) );
  OAI21_X1 U11012 ( .B1(n9781), .B2(n9715), .A(n9705), .ZN(P2_U3479) );
  INV_X1 U11013 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9708) );
  AOI21_X1 U11014 ( .B1(n9707), .B2(n9711), .A(n9706), .ZN(n9782) );
  MUX2_X1 U11015 ( .A(n9708), .B(n9782), .S(n9744), .Z(n9709) );
  OAI21_X1 U11016 ( .B1(n9785), .B2(n9715), .A(n9709), .ZN(P2_U3478) );
  AOI21_X1 U11017 ( .B1(n9712), .B2(n9711), .A(n9710), .ZN(n9786) );
  MUX2_X1 U11018 ( .A(n9713), .B(n9786), .S(n9744), .Z(n9714) );
  OAI21_X1 U11019 ( .B1(n9790), .B2(n9715), .A(n9714), .ZN(P2_U3477) );
  OAI22_X1 U11020 ( .A1(n9719), .A2(n9718), .B1(n9717), .B2(n9716), .ZN(n9720)
         );
  OR2_X1 U11021 ( .A1(n9721), .A2(n9720), .ZN(n9791) );
  MUX2_X1 U11022 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9791), .S(n9744), .Z(
        P2_U3474) );
  NAND3_X1 U11023 ( .A1(n6863), .A2(n8281), .A3(n9722), .ZN(n9723) );
  NAND2_X1 U11024 ( .A1(n6889), .A2(n9723), .ZN(n9731) );
  NAND2_X1 U11025 ( .A1(n9725), .A2(n9724), .ZN(n9728) );
  NAND2_X1 U11026 ( .A1(n9726), .A2(n6257), .ZN(n9727) );
  NAND2_X1 U11027 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  AOI21_X1 U11028 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9736) );
  OR2_X1 U11029 ( .A1(n9732), .A2(n8281), .ZN(n9733) );
  NAND2_X1 U11030 ( .A1(n6885), .A2(n9733), .ZN(n10620) );
  NAND2_X1 U11031 ( .A1(n10620), .A2(n9734), .ZN(n9735) );
  NAND2_X1 U11032 ( .A1(n9736), .A2(n9735), .ZN(n10627) );
  INV_X1 U11033 ( .A(n10627), .ZN(n9742) );
  INV_X1 U11034 ( .A(n9737), .ZN(n9740) );
  AOI22_X1 U11035 ( .A1(n10620), .A2(n9740), .B1(n9739), .B2(n9738), .ZN(n9741) );
  NAND2_X1 U11036 ( .A1(n9742), .A2(n9741), .ZN(n10635) );
  MUX2_X1 U11037 ( .A(n10635), .B(P2_REG1_REG_2__SCAN_IN), .S(n9743), .Z(
        P2_U3461) );
  MUX2_X1 U11038 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9745), .S(n9744), .Z(
        P2_U3459) );
  INV_X1 U11039 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U11040 ( .A1(n9746), .A2(n6261), .ZN(n9748) );
  OR2_X1 U11041 ( .A1(n10652), .A2(n9747), .ZN(n9751) );
  OAI211_X1 U11042 ( .C1(n9749), .C2(n10649), .A(n9748), .B(n9751), .ZN(
        P2_U3458) );
  INV_X1 U11043 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U11044 ( .A1(n9750), .A2(n6261), .ZN(n9752) );
  OAI211_X1 U11045 ( .C1(n9753), .C2(n10649), .A(n9752), .B(n9751), .ZN(
        P2_U3457) );
  MUX2_X1 U11046 ( .A(n9755), .B(n9754), .S(n10649), .Z(n9756) );
  OAI21_X1 U11047 ( .B1(n9757), .B2(n9789), .A(n9756), .ZN(P2_U3453) );
  MUX2_X1 U11048 ( .A(n9759), .B(n9758), .S(n10649), .Z(n9760) );
  OAI21_X1 U11049 ( .B1(n9761), .B2(n9789), .A(n9760), .ZN(P2_U3452) );
  MUX2_X1 U11050 ( .A(n9763), .B(n9762), .S(n10649), .Z(n9764) );
  OAI21_X1 U11051 ( .B1(n9765), .B2(n9789), .A(n9764), .ZN(P2_U3451) );
  INV_X1 U11052 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9767) );
  MUX2_X1 U11053 ( .A(n9767), .B(n9766), .S(n10649), .Z(n9768) );
  OAI21_X1 U11054 ( .B1(n9769), .B2(n9789), .A(n9768), .ZN(P2_U3450) );
  MUX2_X1 U11055 ( .A(n9771), .B(n9770), .S(n10649), .Z(n9772) );
  OAI21_X1 U11056 ( .B1(n9773), .B2(n9789), .A(n9772), .ZN(P2_U3449) );
  MUX2_X1 U11057 ( .A(n9775), .B(n9774), .S(n10649), .Z(n9776) );
  OAI21_X1 U11058 ( .B1(n9777), .B2(n9789), .A(n9776), .ZN(P2_U3448) );
  INV_X1 U11059 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9779) );
  MUX2_X1 U11060 ( .A(n9779), .B(n9778), .S(n10649), .Z(n9780) );
  OAI21_X1 U11061 ( .B1(n9781), .B2(n9789), .A(n9780), .ZN(P2_U3447) );
  INV_X1 U11062 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9783) );
  MUX2_X1 U11063 ( .A(n9783), .B(n9782), .S(n10649), .Z(n9784) );
  OAI21_X1 U11064 ( .B1(n9785), .B2(n9789), .A(n9784), .ZN(P2_U3446) );
  INV_X1 U11065 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9787) );
  MUX2_X1 U11066 ( .A(n9787), .B(n9786), .S(n10649), .Z(n9788) );
  OAI21_X1 U11067 ( .B1(n9790), .B2(n9789), .A(n9788), .ZN(P2_U3444) );
  MUX2_X1 U11068 ( .A(n9791), .B(P2_REG0_REG_15__SCAN_IN), .S(n10652), .Z(
        P2_U3435) );
  INV_X1 U11069 ( .A(n10344), .ZN(n9797) );
  NOR4_X1 U11070 ( .A1(n9793), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9792), .ZN(n9794) );
  AOI21_X1 U11071 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9795), .A(n9794), .ZN(
        n9796) );
  OAI21_X1 U11072 ( .B1(n9797), .B2(n9801), .A(n9796), .ZN(P2_U3264) );
  OAI222_X1 U11073 ( .A1(P2_U3151), .A2(n9802), .B1(n9801), .B2(n9800), .C1(
        n9799), .C2(n9798), .ZN(P2_U3266) );
  MUX2_X1 U11074 ( .A(n9803), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U11075 ( .A(n9862), .ZN(n9806) );
  NOR3_X1 U11076 ( .A1(n9885), .A2(n9880), .A3(n9804), .ZN(n9805) );
  OAI21_X1 U11077 ( .B1(n9806), .B2(n9805), .A(n9922), .ZN(n9811) );
  NOR2_X1 U11078 ( .A1(n9827), .A2(n9887), .ZN(n9807) );
  AOI21_X1 U11079 ( .B1(n9939), .B2(n9865), .A(n9807), .ZN(n10136) );
  OAI22_X1 U11080 ( .A1(n10136), .A2(n10413), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9808), .ZN(n9809) );
  AOI21_X1 U11081 ( .B1(n10143), .B2(n9927), .A(n9809), .ZN(n9810) );
  OAI211_X1 U11082 ( .C1(n10311), .C2(n9931), .A(n9811), .B(n9810), .ZN(
        P1_U3216) );
  NAND2_X1 U11083 ( .A1(n9812), .A2(n9896), .ZN(n9895) );
  XOR2_X1 U11084 ( .A(n9814), .B(n4557), .Z(n9821) );
  INV_X1 U11085 ( .A(n10209), .ZN(n9818) );
  OAI22_X1 U11086 ( .A1(n9826), .A2(n9908), .B1(n9815), .B2(n9887), .ZN(n10201) );
  NAND2_X1 U11087 ( .A1(n10201), .A2(n9916), .ZN(n9816) );
  OAI211_X1 U11088 ( .C1(n10423), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9819)
         );
  AOI21_X1 U11089 ( .B1(n10208), .B2(n10421), .A(n9819), .ZN(n9820) );
  OAI21_X1 U11090 ( .B1(n9821), .B2(n10416), .A(n9820), .ZN(P1_U3219) );
  NAND2_X1 U11091 ( .A1(n9822), .A2(n9823), .ZN(n9824) );
  XOR2_X1 U11092 ( .A(n9825), .B(n9824), .Z(n9832) );
  INV_X1 U11093 ( .A(n10178), .ZN(n9829) );
  OAI22_X1 U11094 ( .A1(n9827), .A2(n9908), .B1(n9826), .B2(n9887), .ZN(n10171) );
  AOI22_X1 U11095 ( .A1(n10171), .A2(n9916), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9828) );
  OAI21_X1 U11096 ( .B1(n10423), .B2(n9829), .A(n9828), .ZN(n9830) );
  AOI21_X1 U11097 ( .B1(n10177), .B2(n10421), .A(n9830), .ZN(n9831) );
  OAI21_X1 U11098 ( .B1(n9832), .B2(n10416), .A(n9831), .ZN(P1_U3223) );
  AOI21_X1 U11099 ( .B1(n4566), .B2(n9833), .A(n9906), .ZN(n9840) );
  OAI22_X1 U11100 ( .A1(n9835), .A2(n9908), .B1(n9834), .B2(n9887), .ZN(n10104) );
  OAI22_X1 U11101 ( .A1(n10109), .A2(n10423), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9836), .ZN(n9838) );
  NOR2_X1 U11102 ( .A1(n10304), .A2(n9931), .ZN(n9837) );
  AOI211_X1 U11103 ( .C1(n9916), .C2(n10104), .A(n9838), .B(n9837), .ZN(n9839)
         );
  OAI21_X1 U11104 ( .B1(n9840), .B2(n10416), .A(n9839), .ZN(P1_U3225) );
  XOR2_X1 U11105 ( .A(n9841), .B(n9842), .Z(n9850) );
  INV_X1 U11106 ( .A(n9843), .ZN(n9846) );
  AOI22_X1 U11107 ( .A1(n9916), .A2(n9844), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9845) );
  OAI21_X1 U11108 ( .B1(n10423), .B2(n9846), .A(n9845), .ZN(n9847) );
  AOI21_X1 U11109 ( .B1(n9848), .B2(n10421), .A(n9847), .ZN(n9849) );
  OAI21_X1 U11110 ( .B1(n9850), .B2(n10416), .A(n9849), .ZN(P1_U3226) );
  XOR2_X1 U11111 ( .A(n9851), .B(n9852), .Z(n9859) );
  AOI21_X1 U11112 ( .B1(n9916), .B2(n9854), .A(n9853), .ZN(n9855) );
  OAI21_X1 U11113 ( .B1(n10423), .B2(n9856), .A(n9855), .ZN(n9857) );
  AOI21_X1 U11114 ( .B1(n10275), .B2(n10421), .A(n9857), .ZN(n9858) );
  OAI21_X1 U11115 ( .B1(n9859), .B2(n10416), .A(n9858), .ZN(P1_U3228) );
  AND3_X1 U11116 ( .A1(n9862), .A2(n9861), .A3(n9860), .ZN(n9863) );
  OAI21_X1 U11117 ( .B1(n9864), .B2(n9863), .A(n9922), .ZN(n9869) );
  NOR2_X1 U11118 ( .A1(n10423), .A2(n10125), .ZN(n9867) );
  AOI22_X1 U11119 ( .A1(n9938), .A2(n9865), .B1(n9940), .B2(n9910), .ZN(n10121) );
  NOR2_X1 U11120 ( .A1(n10121), .A2(n10413), .ZN(n9866) );
  AOI211_X1 U11121 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n9867), 
        .B(n9866), .ZN(n9868) );
  OAI211_X1 U11122 ( .C1(n4881), .C2(n9931), .A(n9869), .B(n9868), .ZN(
        P1_U3229) );
  XNOR2_X1 U11123 ( .A(n9872), .B(n9871), .ZN(n9873) );
  XNOR2_X1 U11124 ( .A(n9870), .B(n9873), .ZN(n9879) );
  OR2_X1 U11125 ( .A1(n9888), .A2(n9908), .ZN(n9875) );
  NAND2_X1 U11126 ( .A1(n6059), .A2(n9910), .ZN(n9874) );
  NAND2_X1 U11127 ( .A1(n9875), .A2(n9874), .ZN(n10186) );
  AOI22_X1 U11128 ( .A1(n10186), .A2(n9916), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9876) );
  OAI21_X1 U11129 ( .B1(n10423), .B2(n10191), .A(n9876), .ZN(n9877) );
  AOI21_X1 U11130 ( .B1(n10197), .B2(n10421), .A(n9877), .ZN(n9878) );
  OAI21_X1 U11131 ( .B1(n9879), .B2(n10416), .A(n9878), .ZN(P1_U3233) );
  INV_X1 U11132 ( .A(n9880), .ZN(n9884) );
  OR2_X1 U11133 ( .A1(n9881), .A2(n9880), .ZN(n9882) );
  AOI22_X1 U11134 ( .A1(n9885), .A2(n9884), .B1(n9883), .B2(n9882), .ZN(n9894)
         );
  OR2_X1 U11135 ( .A1(n9886), .A2(n9908), .ZN(n9890) );
  OR2_X1 U11136 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  NAND2_X1 U11137 ( .A1(n9890), .A2(n9889), .ZN(n10151) );
  AOI22_X1 U11138 ( .A1(n10151), .A2(n9916), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9891) );
  OAI21_X1 U11139 ( .B1(n10423), .B2(n10160), .A(n9891), .ZN(n9892) );
  AOI21_X1 U11140 ( .B1(n10159), .B2(n10421), .A(n9892), .ZN(n9893) );
  OAI21_X1 U11141 ( .B1(n9894), .B2(n10416), .A(n9893), .ZN(P1_U3235) );
  OAI21_X1 U11142 ( .B1(n9896), .B2(n9812), .A(n9895), .ZN(n9897) );
  NAND2_X1 U11143 ( .A1(n9897), .A2(n9922), .ZN(n9903) );
  OAI22_X1 U11144 ( .A1(n10413), .A2(n9899), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9898), .ZN(n9900) );
  AOI21_X1 U11145 ( .B1(n9901), .B2(n9927), .A(n9900), .ZN(n9902) );
  OAI211_X1 U11146 ( .C1(n10330), .C2(n9931), .A(n9903), .B(n9902), .ZN(
        P1_U3238) );
  OAI21_X1 U11147 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  NAND3_X1 U11148 ( .A1(n5064), .A2(n9922), .A3(n9907), .ZN(n9918) );
  OR2_X1 U11149 ( .A1(n9909), .A2(n9908), .ZN(n9912) );
  NAND2_X1 U11150 ( .A1(n9938), .A2(n9910), .ZN(n9911) );
  NAND2_X1 U11151 ( .A1(n9912), .A2(n9911), .ZN(n10089) );
  INV_X1 U11152 ( .A(n10096), .ZN(n9914) );
  OAI22_X1 U11153 ( .A1(n9914), .A2(n10423), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9913), .ZN(n9915) );
  AOI21_X1 U11154 ( .B1(n10089), .B2(n9916), .A(n9915), .ZN(n9917) );
  OAI211_X1 U11155 ( .C1(n10300), .C2(n9931), .A(n9918), .B(n9917), .ZN(
        P1_U3240) );
  OAI21_X1 U11156 ( .B1(n9921), .B2(n9919), .A(n9920), .ZN(n9923) );
  NAND2_X1 U11157 ( .A1(n9923), .A2(n9922), .ZN(n9930) );
  OAI22_X1 U11158 ( .A1(n10413), .A2(n9925), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9924), .ZN(n9926) );
  AOI21_X1 U11159 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9929) );
  OAI211_X1 U11160 ( .C1(n6032), .C2(n9931), .A(n9930), .B(n9929), .ZN(
        P1_U3241) );
  MUX2_X1 U11161 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9932), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U11162 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9933), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U11163 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9934), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U11164 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9935), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11165 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9936), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11166 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9937), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U11167 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9938), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11168 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9939), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U11169 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9940), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U11170 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9941), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11171 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n5021), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11172 ( .A(n9943), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9942), .Z(
        P1_U3574) );
  MUX2_X1 U11173 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n6059), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11174 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9944), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11175 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9945), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11176 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9946), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U11177 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9947), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U11178 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9948), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11179 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9949), .S(P1_U3973), .Z(
        P1_U3567) );
  INV_X1 U11180 ( .A(n9950), .ZN(n9951) );
  MUX2_X1 U11181 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9951), .S(P1_U3973), .Z(
        P1_U3566) );
  INV_X1 U11182 ( .A(n9952), .ZN(n9953) );
  MUX2_X1 U11183 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9953), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11184 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9954), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11185 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9955), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U11186 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9956), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U11187 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9957), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11188 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9958), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U11189 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9959), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U11190 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9960), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U11191 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9961), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11192 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9962), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U11193 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9963), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U11194 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9964), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U11195 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10351) );
  OAI22_X1 U11196 ( .A1(n9966), .A2(n10351), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9965), .ZN(n9967) );
  AOI21_X1 U11197 ( .B1(n9968), .B2(n10022), .A(n9967), .ZN(n9979) );
  MUX2_X1 U11198 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10524), .S(n9969), .Z(n9971) );
  NAND2_X1 U11199 ( .A1(n9971), .A2(n9970), .ZN(n9972) );
  NAND3_X1 U11200 ( .A1(n10033), .A2(n9973), .A3(n9972), .ZN(n9978) );
  OAI211_X1 U11201 ( .C1(n9976), .C2(n9975), .A(n10025), .B(n9974), .ZN(n9977)
         );
  NAND3_X1 U11202 ( .A1(n9979), .A2(n9978), .A3(n9977), .ZN(P1_U3244) );
  AOI22_X1 U11203 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n10021), 
        .B2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9989) );
  XOR2_X1 U11204 ( .A(n9981), .B(n9980), .Z(n9982) );
  AOI22_X1 U11205 ( .A1(n9983), .A2(n10022), .B1(n10033), .B2(n9982), .ZN(
        n9988) );
  OAI211_X1 U11206 ( .C1(n9986), .C2(n9985), .A(n10025), .B(n9984), .ZN(n9987)
         );
  NAND4_X1 U11207 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(
        P1_U3245) );
  NOR2_X1 U11208 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7423), .ZN(n9992) );
  NOR2_X1 U11209 ( .A1(n10007), .A2(n9996), .ZN(n9991) );
  AOI211_X1 U11210 ( .C1(n10021), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9992), .B(
        n9991), .ZN(n10004) );
  OAI211_X1 U11211 ( .C1(n9995), .C2(n9994), .A(n10025), .B(n9993), .ZN(n10003) );
  MUX2_X1 U11212 ( .A(n6670), .B(P1_REG1_REG_3__SCAN_IN), .S(n9996), .Z(n10001) );
  INV_X1 U11213 ( .A(n9997), .ZN(n10000) );
  INV_X1 U11214 ( .A(n9998), .ZN(n9999) );
  OAI211_X1 U11215 ( .C1(n10001), .C2(n10000), .A(n10033), .B(n9999), .ZN(
        n10002) );
  NAND3_X1 U11216 ( .A1(n10004), .A2(n10003), .A3(n10002), .ZN(P1_U3246) );
  INV_X1 U11217 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U11218 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10005), .ZN(n10009) );
  NOR2_X1 U11219 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  AOI211_X1 U11220 ( .C1(n10021), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10009), .B(
        n10008), .ZN(n10020) );
  OAI211_X1 U11221 ( .C1(n10012), .C2(n10011), .A(n10025), .B(n10010), .ZN(
        n10019) );
  INV_X1 U11222 ( .A(n10035), .ZN(n10017) );
  NAND3_X1 U11223 ( .A1(n10015), .A2(n10014), .A3(n10013), .ZN(n10016) );
  NAND3_X1 U11224 ( .A1(n10033), .A2(n10017), .A3(n10016), .ZN(n10018) );
  NAND3_X1 U11225 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(P1_U3248) );
  AND2_X1 U11226 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10410) );
  AOI21_X1 U11227 ( .B1(n10021), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10410), .ZN(
        n10039) );
  NAND2_X1 U11228 ( .A1(n10022), .A2(n10028), .ZN(n10038) );
  INV_X1 U11229 ( .A(n10023), .ZN(n10024) );
  OAI211_X1 U11230 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10037) );
  MUX2_X1 U11231 ( .A(n6676), .B(P1_REG1_REG_6__SCAN_IN), .S(n10028), .Z(
        n10031) );
  INV_X1 U11232 ( .A(n10029), .ZN(n10030) );
  NAND2_X1 U11233 ( .A1(n10031), .A2(n10030), .ZN(n10034) );
  OAI211_X1 U11234 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10036) );
  NAND4_X1 U11235 ( .A1(n10039), .A2(n10038), .A3(n10037), .A4(n10036), .ZN(
        P1_U3249) );
  INV_X1 U11236 ( .A(n10040), .ZN(n10041) );
  NAND2_X1 U11237 ( .A1(n10218), .A2(n10450), .ZN(n10046) );
  AOI21_X1 U11238 ( .B1(n10215), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10044), 
        .ZN(n10045) );
  OAI211_X1 U11239 ( .C1(n4741), .C2(n10456), .A(n10046), .B(n10045), .ZN(
        P1_U3264) );
  NAND2_X1 U11240 ( .A1(n10047), .A2(n10458), .ZN(n10055) );
  INV_X1 U11241 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10048) );
  OAI22_X1 U11242 ( .A1(n10049), .A2(n10190), .B1(n10048), .B2(n8066), .ZN(
        n10052) );
  NOR2_X1 U11243 ( .A1(n10050), .A2(n10194), .ZN(n10051) );
  AOI211_X1 U11244 ( .C1(n10441), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10054) );
  OAI211_X1 U11245 ( .C1(n10056), .C2(n10215), .A(n10055), .B(n10054), .ZN(
        P1_U3356) );
  INV_X1 U11246 ( .A(n10057), .ZN(n10066) );
  NAND2_X1 U11247 ( .A1(n10058), .A2(n10458), .ZN(n10065) );
  AOI22_X1 U11248 ( .A1(n10059), .A2(n10452), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10462), .ZN(n10060) );
  OAI21_X1 U11249 ( .B1(n10061), .B2(n10456), .A(n10060), .ZN(n10062) );
  AOI21_X1 U11250 ( .B1(n10063), .B2(n10450), .A(n10062), .ZN(n10064) );
  OAI211_X1 U11251 ( .C1(n10066), .C2(n10215), .A(n10065), .B(n10064), .ZN(
        P1_U3265) );
  OAI21_X1 U11252 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n10070) );
  NAND2_X1 U11253 ( .A1(n10070), .A2(n10427), .ZN(n10073) );
  INV_X1 U11254 ( .A(n10071), .ZN(n10072) );
  NAND2_X1 U11255 ( .A1(n10073), .A2(n10072), .ZN(n10221) );
  INV_X1 U11256 ( .A(n10221), .ZN(n10086) );
  OAI21_X1 U11257 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n10223) );
  NAND2_X1 U11258 ( .A1(n10223), .A2(n10458), .ZN(n10085) );
  INV_X1 U11259 ( .A(n10077), .ZN(n10078) );
  AOI211_X1 U11260 ( .C1(n10080), .C2(n10079), .A(n10502), .B(n10078), .ZN(
        n10222) );
  AOI22_X1 U11261 ( .A1(n10081), .A2(n10452), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10462), .ZN(n10082) );
  OAI21_X1 U11262 ( .B1(n10296), .B2(n10456), .A(n10082), .ZN(n10083) );
  AOI21_X1 U11263 ( .B1(n10222), .B2(n10450), .A(n10083), .ZN(n10084) );
  OAI211_X1 U11264 ( .C1(n10215), .C2(n10086), .A(n10085), .B(n10084), .ZN(
        P1_U3266) );
  XNOR2_X1 U11265 ( .A(n10088), .B(n10087), .ZN(n10091) );
  INV_X1 U11266 ( .A(n10089), .ZN(n10090) );
  OAI21_X1 U11267 ( .B1(n10091), .B2(n10203), .A(n10090), .ZN(n10226) );
  INV_X1 U11268 ( .A(n10226), .ZN(n10101) );
  XNOR2_X1 U11269 ( .A(n10093), .B(n10092), .ZN(n10228) );
  NAND2_X1 U11270 ( .A1(n10228), .A2(n10458), .ZN(n10100) );
  AOI211_X1 U11271 ( .C1(n10095), .C2(n10110), .A(n10502), .B(n10094), .ZN(
        n10227) );
  AOI22_X1 U11272 ( .A1(n10096), .A2(n10452), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10462), .ZN(n10097) );
  OAI21_X1 U11273 ( .B1(n10300), .B2(n10456), .A(n10097), .ZN(n10098) );
  AOI21_X1 U11274 ( .B1(n10227), .B2(n10450), .A(n10098), .ZN(n10099) );
  OAI211_X1 U11275 ( .C1(n10215), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        P1_U3267) );
  NAND2_X1 U11276 ( .A1(n10119), .A2(n10102), .ZN(n10103) );
  XNOR2_X1 U11277 ( .A(n10103), .B(n10106), .ZN(n10105) );
  AOI21_X1 U11278 ( .B1(n10105), .B2(n10427), .A(n10104), .ZN(n10232) );
  XNOR2_X1 U11279 ( .A(n10107), .B(n10106), .ZN(n10234) );
  NAND2_X1 U11280 ( .A1(n10234), .A2(n10458), .ZN(n10115) );
  INV_X1 U11281 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10108) );
  OAI22_X1 U11282 ( .A1(n10109), .A2(n10190), .B1(n10108), .B2(n8066), .ZN(
        n10112) );
  OAI211_X1 U11283 ( .C1(n10304), .C2(n4599), .A(n10435), .B(n10110), .ZN(
        n10231) );
  NOR2_X1 U11284 ( .A1(n10231), .A2(n10194), .ZN(n10111) );
  AOI211_X1 U11285 ( .C1(n10441), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10114) );
  OAI211_X1 U11286 ( .C1(n10215), .C2(n10232), .A(n10115), .B(n10114), .ZN(
        P1_U3268) );
  NAND2_X1 U11287 ( .A1(n10132), .A2(n10116), .ZN(n10118) );
  NAND2_X1 U11288 ( .A1(n10118), .A2(n10117), .ZN(n10120) );
  NAND3_X1 U11289 ( .A1(n10120), .A2(n10427), .A3(n10119), .ZN(n10122) );
  NAND2_X1 U11290 ( .A1(n10122), .A2(n10121), .ZN(n10237) );
  INV_X1 U11291 ( .A(n10237), .ZN(n10131) );
  XNOR2_X1 U11292 ( .A(n10123), .B(n4796), .ZN(n10239) );
  NAND2_X1 U11293 ( .A1(n10239), .A2(n10458), .ZN(n10130) );
  AOI211_X1 U11294 ( .C1(n10124), .C2(n10140), .A(n10502), .B(n4599), .ZN(
        n10238) );
  INV_X1 U11295 ( .A(n10125), .ZN(n10126) );
  AOI22_X1 U11296 ( .A1(n10126), .A2(n10452), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10462), .ZN(n10127) );
  OAI21_X1 U11297 ( .B1(n4881), .B2(n10456), .A(n10127), .ZN(n10128) );
  AOI21_X1 U11298 ( .B1(n10238), .B2(n10450), .A(n10128), .ZN(n10129) );
  OAI211_X1 U11299 ( .C1(n10215), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        P1_U3269) );
  OAI21_X1 U11300 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10135) );
  NAND2_X1 U11301 ( .A1(n10135), .A2(n10427), .ZN(n10137) );
  NAND2_X1 U11302 ( .A1(n10137), .A2(n10136), .ZN(n10242) );
  INV_X1 U11303 ( .A(n10242), .ZN(n10148) );
  XNOR2_X1 U11304 ( .A(n10139), .B(n10138), .ZN(n10244) );
  NAND2_X1 U11305 ( .A1(n10244), .A2(n10458), .ZN(n10147) );
  INV_X1 U11306 ( .A(n10140), .ZN(n10141) );
  AOI211_X1 U11307 ( .C1(n10142), .C2(n10157), .A(n10502), .B(n10141), .ZN(
        n10243) );
  AOI22_X1 U11308 ( .A1(n10143), .A2(n10452), .B1(n10215), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n10144) );
  OAI21_X1 U11309 ( .B1(n10311), .B2(n10456), .A(n10144), .ZN(n10145) );
  AOI21_X1 U11310 ( .B1(n10243), .B2(n10450), .A(n10145), .ZN(n10146) );
  OAI211_X1 U11311 ( .C1(n10215), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        P1_U3270) );
  XNOR2_X1 U11312 ( .A(n10149), .B(n10154), .ZN(n10150) );
  NAND2_X1 U11313 ( .A1(n10150), .A2(n10427), .ZN(n10153) );
  INV_X1 U11314 ( .A(n10151), .ZN(n10152) );
  NAND2_X1 U11315 ( .A1(n10153), .A2(n10152), .ZN(n10247) );
  INV_X1 U11316 ( .A(n10247), .ZN(n10166) );
  XNOR2_X1 U11317 ( .A(n10155), .B(n10154), .ZN(n10249) );
  NAND2_X1 U11318 ( .A1(n10249), .A2(n10458), .ZN(n10165) );
  INV_X1 U11319 ( .A(n10157), .ZN(n10158) );
  AOI211_X1 U11320 ( .C1(n10159), .C2(n10176), .A(n10502), .B(n10158), .ZN(
        n10248) );
  INV_X1 U11321 ( .A(n10160), .ZN(n10161) );
  AOI22_X1 U11322 ( .A1(n10161), .A2(n10452), .B1(n10215), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n10162) );
  OAI21_X1 U11323 ( .B1(n6206), .B2(n10456), .A(n10162), .ZN(n10163) );
  AOI21_X1 U11324 ( .B1(n10248), .B2(n10450), .A(n10163), .ZN(n10164) );
  OAI211_X1 U11325 ( .C1(n10215), .C2(n10166), .A(n10165), .B(n10164), .ZN(
        P1_U3271) );
  NAND2_X1 U11326 ( .A1(n10167), .A2(n10174), .ZN(n10168) );
  NAND2_X1 U11327 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  NAND2_X1 U11328 ( .A1(n10170), .A2(n10427), .ZN(n10173) );
  INV_X1 U11329 ( .A(n10171), .ZN(n10172) );
  NAND2_X1 U11330 ( .A1(n10173), .A2(n10172), .ZN(n10252) );
  INV_X1 U11331 ( .A(n10252), .ZN(n10183) );
  XNOR2_X1 U11332 ( .A(n10175), .B(n10174), .ZN(n10254) );
  NAND2_X1 U11333 ( .A1(n10254), .A2(n10458), .ZN(n10182) );
  AOI211_X1 U11334 ( .C1(n10177), .C2(n10193), .A(n10502), .B(n10156), .ZN(
        n10253) );
  AOI22_X1 U11335 ( .A1(n10462), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10178), 
        .B2(n10452), .ZN(n10179) );
  OAI21_X1 U11336 ( .B1(n10318), .B2(n10456), .A(n10179), .ZN(n10180) );
  AOI21_X1 U11337 ( .B1(n10253), .B2(n10450), .A(n10180), .ZN(n10181) );
  OAI211_X1 U11338 ( .C1(n10215), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        P1_U3272) );
  INV_X1 U11339 ( .A(n10189), .ZN(n10184) );
  XNOR2_X1 U11340 ( .A(n10185), .B(n10184), .ZN(n10187) );
  AOI21_X1 U11341 ( .B1(n10187), .B2(n10427), .A(n10186), .ZN(n10258) );
  XOR2_X1 U11342 ( .A(n10189), .B(n10188), .Z(n10260) );
  NAND2_X1 U11343 ( .A1(n10260), .A2(n10458), .ZN(n10199) );
  INV_X1 U11344 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10192) );
  OAI22_X1 U11345 ( .A1(n8066), .A2(n10192), .B1(n10191), .B2(n10190), .ZN(
        n10196) );
  OAI211_X1 U11346 ( .C1(n10322), .C2(n4598), .A(n10435), .B(n10193), .ZN(
        n10257) );
  NOR2_X1 U11347 ( .A1(n10257), .A2(n10194), .ZN(n10195) );
  AOI211_X1 U11348 ( .C1(n10441), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10198) );
  OAI211_X1 U11349 ( .C1(n10215), .C2(n10258), .A(n10199), .B(n10198), .ZN(
        P1_U3273) );
  XNOR2_X1 U11350 ( .A(n10200), .B(n10205), .ZN(n10204) );
  INV_X1 U11351 ( .A(n10201), .ZN(n10202) );
  OAI21_X1 U11352 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(n10263) );
  INV_X1 U11353 ( .A(n10263), .ZN(n10214) );
  XNOR2_X1 U11354 ( .A(n10206), .B(n10205), .ZN(n10265) );
  NAND2_X1 U11355 ( .A1(n10265), .A2(n10458), .ZN(n10213) );
  AOI211_X1 U11356 ( .C1(n10208), .C2(n10207), .A(n10502), .B(n4598), .ZN(
        n10264) );
  AOI22_X1 U11357 ( .A1(n10215), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10209), 
        .B2(n10452), .ZN(n10210) );
  OAI21_X1 U11358 ( .B1(n4884), .B2(n10456), .A(n10210), .ZN(n10211) );
  AOI21_X1 U11359 ( .B1(n10264), .B2(n10450), .A(n10211), .ZN(n10212) );
  OAI211_X1 U11360 ( .C1(n10215), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        P1_U3274) );
  INV_X1 U11361 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10219) );
  INV_X1 U11362 ( .A(n10216), .ZN(n10217) );
  NOR2_X1 U11363 ( .A1(n10218), .A2(n10217), .ZN(n10290) );
  MUX2_X1 U11364 ( .A(n10219), .B(n10290), .S(n10537), .Z(n10220) );
  OAI21_X1 U11365 ( .B1(n4741), .B2(n10273), .A(n10220), .ZN(P1_U3552) );
  OAI21_X1 U11366 ( .B1(n10296), .B2(n10273), .A(n10225), .ZN(P1_U3549) );
  INV_X1 U11367 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10229) );
  AOI211_X1 U11368 ( .C1(n10228), .C2(n10520), .A(n10227), .B(n10226), .ZN(
        n10297) );
  MUX2_X1 U11369 ( .A(n10229), .B(n10297), .S(n10537), .Z(n10230) );
  OAI21_X1 U11370 ( .B1(n10300), .B2(n10273), .A(n10230), .ZN(P1_U3548) );
  INV_X1 U11371 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U11372 ( .A1(n10232), .A2(n10231), .ZN(n10233) );
  AOI21_X1 U11373 ( .B1(n10234), .B2(n10520), .A(n10233), .ZN(n10301) );
  MUX2_X1 U11374 ( .A(n10235), .B(n10301), .S(n10537), .Z(n10236) );
  OAI21_X1 U11375 ( .B1(n10304), .B2(n10273), .A(n10236), .ZN(P1_U3547) );
  AOI211_X1 U11376 ( .C1(n10239), .C2(n10520), .A(n10238), .B(n10237), .ZN(
        n10305) );
  MUX2_X1 U11377 ( .A(n10240), .B(n10305), .S(n10537), .Z(n10241) );
  OAI21_X1 U11378 ( .B1(n4881), .B2(n10273), .A(n10241), .ZN(P1_U3546) );
  AOI211_X1 U11379 ( .C1(n10244), .C2(n10520), .A(n10243), .B(n10242), .ZN(
        n10308) );
  MUX2_X1 U11380 ( .A(n10245), .B(n10308), .S(n10537), .Z(n10246) );
  OAI21_X1 U11381 ( .B1(n10311), .B2(n10273), .A(n10246), .ZN(P1_U3545) );
  AOI211_X1 U11382 ( .C1(n10249), .C2(n10520), .A(n10248), .B(n10247), .ZN(
        n10312) );
  MUX2_X1 U11383 ( .A(n10250), .B(n10312), .S(n10537), .Z(n10251) );
  OAI21_X1 U11384 ( .B1(n6206), .B2(n10273), .A(n10251), .ZN(P1_U3544) );
  INV_X1 U11385 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10255) );
  AOI211_X1 U11386 ( .C1(n10254), .C2(n10520), .A(n10253), .B(n10252), .ZN(
        n10315) );
  MUX2_X1 U11387 ( .A(n10255), .B(n10315), .S(n10537), .Z(n10256) );
  OAI21_X1 U11388 ( .B1(n10318), .B2(n10273), .A(n10256), .ZN(P1_U3543) );
  INV_X1 U11389 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U11390 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  AOI21_X1 U11391 ( .B1(n10260), .B2(n10520), .A(n10259), .ZN(n10319) );
  MUX2_X1 U11392 ( .A(n10261), .B(n10319), .S(n10537), .Z(n10262) );
  OAI21_X1 U11393 ( .B1(n10322), .B2(n10273), .A(n10262), .ZN(P1_U3542) );
  AOI211_X1 U11394 ( .C1(n10265), .C2(n10520), .A(n10264), .B(n10263), .ZN(
        n10323) );
  MUX2_X1 U11395 ( .A(n10266), .B(n10323), .S(n10537), .Z(n10267) );
  OAI21_X1 U11396 ( .B1(n4884), .B2(n10273), .A(n10267), .ZN(P1_U3541) );
  AOI211_X1 U11397 ( .C1(n10270), .C2(n10520), .A(n10269), .B(n10268), .ZN(
        n10326) );
  MUX2_X1 U11398 ( .A(n10271), .B(n10326), .S(n10537), .Z(n10272) );
  OAI21_X1 U11399 ( .B1(n10330), .B2(n10273), .A(n10272), .ZN(P1_U3540) );
  AOI21_X1 U11400 ( .B1(n10282), .B2(n10275), .A(n10274), .ZN(n10276) );
  OAI211_X1 U11401 ( .C1(n10278), .C2(n10284), .A(n10277), .B(n10276), .ZN(
        n10331) );
  MUX2_X1 U11402 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10331), .S(n10537), .Z(
        P1_U3539) );
  AOI211_X1 U11403 ( .C1(n10282), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        n10283) );
  OAI21_X1 U11404 ( .B1(n10285), .B2(n10284), .A(n10283), .ZN(n10332) );
  MUX2_X1 U11405 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10332), .S(n10537), .Z(
        P1_U3537) );
  MUX2_X1 U11406 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10286), .S(n10537), .Z(
        P1_U3522) );
  OAI21_X1 U11407 ( .B1(n10289), .B2(n10329), .A(n10288), .ZN(P1_U3521) );
  INV_X1 U11408 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10291) );
  MUX2_X1 U11409 ( .A(n10291), .B(n10290), .S(n10523), .Z(n10292) );
  OAI21_X1 U11410 ( .B1(n4741), .B2(n10329), .A(n10292), .ZN(P1_U3520) );
  INV_X1 U11411 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10294) );
  OAI21_X1 U11412 ( .B1(n10296), .B2(n10329), .A(n10295), .ZN(P1_U3517) );
  MUX2_X1 U11413 ( .A(n10298), .B(n10297), .S(n10523), .Z(n10299) );
  OAI21_X1 U11414 ( .B1(n10300), .B2(n10329), .A(n10299), .ZN(P1_U3516) );
  MUX2_X1 U11415 ( .A(n10302), .B(n10301), .S(n10523), .Z(n10303) );
  OAI21_X1 U11416 ( .B1(n10304), .B2(n10329), .A(n10303), .ZN(P1_U3515) );
  INV_X1 U11417 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10306) );
  MUX2_X1 U11418 ( .A(n10306), .B(n10305), .S(n10523), .Z(n10307) );
  OAI21_X1 U11419 ( .B1(n4881), .B2(n10329), .A(n10307), .ZN(P1_U3514) );
  INV_X1 U11420 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U11421 ( .A(n10309), .B(n10308), .S(n10523), .Z(n10310) );
  OAI21_X1 U11422 ( .B1(n10311), .B2(n10329), .A(n10310), .ZN(P1_U3513) );
  INV_X1 U11423 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10313) );
  MUX2_X1 U11424 ( .A(n10313), .B(n10312), .S(n10523), .Z(n10314) );
  OAI21_X1 U11425 ( .B1(n6206), .B2(n10329), .A(n10314), .ZN(P1_U3512) );
  INV_X1 U11426 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10316) );
  MUX2_X1 U11427 ( .A(n10316), .B(n10315), .S(n10523), .Z(n10317) );
  OAI21_X1 U11428 ( .B1(n10318), .B2(n10329), .A(n10317), .ZN(P1_U3511) );
  MUX2_X1 U11429 ( .A(n10320), .B(n10319), .S(n10523), .Z(n10321) );
  OAI21_X1 U11430 ( .B1(n10322), .B2(n10329), .A(n10321), .ZN(P1_U3510) );
  INV_X1 U11431 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10324) );
  MUX2_X1 U11432 ( .A(n10324), .B(n10323), .S(n10523), .Z(n10325) );
  OAI21_X1 U11433 ( .B1(n4884), .B2(n10329), .A(n10325), .ZN(P1_U3509) );
  INV_X1 U11434 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10327) );
  MUX2_X1 U11435 ( .A(n10327), .B(n10326), .S(n10523), .Z(n10328) );
  OAI21_X1 U11436 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(P1_U3507) );
  MUX2_X1 U11437 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10331), .S(n10523), .Z(
        P1_U3504) );
  MUX2_X1 U11438 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10332), .S(n10523), .Z(
        P1_U3498) );
  MUX2_X1 U11439 ( .A(P1_D_REG_1__SCAN_IN), .B(n10335), .S(n10469), .Z(
        P1_U3440) );
  MUX2_X1 U11440 ( .A(P1_D_REG_0__SCAN_IN), .B(n10336), .S(n10469), .Z(
        P1_U3439) );
  INV_X1 U11441 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10337) );
  NAND3_X1 U11442 ( .A1(n10337), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10340) );
  OAI22_X1 U11443 ( .A1(n10341), .A2(n10340), .B1(n10339), .B2(n10338), .ZN(
        n10342) );
  AOI21_X1 U11444 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10345) );
  INV_X1 U11445 ( .A(n10345), .ZN(P1_U3324) );
  NOR2_X1 U11446 ( .A1(n10346), .A2(n10347), .ZN(n10407) );
  NOR2_X1 U11447 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10403) );
  NOR2_X1 U11448 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10399) );
  INV_X1 U11449 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10395) );
  INV_X1 U11450 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11451 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n10389) );
  NOR2_X1 U11452 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10385) );
  NOR2_X1 U11453 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10378) );
  NOR2_X1 U11454 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10374) );
  NOR2_X1 U11455 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10371) );
  NOR2_X1 U11456 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10369) );
  NOR2_X1 U11457 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10366) );
  NOR2_X1 U11458 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10364) );
  NOR2_X1 U11459 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10360) );
  NAND2_X1 U11460 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10356) );
  INV_X1 U11461 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U11462 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10349), .B2(n10348), .ZN(n10689) );
  NAND2_X1 U11463 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10354) );
  AOI21_X1 U11464 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10653) );
  NAND2_X1 U11465 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10350) );
  NOR2_X1 U11466 ( .A1(n10351), .A2(n10350), .ZN(n10654) );
  NOR2_X1 U11467 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10654), .ZN(n10352) );
  NOR2_X1 U11468 ( .A1(n10653), .A2(n10352), .ZN(n10687) );
  XOR2_X1 U11469 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10686) );
  NAND2_X1 U11470 ( .A1(n10687), .A2(n10686), .ZN(n10353) );
  NAND2_X1 U11471 ( .A1(n10354), .A2(n10353), .ZN(n10688) );
  NAND2_X1 U11472 ( .A1(n10689), .A2(n10688), .ZN(n10355) );
  NAND2_X1 U11473 ( .A1(n10356), .A2(n10355), .ZN(n10691) );
  INV_X1 U11474 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U11475 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n10358), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n10357), .ZN(n10690) );
  NOR2_X1 U11476 ( .A1(n10691), .A2(n10690), .ZN(n10359) );
  NOR2_X1 U11477 ( .A1(n10360), .A2(n10359), .ZN(n10679) );
  INV_X1 U11478 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U11479 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10362), .B1(
        P2_ADDR_REG_5__SCAN_IN), .B2(n10361), .ZN(n10678) );
  NOR2_X1 U11480 ( .A1(n10679), .A2(n10678), .ZN(n10363) );
  NOR2_X1 U11481 ( .A1(n10364), .A2(n10363), .ZN(n10677) );
  XNOR2_X1 U11482 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10676) );
  NOR2_X1 U11483 ( .A1(n10677), .A2(n10676), .ZN(n10365) );
  NOR2_X1 U11484 ( .A1(n10366), .A2(n10365), .ZN(n10683) );
  INV_X1 U11485 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U11486 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10367), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n10596), .ZN(n10682) );
  NOR2_X1 U11487 ( .A1(n10683), .A2(n10682), .ZN(n10368) );
  NOR2_X1 U11488 ( .A1(n10369), .A2(n10368), .ZN(n10685) );
  XNOR2_X1 U11489 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10684) );
  NOR2_X1 U11490 ( .A1(n10685), .A2(n10684), .ZN(n10370) );
  NOR2_X1 U11491 ( .A1(n10371), .A2(n10370), .ZN(n10681) );
  AOI22_X1 U11492 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6713), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10372), .ZN(n10680) );
  NOR2_X1 U11493 ( .A1(n10681), .A2(n10680), .ZN(n10373) );
  NOR2_X1 U11494 ( .A1(n10374), .A2(n10373), .ZN(n10675) );
  INV_X1 U11495 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U11496 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10376), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10375), .ZN(n10674) );
  NOR2_X1 U11497 ( .A1(n10675), .A2(n10674), .ZN(n10377) );
  NOR2_X1 U11498 ( .A1(n10378), .A2(n10377), .ZN(n10673) );
  AOI22_X1 U11499 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n10380), .B1(
        P2_ADDR_REG_11__SCAN_IN), .B2(n10381), .ZN(n10672) );
  NOR2_X1 U11500 ( .A1(n10673), .A2(n10672), .ZN(n10379) );
  AOI21_X1 U11501 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(n10671) );
  INV_X1 U11502 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U11503 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10383), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10382), .ZN(n10670) );
  NOR2_X1 U11504 ( .A1(n10671), .A2(n10670), .ZN(n10384) );
  NOR2_X1 U11505 ( .A1(n10385), .A2(n10384), .ZN(n10669) );
  INV_X1 U11506 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U11507 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n10387), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(n10386), .ZN(n10668) );
  NOR2_X1 U11508 ( .A1(n10669), .A2(n10668), .ZN(n10388) );
  NOR2_X1 U11509 ( .A1(n10389), .A2(n10388), .ZN(n10667) );
  AOI22_X1 U11510 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n10391), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(n10392), .ZN(n10666) );
  NOR2_X1 U11511 ( .A1(n10667), .A2(n10666), .ZN(n10390) );
  AOI21_X1 U11512 ( .B1(n10392), .B2(n10391), .A(n10390), .ZN(n10665) );
  AOI22_X1 U11513 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n10394), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n10395), .ZN(n10664) );
  NOR2_X1 U11514 ( .A1(n10665), .A2(n10664), .ZN(n10393) );
  AOI21_X1 U11515 ( .B1(n10395), .B2(n10394), .A(n10393), .ZN(n10663) );
  INV_X1 U11516 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U11517 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10397), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10396), .ZN(n10662) );
  NOR2_X1 U11518 ( .A1(n10663), .A2(n10662), .ZN(n10398) );
  NOR2_X1 U11519 ( .A1(n10399), .A2(n10398), .ZN(n10661) );
  INV_X1 U11520 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U11521 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10401), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10400), .ZN(n10660) );
  NOR2_X1 U11522 ( .A1(n10661), .A2(n10660), .ZN(n10402) );
  NOR2_X1 U11523 ( .A1(n10403), .A2(n10402), .ZN(n10658) );
  NOR2_X1 U11524 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10658), .ZN(n10405) );
  NAND2_X1 U11525 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10658), .ZN(n10657) );
  OAI21_X1 U11526 ( .B1(n10405), .B2(n10404), .A(n10657), .ZN(n10406) );
  XOR2_X1 U11527 ( .A(n10407), .B(n10406), .Z(ADD_1068_U4) );
  INV_X1 U11528 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U11529 ( .A1(n10652), .A2(n10409), .B1(n10408), .B2(n10649), .ZN(
        P2_U3429) );
  XNOR2_X1 U11530 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U11531 ( .A(n10410), .ZN(n10411) );
  OAI21_X1 U11532 ( .B1(n10413), .B2(n10412), .A(n10411), .ZN(n10420) );
  NAND2_X1 U11533 ( .A1(n10415), .A2(n10414), .ZN(n10417) );
  AOI21_X1 U11534 ( .B1(n10418), .B2(n10417), .A(n10416), .ZN(n10419) );
  AOI211_X1 U11535 ( .C1(n10449), .C2(n10421), .A(n10420), .B(n10419), .ZN(
        n10422) );
  OAI21_X1 U11536 ( .B1(n10424), .B2(n10423), .A(n10422), .ZN(P1_U3239) );
  XNOR2_X1 U11537 ( .A(n10425), .B(n10430), .ZN(n10428) );
  AOI21_X1 U11538 ( .B1(n10428), .B2(n10427), .A(n10426), .ZN(n10516) );
  AOI222_X1 U11539 ( .A1(n10432), .A2(n10441), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n10215), .C1(n10429), .C2(n10452), .ZN(n10439) );
  XNOR2_X1 U11540 ( .A(n10431), .B(n10430), .ZN(n10521) );
  INV_X1 U11541 ( .A(n10432), .ZN(n10518) );
  INV_X1 U11542 ( .A(n10433), .ZN(n10436) );
  OAI211_X1 U11543 ( .C1(n10518), .C2(n10436), .A(n4900), .B(n10435), .ZN(
        n10515) );
  INV_X1 U11544 ( .A(n10515), .ZN(n10437) );
  AOI22_X1 U11545 ( .A1(n10521), .A2(n10458), .B1(n10450), .B2(n10437), .ZN(
        n10438) );
  OAI211_X1 U11546 ( .C1(n10462), .C2(n10516), .A(n10439), .B(n10438), .ZN(
        P1_U3280) );
  AOI222_X1 U11547 ( .A1(n10442), .A2(n10441), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n10215), .C1(n10452), .C2(n10440), .ZN(n10447) );
  AOI22_X1 U11548 ( .A1(n10445), .A2(n10444), .B1(n10450), .B2(n10443), .ZN(
        n10446) );
  OAI211_X1 U11549 ( .C1(n10462), .C2(n10448), .A(n10447), .B(n10446), .ZN(
        P1_U3286) );
  NAND2_X1 U11550 ( .A1(n10451), .A2(n10450), .ZN(n10455) );
  AOI22_X1 U11551 ( .A1(n10462), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10453), 
        .B2(n10452), .ZN(n10454) );
  OAI211_X1 U11552 ( .C1(n4892), .C2(n10456), .A(n10455), .B(n10454), .ZN(
        n10457) );
  AOI21_X1 U11553 ( .B1(n10459), .B2(n10458), .A(n10457), .ZN(n10460) );
  OAI21_X1 U11554 ( .B1(n10462), .B2(n10461), .A(n10460), .ZN(P1_U3287) );
  AND2_X1 U11555 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10470), .ZN(P1_U3294) );
  AND2_X1 U11556 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10470), .ZN(P1_U3295) );
  AND2_X1 U11557 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10470), .ZN(P1_U3296) );
  AND2_X1 U11558 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10470), .ZN(P1_U3297) );
  AND2_X1 U11559 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10470), .ZN(P1_U3298) );
  NOR2_X1 U11560 ( .A1(n10469), .A2(n10463), .ZN(P1_U3299) );
  AND2_X1 U11561 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10470), .ZN(P1_U3300) );
  NOR2_X1 U11562 ( .A1(n10469), .A2(n10464), .ZN(P1_U3301) );
  AND2_X1 U11563 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10470), .ZN(P1_U3302) );
  AND2_X1 U11564 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10470), .ZN(P1_U3303) );
  AND2_X1 U11565 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10470), .ZN(P1_U3304) );
  NOR2_X1 U11566 ( .A1(n10469), .A2(n10465), .ZN(P1_U3305) );
  AND2_X1 U11567 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10470), .ZN(P1_U3306) );
  AND2_X1 U11568 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10470), .ZN(P1_U3307) );
  AND2_X1 U11569 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10470), .ZN(P1_U3308) );
  AND2_X1 U11570 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10470), .ZN(P1_U3309) );
  AND2_X1 U11571 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10470), .ZN(P1_U3310) );
  NOR2_X1 U11572 ( .A1(n10469), .A2(n10466), .ZN(P1_U3311) );
  NOR2_X1 U11573 ( .A1(n10469), .A2(n10467), .ZN(P1_U3312) );
  NOR2_X1 U11574 ( .A1(n10469), .A2(n10468), .ZN(P1_U3313) );
  AND2_X1 U11575 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10470), .ZN(P1_U3314) );
  AND2_X1 U11576 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10470), .ZN(P1_U3315) );
  AND2_X1 U11577 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10470), .ZN(P1_U3316) );
  AND2_X1 U11578 ( .A1(n10470), .A2(P1_D_REG_8__SCAN_IN), .ZN(P1_U3317) );
  AND2_X1 U11579 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10470), .ZN(P1_U3318) );
  AND2_X1 U11580 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10470), .ZN(P1_U3319) );
  AND2_X1 U11581 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10470), .ZN(P1_U3320) );
  AND2_X1 U11582 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10470), .ZN(P1_U3321) );
  AND2_X1 U11583 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10470), .ZN(P1_U3322) );
  AND2_X1 U11584 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10470), .ZN(P1_U3323) );
  OAI21_X1 U11585 ( .B1(n6205), .B2(n10517), .A(n10471), .ZN(n10472) );
  AOI21_X1 U11586 ( .B1(n10473), .B2(n10481), .A(n10472), .ZN(n10475) );
  AND2_X1 U11587 ( .A1(n10475), .A2(n10474), .ZN(n10525) );
  INV_X1 U11588 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U11589 ( .A1(n10523), .A2(n10525), .B1(n10476), .B2(n6596), .ZN(
        P1_U3456) );
  INV_X1 U11590 ( .A(n10477), .ZN(n10479) );
  OAI21_X1 U11591 ( .B1(n10479), .B2(n10517), .A(n10478), .ZN(n10480) );
  AOI21_X1 U11592 ( .B1(n10482), .B2(n10481), .A(n10480), .ZN(n10483) );
  INV_X1 U11593 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U11594 ( .A1(n10523), .A2(n10526), .B1(n10485), .B2(n6596), .ZN(
        P1_U3477) );
  INV_X1 U11595 ( .A(n10486), .ZN(n10489) );
  OAI211_X1 U11596 ( .C1(n10489), .C2(n10517), .A(n10488), .B(n10487), .ZN(
        n10490) );
  AOI21_X1 U11597 ( .B1(n10520), .B2(n10491), .A(n10490), .ZN(n10528) );
  INV_X1 U11598 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U11599 ( .A1(n10523), .A2(n10528), .B1(n10492), .B2(n6596), .ZN(
        P1_U3480) );
  OAI21_X1 U11600 ( .B1(n10494), .B2(n10517), .A(n10493), .ZN(n10495) );
  AOI211_X1 U11601 ( .C1(n10497), .C2(n10520), .A(n10496), .B(n10495), .ZN(
        n10529) );
  INV_X1 U11602 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U11603 ( .A1(n10523), .A2(n10529), .B1(n10498), .B2(n6596), .ZN(
        P1_U3483) );
  NOR2_X1 U11604 ( .A1(n10500), .A2(n10499), .ZN(n10505) );
  OAI22_X1 U11605 ( .A1(n10503), .A2(n10502), .B1(n10501), .B2(n10517), .ZN(
        n10504) );
  NOR3_X1 U11606 ( .A1(n10506), .A2(n10505), .A3(n10504), .ZN(n10531) );
  INV_X1 U11607 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U11608 ( .A1(n10523), .A2(n10531), .B1(n10507), .B2(n6596), .ZN(
        P1_U3486) );
  INV_X1 U11609 ( .A(n10508), .ZN(n10513) );
  OAI211_X1 U11610 ( .C1(n10511), .C2(n10517), .A(n10510), .B(n10509), .ZN(
        n10512) );
  AOI21_X1 U11611 ( .B1(n10513), .B2(n10520), .A(n10512), .ZN(n10533) );
  INV_X1 U11612 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U11613 ( .A1(n10523), .A2(n10533), .B1(n10514), .B2(n6596), .ZN(
        P1_U3489) );
  OAI211_X1 U11614 ( .C1(n10518), .C2(n10517), .A(n10516), .B(n10515), .ZN(
        n10519) );
  AOI21_X1 U11615 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(n10536) );
  INV_X1 U11616 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U11617 ( .A1(n10523), .A2(n10536), .B1(n10522), .B2(n6596), .ZN(
        P1_U3492) );
  AOI22_X1 U11618 ( .A1(n10537), .A2(n10525), .B1(n10524), .B2(n10534), .ZN(
        P1_U3523) );
  AOI22_X1 U11619 ( .A1(n10537), .A2(n10526), .B1(n6680), .B2(n10534), .ZN(
        P1_U3530) );
  AOI22_X1 U11620 ( .A1(n10537), .A2(n10528), .B1(n10527), .B2(n10534), .ZN(
        P1_U3531) );
  AOI22_X1 U11621 ( .A1(n10537), .A2(n10529), .B1(n6724), .B2(n10534), .ZN(
        P1_U3532) );
  AOI22_X1 U11622 ( .A1(n10537), .A2(n10531), .B1(n10530), .B2(n10534), .ZN(
        P1_U3533) );
  AOI22_X1 U11623 ( .A1(n10537), .A2(n10533), .B1(n10532), .B2(n10534), .ZN(
        P1_U3534) );
  AOI22_X1 U11624 ( .A1(n10537), .A2(n10536), .B1(n10535), .B2(n10534), .ZN(
        P1_U3535) );
  INV_X1 U11625 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10655) );
  INV_X1 U11626 ( .A(n10538), .ZN(n10539) );
  AOI21_X1 U11627 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(n10547) );
  AOI211_X1 U11628 ( .C1(n10544), .C2(n10543), .A(n10542), .B(n10561), .ZN(
        n10545) );
  AOI21_X1 U11629 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_U3151), .A(n10545), 
        .ZN(n10546) );
  OAI21_X1 U11630 ( .B1(n10547), .B2(n10615), .A(n10546), .ZN(n10548) );
  AOI21_X1 U11631 ( .B1(n10549), .B2(n10586), .A(n10548), .ZN(n10556) );
  INV_X1 U11632 ( .A(n10550), .ZN(n10551) );
  AOI21_X1 U11633 ( .B1(n10553), .B2(n10552), .A(n10551), .ZN(n10554) );
  OR2_X1 U11634 ( .A1(n10606), .A2(n10554), .ZN(n10555) );
  OAI211_X1 U11635 ( .C1(n10655), .C2(n10597), .A(n10556), .B(n10555), .ZN(
        P2_U3183) );
  INV_X1 U11636 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10568) );
  OAI21_X1 U11637 ( .B1(n10559), .B2(n10558), .A(n10557), .ZN(n10565) );
  AOI211_X1 U11638 ( .C1(n10563), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        n10564) );
  AOI21_X1 U11639 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(n10567) );
  OAI21_X1 U11640 ( .B1(n10597), .B2(n10568), .A(n10567), .ZN(n10569) );
  AOI21_X1 U11641 ( .B1(n10570), .B2(n10586), .A(n10569), .ZN(n10577) );
  INV_X1 U11642 ( .A(n10606), .ZN(n10575) );
  OAI21_X1 U11643 ( .B1(n10573), .B2(n10572), .A(n10571), .ZN(n10574) );
  NAND2_X1 U11644 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  OAI211_X1 U11645 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7106), .A(n10577), .B(
        n10576), .ZN(P2_U3184) );
  AOI21_X1 U11646 ( .B1(n7534), .B2(n10579), .A(n10578), .ZN(n10588) );
  AOI21_X1 U11647 ( .B1(n7535), .B2(n10581), .A(n10580), .ZN(n10582) );
  NOR2_X1 U11648 ( .A1(n10582), .A2(n10615), .ZN(n10583) );
  AOI211_X1 U11649 ( .C1(n10586), .C2(n10585), .A(n10584), .B(n10583), .ZN(
        n10587) );
  OAI21_X1 U11650 ( .B1(n10588), .B2(n10606), .A(n10587), .ZN(n10589) );
  INV_X1 U11651 ( .A(n10589), .ZN(n10595) );
  OAI21_X1 U11652 ( .B1(n10592), .B2(n10591), .A(n10590), .ZN(n10593) );
  NAND2_X1 U11653 ( .A1(n10612), .A2(n10593), .ZN(n10594) );
  OAI211_X1 U11654 ( .C1(n10597), .C2(n10596), .A(n10595), .B(n10594), .ZN(
        P2_U3189) );
  OAI22_X1 U11655 ( .A1(n10598), .A2(n9410), .B1(n10597), .B2(n10387), .ZN(
        n10599) );
  INV_X1 U11656 ( .A(n10599), .ZN(n10619) );
  AOI21_X1 U11657 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(n10616) );
  AOI21_X1 U11658 ( .B1(n10605), .B2(n10604), .A(n10603), .ZN(n10607) );
  OR2_X1 U11659 ( .A1(n10607), .A2(n10606), .ZN(n10614) );
  OAI21_X1 U11660 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(n10611) );
  NAND2_X1 U11661 ( .A1(n10612), .A2(n10611), .ZN(n10613) );
  OAI211_X1 U11662 ( .C1(n10616), .C2(n10615), .A(n10614), .B(n10613), .ZN(
        n10617) );
  INV_X1 U11663 ( .A(n10617), .ZN(n10618) );
  OAI211_X1 U11664 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5469), .A(n10619), .B(
        n10618), .ZN(P2_U3195) );
  INV_X1 U11665 ( .A(n10620), .ZN(n10625) );
  INV_X1 U11666 ( .A(n10621), .ZN(n10624) );
  OAI22_X1 U11667 ( .A1(n10625), .A2(n10624), .B1(n10623), .B2(n10622), .ZN(
        n10626) );
  AOI211_X1 U11668 ( .C1(n10628), .C2(P2_REG3_REG_2__SCAN_IN), .A(n10627), .B(
        n10626), .ZN(n10630) );
  AOI22_X1 U11669 ( .A1(n10632), .A2(n10631), .B1(n10630), .B2(n10629), .ZN(
        P2_U3231) );
  INV_X1 U11670 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U11671 ( .A1(n10652), .A2(n10634), .B1(n10633), .B2(n10649), .ZN(
        P2_U3393) );
  OAI22_X1 U11672 ( .A1(n10649), .A2(P2_REG0_REG_2__SCAN_IN), .B1(n10635), 
        .B2(n10652), .ZN(n10636) );
  INV_X1 U11673 ( .A(n10636), .ZN(P2_U3396) );
  INV_X1 U11674 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U11675 ( .A1(n10652), .A2(n10638), .B1(n10637), .B2(n10649), .ZN(
        P2_U3399) );
  AOI22_X1 U11676 ( .A1(n10652), .A2(n10640), .B1(n10639), .B2(n10649), .ZN(
        P2_U3402) );
  INV_X1 U11677 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U11678 ( .A1(n10652), .A2(n10642), .B1(n10641), .B2(n10649), .ZN(
        P2_U3405) );
  INV_X1 U11679 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U11680 ( .A1(n10652), .A2(n10644), .B1(n10643), .B2(n10649), .ZN(
        P2_U3408) );
  INV_X1 U11681 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U11682 ( .A1(n10652), .A2(n10646), .B1(n10645), .B2(n10649), .ZN(
        P2_U3414) );
  INV_X1 U11683 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U11684 ( .A1(n10652), .A2(n10648), .B1(n10647), .B2(n10649), .ZN(
        P2_U3423) );
  INV_X1 U11685 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U11686 ( .A1(n10652), .A2(n10651), .B1(n10650), .B2(n10649), .ZN(
        P2_U3426) );
  NOR2_X1 U11687 ( .A1(n10654), .A2(n10653), .ZN(n10656) );
  XNOR2_X1 U11688 ( .A(n10656), .B(n10655), .ZN(ADD_1068_U5) );
  XOR2_X1 U11689 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11690 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10658), .A(n10657), 
        .ZN(n10659) );
  XNOR2_X1 U11691 ( .A(n10659), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  XNOR2_X1 U11692 ( .A(n10661), .B(n10660), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11693 ( .A(n10663), .B(n10662), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11694 ( .A(n10665), .B(n10664), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11695 ( .A(n10667), .B(n10666), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11696 ( .A(n10669), .B(n10668), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11697 ( .A(n10671), .B(n10670), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11698 ( .A(n10673), .B(n10672), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11699 ( .A(n10675), .B(n10674), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11700 ( .A(n10677), .B(n10676), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11701 ( .A(n10679), .B(n10678), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11702 ( .A(n10681), .B(n10680), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11703 ( .A(n10683), .B(n10682), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11704 ( .A(n10685), .B(n10684), .ZN(ADD_1068_U48) );
  XOR2_X1 U11705 ( .A(n10687), .B(n10686), .Z(ADD_1068_U54) );
  XOR2_X1 U11706 ( .A(n10689), .B(n10688), .Z(ADD_1068_U53) );
  XNOR2_X1 U11707 ( .A(n10691), .B(n10690), .ZN(ADD_1068_U52) );
  OAI21_X1 U6339 ( .B1(n4693), .B2(n9833), .A(n4688), .ZN(n9906) );
  AOI21_X1 U5044 ( .B1(n9880), .B2(n4690), .A(n4689), .ZN(n4688) );
  INV_X1 U5056 ( .A(n5891), .ZN(n7427) );
  NAND2_X1 U5078 ( .A1(n5219), .A2(n5218), .ZN(n5566) );
  XNOR2_X1 U5236 ( .A(n9520), .B(n9523), .ZN(n9535) );
  CLKBUF_X1 U5996 ( .A(n6277), .Z(n8822) );
  CLKBUF_X1 U6340 ( .A(n6267), .Z(n4526) );
endmodule

