

module b20_C_SARLock_k_64_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173;

  INV_X4 U4801 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  CLKBUF_X2 U4802 ( .A(n6305), .Z(n4295) );
  CLKBUF_X3 U4803 ( .A(n6310), .Z(n4294) );
  CLKBUF_X1 U4804 ( .A(n5658), .Z(n5682) );
  INV_X1 U4805 ( .A(n5625), .ZN(n5614) );
  INV_X1 U4806 ( .A(n5625), .ZN(n5609) );
  INV_X1 U4807 ( .A(n7121), .ZN(n5500) );
  AND2_X1 U4808 ( .A1(n4845), .A2(n5568), .ZN(n4644) );
  INV_X2 U4809 ( .A(n5605), .ZN(n5834) );
  INV_X1 U4810 ( .A(n6842), .ZN(n5949) );
  BUF_X1 U4811 ( .A(n5272), .Z(n7124) );
  INV_X1 U4812 ( .A(n8256), .ZN(n8264) );
  NAND2_X1 U4813 ( .A1(n4907), .A2(n4906), .ZN(n5134) );
  NAND2_X2 U4814 ( .A1(n7731), .A2(n6364), .ZN(n6416) );
  XNOR2_X1 U4815 ( .A(n4900), .B(SI_5_), .ZN(n5074) );
  XNOR2_X1 U4816 ( .A(n5298), .B(n5470), .ZN(n8609) );
  XNOR2_X1 U4817 ( .A(n5585), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6364) );
  AND3_X2 U4819 ( .A1(n4645), .A2(n4490), .A3(n4644), .ZN(n5954) );
  NAND2_X2 U4820 ( .A1(n8339), .A2(n5513), .ZN(n6377) );
  NOR2_X1 U4821 ( .A1(n7977), .A2(n7978), .ZN(n7982) );
  XNOR2_X2 U4822 ( .A(n9094), .B(n9090), .ZN(n9231) );
  NAND2_X2 U4823 ( .A1(n4614), .A2(n4615), .ZN(n8654) );
  XNOR2_X2 U4824 ( .A(n5087), .B(n5086), .ZN(n6391) );
  NAND2_X1 U4825 ( .A1(n4447), .A2(n4896), .ZN(n5087) );
  OAI211_X2 U4826 ( .C1(n6416), .C2(n6457), .A(n5674), .B(n5673), .ZN(n7336)
         );
  AOI22_X1 U4827 ( .A1(n6084), .A2(n6310), .B1(n6311), .B2(n6085), .ZN(n6090)
         );
  INV_X1 U4828 ( .A(n6078), .ZN(n6310) );
  NAND4_X4 U4829 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n5481)
         );
  CLKBUF_X1 U4830 ( .A(n6364), .Z(n4296) );
  NAND2_X2 U4831 ( .A1(n5831), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5832) );
  AND2_X1 U4832 ( .A1(n4430), .A2(n4428), .ZN(n8339) );
  NAND2_X1 U4833 ( .A1(n6022), .A2(n6021), .ZN(n9471) );
  AND3_X1 U4834 ( .A1(n4673), .A2(n4321), .A3(n4672), .ZN(n7108) );
  NAND2_X2 U4835 ( .A1(n8104), .A2(n8107), .ZN(n6777) );
  NAND4_X1 U4836 ( .A1(n5059), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n8475)
         );
  INV_X1 U4837 ( .A(n6298), .ZN(n6308) );
  INV_X1 U4838 ( .A(n6084), .ZN(n5992) );
  OR2_X1 U4839 ( .A1(n5272), .A2(n6554), .ZN(n5013) );
  BUF_X1 U4840 ( .A(n5039), .Z(n5211) );
  NAND2_X2 U4841 ( .A1(n5007), .A2(n5006), .ZN(n7121) );
  CLKBUF_X2 U4842 ( .A(n5034), .Z(n5506) );
  INV_X2 U4843 ( .A(n8609), .ZN(n8622) );
  XNOR2_X1 U4844 ( .A(n4519), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8610) );
  INV_X4 U4845 ( .A(n6388), .ZN(n6389) );
  AOI21_X1 U4846 ( .B1(n4560), .B2(n4756), .A(n4559), .ZN(n8317) );
  AOI21_X1 U4847 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8053) );
  NAND2_X1 U4848 ( .A1(n4765), .A2(n4763), .ZN(n9241) );
  OAI21_X1 U4849 ( .B1(n7982), .B2(n4476), .A(n7987), .ZN(n8042) );
  XNOR2_X1 U4850 ( .A(n9386), .B(n9392), .ZN(n9738) );
  NAND2_X1 U4851 ( .A1(n4781), .A2(n4779), .ZN(n8926) );
  AND2_X1 U4852 ( .A1(n4616), .A2(n4320), .ZN(n8663) );
  OR2_X1 U4853 ( .A1(n9382), .A2(n9383), .ZN(n9385) );
  OR2_X2 U4854 ( .A1(n6264), .A2(n9113), .ZN(n9116) );
  NAND2_X1 U4855 ( .A1(n4842), .A2(n4841), .ZN(n4840) );
  AOI21_X1 U4856 ( .B1(n4397), .B2(n4473), .A(n7948), .ZN(n7960) );
  OR2_X1 U4857 ( .A1(n8768), .A2(n4448), .ZN(n4450) );
  OAI21_X2 U4858 ( .B1(n7341), .B2(n5176), .A(n5175), .ZN(n7368) );
  OAI21_X1 U4859 ( .B1(n7050), .B2(n5709), .A(n8006), .ZN(n7358) );
  OR2_X1 U4860 ( .A1(n9784), .A2(n9274), .ZN(n6010) );
  AND2_X1 U4861 ( .A1(n7217), .A2(n7863), .ZN(n7219) );
  NAND2_X1 U4862 ( .A1(n4830), .A2(n4829), .ZN(n7217) );
  NOR2_X1 U4863 ( .A1(n6846), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U4864 ( .A1(n5204), .A2(n4928), .ZN(n4746) );
  INV_X2 U4865 ( .A(n8767), .ZN(n8780) );
  NAND2_X2 U4866 ( .A1(n6957), .A2(n9978), .ZN(n9984) );
  OAI211_X1 U4867 ( .C1(n5506), .C2(n6585), .A(n5077), .B(n5076), .ZN(n10081)
         );
  AND3_X1 U4868 ( .A1(n5095), .A2(n5094), .A3(n5093), .ZN(n10076) );
  NAND4_X2 U4869 ( .A1(n5070), .A2(n5069), .A3(n5068), .A4(n5067), .ZN(n8474)
         );
  NAND4_X1 U4870 ( .A1(n5044), .A2(n5043), .A3(n5042), .A4(n5041), .ZN(n8476)
         );
  NAND4_X1 U4871 ( .A1(n4861), .A2(n5029), .A3(n5028), .A4(n5027), .ZN(n6783)
         );
  AND3_X1 U4872 ( .A1(n5052), .A2(n5051), .A3(n5050), .ZN(n6916) );
  NAND3_X1 U4873 ( .A1(n4445), .A2(n4899), .A3(n4444), .ZN(n5075) );
  INV_X2 U4874 ( .A(n8103), .ZN(n8252) );
  AOI21_X1 U4875 ( .B1(n4303), .B2(n4728), .A(n4341), .ZN(n4723) );
  INV_X2 U4876 ( .A(n5703), .ZN(n6345) );
  INV_X2 U4877 ( .A(n5038), .ZN(n7119) );
  NAND2_X1 U4878 ( .A1(n9330), .A2(n7837), .ZN(n9983) );
  NAND2_X1 U4879 ( .A1(n6416), .A2(n6389), .ZN(n5703) );
  MUX2_X1 U4880 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9801), .S(n6416), .Z(n7024) );
  AND2_X1 U4881 ( .A1(n5965), .A2(n5964), .ZN(n5967) );
  XNOR2_X1 U4882 ( .A(n5473), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6643) );
  AND2_X1 U4883 ( .A1(n5957), .A2(n4315), .ZN(n5964) );
  NAND2_X1 U4884 ( .A1(n5594), .A2(n5593), .ZN(n7731) );
  AND2_X2 U4885 ( .A1(n5578), .A2(n5579), .ZN(n5645) );
  NAND2_X1 U4886 ( .A1(n8897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5002) );
  INV_X1 U4887 ( .A(n8342), .ZN(n5006) );
  INV_X2 U4888 ( .A(n8610), .ZN(n8318) );
  XNOR2_X1 U4889 ( .A(n5005), .B(n5004), .ZN(n8342) );
  XNOR2_X1 U4890 ( .A(n5575), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U4891 ( .A1(n5818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U4892 ( .A(n4894), .B(SI_3_), .ZN(n5062) );
  OR2_X1 U4893 ( .A1(n5000), .A2(n5147), .ZN(n4976) );
  NAND2_X1 U4894 ( .A1(n4648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U4895 ( .A1(n5529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4519) );
  OAI21_X1 U4896 ( .B1(n6357), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4888), .ZN(
        n4889) );
  AND2_X2 U4897 ( .A1(n4812), .A2(n4814), .ZN(n4975) );
  INV_X1 U4898 ( .A(n5163), .ZN(n4814) );
  NAND2_X1 U4899 ( .A1(n4704), .A2(n4317), .ZN(n6579) );
  AND2_X1 U4900 ( .A1(n4862), .A2(n4846), .ZN(n4845) );
  AND2_X1 U4901 ( .A1(n4313), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U4902 ( .A1(n4496), .A2(n4879), .ZN(n4501) );
  NAND2_X1 U4903 ( .A1(n4881), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4502) );
  AND2_X1 U4904 ( .A1(n5595), .A2(n5596), .ZN(n5652) );
  AND3_X1 U4905 ( .A1(n9020), .A2(n9019), .A3(n5474), .ZN(n4970) );
  AND4_X1 U4906 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5630), .ZN(n5567)
         );
  NAND2_X1 U4907 ( .A1(n4498), .A2(n4497), .ZN(n4496) );
  AND2_X1 U4908 ( .A1(n4961), .A2(n4966), .ZN(n4697) );
  INV_X1 U4909 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5829) );
  INV_X1 U4910 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5816) );
  NOR2_X1 U4911 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4962) );
  NOR2_X1 U4912 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5563) );
  NOR2_X1 U4913 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4963) );
  NOR2_X1 U4914 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4964) );
  NOR2_X1 U4915 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5562) );
  NOR2_X1 U4916 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5561) );
  NOR2_X1 U4917 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5564) );
  NOR2_X1 U4918 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5281) );
  INV_X1 U4919 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5474) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5595) );
  INV_X1 U4921 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5596) );
  INV_X4 U4922 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4923 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4879) );
  INV_X1 U4924 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4498) );
  NAND4_X2 U4925 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n6084)
         );
  NAND2_X2 U4926 ( .A1(n5008), .A2(n5006), .ZN(n5039) );
  AOI21_X2 U4927 ( .B1(n9195), .B2(n6191), .A(n4877), .ZN(n6198) );
  INV_X2 U4928 ( .A(n6035), .ZN(n9330) );
  AOI211_X2 U4929 ( .C1(n9766), .C2(n9260), .A(n9100), .B(n9099), .ZN(n9101)
         );
  AOI21_X2 U4930 ( .B1(n4587), .B2(n4589), .A(n4343), .ZN(n6909) );
  NAND2_X1 U4931 ( .A1(n5007), .A2(n8342), .ZN(n5038) );
  OAI222_X1 U4932 ( .A1(n5007), .A2(P2_U3151), .B1(n8907), .B2(n8906), .C1(
        n8905), .C2(n8904), .ZN(P2_U3265) );
  NAND2_X1 U4933 ( .A1(n5025), .A2(n6648), .ZN(n8104) );
  NAND2_X1 U4934 ( .A1(n6073), .A2(n7985), .ZN(n6075) );
  AND2_X1 U4935 ( .A1(n5571), .A2(n5572), .ZN(n4860) );
  INV_X1 U4936 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5572) );
  AOI21_X1 U4937 ( .B1(n4742), .B2(n4741), .A(n4740), .ZN(n4739) );
  NAND2_X1 U4938 ( .A1(n4458), .A2(n4457), .ZN(n5314) );
  AOI21_X1 U4939 ( .B1(n4460), .B2(n4462), .A(SI_20_), .ZN(n4457) );
  NAND2_X1 U4940 ( .A1(n5265), .A2(n4460), .ZN(n4458) );
  OAI21_X1 U4941 ( .B1(n5265), .B2(n4462), .A(n4460), .ZN(n5313) );
  INV_X1 U4942 ( .A(n5128), .ZN(n4904) );
  INV_X1 U4943 ( .A(n8465), .ZN(n7694) );
  NAND2_X1 U4944 ( .A1(n5495), .A2(n5494), .ZN(n8310) );
  OR2_X1 U4945 ( .A1(n8636), .A2(n8643), .ZN(n5494) );
  OR2_X1 U4946 ( .A1(n5277), .A2(n8391), .ZN(n4869) );
  NOR2_X1 U4947 ( .A1(n4354), .A2(n4780), .ZN(n4779) );
  INV_X1 U4948 ( .A(n8928), .ZN(n4780) );
  NAND2_X1 U4949 ( .A1(n4410), .A2(n4409), .ZN(n4408) );
  NAND2_X1 U4950 ( .A1(n4545), .A2(n8236), .ZN(n4544) );
  OR2_X1 U4951 ( .A1(n9736), .A2(n6030), .ZN(n7952) );
  AND2_X1 U4952 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  AOI21_X1 U4953 ( .B1(n4658), .B2(n4660), .A(n4657), .ZN(n4656) );
  INV_X1 U4954 ( .A(n4661), .ZN(n4658) );
  INV_X1 U4955 ( .A(n4660), .ZN(n4659) );
  AND2_X1 U4956 ( .A1(n8312), .A2(n8270), .ZN(n4750) );
  NAND2_X1 U4957 ( .A1(n6698), .A2(n6580), .ZN(n6581) );
  NAND2_X1 U4958 ( .A1(n4567), .A2(n4566), .ZN(n6796) );
  AOI21_X1 U4959 ( .B1(n4568), .B2(n4570), .A(n4319), .ZN(n4566) );
  NAND2_X1 U4960 ( .A1(n4700), .A2(n8538), .ZN(n4699) );
  OR2_X1 U4961 ( .A1(n4718), .A2(n4720), .ZN(n4715) );
  NAND2_X1 U4962 ( .A1(n4718), .A2(n4382), .ZN(n4716) );
  NAND2_X1 U4963 ( .A1(n8879), .A2(n8740), .ZN(n4603) );
  OR2_X1 U4964 ( .A1(n8873), .A2(n8730), .ZN(n8219) );
  OR2_X1 U4965 ( .A1(n8891), .A2(n8391), .ZN(n8203) );
  OR2_X1 U4966 ( .A1(n8174), .A2(n8466), .ZN(n8177) );
  INV_X1 U4967 ( .A(n8610), .ZN(n6596) );
  OR2_X1 U4968 ( .A1(n9340), .A2(n9264), .ZN(n7983) );
  AND2_X1 U4969 ( .A1(n9340), .A2(n9264), .ZN(n7986) );
  OR2_X1 U4970 ( .A1(n9655), .A2(n5933), .ZN(n7963) );
  NAND2_X1 U4971 ( .A1(n9736), .A2(n6030), .ZN(n7954) );
  OR2_X1 U4972 ( .A1(n9224), .A2(n5736), .ZN(n7889) );
  OR2_X1 U4973 ( .A1(n7812), .A2(n5708), .ZN(n8006) );
  NAND2_X1 U4974 ( .A1(n6349), .A2(n6348), .ZN(n9363) );
  OR2_X1 U4975 ( .A1(n9741), .A2(n9426), .ZN(n7958) );
  OR2_X1 U4976 ( .A1(n9202), .A2(n9276), .ZN(n6006) );
  NAND2_X1 U4977 ( .A1(n4722), .A2(n5444), .ZN(n5456) );
  NAND2_X1 U4978 ( .A1(n5443), .A2(n5442), .ZN(n4722) );
  OAI21_X1 U4979 ( .B1(n5313), .B2(n5312), .A(n5311), .ZN(n5315) );
  INV_X1 U4980 ( .A(n4847), .ZN(n4846) );
  INV_X1 U4981 ( .A(n4950), .ZN(n4468) );
  NAND2_X1 U4982 ( .A1(n4944), .A2(n4943), .ZN(n5265) );
  NAND2_X1 U4983 ( .A1(n4403), .A2(n4926), .ZN(n5204) );
  NAND2_X1 U4984 ( .A1(n4925), .A2(SI_12_), .ZN(n4926) );
  NAND2_X1 U4985 ( .A1(n4400), .A2(n4398), .ZN(n4403) );
  XNOR2_X1 U4986 ( .A(n4929), .B(SI_13_), .ZN(n5203) );
  XNOR2_X1 U4987 ( .A(n4924), .B(SI_12_), .ZN(n5189) );
  NAND2_X1 U4988 ( .A1(n4732), .A2(n4734), .ZN(n5129) );
  AOI21_X1 U4989 ( .B1(n5110), .B2(n4735), .A(n4339), .ZN(n4734) );
  OAI21_X1 U4990 ( .B1(n8368), .B2(n4651), .A(n4649), .ZN(n8077) );
  AOI21_X1 U4991 ( .B1(n8073), .B2(n4650), .A(n4356), .ZN(n4649) );
  INV_X1 U4992 ( .A(n8073), .ZN(n4651) );
  NAND4_X1 U4993 ( .A1(n5016), .A2(n5015), .A3(n5014), .A4(n5013), .ZN(n6625)
         );
  OR2_X1 U4994 ( .A1(n5038), .A2(n5012), .ZN(n5016) );
  NOR2_X1 U4995 ( .A1(n4527), .A2(n6939), .ZN(n4526) );
  INV_X1 U4996 ( .A(n10053), .ZN(n4524) );
  OR2_X1 U4997 ( .A1(n5353), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5373) );
  NOR2_X1 U4998 ( .A1(n4328), .A2(n4588), .ZN(n4587) );
  INV_X1 U4999 ( .A(n5053), .ZN(n4588) );
  NAND2_X1 U5000 ( .A1(n6625), .A2(n10067), .ZN(n8107) );
  NAND2_X1 U5001 ( .A1(n8104), .A2(n6778), .ZN(n8108) );
  OR2_X1 U5002 ( .A1(n6783), .A2(n7772), .ZN(n6778) );
  AOI21_X1 U5003 ( .B1(n4305), .B2(n4437), .A(n4433), .ZN(n4432) );
  NAND2_X1 U5004 ( .A1(n4437), .A2(n4435), .ZN(n4434) );
  AOI21_X1 U5005 ( .B1(n4297), .B2(n4300), .A(n4342), .ZN(n4615) );
  OR2_X1 U5006 ( .A1(n8867), .A2(n8692), .ZN(n8222) );
  AND2_X1 U5007 ( .A1(n8760), .A2(n8462), .ZN(n5294) );
  OR2_X1 U5008 ( .A1(n8817), .A2(n8729), .ZN(n8211) );
  INV_X1 U5009 ( .A(n8253), .ZN(n5299) );
  AND2_X1 U5010 ( .A1(n4816), .A2(n4972), .ZN(n4813) );
  NOR2_X1 U5011 ( .A1(n7388), .A2(n4795), .ZN(n4794) );
  INV_X1 U5012 ( .A(n6149), .ZN(n4795) );
  AOI21_X1 U5013 ( .B1(n4766), .B2(n4767), .A(n4764), .ZN(n4763) );
  INV_X1 U5014 ( .A(n9242), .ZN(n4764) );
  NAND2_X1 U5015 ( .A1(n9351), .A2(n7963), .ZN(n9348) );
  XNOR2_X1 U5016 ( .A(n9363), .B(n9265), .ZN(n9353) );
  OR2_X1 U5017 ( .A1(n5917), .A2(n5916), .ZN(n9364) );
  AOI21_X1 U5018 ( .B1(n4836), .B2(n4838), .A(n4362), .ZN(n4834) );
  INV_X1 U5019 ( .A(n4836), .ZN(n4835) );
  NAND2_X1 U5020 ( .A1(n9437), .A2(n5890), .ZN(n9436) );
  INV_X1 U5021 ( .A(n9471), .ZN(n4842) );
  OR2_X1 U5022 ( .A1(n9723), .A2(n6007), .ZN(n8014) );
  NAND2_X1 U5023 ( .A1(n6837), .A2(n7995), .ZN(n5623) );
  AND2_X1 U5024 ( .A1(n5987), .A2(n9790), .ZN(n6368) );
  AND2_X1 U5025 ( .A1(n5574), .A2(n4860), .ZN(n4647) );
  NOR2_X1 U5026 ( .A1(n5346), .A2(n4745), .ZN(n4744) );
  INV_X1 U5027 ( .A(n5328), .ZN(n4745) );
  AND2_X1 U5028 ( .A1(n5365), .A2(n5351), .ZN(n5363) );
  INV_X1 U5029 ( .A(n8664), .ZN(n8644) );
  NAND2_X1 U5030 ( .A1(n4686), .A2(n4689), .ZN(n8400) );
  AOI22_X1 U5031 ( .A1(n4298), .A2(n8388), .B1(n8463), .B2(n4690), .ZN(n4689)
         );
  OR2_X1 U5032 ( .A1(n5510), .A2(n7198), .ZN(n4430) );
  AOI21_X1 U5033 ( .B1(n5509), .B2(n8769), .A(n4429), .ZN(n4428) );
  INV_X1 U5034 ( .A(n5508), .ZN(n4429) );
  NAND2_X1 U5035 ( .A1(n6100), .A2(n6099), .ZN(n6810) );
  NOR2_X1 U5036 ( .A1(n6360), .A2(n9617), .ZN(n9336) );
  NAND2_X1 U5037 ( .A1(n4388), .A2(n8120), .ZN(n8140) );
  OAI21_X1 U5038 ( .B1(n8118), .B2(n8119), .A(n8117), .ZN(n4388) );
  AND2_X1 U5039 ( .A1(n8152), .A2(n8146), .ZN(n8129) );
  OAI21_X1 U5040 ( .B1(n8166), .B2(n8291), .A(n8165), .ZN(n8167) );
  MUX2_X1 U5041 ( .A(n8155), .B(n8154), .S(n8264), .Z(n8166) );
  INV_X1 U5042 ( .A(n8185), .ZN(n4540) );
  OAI21_X1 U5043 ( .B1(n8185), .B2(n4539), .A(n8295), .ZN(n4538) );
  NAND2_X1 U5044 ( .A1(n8210), .A2(n8264), .ZN(n4557) );
  INV_X1 U5045 ( .A(n7906), .ZN(n4406) );
  NAND2_X1 U5046 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  INV_X1 U5047 ( .A(n8218), .ZN(n4552) );
  INV_X1 U5048 ( .A(n5296), .ZN(n4463) );
  NAND2_X1 U5049 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  OAI21_X1 U5050 ( .B1(n7960), .B2(n7959), .A(n4472), .ZN(n4396) );
  NAND2_X1 U5051 ( .A1(n9353), .A2(n4316), .ZN(n4417) );
  INV_X1 U5052 ( .A(n9408), .ZN(n6030) );
  NOR2_X1 U5053 ( .A1(n9655), .A2(n9736), .ZN(n4495) );
  INV_X1 U5054 ( .A(n9529), .ZN(n4629) );
  NAND2_X1 U5055 ( .A1(n5460), .A2(n5459), .ZN(n6338) );
  NAND2_X1 U5056 ( .A1(n5456), .A2(n5455), .ZN(n5460) );
  OAI211_X1 U5057 ( .C1(n4502), .C2(P1_DATAO_REG_8__SCAN_IN), .A(n4500), .B(
        n4499), .ZN(n4910) );
  INV_X1 U5058 ( .A(n4668), .ZN(n4665) );
  NAND2_X1 U5059 ( .A1(n6612), .A2(n6571), .ZN(n6572) );
  NAND2_X1 U5060 ( .A1(n4394), .A2(n4393), .ZN(n6573) );
  INV_X1 U5061 ( .A(n6572), .ZN(n4394) );
  OR2_X1 U5062 ( .A1(n7708), .A2(n7707), .ZN(n7710) );
  NAND2_X1 U5063 ( .A1(n4510), .A2(n8486), .ZN(n4507) );
  OR2_X1 U5064 ( .A1(n7718), .A2(n4508), .ZN(n4506) );
  NAND2_X1 U5065 ( .A1(n4510), .A2(n4509), .ZN(n4508) );
  INV_X1 U5066 ( .A(n7719), .ZN(n4509) );
  NOR2_X1 U5067 ( .A1(n8613), .A2(n8758), .ZN(n4721) );
  OR2_X1 U5068 ( .A1(n8829), .A2(n8774), .ZN(n8198) );
  NAND2_X1 U5069 ( .A1(n4805), .A2(n8287), .ZN(n4455) );
  INV_X1 U5070 ( .A(n8143), .ZN(n4805) );
  AND2_X1 U5071 ( .A1(n8126), .A2(n7099), .ZN(n8131) );
  INV_X1 U5072 ( .A(n8146), .ZN(n4802) );
  OR2_X1 U5073 ( .A1(n8454), .A2(n8792), .ZN(n8242) );
  INV_X1 U5074 ( .A(n8851), .ZN(n5399) );
  NOR2_X1 U5075 ( .A1(n4443), .A2(n8271), .ZN(n4440) );
  INV_X1 U5076 ( .A(n8234), .ZN(n4443) );
  OR2_X1 U5077 ( .A1(n8851), .A2(n8080), .ZN(n8234) );
  NAND2_X1 U5078 ( .A1(n8851), .A2(n8080), .ZN(n8235) );
  NAND2_X1 U5079 ( .A1(n4344), .A2(n4613), .ZN(n4611) );
  NOR2_X1 U5080 ( .A1(n5201), .A2(n4610), .ZN(n4609) );
  INV_X1 U5081 ( .A(n5188), .ZN(n4610) );
  NOR2_X1 U5082 ( .A1(n4777), .A2(n4773), .ZN(n4772) );
  INV_X1 U5083 ( .A(n6211), .ZN(n4773) );
  INV_X1 U5084 ( .A(n9167), .ZN(n4777) );
  INV_X1 U5085 ( .A(n6216), .ZN(n4776) );
  AOI22_X1 U5086 ( .A1(n9288), .A2(n6311), .B1(n6101), .B2(n7024), .ZN(n6082)
         );
  NOR2_X1 U5087 ( .A1(n6267), .A2(n4791), .ZN(n4790) );
  INV_X1 U5088 ( .A(n6265), .ZN(n4791) );
  INV_X1 U5089 ( .A(n5712), .ZN(n5739) );
  NOR2_X1 U5090 ( .A1(n9363), .A2(n4494), .ZN(n4493) );
  INV_X1 U5091 ( .A(n4495), .ZN(n4494) );
  OR2_X1 U5092 ( .A1(n9671), .A2(n9410), .ZN(n7957) );
  NOR2_X1 U5093 ( .A1(n9504), .A2(n9752), .ZN(n9455) );
  NOR2_X1 U5094 ( .A1(n9521), .A2(n9766), .ZN(n4483) );
  OR2_X1 U5095 ( .A1(n9521), .A2(n9501), .ZN(n9492) );
  NAND2_X1 U5096 ( .A1(n9530), .A2(n9529), .ZN(n4633) );
  AOI21_X1 U5097 ( .B1(n4854), .B2(n7210), .A(n9954), .ZN(n4852) );
  INV_X1 U5098 ( .A(n4854), .ZN(n4853) );
  INV_X1 U5099 ( .A(n7854), .ZN(n4624) );
  OR2_X1 U5100 ( .A1(n9159), .A2(n6874), .ZN(n4486) );
  NAND2_X1 U5101 ( .A1(n9406), .A2(n9407), .ZN(n9405) );
  AND2_X1 U5102 ( .A1(n9680), .A2(n9475), .ZN(n6024) );
  OAI21_X1 U5103 ( .B1(n4866), .B2(n4827), .A(n6016), .ZN(n4826) );
  NAND2_X1 U5104 ( .A1(n6813), .A2(n6874), .ZN(n7852) );
  NAND2_X1 U5105 ( .A1(n8001), .A2(n7854), .ZN(n7842) );
  AND2_X1 U5106 ( .A1(n7027), .A2(n5949), .ZN(n6859) );
  AND2_X1 U5107 ( .A1(n5570), .A2(n4489), .ZN(n4490) );
  NAND2_X1 U5108 ( .A1(n5422), .A2(n5421), .ZN(n5443) );
  AND4_X1 U5109 ( .A1(n4645), .A2(n4644), .A3(n4490), .A4(n4860), .ZN(n5586)
         );
  NAND2_X1 U5110 ( .A1(n4301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5937) );
  INV_X1 U5111 ( .A(n4465), .ZN(n4464) );
  OAI21_X1 U5112 ( .B1(n4470), .B2(n4466), .A(n4953), .ZN(n4465) );
  NAND2_X1 U5113 ( .A1(n4940), .A2(n4939), .ZN(n5249) );
  NAND2_X1 U5114 ( .A1(n4923), .A2(n4922), .ZN(n5177) );
  NAND2_X1 U5115 ( .A1(n4912), .A2(n4913), .ZN(n5133) );
  XNOR2_X1 U5116 ( .A(n4905), .B(SI_7_), .ZN(n5128) );
  INV_X1 U5117 ( .A(SI_6_), .ZN(n9033) );
  OAI21_X1 U5118 ( .B1(n6388), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4454), .ZN(
        n4884) );
  NAND2_X1 U5119 ( .A1(n6388), .A2(n6398), .ZN(n4454) );
  NOR2_X1 U5120 ( .A1(n8066), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5121 ( .A1(n8065), .A2(n4332), .ZN(n4660) );
  NOR2_X1 U5122 ( .A1(n4670), .A2(n7543), .ZN(n4668) );
  AND2_X1 U5123 ( .A1(n8159), .A2(n8157), .ZN(n7536) );
  OR2_X1 U5124 ( .A1(n8400), .A2(n8401), .ZN(n8399) );
  OR2_X1 U5125 ( .A1(n6820), .A2(n4676), .ZN(n4673) );
  OR2_X1 U5126 ( .A1(n7080), .A2(n6821), .ZN(n4676) );
  OR2_X1 U5127 ( .A1(n7079), .A2(n8474), .ZN(n4674) );
  OR2_X1 U5128 ( .A1(n7080), .A2(n4677), .ZN(n4675) );
  NOR2_X1 U5129 ( .A1(n8085), .A2(n8409), .ZN(n4871) );
  NAND2_X1 U5130 ( .A1(n8269), .A2(n8268), .ZN(n4561) );
  NAND2_X1 U5131 ( .A1(n4753), .A2(n4330), .ZN(n4752) );
  AND2_X1 U5132 ( .A1(n7128), .A2(n7127), .ZN(n8628) );
  AND2_X1 U5133 ( .A1(n5453), .A2(n5452), .ZN(n8643) );
  XNOR2_X1 U5134 ( .A(n6555), .B(n6695), .ZN(n6689) );
  OAI21_X1 U5135 ( .B1(n6579), .B2(n6678), .A(n4571), .ZN(n6700) );
  NAND2_X1 U5136 ( .A1(n6579), .A2(n6678), .ZN(n4571) );
  OAI21_X1 U5137 ( .B1(n6579), .B2(n5040), .A(n4395), .ZN(n6703) );
  NAND2_X1 U5138 ( .A1(n6579), .A2(n5040), .ZN(n4395) );
  OR2_X1 U5139 ( .A1(n6581), .A2(n6720), .ZN(n6582) );
  OR2_X1 U5140 ( .A1(n6734), .A2(n6733), .ZN(n4514) );
  OR2_X1 U5141 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  AOI21_X1 U5142 ( .B1(n6589), .B2(n4569), .A(n4380), .ZN(n4568) );
  INV_X1 U5143 ( .A(n6589), .ZN(n4570) );
  NAND2_X1 U5144 ( .A1(n6736), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6735) );
  OR2_X1 U5145 ( .A1(n6796), .A2(n6939), .ZN(n6797) );
  AOI21_X1 U5146 ( .B1(n4524), .B2(n4526), .A(n6930), .ZN(n4521) );
  INV_X1 U5147 ( .A(n7147), .ZN(n4710) );
  NAND2_X1 U5148 ( .A1(n6946), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U5149 ( .A1(n4586), .A2(n7508), .ZN(n4585) );
  NAND2_X1 U5150 ( .A1(n4585), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4584) );
  NOR2_X1 U5151 ( .A1(n7509), .A2(n7510), .ZN(n7511) );
  OR2_X1 U5152 ( .A1(n7511), .A2(n7512), .ZN(n4503) );
  AND2_X1 U5153 ( .A1(n7492), .A2(n7519), .ZN(n7632) );
  NOR2_X1 U5154 ( .A1(n7494), .A2(n7506), .ZN(n7631) );
  NAND2_X1 U5155 ( .A1(n4712), .A2(n4711), .ZN(n7703) );
  INV_X1 U5156 ( .A(n7634), .ZN(n4711) );
  NAND2_X1 U5157 ( .A1(n4582), .A2(n7725), .ZN(n4580) );
  INV_X1 U5158 ( .A(n7710), .ZN(n4582) );
  OR2_X1 U5159 ( .A1(n8537), .A2(n8536), .ZN(n4700) );
  INV_X1 U5160 ( .A(n4699), .ZN(n8560) );
  NOR2_X1 U5161 ( .A1(n8577), .A2(n8578), .ZN(n8581) );
  NOR2_X1 U5162 ( .A1(n8454), .A2(n8773), .ZN(n6045) );
  NOR2_X1 U5163 ( .A1(n8643), .A2(n8775), .ZN(n8646) );
  NAND2_X1 U5164 ( .A1(n5391), .A2(n5390), .ZN(n5410) );
  NAND2_X1 U5165 ( .A1(n5320), .A2(n5319), .ZN(n5337) );
  OR2_X1 U5166 ( .A1(n5287), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5304) );
  AND2_X1 U5167 ( .A1(n4419), .A2(n4421), .ZN(n7610) );
  INV_X1 U5168 ( .A(n4422), .ZN(n4421) );
  OAI21_X1 U5169 ( .B1(n4427), .B2(n4423), .A(n8187), .ZN(n4422) );
  AND4_X1 U5170 ( .A1(n5276), .A2(n5275), .A3(n5274), .A4(n5273), .ZN(n8391)
         );
  NAND2_X1 U5171 ( .A1(n4991), .A2(n4990), .ZN(n5223) );
  INV_X1 U5172 ( .A(n5209), .ZN(n4991) );
  OR2_X1 U5173 ( .A1(n7368), .A2(n7536), .ZN(n7369) );
  OR2_X1 U5174 ( .A1(n5169), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5182) );
  OR2_X1 U5175 ( .A1(n10106), .A2(n7418), .ZN(n8130) );
  AND4_X1 U5176 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n7537)
         );
  INV_X1 U5177 ( .A(n8470), .ZN(n7418) );
  NAND2_X1 U5178 ( .A1(n4617), .A2(n5132), .ZN(n7101) );
  NAND2_X1 U5179 ( .A1(n7038), .A2(n5483), .ZN(n4617) );
  AND2_X1 U5180 ( .A1(n8113), .A2(n8107), .ZN(n4806) );
  INV_X1 U5181 ( .A(n8119), .ZN(n8279) );
  NAND2_X1 U5182 ( .A1(n8242), .A2(n8243), .ZN(n8641) );
  NAND2_X1 U5183 ( .A1(n8234), .A2(n8235), .ZN(n8670) );
  OR2_X1 U5184 ( .A1(n8677), .A2(n4300), .ZN(n4616) );
  NAND2_X1 U5185 ( .A1(n4819), .A2(n4334), .ZN(n8675) );
  INV_X1 U5186 ( .A(n8274), .ZN(n4820) );
  AND2_X1 U5187 ( .A1(n5379), .A2(n5378), .ZN(n8693) );
  OR2_X1 U5188 ( .A1(n8274), .A2(n8273), .ZN(n8689) );
  NAND2_X1 U5189 ( .A1(n4594), .A2(n4591), .ZN(n8705) );
  INV_X1 U5190 ( .A(n4592), .ZN(n4591) );
  OAI22_X1 U5191 ( .A1(n4593), .A2(n8716), .B1(n8873), .B2(n8706), .ZN(n4592)
         );
  NAND2_X1 U5192 ( .A1(n4598), .A2(n4603), .ZN(n4597) );
  INV_X1 U5193 ( .A(n4601), .ZN(n4598) );
  NAND2_X1 U5194 ( .A1(n4603), .A2(n4600), .ZN(n4599) );
  AND2_X1 U5195 ( .A1(n8219), .A2(n8220), .ZN(n8716) );
  AND2_X1 U5196 ( .A1(n8217), .A2(n8713), .ZN(n8727) );
  NAND2_X1 U5197 ( .A1(n4450), .A2(n4451), .ZN(n8743) );
  NAND2_X1 U5198 ( .A1(n8743), .A2(n8742), .ZN(n8741) );
  NAND2_X1 U5199 ( .A1(n5301), .A2(n5300), .ZN(n8817) );
  AND4_X1 U5200 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8776)
         );
  INV_X1 U5201 ( .A(n8750), .ZN(n8773) );
  OR2_X1 U5202 ( .A1(n8256), .A2(n6662), .ZN(n8775) );
  NOR2_X1 U5203 ( .A1(n8183), .A2(n4426), .ZN(n4425) );
  INV_X1 U5204 ( .A(n5489), .ZN(n4426) );
  NAND2_X1 U5205 ( .A1(n5208), .A2(n5207), .ZN(n8174) );
  AND2_X1 U5206 ( .A1(n8264), .A2(n6662), .ZN(n8750) );
  INV_X1 U5207 ( .A(n8775), .ZN(n8752) );
  NOR2_X1 U5208 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4811) );
  INV_X1 U5209 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5004) );
  NOR2_X1 U5210 ( .A1(n5049), .A2(n4965), .ZN(n5148) );
  OR2_X1 U5211 ( .A1(n5088), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U5212 ( .A1(n4564), .A2(n4563), .ZN(n5088) );
  INV_X1 U5213 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4563) );
  INV_X1 U5214 ( .A(n5049), .ZN(n4564) );
  NAND2_X1 U5215 ( .A1(n5047), .A2(n4961), .ZN(n5049) );
  NAND2_X1 U5216 ( .A1(n5147), .A2(n4961), .ZN(n4703) );
  INV_X1 U5217 ( .A(n6267), .ZN(n4787) );
  NAND2_X1 U5218 ( .A1(n7468), .A2(n6345), .ZN(n4477) );
  NAND2_X1 U5219 ( .A1(n5786), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5797) );
  INV_X1 U5220 ( .A(n9285), .ZN(n6872) );
  NAND2_X1 U5221 ( .A1(n6141), .A2(n4797), .ZN(n4796) );
  AND2_X1 U5222 ( .A1(n4318), .A2(n6140), .ZN(n4797) );
  INV_X1 U5223 ( .A(n9844), .ZN(n4761) );
  NAND2_X1 U5224 ( .A1(n4345), .A2(n4770), .ZN(n4766) );
  OR2_X1 U5225 ( .A1(n9176), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U5226 ( .A1(n4770), .A2(n6283), .ZN(n4767) );
  CLKBUF_X1 U5227 ( .A(n9143), .Z(n9144) );
  NOR2_X1 U5228 ( .A1(n7983), .A2(n7984), .ZN(n4476) );
  OR3_X1 U5229 ( .A1(n8036), .A2(n7986), .A3(n7834), .ZN(n7979) );
  NAND2_X1 U5230 ( .A1(n5645), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5613) );
  NOR2_X1 U5231 ( .A1(n9445), .A2(n9671), .ZN(n9428) );
  INV_X1 U5232 ( .A(n9266), .ZN(n9426) );
  OR2_X1 U5233 ( .A1(n9676), .A2(n9425), .ZN(n7777) );
  INV_X1 U5234 ( .A(n9423), .ZN(n5901) );
  NAND2_X1 U5235 ( .A1(n5878), .A2(n9461), .ZN(n9437) );
  NAND2_X1 U5236 ( .A1(n9551), .A2(n4481), .ZN(n9504) );
  NOR2_X1 U5237 ( .A1(n9757), .A2(n4482), .ZN(n4481) );
  INV_X1 U5238 ( .A(n4483), .ZN(n4482) );
  AND2_X1 U5239 ( .A1(n5815), .A2(n8019), .ZN(n4626) );
  OAI21_X1 U5240 ( .B1(n5778), .B2(n4642), .A(n4640), .ZN(n9577) );
  AOI21_X1 U5241 ( .B1(n4643), .B2(n9611), .A(n4641), .ZN(n4640) );
  INV_X1 U5242 ( .A(n4643), .ZN(n4642) );
  INV_X1 U5243 ( .A(n7905), .ZN(n4641) );
  INV_X1 U5244 ( .A(n6012), .ZN(n9576) );
  AND2_X1 U5245 ( .A1(n9592), .A2(n8014), .ZN(n4643) );
  NAND2_X1 U5246 ( .A1(n5778), .A2(n5777), .ZN(n9608) );
  OR2_X1 U5247 ( .A1(n7449), .A2(n9130), .ZN(n7567) );
  NOR2_X1 U5248 ( .A1(n7567), .A2(n9202), .ZN(n9616) );
  OR2_X1 U5249 ( .A1(n9130), .A2(n5751), .ZN(n7890) );
  INV_X1 U5250 ( .A(n4634), .ZN(n4635) );
  OAI21_X1 U5251 ( .B1(n5737), .B2(n4639), .A(n7820), .ZN(n4634) );
  OR2_X1 U5252 ( .A1(n7358), .A2(n7811), .ZN(n7403) );
  AOI21_X1 U5253 ( .B1(n7808), .B2(n4832), .A(n4337), .ZN(n4829) );
  NAND2_X1 U5254 ( .A1(n4831), .A2(n7089), .ZN(n4830) );
  NAND2_X1 U5255 ( .A1(n7089), .A2(n7088), .ZN(n7087) );
  INV_X1 U5256 ( .A(n9995), .ZN(n9595) );
  NOR2_X1 U5257 ( .A1(n9288), .A2(n9976), .ZN(n7802) );
  AOI21_X1 U5258 ( .B1(n4839), .B2(n6023), .A(n4837), .ZN(n4836) );
  INV_X1 U5259 ( .A(n9454), .ZN(n4837) );
  OR2_X1 U5260 ( .A1(n9757), .A2(n9268), .ZN(n6021) );
  NAND2_X1 U5261 ( .A1(n6748), .A2(n6345), .ZN(n4413) );
  INV_X1 U5262 ( .A(n6416), .ZN(n5833) );
  OR2_X1 U5263 ( .A1(n9130), .A2(n9277), .ZN(n6005) );
  NAND2_X1 U5264 ( .A1(n7855), .A2(n7852), .ZN(n7801) );
  AND2_X1 U5265 ( .A1(n5960), .A2(n5966), .ZN(n6410) );
  XNOR2_X1 U5266 ( .A(n5576), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5579) );
  INV_X1 U5267 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5573) );
  NOR2_X1 U5268 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5591) );
  XNOR2_X1 U5269 ( .A(n5456), .B(n5455), .ZN(n7729) );
  OAI21_X1 U5270 ( .B1(n4860), .B2(n9791), .A(n5584), .ZN(n4859) );
  XNOR2_X1 U5271 ( .A(n5420), .B(n5419), .ZN(n7680) );
  XNOR2_X1 U5272 ( .A(n5401), .B(n5400), .ZN(n7629) );
  INV_X1 U5273 ( .A(n5345), .ZN(n4743) );
  OAI21_X1 U5274 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(n5347) );
  XNOR2_X1 U5275 ( .A(n5937), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U5276 ( .A1(n4645), .A2(n4644), .ZN(n5938) );
  NAND2_X1 U5277 ( .A1(n4469), .A2(n4950), .ZN(n5279) );
  NAND2_X1 U5278 ( .A1(n4471), .A2(n4470), .ZN(n4469) );
  INV_X1 U5279 ( .A(n5265), .ZN(n4471) );
  XNOR2_X1 U5280 ( .A(n5217), .B(n5216), .ZN(n6748) );
  NAND2_X1 U5281 ( .A1(n4746), .A2(n4930), .ZN(n5217) );
  NAND2_X1 U5282 ( .A1(n4400), .A2(n4923), .ZN(n5190) );
  NAND2_X1 U5283 ( .A1(n4724), .A2(n4725), .ZN(n5162) );
  OR2_X1 U5284 ( .A1(n5134), .A2(n4728), .ZN(n4724) );
  XNOR2_X1 U5285 ( .A(n4903), .B(n9033), .ZN(n5110) );
  NAND2_X1 U5286 ( .A1(n5086), .A2(n4446), .ZN(n4444) );
  INV_X1 U5287 ( .A(n5506), .ZN(n6382) );
  AND4_X1 U5288 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n7113)
         );
  NAND2_X1 U5289 ( .A1(n4685), .A2(n8089), .ZN(n8344) );
  AND2_X1 U5290 ( .A1(n5343), .A2(n5342), .ZN(n8692) );
  XNOR2_X1 U5291 ( .A(n8077), .B(n8075), .ZN(n8352) );
  AND3_X1 U5292 ( .A1(n5011), .A2(n5010), .A3(n5009), .ZN(n8740) );
  AOI21_X1 U5293 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4679) );
  INV_X1 U5294 ( .A(n8092), .ZN(n4680) );
  INV_X1 U5295 ( .A(n8448), .ZN(n4681) );
  AND2_X1 U5296 ( .A1(n5359), .A2(n5358), .ZN(n8430) );
  AND3_X1 U5297 ( .A1(n5309), .A2(n5308), .A3(n5307), .ZN(n8729) );
  AOI22_X1 U5298 ( .A1(n7689), .A2(n7688), .B1(n7694), .B2(n7687), .ZN(n7692)
         );
  NAND2_X1 U5299 ( .A1(n5416), .A2(n5415), .ZN(n8664) );
  INV_X1 U5300 ( .A(n8693), .ZN(n8665) );
  INV_X1 U5301 ( .A(n8430), .ZN(n8707) );
  INV_X1 U5302 ( .A(n8692), .ZN(n8718) );
  NAND2_X1 U5303 ( .A1(n7119), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5059) );
  OR2_X1 U5304 ( .A1(n5272), .A2(n7769), .ZN(n5029) );
  AOI21_X1 U5305 ( .B1(n6734), .B2(n4311), .A(n4511), .ZN(n6794) );
  INV_X1 U5306 ( .A(n4512), .ZN(n4511) );
  AOI21_X1 U5307 ( .B1(n4311), .B2(n6733), .A(n6790), .ZN(n4512) );
  NOR2_X1 U5308 ( .A1(n7138), .A2(n7137), .ZN(n7509) );
  OR2_X1 U5309 ( .A1(n7631), .A2(n7632), .ZN(n4712) );
  INV_X1 U5310 ( .A(n7703), .ZN(n7702) );
  AND3_X1 U5311 ( .A1(n4580), .A2(n8492), .A3(P2_REG1_REG_13__SCAN_IN), .ZN(
        n8493) );
  NOR2_X1 U5312 ( .A1(n8597), .A2(n8598), .ZN(n8601) );
  NOR2_X1 U5313 ( .A1(n8604), .A2(n4386), .ZN(n4385) );
  NOR2_X1 U5314 ( .A1(n4387), .A2(n8618), .ZN(n4386) );
  OAI21_X1 U5315 ( .B1(n4532), .B2(n10055), .A(n4529), .ZN(n4528) );
  XNOR2_X1 U5316 ( .A(n4534), .B(n4533), .ZN(n4532) );
  AOI21_X1 U5317 ( .B1(n8621), .B2(n10060), .A(n4530), .ZN(n4529) );
  INV_X1 U5318 ( .A(n8615), .ZN(n4533) );
  NAND2_X1 U5319 ( .A1(n5462), .A2(n5461), .ZN(n8337) );
  NAND2_X1 U5320 ( .A1(n4979), .A2(n4978), .ZN(n8734) );
  NAND2_X1 U5321 ( .A1(n5512), .A2(n10082), .ZN(n5513) );
  AOI21_X1 U5322 ( .B1(n7468), .B2(n8252), .A(n5352), .ZN(n8861) );
  AND2_X1 U5323 ( .A1(n4975), .A2(n4810), .ZN(n5000) );
  OR2_X1 U5324 ( .A1(n5471), .A2(n5147), .ZN(n5298) );
  NAND2_X1 U5325 ( .A1(n4477), .A2(n5870), .ZN(n9680) );
  NAND2_X1 U5326 ( .A1(n9241), .A2(n6304), .ZN(n6319) );
  AOI21_X1 U5327 ( .B1(n9094), .B2(n6254), .A(n6253), .ZN(n6264) );
  INV_X1 U5328 ( .A(n9856), .ZN(n9247) );
  AOI21_X1 U5329 ( .B1(n9651), .B2(n9637), .A(n9368), .ZN(n9369) );
  AOI21_X1 U5330 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9350) );
  NAND2_X1 U5331 ( .A1(n9360), .A2(n9648), .ZN(n9371) );
  INV_X1 U5332 ( .A(n9741), .ZN(n9404) );
  INV_X1 U5333 ( .A(n9752), .ZN(n9485) );
  INV_X1 U5334 ( .A(n9757), .ZN(n9508) );
  OR2_X1 U5335 ( .A1(n6324), .A2(n8047), .ZN(n9978) );
  OR2_X1 U5336 ( .A1(n5703), .A2(n6399), .ZN(n5607) );
  XNOR2_X1 U5337 ( .A(n9349), .B(n7832), .ZN(n9660) );
  NAND2_X1 U5338 ( .A1(n6358), .A2(n6416), .ZN(n9340) );
  NAND2_X1 U5339 ( .A1(n5602), .A2(n5601), .ZN(n6842) );
  AND2_X1 U5340 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  OR2_X1 U5341 ( .A1(n6416), .A2(n6538), .ZN(n5599) );
  AOI21_X1 U5342 ( .B1(n8105), .B2(n8104), .A(n4389), .ZN(n8111) );
  INV_X1 U5343 ( .A(n8107), .ZN(n4389) );
  NAND2_X1 U5344 ( .A1(n4543), .A2(n4542), .ZN(n8149) );
  NAND2_X1 U5345 ( .A1(n8129), .A2(n8256), .ZN(n4543) );
  AND2_X1 U5346 ( .A1(n8198), .A2(n8187), .ZN(n4541) );
  INV_X1 U5347 ( .A(n4538), .ZN(n4537) );
  NAND2_X1 U5348 ( .A1(n7990), .A2(n7975), .ZN(n4411) );
  NAND2_X1 U5349 ( .A1(n7898), .A2(n7897), .ZN(n4412) );
  NOR2_X1 U5350 ( .A1(n7902), .A2(n8016), .ZN(n4409) );
  NAND2_X1 U5351 ( .A1(n4555), .A2(n4324), .ZN(n4554) );
  INV_X1 U5352 ( .A(n8216), .ZN(n4556) );
  NOR2_X1 U5353 ( .A1(n8704), .A2(n8221), .ZN(n4550) );
  INV_X1 U5354 ( .A(n7910), .ZN(n4404) );
  NAND2_X1 U5355 ( .A1(n4407), .A2(n4406), .ZN(n4405) );
  NAND2_X1 U5356 ( .A1(n4549), .A2(n4548), .ZN(n4547) );
  NOR2_X1 U5357 ( .A1(n8228), .A2(n8264), .ZN(n4548) );
  AOI21_X1 U5358 ( .B1(n8233), .B2(n8264), .A(n8670), .ZN(n4546) );
  AND2_X1 U5359 ( .A1(n7958), .A2(n7957), .ZN(n4472) );
  NOR2_X1 U5360 ( .A1(n7943), .A2(n9438), .ZN(n4473) );
  AND2_X1 U5361 ( .A1(n9951), .A2(n6000), .ZN(n7866) );
  NAND2_X1 U5362 ( .A1(n8246), .A2(n4747), .ZN(n4748) );
  INV_X1 U5363 ( .A(n8250), .ZN(n4747) );
  INV_X1 U5364 ( .A(n8487), .ZN(n4510) );
  AND2_X1 U5365 ( .A1(n8582), .A2(n4504), .ZN(n8585) );
  NAND2_X1 U5366 ( .A1(n8583), .A2(n8596), .ZN(n4504) );
  NAND2_X1 U5367 ( .A1(n7536), .A2(n5188), .ZN(n4612) );
  INV_X1 U5368 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4966) );
  INV_X1 U5369 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9013) );
  INV_X1 U5370 ( .A(n5990), .ZN(n7806) );
  NOR2_X1 U5371 ( .A1(n9784), .A2(n9723), .ZN(n4480) );
  INV_X1 U5372 ( .A(n4744), .ZN(n4741) );
  INV_X1 U5373 ( .A(n5363), .ZN(n4740) );
  AOI21_X1 U5374 ( .B1(n4464), .B2(n4329), .A(n4461), .ZN(n4460) );
  INV_X1 U5375 ( .A(n4959), .ZN(n4461) );
  NAND2_X1 U5376 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  AND2_X1 U5377 ( .A1(n5234), .A2(n5232), .ZN(n4936) );
  NOR2_X1 U5378 ( .A1(n4927), .A2(n4399), .ZN(n4398) );
  INV_X1 U5379 ( .A(n4923), .ZN(n4399) );
  INV_X1 U5380 ( .A(n5189), .ZN(n4927) );
  AND2_X1 U5381 ( .A1(n4874), .A2(n4475), .ZN(n4729) );
  NAND2_X1 U5382 ( .A1(n4474), .A2(n4913), .ZN(n4475) );
  INV_X1 U5383 ( .A(n4912), .ZN(n4474) );
  NAND2_X1 U5384 ( .A1(n4914), .A2(n8998), .ZN(n4917) );
  NOR2_X1 U5385 ( .A1(n4733), .A2(n4731), .ZN(n4730) );
  INV_X1 U5386 ( .A(n5110), .ZN(n4731) );
  INV_X1 U5387 ( .A(n4902), .ZN(n4735) );
  INV_X1 U5388 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4497) );
  OR2_X1 U5389 ( .A1(n8425), .A2(n8692), .ZN(n8073) );
  INV_X1 U5390 ( .A(n8072), .ZN(n4650) );
  NOR2_X1 U5391 ( .A1(n8246), .A2(n8247), .ZN(n8251) );
  NAND2_X1 U5392 ( .A1(n8270), .A2(n4755), .ZN(n4754) );
  INV_X1 U5393 ( .A(n8310), .ZN(n4755) );
  NOR3_X1 U5394 ( .A1(n4800), .A2(n8316), .A3(n4799), .ZN(n4798) );
  NOR2_X1 U5395 ( .A1(n8307), .A2(n8838), .ZN(n4800) );
  NAND2_X1 U5396 ( .A1(n8838), .A2(n8460), .ZN(n8312) );
  NAND2_X1 U5397 ( .A1(n7703), .A2(n4873), .ZN(n7704) );
  INV_X1 U5398 ( .A(n8496), .ZN(n4581) );
  OR2_X1 U5399 ( .A1(n8509), .A2(n8508), .ZN(n8510) );
  AND2_X1 U5400 ( .A1(n4699), .A2(n4698), .ZN(n8595) );
  NAND2_X1 U5401 ( .A1(n8561), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4698) );
  OR2_X1 U5402 ( .A1(n8760), .A2(n8776), .ZN(n8204) );
  OR2_X1 U5403 ( .A1(n4425), .A2(n8184), .ZN(n4423) );
  INV_X1 U5404 ( .A(n8196), .ZN(n4427) );
  OR2_X1 U5405 ( .A1(n4427), .A2(n8184), .ZN(n4424) );
  NAND2_X1 U5406 ( .A1(n10106), .A2(n7418), .ZN(n8152) );
  NAND2_X1 U5407 ( .A1(n4983), .A2(n4982), .ZN(n5103) );
  INV_X1 U5408 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4982) );
  INV_X1 U5409 ( .A(n5080), .ZN(n4983) );
  NAND2_X1 U5410 ( .A1(n6676), .A2(n8119), .ZN(n4589) );
  NAND2_X1 U5411 ( .A1(n8622), .A2(n5511), .ZN(n6644) );
  NAND2_X1 U5412 ( .A1(n4597), .A2(n4599), .ZN(n4593) );
  NOR2_X1 U5413 ( .A1(n4596), .A2(n8716), .ZN(n4595) );
  INV_X1 U5414 ( .A(n4597), .ZN(n4596) );
  NAND2_X1 U5415 ( .A1(n4818), .A2(n4600), .ZN(n4817) );
  AOI21_X1 U5416 ( .B1(n4807), .B2(n4453), .A(n4452), .ZN(n4451) );
  INV_X1 U5417 ( .A(n8203), .ZN(n4453) );
  INV_X1 U5418 ( .A(n8204), .ZN(n4452) );
  INV_X1 U5419 ( .A(n4807), .ZN(n4448) );
  OR2_X1 U5420 ( .A1(n10117), .A2(n7537), .ZN(n8159) );
  NAND2_X1 U5421 ( .A1(n4975), .A2(n4974), .ZN(n5529) );
  INV_X2 U5422 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U5423 ( .A1(n5218), .A2(n9020), .ZN(n5283) );
  NAND3_X1 U5424 ( .A1(n4964), .A2(n4963), .A3(n4962), .ZN(n4965) );
  NAND2_X1 U5425 ( .A1(n4789), .A2(n4783), .ZN(n4782) );
  INV_X1 U5426 ( .A(n4790), .ZN(n4783) );
  NOR2_X1 U5427 ( .A1(n5838), .A2(n5837), .ZN(n5846) );
  INV_X1 U5428 ( .A(n9220), .ZN(n4760) );
  AOI21_X1 U5429 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n7974) );
  AND2_X1 U5430 ( .A1(n7969), .A2(n7970), .ZN(n4414) );
  AOI21_X1 U5431 ( .B1(n7966), .B2(n7975), .A(n4417), .ZN(n4416) );
  NAND2_X1 U5432 ( .A1(n7830), .A2(n7954), .ZN(n4621) );
  INV_X1 U5433 ( .A(n7954), .ZN(n4622) );
  INV_X1 U5434 ( .A(n5883), .ZN(n5882) );
  INV_X1 U5435 ( .A(n5745), .ZN(n5743) );
  INV_X1 U5436 ( .A(n7889), .ZN(n4639) );
  AND2_X1 U5437 ( .A1(n5951), .A2(n4456), .ZN(n7352) );
  NAND2_X1 U5438 ( .A1(n5695), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5683) );
  INV_X1 U5439 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5675) );
  NOR2_X1 U5440 ( .A1(n5683), .A2(n5675), .ZN(n5677) );
  AND2_X1 U5441 ( .A1(n7808), .A2(n7088), .ZN(n4831) );
  INV_X1 U5442 ( .A(n5998), .ZN(n4832) );
  NAND2_X1 U5443 ( .A1(n6035), .A2(n8049), .ZN(n6072) );
  AOI21_X1 U5444 ( .B1(n4299), .B2(n4622), .A(n7967), .ZN(n4618) );
  NAND2_X1 U5445 ( .A1(n9420), .A2(n7956), .ZN(n9406) );
  OR2_X1 U5446 ( .A1(n9444), .A2(n9676), .ZN(n9445) );
  AND2_X1 U5447 ( .A1(n5863), .A2(n4628), .ZN(n4627) );
  NAND2_X1 U5448 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U5449 ( .A1(n4633), .A2(n4630), .ZN(n9493) );
  NAND2_X1 U5450 ( .A1(n9556), .A2(n6015), .ZN(n4828) );
  AND2_X1 U5451 ( .A1(n9616), .A2(n4478), .ZN(n9567) );
  AND2_X1 U5452 ( .A1(n4302), .A2(n9570), .ZN(n4478) );
  NAND2_X1 U5453 ( .A1(n9616), .A2(n4302), .ZN(n9581) );
  NAND2_X1 U5454 ( .A1(n9616), .A2(n4480), .ZN(n9598) );
  NOR2_X1 U5455 ( .A1(n6085), .A2(n7024), .ZN(n7027) );
  OAI21_X1 U5456 ( .B1(n6341), .B2(n6340), .A(n6339), .ZN(n6352) );
  OR2_X1 U5457 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  XNOR2_X1 U5458 ( .A(n6338), .B(n6337), .ZN(n6341) );
  AND2_X1 U5459 ( .A1(n5421), .A2(n5407), .ZN(n5419) );
  INV_X1 U5460 ( .A(n5264), .ZN(n4470) );
  NAND2_X1 U5461 ( .A1(n5569), .A2(n4848), .ZN(n4847) );
  INV_X1 U5462 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5569) );
  INV_X1 U5463 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4848) );
  INV_X1 U5464 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U5465 ( .A1(n4931), .A2(n9004), .ZN(n5232) );
  INV_X1 U5466 ( .A(n5203), .ZN(n4928) );
  NAND3_X1 U5467 ( .A1(n4402), .A2(n4723), .A3(n4401), .ZN(n4400) );
  AND2_X1 U5468 ( .A1(n5711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5712) );
  AOI21_X1 U5469 ( .B1(n4729), .B2(n4727), .A(n4726), .ZN(n4725) );
  INV_X1 U5470 ( .A(n4913), .ZN(n4727) );
  INV_X1 U5471 ( .A(n4917), .ZN(n4726) );
  INV_X1 U5472 ( .A(n4729), .ZN(n4728) );
  OR3_X1 U5473 ( .A1(n5669), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n5710) );
  INV_X1 U5474 ( .A(n4896), .ZN(n4446) );
  OAI21_X1 U5475 ( .B1(n6389), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4893), .ZN(
        n4894) );
  INV_X1 U5476 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4880) );
  AND2_X1 U5477 ( .A1(n8415), .A2(n8063), .ZN(n8360) );
  INV_X1 U5478 ( .A(n8089), .ZN(n4684) );
  XNOR2_X1 U5479 ( .A(n8249), .B(n8461), .ZN(n8302) );
  NOR2_X1 U5480 ( .A1(n7541), .A2(n7540), .ZN(n4670) );
  NAND2_X1 U5481 ( .A1(n7422), .A2(n4671), .ZN(n4669) );
  NOR2_X1 U5482 ( .A1(n4688), .A2(n4360), .ZN(n4687) );
  INV_X1 U5483 ( .A(n7691), .ZN(n4688) );
  AOI21_X1 U5484 ( .B1(n4656), .B2(n4659), .A(n4654), .ZN(n4653) );
  INV_X1 U5485 ( .A(n8416), .ZN(n4654) );
  NAND2_X1 U5486 ( .A1(n4309), .A2(n4671), .ZN(n4666) );
  NAND2_X1 U5487 ( .A1(n4309), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5488 ( .A1(n6699), .A2(n6700), .ZN(n6698) );
  AND2_X1 U5489 ( .A1(n6609), .A2(n6569), .ZN(n6724) );
  NAND2_X1 U5490 ( .A1(n4392), .A2(n4391), .ZN(n6569) );
  NAND2_X1 U5491 ( .A1(n6724), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U5492 ( .A1(n6722), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6721) );
  AOI21_X1 U5493 ( .B1(n6574), .B2(n4708), .A(n4383), .ZN(n4707) );
  NAND2_X1 U5494 ( .A1(n4381), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6737) );
  INV_X1 U5495 ( .A(n6564), .ZN(n4513) );
  OAI21_X1 U5496 ( .B1(n4575), .B2(n6797), .A(n4574), .ZN(n10046) );
  AOI21_X1 U5497 ( .B1(n10043), .B2(n4576), .A(n4378), .ZN(n4574) );
  OAI21_X1 U5498 ( .B1(n7140), .B2(n7142), .A(n4565), .ZN(n7497) );
  OR2_X1 U5499 ( .A1(n7632), .A2(n7493), .ZN(n7494) );
  NOR2_X1 U5500 ( .A1(n7492), .A2(n7519), .ZN(n7493) );
  OR2_X1 U5501 ( .A1(n6636), .A2(n6380), .ZN(n6591) );
  AND2_X1 U5502 ( .A1(n4503), .A2(n4374), .ZN(n7641) );
  NOR2_X1 U5503 ( .A1(n7641), .A2(n7642), .ZN(n7716) );
  AND2_X1 U5504 ( .A1(n4584), .A2(n4312), .ZN(n7648) );
  NOR2_X1 U5505 ( .A1(n7718), .A2(n7719), .ZN(n8485) );
  OR2_X1 U5506 ( .A1(n7704), .A2(n7709), .ZN(n4701) );
  AND2_X1 U5507 ( .A1(n4506), .A2(n4375), .ZN(n8517) );
  OR2_X1 U5508 ( .A1(n8510), .A2(n8534), .ZN(n4572) );
  NAND3_X1 U5509 ( .A1(n4572), .A2(P2_REG1_REG_15__SCAN_IN), .A3(n8528), .ZN(
        n4573) );
  AOI21_X1 U5510 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8561), .A(n8556), .ZN(
        n8576) );
  NAND2_X1 U5511 ( .A1(n4505), .A2(n8566), .ZN(n8571) );
  OR2_X1 U5512 ( .A1(n8567), .A2(n8568), .ZN(n4505) );
  NAND2_X1 U5513 ( .A1(n8571), .A2(n8570), .ZN(n8582) );
  INV_X1 U5514 ( .A(n8605), .ZN(n4387) );
  NAND2_X1 U5515 ( .A1(n4718), .A2(n8619), .ZN(n4717) );
  NAND2_X1 U5516 ( .A1(n4716), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5517 ( .A1(n10047), .A2(n8622), .ZN(n4531) );
  OAI21_X1 U5518 ( .B1(n8614), .B2(n8613), .A(n8612), .ZN(n4534) );
  INV_X1 U5519 ( .A(n5463), .ZN(n8332) );
  INV_X1 U5520 ( .A(n5431), .ZN(n5430) );
  OR2_X1 U5521 ( .A1(n5447), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5463) );
  OR2_X1 U5522 ( .A1(n5410), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U5523 ( .A1(n5372), .A2(n9001), .ZN(n5392) );
  OR2_X1 U5524 ( .A1(n5337), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5353) );
  OR2_X1 U5525 ( .A1(n5306), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5321) );
  NOR2_X1 U5526 ( .A1(n8763), .A2(n4808), .ZN(n4807) );
  INV_X1 U5527 ( .A(n8191), .ZN(n4808) );
  NAND2_X1 U5528 ( .A1(n8768), .A2(n8203), .ZN(n4809) );
  NAND2_X1 U5529 ( .A1(n4995), .A2(n4994), .ZN(n5287) );
  INV_X1 U5530 ( .A(n5270), .ZN(n4995) );
  NAND2_X1 U5531 ( .A1(n4993), .A2(n4992), .ZN(n5256) );
  OR2_X1 U5532 ( .A1(n5256), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5270) );
  AND4_X1 U5533 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n8392)
         );
  OR2_X1 U5534 ( .A1(n5223), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U5535 ( .A1(n4989), .A2(n4988), .ZN(n5209) );
  INV_X1 U5536 ( .A(n5195), .ZN(n4989) );
  OR2_X1 U5537 ( .A1(n5182), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5195) );
  AND2_X1 U5538 ( .A1(n5486), .A2(n8130), .ZN(n4821) );
  INV_X1 U5539 ( .A(n7536), .ZN(n8291) );
  NAND2_X1 U5540 ( .A1(n4987), .A2(n4986), .ZN(n5169) );
  INV_X1 U5541 ( .A(n5152), .ZN(n4987) );
  NAND2_X1 U5542 ( .A1(n4803), .A2(n4801), .ZN(n7192) );
  AOI21_X1 U5543 ( .B1(n4804), .B2(n5483), .A(n4802), .ZN(n4801) );
  OR2_X1 U5544 ( .A1(n5139), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5152) );
  OR2_X1 U5545 ( .A1(n5103), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U5546 ( .A1(n4985), .A2(n4984), .ZN(n5139) );
  INV_X1 U5547 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n4984) );
  INV_X1 U5548 ( .A(n5118), .ZN(n4985) );
  NAND2_X1 U5549 ( .A1(n5482), .A2(n8143), .ZN(n7036) );
  NAND2_X1 U5550 ( .A1(n4981), .A2(n4980), .ZN(n5080) );
  INV_X1 U5551 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4980) );
  OR2_X1 U5552 ( .A1(n7764), .A2(n5498), .ZN(n7198) );
  NAND2_X1 U5553 ( .A1(n6674), .A2(n8112), .ZN(n7064) );
  INV_X1 U5554 ( .A(n6403), .ZN(n6666) );
  OR2_X1 U5555 ( .A1(n8628), .A2(n8627), .ZN(n8833) );
  NAND2_X1 U5556 ( .A1(n8640), .A2(n8243), .ZN(n5492) );
  INV_X1 U5557 ( .A(n4440), .ZN(n4439) );
  AOI21_X1 U5558 ( .B1(n4442), .B2(n4440), .A(n4438), .ZN(n4437) );
  INV_X1 U5559 ( .A(n8235), .ZN(n4438) );
  AND2_X1 U5560 ( .A1(n4435), .A2(n8237), .ZN(n8655) );
  AND3_X1 U5561 ( .A1(n5325), .A2(n5324), .A3(n5323), .ZN(n8730) );
  NOR2_X1 U5562 ( .A1(n8727), .A2(n4605), .ZN(n4601) );
  OR2_X1 U5563 ( .A1(n8737), .A2(n8742), .ZN(n4602) );
  NOR2_X1 U5564 ( .A1(n4608), .A2(n4611), .ZN(n4607) );
  INV_X1 U5565 ( .A(n8292), .ZN(n4608) );
  NAND2_X1 U5566 ( .A1(n4606), .A2(n4611), .ZN(n7457) );
  NAND2_X1 U5567 ( .A1(n7368), .A2(n4609), .ZN(n4606) );
  AND2_X1 U5568 ( .A1(n6636), .A2(n6753), .ZN(n6403) );
  AND2_X1 U5569 ( .A1(n4974), .A2(n4977), .ZN(n4810) );
  NAND2_X1 U5570 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  AND2_X1 U5571 ( .A1(n4692), .A2(n5470), .ZN(n4691) );
  NOR2_X1 U5572 ( .A1(n4693), .A2(n5282), .ZN(n4692) );
  NAND2_X1 U5573 ( .A1(n4694), .A2(n9020), .ZN(n4693) );
  INV_X1 U5574 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4694) );
  OR2_X1 U5575 ( .A1(n5866), .A2(n9208), .ZN(n5872) );
  NAND2_X1 U5576 ( .A1(n5871), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5883) );
  INV_X1 U5577 ( .A(n5872), .ZN(n5871) );
  OR2_X1 U5578 ( .A1(n5858), .A2(n9117), .ZN(n5866) );
  AND2_X1 U5579 ( .A1(n6248), .A2(n6249), .ZN(n9111) );
  AOI21_X1 U5580 ( .B1(n4776), .B2(n9167), .A(n4775), .ZN(n4774) );
  INV_X1 U5581 ( .A(n6226), .ZN(n4775) );
  NAND2_X1 U5582 ( .A1(n9175), .A2(n9176), .ZN(n9174) );
  NAND2_X1 U5583 ( .A1(n9123), .A2(n9124), .ZN(n9195) );
  OR2_X1 U5584 ( .A1(n5717), .A2(n9064), .ZN(n5729) );
  AND2_X1 U5585 ( .A1(n5693), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5695) );
  AND3_X1 U5586 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5693) );
  AND2_X1 U5587 ( .A1(n6413), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6384) );
  AND2_X1 U5588 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NOR2_X1 U5589 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5565) );
  NOR2_X1 U5590 ( .A1(n7973), .A2(n4492), .ZN(n4491) );
  INV_X1 U5591 ( .A(n4493), .ZN(n4492) );
  NAND2_X1 U5592 ( .A1(n4620), .A2(n7954), .ZN(n5934) );
  AND2_X1 U5593 ( .A1(n9428), .A2(n9404), .ZN(n9387) );
  AND2_X1 U5594 ( .A1(n9766), .A2(n9270), .ZN(n6018) );
  AND2_X1 U5595 ( .A1(n9567), .A2(n9556), .ZN(n9551) );
  NAND2_X1 U5596 ( .A1(n9542), .A2(n5828), .ZN(n9546) );
  INV_X1 U5597 ( .A(n5809), .ZN(n5807) );
  NAND2_X1 U5598 ( .A1(n7441), .A2(n7440), .ZN(n7439) );
  NAND2_X1 U5599 ( .A1(n7353), .A2(n7488), .ZN(n7449) );
  NAND2_X1 U5600 ( .A1(n7396), .A2(n7817), .ZN(n7395) );
  NAND2_X1 U5601 ( .A1(n7403), .A2(n5737), .ZN(n7405) );
  NAND2_X1 U5602 ( .A1(n8003), .A2(n8002), .ZN(n5709) );
  AOI21_X1 U5603 ( .B1(n4852), .B2(n4853), .A(n4336), .ZN(n4849) );
  NAND2_X1 U5604 ( .A1(n4487), .A2(n4484), .ZN(n7227) );
  NOR2_X1 U5605 ( .A1(n4486), .A2(n4485), .ZN(n4484) );
  NOR2_X1 U5606 ( .A1(n6873), .A2(n4379), .ZN(n7228) );
  NAND2_X1 U5607 ( .A1(n4625), .A2(n7852), .ZN(n7092) );
  OAI21_X1 U5608 ( .B1(n8001), .B2(n7845), .A(n4338), .ZN(n4625) );
  NAND2_X1 U5609 ( .A1(n4624), .A2(n7997), .ZN(n4623) );
  NAND2_X1 U5610 ( .A1(n4487), .A2(n4488), .ZN(n7090) );
  INV_X1 U5611 ( .A(n4486), .ZN(n4488) );
  INV_X1 U5612 ( .A(n9617), .ZN(n9966) );
  AND2_X1 U5613 ( .A1(n6504), .A2(n6414), .ZN(n9465) );
  OR2_X1 U5614 ( .A1(n9727), .A2(n7993), .ZN(n6324) );
  INV_X1 U5615 ( .A(n9348), .ZN(n7832) );
  AND2_X1 U5616 ( .A1(n7958), .A2(n7962), .ZN(n9407) );
  AND2_X1 U5617 ( .A1(n7776), .A2(n9462), .ZN(n9474) );
  NAND2_X1 U5618 ( .A1(n5845), .A2(n5844), .ZN(n9521) );
  OAI22_X1 U5619 ( .A1(n9559), .A2(n4823), .B1(n4825), .B2(n4822), .ZN(n9528)
         );
  NAND2_X1 U5620 ( .A1(n4828), .A2(n6014), .ZN(n4823) );
  INV_X1 U5621 ( .A(n4828), .ZN(n4822) );
  INV_X1 U5622 ( .A(n4826), .ZN(n4825) );
  AND2_X1 U5623 ( .A1(n7919), .A2(n7989), .ZN(n9529) );
  NAND2_X1 U5624 ( .A1(n5820), .A2(n5819), .ZN(n9703) );
  AOI21_X1 U5625 ( .B1(n9607), .B2(n6009), .A(n6008), .ZN(n9590) );
  NAND2_X1 U5626 ( .A1(n8013), .A2(n8010), .ZN(n7883) );
  NAND2_X1 U5627 ( .A1(n7842), .A2(n7997), .ZN(n6869) );
  AND2_X1 U5628 ( .A1(n6037), .A2(n6068), .ZN(n9724) );
  INV_X1 U5629 ( .A(n6085), .ZN(n5991) );
  XNOR2_X1 U5630 ( .A(n6352), .B(n6351), .ZN(n8326) );
  XNOR2_X1 U5631 ( .A(n6341), .B(SI_29_), .ZN(n8340) );
  XNOR2_X1 U5632 ( .A(n5443), .B(n5442), .ZN(n7700) );
  OR2_X1 U5633 ( .A1(n5586), .A2(n9791), .ZN(n5959) );
  NAND2_X1 U5634 ( .A1(n5936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U5635 ( .A1(n4459), .A2(n4464), .ZN(n5297) );
  NAND2_X1 U5636 ( .A1(n5265), .A2(n4467), .ZN(n4459) );
  XNOR2_X1 U5637 ( .A(n4562), .B(n4874), .ZN(n6418) );
  OAI21_X1 U5638 ( .B1(n5134), .B2(n5133), .A(n4913), .ZN(n4562) );
  XNOR2_X1 U5639 ( .A(n4897), .B(SI_4_), .ZN(n5086) );
  AND2_X1 U5640 ( .A1(n5131), .A2(n5130), .ZN(n10093) );
  NAND2_X1 U5641 ( .A1(n4685), .A2(n4682), .ZN(n8345) );
  NAND2_X1 U5642 ( .A1(n8399), .A2(n4661), .ZN(n4655) );
  NAND2_X1 U5643 ( .A1(n4669), .A2(n4667), .ZN(n7544) );
  INV_X1 U5644 ( .A(n4670), .ZN(n4667) );
  NAND2_X1 U5645 ( .A1(n8056), .A2(n4868), .ZN(n8390) );
  OR2_X1 U5646 ( .A1(n6820), .A2(n6821), .ZN(n4678) );
  NAND2_X1 U5647 ( .A1(n8368), .A2(n8072), .ZN(n8427) );
  AND2_X1 U5648 ( .A1(n5286), .A2(n5285), .ZN(n8823) );
  NAND2_X1 U5649 ( .A1(n8399), .A2(n8436), .ZN(n8358) );
  INV_X1 U5650 ( .A(n7082), .ZN(n4672) );
  NAND2_X1 U5651 ( .A1(n4321), .A2(n4673), .ZN(n7081) );
  AND2_X1 U5652 ( .A1(n6656), .A2(n6655), .ZN(n8458) );
  OR2_X1 U5653 ( .A1(n4878), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U5654 ( .A1(n7692), .A2(n7691), .ZN(n8056) );
  INV_X1 U5655 ( .A(n8458), .ZN(n8439) );
  AND2_X1 U5656 ( .A1(n8306), .A2(n4757), .ZN(n4756) );
  NAND2_X1 U5657 ( .A1(n4752), .A2(n4304), .ZN(n4559) );
  AND2_X1 U5658 ( .A1(n4313), .A2(n4816), .ZN(n4815) );
  INV_X1 U5659 ( .A(n8643), .ZN(n8461) );
  INV_X1 U5660 ( .A(n7113), .ZN(n8473) );
  CLKBUF_X1 U5661 ( .A(n6625), .Z(n8477) );
  OR2_X1 U5662 ( .A1(n6591), .A2(P2_U3151), .ZN(n8588) );
  OAI22_X1 U5663 ( .A1(n6697), .A2(n6696), .B1(n6709), .B2(n6558), .ZN(n6718)
         );
  NOR2_X1 U5664 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  INV_X1 U5665 ( .A(n6624), .ZN(n4517) );
  INV_X1 U5666 ( .A(n6560), .ZN(n4518) );
  NAND2_X1 U5667 ( .A1(n4514), .A2(n4515), .ZN(n6563) );
  AND2_X1 U5668 ( .A1(n4514), .A2(n4311), .ZN(n6791) );
  OAI21_X1 U5669 ( .B1(n6736), .B2(n4570), .A(n4568), .ZN(n6795) );
  NAND2_X1 U5670 ( .A1(n4377), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10044) );
  AND2_X1 U5671 ( .A1(n4525), .A2(n4524), .ZN(n10052) );
  OR2_X1 U5672 ( .A1(n6925), .A2(n4526), .ZN(n4525) );
  XNOR2_X1 U5673 ( .A(n7139), .B(n7134), .ZN(n6936) );
  NAND2_X1 U5674 ( .A1(n6936), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7141) );
  AND2_X1 U5675 ( .A1(n4523), .A2(n4522), .ZN(n7132) );
  AND2_X1 U5676 ( .A1(n7148), .A2(n7147), .ZN(n7152) );
  NAND2_X1 U5677 ( .A1(n4312), .A2(n4585), .ZN(n7501) );
  INV_X1 U5678 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5679 ( .A(n4503), .ZN(n7640) );
  NAND2_X1 U5680 ( .A1(n4701), .A2(n8478), .ZN(n7705) );
  AND2_X1 U5681 ( .A1(n4702), .A2(n8478), .ZN(n8482) );
  NOR2_X1 U5682 ( .A1(n8482), .A2(n8481), .ZN(n8502) );
  INV_X1 U5683 ( .A(n8493), .ZN(n4578) );
  INV_X1 U5684 ( .A(n4700), .ZN(n8540) );
  AND2_X1 U5685 ( .A1(n8528), .A2(n4573), .ZN(n8531) );
  XNOR2_X1 U5686 ( .A(n8576), .B(n8596), .ZN(n8557) );
  NOR2_X1 U5687 ( .A1(n8557), .A2(n8824), .ZN(n8577) );
  XNOR2_X1 U5688 ( .A(n8310), .B(n8248), .ZN(n5510) );
  NAND2_X1 U5689 ( .A1(n6048), .A2(n6047), .ZN(n8633) );
  NOR2_X1 U5690 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  NAND2_X1 U5691 ( .A1(n6044), .A2(n8769), .ZN(n6048) );
  OAI21_X1 U5692 ( .B1(n8648), .B2(n8738), .A(n8647), .ZN(n8794) );
  NOR2_X1 U5693 ( .A1(n8644), .A2(n8773), .ZN(n8645) );
  AOI21_X1 U5694 ( .B1(n5879), .B2(n8252), .A(n5371), .ZN(n8683) );
  NAND2_X1 U5695 ( .A1(n4809), .A2(n4807), .ZN(n8761) );
  INV_X1 U5696 ( .A(n8823), .ZN(n8760) );
  NAND2_X1 U5697 ( .A1(n5255), .A2(n5254), .ZN(n8829) );
  NAND2_X1 U5698 ( .A1(n7369), .A2(n5188), .ZN(n7433) );
  NAND2_X1 U5699 ( .A1(n5194), .A2(n5193), .ZN(n8169) );
  NAND2_X1 U5700 ( .A1(n7191), .A2(n8130), .ZN(n7340) );
  NAND2_X1 U5701 ( .A1(n4418), .A2(n5137), .ZN(n7244) );
  NAND2_X1 U5702 ( .A1(n6408), .A2(n8252), .ZN(n4418) );
  INV_X1 U5703 ( .A(n8698), .ZN(n8785) );
  AND2_X1 U5704 ( .A1(n8108), .A2(n8107), .ZN(n6675) );
  OR2_X1 U5705 ( .A1(n6667), .A2(n6666), .ZN(n8756) );
  XNOR2_X1 U5706 ( .A(n6050), .B(n6042), .ZN(n8639) );
  NOR2_X1 U5707 ( .A1(n8794), .A2(n8793), .ZN(n8839) );
  AND2_X1 U5708 ( .A1(n8792), .A2(n10118), .ZN(n8793) );
  NAND2_X1 U5709 ( .A1(n5409), .A2(n5408), .ZN(n8845) );
  NAND2_X1 U5710 ( .A1(n7680), .A2(n8252), .ZN(n5409) );
  XOR2_X1 U5711 ( .A(n8653), .B(n8655), .Z(n8848) );
  OAI21_X1 U5712 ( .B1(n8675), .B2(n4439), .A(n4437), .ZN(n8653) );
  NAND2_X1 U5713 ( .A1(n5389), .A2(n5388), .ZN(n8851) );
  NAND2_X1 U5714 ( .A1(n7629), .A2(n8252), .ZN(n5389) );
  NAND2_X1 U5715 ( .A1(n4616), .A2(n4297), .ZN(n8662) );
  INV_X1 U5716 ( .A(n8683), .ZN(n8856) );
  CLKBUF_X1 U5717 ( .A(n8677), .Z(n8678) );
  NAND2_X1 U5718 ( .A1(n4819), .A2(n8222), .ZN(n8688) );
  NAND2_X1 U5719 ( .A1(n5336), .A2(n5335), .ZN(n8867) );
  NAND2_X1 U5720 ( .A1(n5318), .A2(n5317), .ZN(n8873) );
  NAND2_X1 U5721 ( .A1(n4590), .A2(n4597), .ZN(n8717) );
  OR2_X1 U5722 ( .A1(n8737), .A2(n4599), .ZN(n4590) );
  NAND2_X1 U5723 ( .A1(n8741), .A2(n4818), .ZN(n8714) );
  INV_X1 U5724 ( .A(n8734), .ZN(n8879) );
  NAND2_X1 U5725 ( .A1(n8741), .A2(n8211), .ZN(n8725) );
  NAND2_X1 U5726 ( .A1(n5269), .A2(n5268), .ZN(n8891) );
  AND2_X1 U5727 ( .A1(n8779), .A2(n8778), .ZN(n8888) );
  NAND2_X1 U5728 ( .A1(n5239), .A2(n5238), .ZN(n7690) );
  NAND2_X1 U5729 ( .A1(n5490), .A2(n4425), .ZN(n4420) );
  NAND2_X1 U5730 ( .A1(n5222), .A2(n5221), .ZN(n7677) );
  INV_X1 U5731 ( .A(n8878), .ZN(n8890) );
  NAND2_X1 U5732 ( .A1(n5490), .A2(n5489), .ZN(n7614) );
  NAND2_X1 U5733 ( .A1(n5003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5005) );
  INV_X1 U5734 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8991) );
  INV_X1 U5735 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6420) );
  INV_X1 U5736 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U5737 ( .A1(n5049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U5738 ( .A1(n5048), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U5739 ( .A1(n5021), .A2(n5020), .ZN(n6695) );
  AND2_X1 U5740 ( .A1(n4784), .A2(n4785), .ZN(n8927) );
  AOI21_X1 U5741 ( .B1(n9116), .B2(n4788), .A(n4354), .ZN(n4784) );
  AND2_X1 U5742 ( .A1(n6163), .A2(n6165), .ZN(n9843) );
  NOR2_X1 U5743 ( .A1(n6333), .A2(n9262), .ZN(n6320) );
  NAND2_X1 U5744 ( .A1(n5742), .A2(n5741), .ZN(n9130) );
  NAND2_X1 U5745 ( .A1(n9174), .A2(n6283), .ZN(n9133) );
  NAND2_X1 U5746 ( .A1(n9165), .A2(n9167), .ZN(n9166) );
  NAND2_X1 U5747 ( .A1(n9144), .A2(n6211), .ZN(n4778) );
  NAND2_X1 U5748 ( .A1(n6109), .A2(n6108), .ZN(n6845) );
  INV_X1 U5749 ( .A(n4785), .ZN(n9205) );
  NAND2_X1 U5750 ( .A1(n9116), .A2(n6265), .ZN(n4786) );
  NAND2_X1 U5751 ( .A1(n5727), .A2(n5726), .ZN(n9224) );
  NAND2_X1 U5752 ( .A1(n4762), .A2(n4766), .ZN(n9243) );
  OR2_X1 U5753 ( .A1(n9175), .A2(n4767), .ZN(n4762) );
  AND2_X1 U5754 ( .A1(n6329), .A2(n8052), .ZN(n9856) );
  INV_X1 U5755 ( .A(n8040), .ZN(n8041) );
  AOI21_X1 U5756 ( .B1(n7838), .B2(n6035), .A(n7837), .ZN(n8045) );
  INV_X1 U5757 ( .A(n6034), .ZN(n8049) );
  NAND2_X1 U5758 ( .A1(n5924), .A2(n5923), .ZN(n9408) );
  NAND4_X1 U5759 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n9285)
         );
  NAND4_X1 U5760 ( .A1(n5583), .A2(n5582), .A3(n5581), .A4(n5580), .ZN(n9286)
         );
  NAND2_X1 U5761 ( .A1(n5658), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5610) );
  NAND4_X1 U5762 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n9288)
         );
  NAND2_X1 U5763 ( .A1(n5892), .A2(n5891), .ZN(n9671) );
  NAND2_X1 U5764 ( .A1(n7629), .A2(n6345), .ZN(n5892) );
  NAND2_X1 U5765 ( .A1(n9436), .A2(n7777), .ZN(n9422) );
  XNOR2_X1 U5766 ( .A(n9419), .B(n5901), .ZN(n9673) );
  INV_X1 U5767 ( .A(n9680), .ZN(n9460) );
  NAND2_X1 U5768 ( .A1(n4840), .A2(n4843), .ZN(n9453) );
  NAND2_X1 U5769 ( .A1(n5804), .A2(n8019), .ZN(n9561) );
  NAND2_X1 U5770 ( .A1(n9608), .A2(n4643), .ZN(n9591) );
  AND2_X1 U5771 ( .A1(n9608), .A2(n8014), .ZN(n9593) );
  NAND2_X1 U5772 ( .A1(n7219), .A2(n4855), .ZN(n4851) );
  INV_X1 U5773 ( .A(n7336), .ZN(n7257) );
  AND2_X1 U5774 ( .A1(n4856), .A2(n4855), .ZN(n7202) );
  OR2_X1 U5775 ( .A1(n7219), .A2(n4864), .ZN(n4856) );
  NAND2_X1 U5776 ( .A1(n7047), .A2(n7808), .ZN(n7046) );
  NAND2_X1 U5777 ( .A1(n7087), .A2(n5998), .ZN(n7047) );
  INV_X1 U5778 ( .A(n9637), .ZN(n9970) );
  NAND2_X1 U5779 ( .A1(n5926), .A2(n5925), .ZN(n9655) );
  NAND2_X1 U5780 ( .A1(n5716), .A2(n5715), .ZN(n7379) );
  NOR3_X1 U5781 ( .A1(n9652), .A2(n9651), .A3(n9650), .ZN(n9653) );
  NAND2_X1 U5782 ( .A1(n9385), .A2(n9384), .ZN(n9386) );
  NAND2_X1 U5783 ( .A1(n5903), .A2(n5902), .ZN(n9741) );
  XOR2_X1 U5784 ( .A(n9407), .B(n9382), .Z(n9743) );
  NAND2_X1 U5785 ( .A1(n9471), .A2(n4839), .ZN(n4833) );
  NAND2_X1 U5786 ( .A1(n5865), .A2(n5864), .ZN(n9752) );
  NAND2_X1 U5787 ( .A1(n5855), .A2(n5854), .ZN(n9757) );
  NAND2_X1 U5788 ( .A1(n4824), .A2(n6014), .ZN(n9541) );
  NAND2_X1 U5789 ( .A1(n9559), .A2(n4866), .ZN(n4824) );
  NAND2_X1 U5790 ( .A1(n5755), .A2(n5754), .ZN(n9202) );
  INV_X1 U5791 ( .A(n6874), .ZN(n6965) );
  AND2_X1 U5792 ( .A1(n10030), .A2(n9724), .ZN(n9785) );
  INV_X1 U5793 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5794 ( .A1(n5589), .A2(n5588), .ZN(n5594) );
  NOR2_X1 U5795 ( .A1(n5573), .A2(n9791), .ZN(n5588) );
  INV_X1 U5796 ( .A(n4859), .ZN(n4858) );
  OR2_X1 U5797 ( .A1(n5954), .A2(n9791), .ZN(n4857) );
  NAND2_X1 U5798 ( .A1(n4738), .A2(n4742), .ZN(n5364) );
  NAND2_X1 U5799 ( .A1(n5330), .A2(n4744), .ZN(n4738) );
  INV_X1 U5800 ( .A(n7993), .ZN(n7803) );
  INV_X1 U5801 ( .A(n5962), .ZN(n7837) );
  INV_X1 U5802 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U5803 ( .A1(n4736), .A2(n4902), .ZN(n5111) );
  NAND2_X1 U5804 ( .A1(n5075), .A2(n5074), .ZN(n4736) );
  INV_X1 U5805 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9027) );
  INV_X1 U5806 ( .A(n4712), .ZN(n7635) );
  OR2_X1 U5807 ( .A1(n8603), .A2(n4384), .ZN(P2_U3200) );
  OAI21_X1 U5808 ( .B1(n8606), .B2(n8624), .A(n4385), .ZN(n4384) );
  XNOR2_X1 U5809 ( .A(n8601), .B(n4719), .ZN(n8602) );
  INV_X1 U5810 ( .A(n4528), .ZN(n8623) );
  NOR2_X1 U5811 ( .A1(n5558), .A2(n4872), .ZN(n5559) );
  OAI21_X1 U5812 ( .B1(n6377), .B2(n10121), .A(n4863), .ZN(n6379) );
  AOI21_X1 U5813 ( .B1(n9371), .B2(n9984), .A(n9370), .ZN(n9372) );
  INV_X1 U5814 ( .A(n9369), .ZN(n9370) );
  OR2_X1 U5815 ( .A1(n9340), .A2(n9715), .ZN(n6371) );
  MUX2_X1 U5816 ( .A(n6370), .B(n6373), .S(n10042), .Z(n6372) );
  OR2_X1 U5817 ( .A1(n9340), .A2(n9781), .ZN(n6375) );
  MUX2_X1 U5818 ( .A(n6374), .B(n6373), .S(n10030), .Z(n6376) );
  INV_X1 U5819 ( .A(n5989), .ZN(n6041) );
  AND2_X1 U5820 ( .A1(n8670), .A2(n4320), .ZN(n4297) );
  OR2_X1 U5821 ( .A1(n8463), .A2(n4690), .ZN(n4298) );
  INV_X2 U5822 ( .A(n5731), .ZN(n5696) );
  AND2_X1 U5823 ( .A1(n8327), .A2(n5577), .ZN(n5635) );
  AND2_X1 U5824 ( .A1(n7832), .A2(n4621), .ZN(n4299) );
  INV_X1 U5825 ( .A(n7210), .ZN(n4855) );
  AND2_X1 U5826 ( .A1(n8683), .A2(n8693), .ZN(n4300) );
  NAND3_X1 U5827 ( .A1(n4645), .A2(n4644), .A3(n4489), .ZN(n4301) );
  AND2_X1 U5828 ( .A1(n4480), .A2(n4479), .ZN(n4302) );
  AND2_X1 U5829 ( .A1(n4725), .A2(n5161), .ZN(n4303) );
  NAND2_X1 U5830 ( .A1(n8270), .A2(n8261), .ZN(n8247) );
  NAND2_X1 U5831 ( .A1(n4602), .A2(n4604), .ZN(n8726) );
  NAND2_X1 U5832 ( .A1(n5437), .A2(n5436), .ZN(n8656) );
  INV_X1 U5833 ( .A(n8656), .ZN(n8454) );
  NAND2_X1 U5834 ( .A1(n4814), .A2(n4815), .ZN(n5478) );
  INV_X1 U5835 ( .A(n4975), .ZN(n5516) );
  INV_X1 U5836 ( .A(n9784), .ZN(n9601) );
  NAND2_X1 U5837 ( .A1(n5785), .A2(n5784), .ZN(n9784) );
  NAND2_X1 U5838 ( .A1(n8316), .A2(n5511), .ZN(n4304) );
  AND2_X1 U5839 ( .A1(n4439), .A2(n4435), .ZN(n4305) );
  AOI21_X1 U5840 ( .B1(n8675), .B2(n8231), .A(n8271), .ZN(n4436) );
  AND2_X1 U5841 ( .A1(n4647), .A2(n4646), .ZN(n4306) );
  AND2_X1 U5842 ( .A1(n8217), .A2(n8211), .ZN(n4818) );
  AND4_X1 U5843 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n8774)
         );
  NAND2_X1 U5844 ( .A1(n4645), .A2(n5568), .ZN(n5779) );
  AND2_X1 U5845 ( .A1(n9551), .A2(n4483), .ZN(n4307) );
  NAND2_X1 U5846 ( .A1(n5668), .A2(n5667), .ZN(n9959) );
  INV_X1 U5847 ( .A(n9959), .ZN(n4456) );
  AND2_X1 U5848 ( .A1(n4581), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4308) );
  INV_X1 U5849 ( .A(n6650), .ZN(n7534) );
  NAND2_X1 U5850 ( .A1(n7584), .A2(n8467), .ZN(n4309) );
  NAND2_X1 U5851 ( .A1(n9116), .A2(n4790), .ZN(n4785) );
  OR2_X1 U5852 ( .A1(n4696), .A2(n4965), .ZN(n4310) );
  OAI211_X1 U5853 ( .C1(n6416), .C2(n6469), .A(n5705), .B(n5704), .ZN(n9634)
         );
  NAND2_X1 U5854 ( .A1(n4633), .A2(n7989), .ZN(n7781) );
  AND2_X1 U5855 ( .A1(n4513), .A2(n4515), .ZN(n4311) );
  NAND2_X1 U5856 ( .A1(n7500), .A2(n7519), .ZN(n4312) );
  AND4_X1 U5857 ( .A1(n4971), .A2(n4970), .A3(n4969), .A4(n5281), .ZN(n4313)
         );
  AND2_X1 U5858 ( .A1(n4655), .A2(n4660), .ZN(n4314) );
  NAND2_X1 U5859 ( .A1(n5954), .A2(n5571), .ZN(n4315) );
  INV_X1 U5860 ( .A(n8308), .ZN(n4799) );
  NAND2_X1 U5861 ( .A1(n7967), .A2(n7984), .ZN(n4316) );
  AND2_X1 U5862 ( .A1(n5049), .A2(n4703), .ZN(n4317) );
  INV_X1 U5863 ( .A(n8080), .ZN(n8680) );
  NAND2_X1 U5864 ( .A1(n7251), .A2(n6147), .ZN(n4318) );
  AND2_X1 U5865 ( .A1(n8327), .A2(n5579), .ZN(n5658) );
  AND2_X1 U5866 ( .A1(n6798), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4319) );
  AOI21_X1 U5867 ( .B1(n8378), .B2(n8086), .A(n4870), .ZN(n8447) );
  XNOR2_X1 U5868 ( .A(n5134), .B(n5133), .ZN(n6408) );
  NAND2_X1 U5869 ( .A1(n8856), .A2(n8665), .ZN(n4320) );
  NAND2_X1 U5870 ( .A1(n6029), .A2(n6028), .ZN(n9382) );
  NAND2_X1 U5871 ( .A1(n4833), .A2(n4836), .ZN(n9435) );
  AND2_X1 U5872 ( .A1(n4675), .A2(n4674), .ZN(n4321) );
  AND2_X1 U5873 ( .A1(n9475), .A2(n5870), .ZN(n4322) );
  NAND2_X1 U5874 ( .A1(n7952), .A2(n7954), .ZN(n7830) );
  INV_X1 U5875 ( .A(n9280), .ZN(n9957) );
  INV_X1 U5876 ( .A(n8180), .ZN(n4539) );
  OR2_X1 U5877 ( .A1(n10106), .A2(n8470), .ZN(n4323) );
  OR2_X1 U5878 ( .A1(n7690), .A2(n8392), .ZN(n8187) );
  OR2_X1 U5879 ( .A1(n8215), .A2(n8264), .ZN(n4324) );
  AND2_X1 U5880 ( .A1(n4786), .A2(n6267), .ZN(n4325) );
  OAI21_X1 U5881 ( .B1(n9471), .B2(n4835), .A(n4834), .ZN(n9417) );
  INV_X1 U5882 ( .A(n9611), .ZN(n5777) );
  NOR2_X1 U5883 ( .A1(n8581), .A2(n8580), .ZN(n4326) );
  AND2_X1 U5884 ( .A1(n8211), .A2(n8212), .ZN(n8742) );
  INV_X1 U5885 ( .A(n8742), .ZN(n4600) );
  AND2_X1 U5886 ( .A1(n4840), .A2(n4839), .ZN(n4327) );
  NOR2_X1 U5887 ( .A1(n8475), .A2(n7062), .ZN(n4328) );
  NAND2_X1 U5888 ( .A1(n4413), .A2(n5770), .ZN(n9723) );
  AND2_X1 U5889 ( .A1(n8845), .A2(n8644), .ZN(n8238) );
  INV_X1 U5890 ( .A(n8238), .ZN(n4435) );
  NAND2_X1 U5891 ( .A1(n4778), .A2(n6216), .ZN(n9165) );
  AND2_X1 U5892 ( .A1(n4466), .A2(n4463), .ZN(n4329) );
  NOR2_X1 U5893 ( .A1(n8315), .A2(n8314), .ZN(n4330) );
  INV_X1 U5894 ( .A(n7973), .ZN(n9732) );
  NAND2_X1 U5895 ( .A1(n6347), .A2(n6346), .ZN(n7973) );
  INV_X1 U5896 ( .A(n9766), .ZN(n9535) );
  NAND2_X1 U5897 ( .A1(n5836), .A2(n5835), .ZN(n9766) );
  OR2_X1 U5898 ( .A1(n5360), .A2(n8707), .ZN(n4331) );
  INV_X1 U5899 ( .A(n8271), .ZN(n4441) );
  NAND2_X1 U5900 ( .A1(n8255), .A2(n8254), .ZN(n8311) );
  INV_X1 U5901 ( .A(n8311), .ZN(n8838) );
  NAND2_X1 U5902 ( .A1(n5806), .A2(n5805), .ZN(n9775) );
  NAND2_X1 U5903 ( .A1(n8437), .A2(n8360), .ZN(n4332) );
  AND2_X1 U5904 ( .A1(n7107), .A2(n8473), .ZN(n4333) );
  XNOR2_X1 U5905 ( .A(n4918), .B(SI_10_), .ZN(n5161) );
  INV_X1 U5906 ( .A(n4605), .ZN(n4604) );
  AND2_X1 U5907 ( .A1(n4820), .A2(n8222), .ZN(n4334) );
  NAND2_X1 U5908 ( .A1(n9655), .A2(n5933), .ZN(n9351) );
  AND2_X1 U5909 ( .A1(n4602), .A2(n4601), .ZN(n4335) );
  INV_X1 U5910 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4961) );
  INV_X1 U5911 ( .A(n9736), .ZN(n9391) );
  NAND2_X1 U5912 ( .A1(n5915), .A2(n5914), .ZN(n9736) );
  NOR2_X1 U5913 ( .A1(n9959), .A2(n9279), .ZN(n4336) );
  INV_X1 U5914 ( .A(n5201), .ZN(n4613) );
  INV_X1 U5915 ( .A(n4844), .ZN(n4843) );
  NOR2_X1 U5916 ( .A1(n9118), .A2(n9485), .ZN(n4844) );
  AND2_X1 U5917 ( .A1(n7163), .A2(n5999), .ZN(n4337) );
  AND2_X1 U5918 ( .A1(n4623), .A2(n7855), .ZN(n4338) );
  AND2_X1 U5919 ( .A1(n4903), .A2(SI_6_), .ZN(n4339) );
  OR2_X1 U5920 ( .A1(n5934), .A2(n7832), .ZN(n4340) );
  AND2_X1 U5921 ( .A1(n4919), .A2(SI_10_), .ZN(n4341) );
  AND2_X1 U5922 ( .A1(n5399), .A2(n8080), .ZN(n4342) );
  AND2_X1 U5923 ( .A1(n8475), .A2(n7062), .ZN(n4343) );
  OR2_X1 U5924 ( .A1(n8337), .A2(n8097), .ZN(n8270) );
  NAND2_X1 U5925 ( .A1(n4612), .A2(n5202), .ZN(n4344) );
  NAND2_X1 U5926 ( .A1(n9134), .A2(n4768), .ZN(n4345) );
  AND2_X1 U5927 ( .A1(n8198), .A2(n8195), .ZN(n8275) );
  OR2_X1 U5928 ( .A1(n8845), .A2(n8644), .ZN(n8237) );
  INV_X1 U5929 ( .A(n8237), .ZN(n4433) );
  AND2_X1 U5930 ( .A1(n8292), .A2(n4609), .ZN(n4346) );
  AND2_X1 U5931 ( .A1(n4451), .A2(n4818), .ZN(n4347) );
  AND2_X1 U5932 ( .A1(n4974), .A2(n4811), .ZN(n4348) );
  AND2_X1 U5933 ( .A1(n4865), .A2(n6028), .ZN(n4349) );
  INV_X1 U5934 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4390) );
  AND2_X1 U5935 ( .A1(n8215), .A2(n4817), .ZN(n4350) );
  AND2_X1 U5936 ( .A1(n4934), .A2(n4930), .ZN(n4351) );
  AND2_X1 U5937 ( .A1(n5901), .A2(n7777), .ZN(n4352) );
  NAND2_X1 U5938 ( .A1(n8510), .A2(n8534), .ZN(n8528) );
  AND2_X1 U5939 ( .A1(n5262), .A2(n5246), .ZN(n4353) );
  INV_X1 U5940 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4489) );
  OR2_X1 U5941 ( .A1(n8734), .A2(n8740), .ZN(n8217) );
  INV_X1 U5942 ( .A(n4631), .ZN(n4630) );
  OR2_X1 U5943 ( .A1(n5853), .A2(n4632), .ZN(n4631) );
  INV_X1 U5944 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4816) );
  INV_X1 U5945 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4569) );
  INV_X1 U5946 ( .A(n6585), .ZN(n4393) );
  INV_X1 U5947 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n4576) );
  AND2_X1 U5948 ( .A1(n9616), .A2(n9623), .ZN(n9597) );
  INV_X1 U5949 ( .A(n5635), .ZN(n5731) );
  AND2_X1 U5950 ( .A1(n4787), .A2(n9206), .ZN(n4354) );
  NOR2_X1 U5951 ( .A1(n5779), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U5952 ( .A1(n5881), .A2(n5880), .ZN(n9676) );
  OR3_X1 U5953 ( .A1(n6333), .A2(n9262), .A3(n4875), .ZN(n4355) );
  INV_X1 U5954 ( .A(n7989), .ZN(n4632) );
  NAND2_X1 U5955 ( .A1(n4420), .A2(n7613), .ZN(n7658) );
  INV_X1 U5956 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4708) );
  INV_X1 U5957 ( .A(n4868), .ZN(n4690) );
  AND2_X1 U5958 ( .A1(n8425), .A2(n8692), .ZN(n4356) );
  NAND2_X1 U5959 ( .A1(n9551), .A2(n9535), .ZN(n9520) );
  OR2_X1 U5960 ( .A1(n6378), .A2(n8878), .ZN(n4357) );
  AND2_X1 U5961 ( .A1(n4580), .A2(n8492), .ZN(n4358) );
  AND2_X1 U5962 ( .A1(n4572), .A2(n8528), .ZN(n4359) );
  INV_X1 U5963 ( .A(n6023), .ZN(n4841) );
  INV_X1 U5964 ( .A(n4839), .ZN(n4838) );
  NOR2_X1 U5965 ( .A1(n6024), .A2(n4844), .ZN(n4839) );
  NAND2_X1 U5966 ( .A1(n4809), .A2(n8191), .ZN(n8762) );
  INV_X1 U5967 ( .A(n4467), .ZN(n4466) );
  NOR2_X1 U5968 ( .A1(n4954), .A2(n4468), .ZN(n4467) );
  INV_X1 U5969 ( .A(n6014), .ZN(n4827) );
  INV_X1 U5970 ( .A(n8231), .ZN(n4442) );
  AND2_X1 U5971 ( .A1(n8272), .A2(n8674), .ZN(n8231) );
  NOR2_X1 U5972 ( .A1(n8388), .A2(n8463), .ZN(n4360) );
  AND2_X1 U5973 ( .A1(n4578), .A2(n8492), .ZN(n4361) );
  INV_X1 U5974 ( .A(n6283), .ZN(n4769) );
  OR2_X1 U5975 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  AND2_X1 U5976 ( .A1(n9676), .A2(n9466), .ZN(n4362) );
  OR2_X1 U5977 ( .A1(n5283), .A2(n5282), .ZN(n4363) );
  INV_X1 U5978 ( .A(n4789), .ZN(n4788) );
  NAND2_X1 U5979 ( .A1(n9206), .A2(n6265), .ZN(n4789) );
  AND2_X1 U5980 ( .A1(n6165), .A2(n9844), .ZN(n4364) );
  AOI21_X1 U5981 ( .B1(n4744), .B2(n5329), .A(n4743), .ZN(n4742) );
  NAND2_X1 U5982 ( .A1(n5428), .A2(n5427), .ZN(n8792) );
  INV_X1 U5983 ( .A(n8792), .ZN(n5438) );
  OR2_X1 U5984 ( .A1(n9508), .A2(n9477), .ZN(n4365) );
  NOR2_X1 U5985 ( .A1(n8485), .A2(n8486), .ZN(n4366) );
  NOR2_X1 U5986 ( .A1(n7142), .A2(n6931), .ZN(n4367) );
  AND2_X1 U5987 ( .A1(n4669), .A2(n4668), .ZN(n4368) );
  INV_X1 U5988 ( .A(n8249), .ZN(n8636) );
  AND2_X1 U5989 ( .A1(n5446), .A2(n5445), .ZN(n8249) );
  INV_X1 U5990 ( .A(n4683), .ZN(n4682) );
  OR2_X1 U5991 ( .A1(n8343), .A2(n4684), .ZN(n4683) );
  AND2_X1 U5992 ( .A1(n6062), .A2(n6061), .ZN(n10121) );
  NAND2_X1 U5993 ( .A1(n5796), .A2(n5795), .ZN(n9583) );
  INV_X1 U5994 ( .A(n9583), .ZN(n4479) );
  AND2_X1 U5995 ( .A1(n7352), .A2(n9850), .ZN(n7353) );
  NAND2_X1 U5996 ( .A1(n7036), .A2(n8287), .ZN(n7035) );
  NOR2_X1 U5997 ( .A1(n6873), .A2(n6874), .ZN(n4369) );
  INV_X1 U5998 ( .A(n8436), .ZN(n4662) );
  AND2_X1 U5999 ( .A1(n4851), .A2(n4854), .ZN(n4370) );
  INV_X1 U6000 ( .A(n8415), .ZN(n4657) );
  AOI21_X1 U6001 ( .B1(n5737), .B2(n7811), .A(n4639), .ZN(n4638) );
  NAND2_X1 U6002 ( .A1(n4796), .A2(n6149), .ZN(n7385) );
  NAND2_X1 U6003 ( .A1(n9157), .A2(n9156), .ZN(n9155) );
  NAND2_X1 U6004 ( .A1(n8484), .A2(n8505), .ZN(n4371) );
  AND2_X1 U6005 ( .A1(n4583), .A2(n4312), .ZN(n4372) );
  INV_X1 U6006 ( .A(n5951), .ZN(n9965) );
  NOR2_X1 U6007 ( .A1(n7227), .A2(n7336), .ZN(n5951) );
  AND2_X1 U6008 ( .A1(n4678), .A2(n4677), .ZN(n4373) );
  NAND2_X1 U6009 ( .A1(n7507), .A2(n7508), .ZN(n4374) );
  AND2_X1 U6010 ( .A1(n4507), .A2(n4371), .ZN(n4375) );
  AND2_X1 U6011 ( .A1(n7141), .A2(n7140), .ZN(n4376) );
  AND2_X1 U6012 ( .A1(n6797), .A2(n10043), .ZN(n4377) );
  INV_X1 U6013 ( .A(n8769), .ZN(n8738) );
  NAND2_X1 U6014 ( .A1(n8314), .A2(n6055), .ZN(n8769) );
  XOR2_X1 U6015 ( .A(n10048), .B(P2_REG1_REG_8__SCAN_IN), .Z(n4378) );
  NAND2_X1 U6016 ( .A1(n6034), .A2(n9330), .ZN(n7984) );
  OR2_X1 U6017 ( .A1(n4486), .A2(n9634), .ZN(n4379) );
  INV_X1 U6018 ( .A(n8600), .ZN(n4719) );
  XOR2_X1 U6019 ( .A(n6798), .B(n6588), .Z(n4380) );
  NAND2_X1 U6020 ( .A1(n4589), .A2(n5053), .ZN(n7057) );
  AND2_X1 U6021 ( .A1(n6573), .A2(n6574), .ZN(n4381) );
  INV_X1 U6022 ( .A(n6873), .ZN(n4487) );
  NAND2_X1 U6023 ( .A1(n7021), .A2(n5990), .ZN(n7020) );
  INV_X1 U6024 ( .A(n8619), .ZN(n4720) );
  OR2_X1 U6025 ( .A1(n4719), .A2(n4720), .ZN(n4382) );
  INV_X1 U6026 ( .A(n6720), .ZN(n4391) );
  XOR2_X1 U6027 ( .A(n6798), .B(n6901), .Z(n4383) );
  INV_X1 U6028 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6029 ( .A1(n7350), .A2(n6003), .ZN(n7396) );
  INV_X1 U6030 ( .A(n5074), .ZN(n4733) );
  NAND2_X1 U6031 ( .A1(n4850), .A2(n4849), .ZN(n7351) );
  AOI21_X1 U6032 ( .B1(n9528), .B2(n6019), .A(n6018), .ZN(n9514) );
  NAND2_X1 U6033 ( .A1(n9217), .A2(n9219), .ZN(n9123) );
  NAND2_X1 U6034 ( .A1(n6847), .A2(n6117), .ZN(n6124) );
  NAND2_X2 U6035 ( .A1(n8926), .A2(n8930), .ZN(n9175) );
  NAND2_X2 U6036 ( .A1(n6162), .A2(n6161), .ZN(n6165) );
  XNOR2_X2 U6037 ( .A(n6088), .B(n6298), .ZN(n6089) );
  OR2_X1 U6038 ( .A1(n7850), .A2(n7849), .ZN(n7874) );
  NAND2_X1 U6039 ( .A1(n5623), .A2(n5994), .ZN(n8001) );
  NAND2_X1 U6040 ( .A1(n4408), .A2(n7907), .ZN(n4407) );
  NAND2_X1 U6041 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  NAND2_X1 U6042 ( .A1(n4405), .A2(n4404), .ZN(n7917) );
  AOI211_X1 U6043 ( .C1(n7972), .C2(n7983), .A(n7971), .B(n7986), .ZN(n7978)
         );
  NAND2_X1 U6044 ( .A1(n7968), .A2(n7984), .ZN(n4415) );
  XNOR2_X1 U6045 ( .A(n8595), .B(n8596), .ZN(n8562) );
  NAND2_X1 U6046 ( .A1(n6702), .A2(n6703), .ZN(n6701) );
  INV_X1 U6047 ( .A(n6568), .ZN(n4392) );
  NAND2_X1 U6048 ( .A1(n4706), .A2(n4707), .ZN(n6800) );
  AOI21_X1 U6049 ( .B1(n8598), .B2(n4719), .A(n4721), .ZN(n4718) );
  NAND2_X1 U6050 ( .A1(n8150), .A2(n8149), .ZN(n8153) );
  NAND2_X1 U6051 ( .A1(n4554), .A2(n8219), .ZN(n4553) );
  NAND2_X1 U6052 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U6053 ( .A1(n8209), .A2(n8256), .ZN(n4558) );
  NAND2_X1 U6054 ( .A1(n8197), .A2(n4541), .ZN(n8188) );
  NAND2_X1 U6055 ( .A1(n4561), .A2(n5511), .ZN(n4560) );
  NAND2_X1 U6056 ( .A1(n4544), .A2(n8655), .ZN(n8241) );
  NAND2_X1 U6057 ( .A1(n4551), .A2(n4550), .ZN(n8227) );
  NAND2_X1 U6058 ( .A1(n4749), .A2(n8260), .ZN(n8269) );
  NAND2_X1 U6059 ( .A1(n8230), .A2(n8229), .ZN(n4549) );
  MUX2_X1 U6060 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8908), .S(n5506), .Z(n7760) );
  NAND2_X1 U6061 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  XNOR2_X2 U6062 ( .A(n5832), .B(n4390), .ZN(n6035) );
  NAND2_X1 U6063 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U6064 ( .A1(n6109), .A2(n4792), .ZN(n6847) );
  OAI21_X1 U6065 ( .B1(n4759), .B2(n6163), .A(n4758), .ZN(n9217) );
  NOR2_X1 U6066 ( .A1(n8506), .A2(n8513), .ZN(n8537) );
  AOI21_X1 U6067 ( .B1(n4396), .B2(n7962), .A(n7961), .ZN(n7965) );
  NAND2_X1 U6068 ( .A1(n7944), .A2(n7945), .ZN(n4397) );
  NAND2_X1 U6069 ( .A1(n5134), .A2(n4303), .ZN(n4402) );
  NAND2_X1 U6070 ( .A1(n4723), .A2(n4402), .ZN(n5178) );
  INV_X1 U6071 ( .A(n5177), .ZN(n4401) );
  NAND3_X1 U6072 ( .A1(n5063), .A2(n5062), .A3(n5086), .ZN(n4445) );
  MUX2_X1 U6073 ( .A(n6386), .B(n6390), .S(n6388), .Z(n4897) );
  OR2_X1 U6074 ( .A1(n5490), .A2(n4424), .ZN(n4419) );
  INV_X1 U6075 ( .A(n8675), .ZN(n4431) );
  OAI21_X1 U6076 ( .B1(n4431), .B2(n4434), .A(n4432), .ZN(n8640) );
  NAND2_X1 U6077 ( .A1(n5063), .A2(n5062), .ZN(n4447) );
  NAND2_X1 U6078 ( .A1(n4449), .A2(n4350), .ZN(n5491) );
  NAND2_X1 U6079 ( .A1(n4347), .A2(n4450), .ZN(n4449) );
  NAND2_X4 U6080 ( .A1(n4501), .A2(n4502), .ZN(n6388) );
  AND2_X1 U6081 ( .A1(n4455), .A2(n8131), .ZN(n4804) );
  NAND2_X1 U6082 ( .A1(n4477), .A2(n4322), .ZN(n7940) );
  NAND2_X1 U6083 ( .A1(n10014), .A2(n5999), .ZN(n4485) );
  AND2_X1 U6084 ( .A1(n9387), .A2(n4493), .ZN(n9361) );
  NAND2_X1 U6085 ( .A1(n9387), .A2(n4491), .ZN(n9341) );
  NAND2_X1 U6086 ( .A1(n9387), .A2(n4495), .ZN(n9362) );
  NAND2_X1 U6087 ( .A1(n9387), .A2(n9391), .ZN(n9388) );
  NAND3_X1 U6088 ( .A1(n4496), .A2(n4879), .A3(n4908), .ZN(n4500) );
  NAND3_X1 U6089 ( .A1(n4501), .A2(n4502), .A3(n6409), .ZN(n4499) );
  NAND2_X1 U6090 ( .A1(n4506), .A2(n4507), .ZN(n8516) );
  OR2_X1 U6091 ( .A1(n6562), .A2(n4393), .ZN(n4515) );
  NOR2_X1 U6092 ( .A1(n6603), .A2(n4516), .ZN(n6734) );
  NAND2_X1 U6093 ( .A1(n6925), .A2(n4524), .ZN(n4520) );
  NAND2_X1 U6094 ( .A1(n4520), .A2(n4521), .ZN(n4523) );
  INV_X1 U6095 ( .A(n4525), .ZN(n10054) );
  INV_X1 U6096 ( .A(n4523), .ZN(n6934) );
  INV_X1 U6097 ( .A(n6933), .ZN(n4522) );
  INV_X1 U6098 ( .A(n6926), .ZN(n4527) );
  NAND3_X1 U6099 ( .A1(n8616), .A2(n8617), .A3(n4531), .ZN(n4530) );
  INV_X1 U6100 ( .A(n8182), .ZN(n4536) );
  NAND2_X1 U6101 ( .A1(n8181), .A2(n4540), .ZN(n4535) );
  OAI21_X1 U6102 ( .B1(n4536), .B2(n4535), .A(n4537), .ZN(n8197) );
  NAND3_X1 U6103 ( .A1(n8130), .A2(n8126), .A3(n8264), .ZN(n4542) );
  NAND3_X1 U6104 ( .A1(n4558), .A2(n4557), .A3(n4556), .ZN(n4555) );
  MUX2_X1 U6105 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6388), .Z(n4903) );
  NOR2_X4 U6106 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5047) );
  NAND2_X1 U6107 ( .A1(n6936), .A2(n4367), .ZN(n4565) );
  NAND2_X1 U6108 ( .A1(n6736), .A2(n4568), .ZN(n4567) );
  INV_X1 U6109 ( .A(n4573), .ZN(n8529) );
  INV_X1 U6110 ( .A(n10043), .ZN(n4575) );
  NAND2_X1 U6111 ( .A1(n8494), .A2(n4581), .ZN(n4577) );
  NAND2_X1 U6112 ( .A1(n4579), .A2(n4577), .ZN(n8509) );
  NAND3_X1 U6113 ( .A1(n4580), .A2(n8492), .A3(n4308), .ZN(n4579) );
  INV_X1 U6114 ( .A(n7500), .ZN(n4586) );
  NAND2_X1 U6115 ( .A1(n8737), .A2(n4595), .ZN(n4594) );
  NOR2_X1 U6116 ( .A1(n8367), .A2(n8729), .ZN(n4605) );
  AOI21_X1 U6117 ( .B1(n7368), .B2(n4346), .A(n4607), .ZN(n7456) );
  NAND2_X1 U6118 ( .A1(n8677), .A2(n4297), .ZN(n4614) );
  NAND2_X1 U6119 ( .A1(n7606), .A2(n5263), .ZN(n8772) );
  NAND2_X1 U6120 ( .A1(n5247), .A2(n4353), .ZN(n7606) );
  NAND2_X1 U6121 ( .A1(n5247), .A2(n5246), .ZN(n7604) );
  OAI21_X2 U6122 ( .B1(n7101), .B2(n5145), .A(n5146), .ZN(n7194) );
  OAI21_X1 U6123 ( .B1(n9393), .B2(n4622), .A(n4299), .ZN(n9352) );
  NAND2_X1 U6124 ( .A1(n4619), .A2(n4618), .ZN(n9355) );
  NAND2_X1 U6125 ( .A1(n9393), .A2(n4299), .ZN(n4619) );
  NAND2_X1 U6126 ( .A1(n9393), .A2(n9392), .ZN(n4620) );
  NAND2_X1 U6127 ( .A1(n5804), .A2(n4626), .ZN(n9542) );
  OAI21_X1 U6128 ( .B1(n9530), .B2(n4631), .A(n4627), .ZN(n9496) );
  OAI21_X1 U6129 ( .B1(n7358), .B2(n4636), .A(n4635), .ZN(n7442) );
  INV_X1 U6130 ( .A(n4638), .ZN(n4636) );
  NAND2_X1 U6131 ( .A1(n4637), .A2(n4638), .ZN(n7443) );
  NAND2_X1 U6132 ( .A1(n7358), .A2(n5737), .ZN(n4637) );
  NAND2_X1 U6133 ( .A1(n9436), .A2(n4352), .ZN(n9420) );
  INV_X2 U6134 ( .A(n5768), .ZN(n4645) );
  NAND2_X1 U6135 ( .A1(n5954), .A2(n4647), .ZN(n5590) );
  NAND2_X1 U6136 ( .A1(n5954), .A2(n4306), .ZN(n4648) );
  NAND2_X1 U6137 ( .A1(n8770), .A2(n4869), .ZN(n8749) );
  NAND2_X1 U6138 ( .A1(n5160), .A2(n5159), .ZN(n7341) );
  AOI22_X1 U6139 ( .A1(n8654), .A2(n5418), .B1(n5417), .B2(n8644), .ZN(n8642)
         );
  NAND2_X1 U6140 ( .A1(n5102), .A2(n5101), .ZN(n6899) );
  NAND2_X1 U6141 ( .A1(n8703), .A2(n5344), .ZN(n8690) );
  NAND2_X1 U6142 ( .A1(n8772), .A2(n8771), .ZN(n8770) );
  NOR2_X1 U6143 ( .A1(n8545), .A2(n8544), .ZN(n8567) );
  NOR3_X1 U6144 ( .A1(n6717), .A2(n6605), .A3(n6604), .ZN(n6603) );
  NOR2_X1 U6145 ( .A1(n8585), .A2(n8584), .ZN(n8614) );
  NOR2_X1 U6146 ( .A1(n8517), .A2(n8518), .ZN(n8544) );
  INV_X4 U6147 ( .A(n6388), .ZN(n6357) );
  NAND2_X1 U6148 ( .A1(n7014), .A2(n5622), .ZN(n6837) );
  NAND2_X1 U6149 ( .A1(n7806), .A2(n7802), .ZN(n7014) );
  XNOR2_X1 U6150 ( .A(n9355), .B(n9354), .ZN(n9358) );
  NAND2_X1 U6151 ( .A1(n9473), .A2(n9474), .ZN(n9472) );
  OR2_X1 U6152 ( .A1(n8253), .A2(n6398), .ZN(n5024) );
  NAND2_X2 U6153 ( .A1(n6416), .A2(n6388), .ZN(n5605) );
  NAND3_X2 U6154 ( .A1(n5024), .A2(n5023), .A3(n5022), .ZN(n6648) );
  INV_X1 U6155 ( .A(n6648), .ZN(n10067) );
  NAND2_X1 U6156 ( .A1(n8399), .A2(n4656), .ZN(n4652) );
  NAND2_X1 U6157 ( .A1(n4652), .A2(n4653), .ZN(n8417) );
  INV_X1 U6158 ( .A(n7422), .ZN(n4663) );
  OAI21_X1 U6159 ( .B1(n4663), .B2(n4666), .A(n4664), .ZN(n7585) );
  NAND2_X1 U6160 ( .A1(n7422), .A2(n7421), .ZN(n7542) );
  NOR2_X1 U6161 ( .A1(n7540), .A2(n7420), .ZN(n4671) );
  INV_X1 U6162 ( .A(n4678), .ZN(n6887) );
  NAND2_X1 U6163 ( .A1(n6888), .A2(n6893), .ZN(n4677) );
  OAI21_X1 U6164 ( .B1(n8447), .B2(n4683), .A(n4679), .ZN(n8094) );
  NAND2_X1 U6165 ( .A1(n8447), .A2(n8448), .ZN(n4685) );
  NAND2_X1 U6166 ( .A1(n7692), .A2(n4687), .ZN(n4686) );
  AND2_X1 U6167 ( .A1(n5218), .A2(n4692), .ZN(n5471) );
  NAND2_X1 U6168 ( .A1(n5218), .A2(n4691), .ZN(n5472) );
  INV_X1 U6169 ( .A(n4965), .ZN(n4695) );
  NAND3_X1 U6170 ( .A1(n4695), .A2(n5047), .A3(n4697), .ZN(n5163) );
  NAND3_X1 U6171 ( .A1(n4697), .A2(n5047), .A3(n4816), .ZN(n4696) );
  NAND3_X1 U6172 ( .A1(n4701), .A2(n8478), .A3(P2_REG2_REG_13__SCAN_IN), .ZN(
        n4702) );
  INV_X1 U6173 ( .A(n4702), .ZN(n8479) );
  NAND2_X1 U6174 ( .A1(n7704), .A2(n7709), .ZN(n8478) );
  INV_X1 U6175 ( .A(n6573), .ZN(n4705) );
  NAND2_X1 U6176 ( .A1(n4705), .A2(n6574), .ZN(n4706) );
  OAI21_X1 U6177 ( .B1(n6946), .B2(n4710), .A(n4709), .ZN(n7490) );
  AOI21_X1 U6178 ( .B1(n7147), .B2(n6932), .A(n7151), .ZN(n4709) );
  OAI211_X1 U6179 ( .C1(n4717), .C2(n8597), .A(n4714), .B(n4713), .ZN(n8621)
         );
  NAND3_X1 U6180 ( .A1(n8597), .A2(n4719), .A3(n4720), .ZN(n4713) );
  NAND2_X1 U6181 ( .A1(n5075), .A2(n4730), .ZN(n4732) );
  NAND2_X1 U6182 ( .A1(n5315), .A2(n5314), .ZN(n5330) );
  NAND2_X1 U6183 ( .A1(n4737), .A2(n4739), .ZN(n5366) );
  NAND3_X1 U6184 ( .A1(n5315), .A2(n5314), .A3(n4742), .ZN(n4737) );
  NAND2_X1 U6185 ( .A1(n4746), .A2(n4351), .ZN(n5233) );
  NAND2_X1 U6186 ( .A1(n8248), .A2(n4748), .ZN(n8267) );
  NAND3_X1 U6187 ( .A1(n4748), .A2(n8248), .A3(n8249), .ZN(n4751) );
  INV_X1 U6188 ( .A(n8247), .ZN(n8248) );
  NAND3_X1 U6189 ( .A1(n4751), .A2(n8265), .A3(n4750), .ZN(n4749) );
  NAND2_X1 U6190 ( .A1(n4798), .A2(n4754), .ZN(n4753) );
  NAND2_X1 U6191 ( .A1(n8307), .A2(n8628), .ZN(n4757) );
  AND2_X2 U6192 ( .A1(n6069), .A2(n7030), .ZN(n6070) );
  OR2_X2 U6193 ( .A1(n9983), .A2(n7803), .ZN(n7030) );
  INV_X1 U6194 ( .A(n6165), .ZN(n4759) );
  AOI21_X2 U6195 ( .B1(n6165), .B2(n4761), .A(n4760), .ZN(n4758) );
  NAND2_X1 U6196 ( .A1(n9842), .A2(n6165), .ZN(n9218) );
  NAND2_X1 U6197 ( .A1(n4364), .A2(n6163), .ZN(n9842) );
  NAND2_X1 U6198 ( .A1(n9175), .A2(n4766), .ZN(n4765) );
  NAND2_X1 U6199 ( .A1(n6289), .A2(n6288), .ZN(n4770) );
  NAND2_X1 U6200 ( .A1(n9143), .A2(n4772), .ZN(n4771) );
  NAND2_X2 U6201 ( .A1(n4771), .A2(n4774), .ZN(n9094) );
  NAND2_X1 U6202 ( .A1(n9116), .A2(n4782), .ZN(n4781) );
  INV_X1 U6203 ( .A(n6108), .ZN(n4793) );
  NAND2_X1 U6204 ( .A1(n4796), .A2(n4794), .ZN(n7386) );
  NAND2_X1 U6205 ( .A1(n6141), .A2(n6140), .ZN(n7249) );
  OAI21_X2 U6206 ( .B1(n5779), .B2(n4847), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5817) );
  NAND2_X1 U6207 ( .A1(n5482), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U6208 ( .A1(n8112), .A2(n8113), .ZN(n8119) );
  NAND3_X1 U6209 ( .A1(n8112), .A2(n4806), .A3(n8108), .ZN(n6674) );
  NAND2_X1 U6210 ( .A1(n4975), .A2(n4348), .ZN(n5003) );
  NAND3_X1 U6211 ( .A1(n5007), .A2(n5006), .A3(P2_REG1_REG_2__SCAN_IN), .ZN(
        n5044) );
  XNOR2_X2 U6212 ( .A(n5002), .B(n8898), .ZN(n5007) );
  NAND2_X1 U6213 ( .A1(n8702), .A2(n8225), .ZN(n4819) );
  NAND2_X1 U6214 ( .A1(n7366), .A2(n8161), .ZN(n5487) );
  NAND2_X1 U6215 ( .A1(n7191), .A2(n4821), .ZN(n7366) );
  XNOR2_X2 U6216 ( .A(n6085), .B(n5992), .ZN(n5990) );
  NAND2_X2 U6217 ( .A1(n5608), .A2(n5607), .ZN(n6085) );
  NAND2_X1 U6218 ( .A1(n6029), .A2(n4349), .ZN(n9346) );
  NAND2_X1 U6219 ( .A1(n9346), .A2(n9345), .ZN(n9349) );
  NAND2_X1 U6220 ( .A1(n7219), .A2(n4852), .ZN(n4850) );
  AOI21_X2 U6221 ( .B1(n4855), .B2(n4864), .A(n6002), .ZN(n4854) );
  INV_X1 U6222 ( .A(n4856), .ZN(n7203) );
  NAND2_X1 U6223 ( .A1(n4857), .A2(n4858), .ZN(n5585) );
  NAND2_X1 U6224 ( .A1(n5158), .A2(n4323), .ZN(n5160) );
  XNOR2_X1 U6225 ( .A(n6043), .B(n6042), .ZN(n6044) );
  OAI21_X1 U6226 ( .B1(n9660), .B2(n9787), .A(n6038), .ZN(n6039) );
  INV_X1 U6227 ( .A(n5590), .ZN(n5592) );
  INV_X1 U6228 ( .A(n6319), .ZN(n8910) );
  NAND2_X1 U6229 ( .A1(n5586), .A2(n5587), .ZN(n5589) );
  XOR2_X1 U6230 ( .A(n8640), .B(n8641), .Z(n8842) );
  INV_X1 U6231 ( .A(n5510), .ZN(n5512) );
  INV_X1 U6232 ( .A(n5007), .ZN(n5008) );
  XNOR2_X1 U6233 ( .A(n5959), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5966) );
  AOI21_X2 U6234 ( .B1(n8749), .B2(n5295), .A(n5294), .ZN(n8737) );
  NAND2_X1 U6235 ( .A1(n8705), .A2(n8704), .ZN(n8703) );
  OR2_X1 U6236 ( .A1(n5038), .A2(n5026), .ZN(n4861) );
  AND3_X1 U6237 ( .A1(n5816), .A2(n5829), .A3(n4390), .ZN(n4862) );
  AND2_X1 U6238 ( .A1(n6774), .A2(n7416), .ZN(n10082) );
  OR2_X1 U6239 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(n10119), .ZN(n4863) );
  AND2_X1 U6240 ( .A1(n6001), .A2(n10014), .ZN(n4864) );
  NOR2_X1 U6241 ( .A1(n9383), .A2(n4876), .ZN(n4865) );
  OR2_X1 U6242 ( .A1(n9570), .A2(n6013), .ZN(n4866) );
  OR2_X1 U6243 ( .A1(n9601), .A2(n7901), .ZN(n4867) );
  OR2_X1 U6244 ( .A1(n8055), .A2(n8392), .ZN(n4868) );
  AND2_X1 U6245 ( .A1(n10133), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4872) );
  NAND2_X1 U6246 ( .A1(n7706), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4873) );
  INV_X1 U6247 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6396) );
  XNOR2_X1 U6248 ( .A(n5969), .B(n5968), .ZN(n6034) );
  AND2_X1 U6249 ( .A1(n4917), .A2(n4916), .ZN(n4874) );
  INV_X1 U6250 ( .A(n8156), .ZN(n5486) );
  OR2_X1 U6251 ( .A1(n6316), .A2(n6315), .ZN(n4875) );
  INV_X1 U6252 ( .A(n6814), .ZN(n5950) );
  INV_X1 U6253 ( .A(n8275), .ZN(n5262) );
  XNOR2_X1 U6254 ( .A(n5381), .B(n5380), .ZN(n5879) );
  INV_X1 U6255 ( .A(n8302), .ZN(n6042) );
  INV_X1 U6256 ( .A(n6538), .ZN(n5598) );
  INV_X1 U6257 ( .A(n5579), .ZN(n5577) );
  NOR2_X1 U6258 ( .A1(n6031), .A2(n7830), .ZN(n4876) );
  NOR2_X1 U6259 ( .A1(n6190), .A2(n9197), .ZN(n4877) );
  NOR2_X1 U6260 ( .A1(n8082), .A2(n8382), .ZN(n4878) );
  INV_X1 U6261 ( .A(n8861), .ZN(n5360) );
  MUX2_X1 U6262 ( .A(n8111), .B(n8110), .S(n8256), .Z(n8118) );
  AND2_X1 U6263 ( .A1(n8146), .A2(n8145), .ZN(n8147) );
  NOR2_X1 U6264 ( .A1(n8460), .A2(n8264), .ZN(n8258) );
  NOR2_X1 U6265 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  OR2_X1 U6266 ( .A1(n7532), .A2(n8469), .ZN(n5175) );
  INV_X1 U6267 ( .A(n6625), .ZN(n5025) );
  NOR2_X1 U6268 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  NAND2_X1 U6269 ( .A1(n8305), .A2(n5496), .ZN(n8306) );
  INV_X1 U6270 ( .A(n7490), .ZN(n7150) );
  INV_X1 U6271 ( .A(n5392), .ZN(n5391) );
  OR2_X1 U6272 ( .A1(n8867), .A2(n8718), .ZN(n5344) );
  NAND2_X1 U6273 ( .A1(n5117), .A2(n5116), .ZN(n7038) );
  OR2_X1 U6274 ( .A1(n8049), .A2(n6068), .ZN(n6069) );
  INV_X1 U6275 ( .A(n5788), .ZN(n5786) );
  INV_X1 U6276 ( .A(n9353), .ZN(n9354) );
  NAND2_X1 U6277 ( .A1(n6872), .A2(n6814), .ZN(n7997) );
  INV_X1 U6278 ( .A(n5216), .ZN(n4934) );
  OR2_X1 U6279 ( .A1(n5710), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5711) );
  INV_X1 U6280 ( .A(n5304), .ZN(n4997) );
  INV_X1 U6281 ( .A(n8472), .ZN(n7237) );
  XNOR2_X1 U6282 ( .A(n6940), .B(n6927), .ZN(n6938) );
  NAND2_X1 U6283 ( .A1(n5430), .A2(n5429), .ZN(n5447) );
  INV_X1 U6284 ( .A(n5321), .ZN(n5320) );
  INV_X1 U6285 ( .A(n8285), .ZN(n5484) );
  AND2_X1 U6286 ( .A1(n8136), .A2(n8121), .ZN(n8278) );
  OR2_X1 U6287 ( .A1(n6772), .A2(n6632), .ZN(n6639) );
  INV_X1 U6288 ( .A(n6118), .ZN(n6295) );
  OR2_X1 U6289 ( .A1(n5894), .A2(n5893), .ZN(n5906) );
  NAND2_X1 U6290 ( .A1(n5882), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6291 ( .A1(n5743), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5758) );
  INV_X1 U6292 ( .A(n9340), .ZN(n6359) );
  OR2_X1 U6293 ( .A1(n4876), .A2(n6033), .ZN(n9345) );
  NAND2_X1 U6294 ( .A1(n5834), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U6295 ( .A1(n4920), .A2(n9008), .ZN(n4923) );
  NAND2_X1 U6296 ( .A1(n4910), .A2(n4909), .ZN(n4913) );
  NAND2_X1 U6297 ( .A1(n6389), .A2(n9028), .ZN(n4893) );
  NAND2_X1 U6298 ( .A1(n4997), .A2(n4996), .ZN(n5306) );
  NAND2_X1 U6299 ( .A1(n7236), .A2(n7237), .ZN(n7238) );
  OR2_X1 U6300 ( .A1(n8071), .A2(n8706), .ZN(n8072) );
  OR2_X1 U6301 ( .A1(n6664), .A2(n6663), .ZN(n8429) );
  INV_X1 U6302 ( .A(n5039), .ZN(n5464) );
  OR2_X1 U6303 ( .A1(n5211), .A2(n6908), .ZN(n5083) );
  OR2_X1 U6304 ( .A1(P2_U3150), .A2(n6592), .ZN(n8594) );
  NOR2_X1 U6305 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  INV_X1 U6306 ( .A(n5483), .ZN(n8287) );
  NAND2_X1 U6307 ( .A1(n8792), .A2(n8454), .ZN(n8243) );
  INV_X1 U6308 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5089) );
  OR2_X1 U6309 ( .A1(n5771), .A2(n8922), .ZN(n5788) );
  OR2_X1 U6310 ( .A1(n5797), .A2(n9150), .ZN(n5809) );
  NAND2_X1 U6311 ( .A1(n5807), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5822) );
  OR2_X1 U6312 ( .A1(n5729), .A2(n5728), .ZN(n5745) );
  OR2_X1 U6313 ( .A1(n5822), .A2(n5821), .ZN(n5838) );
  AND2_X1 U6314 ( .A1(n9364), .A2(n5918), .ZN(n9389) );
  INV_X1 U6315 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9064) );
  INV_X1 U6316 ( .A(n9466), .ZN(n9425) );
  AND2_X1 U6317 ( .A1(n5961), .A2(n6411), .ZN(n6954) );
  NAND2_X1 U6318 ( .A1(n9655), .A2(n9785), .ZN(n6038) );
  OR2_X1 U6319 ( .A1(n9521), .A2(n9269), .ZN(n6020) );
  OR2_X1 U6320 ( .A1(n9775), .A2(n9272), .ZN(n6014) );
  NOR2_X1 U6321 ( .A1(n9723), .A2(n9275), .ZN(n6008) );
  AND2_X1 U6322 ( .A1(n5940), .A2(n7985), .ZN(n9995) );
  AND2_X1 U6323 ( .A1(n5402), .A2(n5387), .ZN(n5400) );
  NAND2_X1 U6324 ( .A1(n5232), .A2(n4933), .ZN(n5216) );
  INV_X1 U6325 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5630) );
  AOI22_X1 U6326 ( .A1(n6760), .A2(n6761), .B1(n6756), .B2(n6651), .ZN(n6658)
         );
  AOI22_X1 U6327 ( .A1(n7321), .A2(n7320), .B1(n7319), .B2(n7318), .ZN(n7323)
         );
  INV_X1 U6328 ( .A(n8453), .ZN(n8420) );
  INV_X1 U6329 ( .A(n8404), .ZN(n8450) );
  AND2_X1 U6330 ( .A1(n5398), .A2(n5397), .ZN(n8080) );
  AND2_X1 U6331 ( .A1(n8177), .A2(n8176), .ZN(n8292) );
  OR2_X1 U6332 ( .A1(n10108), .A2(n6774), .ZN(n8682) );
  AND2_X1 U6333 ( .A1(n6634), .A2(n6056), .ZN(n6773) );
  NAND2_X1 U6334 ( .A1(n8222), .A2(n8225), .ZN(n8704) );
  NAND2_X1 U6335 ( .A1(n8277), .A2(n7416), .ZN(n10108) );
  AND2_X1 U6336 ( .A1(n7198), .A2(n10102), .ZN(n10113) );
  INV_X1 U6337 ( .A(n10108), .ZN(n10118) );
  INV_X1 U6338 ( .A(n10113), .ZN(n10080) );
  INV_X1 U6339 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5125) );
  INV_X1 U6340 ( .A(n9262), .ZN(n9852) );
  NAND2_X1 U6341 ( .A1(n7981), .A2(n9330), .ZN(n8044) );
  OR2_X1 U6342 ( .A1(n9245), .A2(n5908), .ZN(n5913) );
  INV_X1 U6343 ( .A(n9837), .ZN(n9943) );
  OR2_X1 U6344 ( .A1(n9680), .A2(n9475), .ZN(n9454) );
  AND2_X1 U6345 ( .A1(n7865), .A2(n9951), .ZN(n7210) );
  AND2_X1 U6346 ( .A1(n9984), .A2(n6035), .ZN(n9637) );
  NOR2_X1 U6347 ( .A1(n9380), .A2(n9374), .ZN(n9656) );
  AND2_X1 U6348 ( .A1(n10042), .A2(n9724), .ZN(n9719) );
  INV_X1 U6349 ( .A(n7830), .ZN(n9392) );
  OR2_X1 U6350 ( .A1(n7984), .A2(n5962), .ZN(n9727) );
  NAND2_X1 U6351 ( .A1(n6958), .A2(n9727), .ZN(n10026) );
  AND2_X1 U6352 ( .A1(n5985), .A2(n6955), .ZN(n6369) );
  XNOR2_X1 U6353 ( .A(n5364), .B(n5363), .ZN(n7468) );
  AND2_X1 U6354 ( .A1(n5714), .A2(n5724), .ZN(n6487) );
  AND2_X1 U6355 ( .A1(n6754), .A2(n8324), .ZN(n8404) );
  OR2_X1 U6356 ( .A1(n6664), .A2(n6662), .ZN(n8453) );
  AND2_X1 U6357 ( .A1(n7128), .A2(n5468), .ZN(n8097) );
  AOI211_X1 U6358 ( .C1(n8785), .C2(n8337), .A(n8336), .B(n8335), .ZN(n8338)
         );
  AND2_X1 U6359 ( .A1(n6779), .A2(n8756), .ZN(n8767) );
  OR2_X1 U6360 ( .A1(n8767), .A2(n6776), .ZN(n8788) );
  INV_X1 U6361 ( .A(n10135), .ZN(n10133) );
  OR2_X1 U6362 ( .A1(n10121), .A2(n10108), .ZN(n8878) );
  OR2_X1 U6363 ( .A1(n10121), .A2(n10113), .ZN(n8894) );
  AND2_X1 U6364 ( .A1(n6642), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6753) );
  INV_X1 U6365 ( .A(n6643), .ZN(n8277) );
  INV_X1 U6366 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6425) );
  INV_X1 U6367 ( .A(n9723), .ZN(n9623) );
  NAND2_X1 U6368 ( .A1(n8910), .A2(n6320), .ZN(n6335) );
  INV_X1 U6369 ( .A(n9676), .ZN(n9450) );
  INV_X1 U6370 ( .A(n9703), .ZN(n9556) );
  NAND2_X1 U6371 ( .A1(n5900), .A2(n5899), .ZN(n9267) );
  NAND2_X1 U6372 ( .A1(n9984), .A2(n6959), .ZN(n9606) );
  INV_X1 U6373 ( .A(n10042), .ZN(n10039) );
  INV_X1 U6374 ( .A(n6039), .ZN(n6040) );
  INV_X1 U6375 ( .A(n9785), .ZN(n9781) );
  INV_X1 U6376 ( .A(n10030), .ZN(n10028) );
  INV_X1 U6377 ( .A(n9992), .ZN(n9993) );
  INV_X1 U6378 ( .A(n5964), .ZN(n7555) );
  INV_X1 U6379 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6423) );
  INV_X1 U6380 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6409) );
  INV_X1 U6381 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U6382 ( .A1(n6053), .A2(n6052), .ZN(P2_U3487) );
  NAND2_X1 U6383 ( .A1(n6066), .A2(n6065), .ZN(P2_U3455) );
  NAND2_X1 U6384 ( .A1(n6041), .A2(n6040), .ZN(P1_U3518) );
  NAND2_X1 U6385 ( .A1(n4880), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4881) );
  INV_X1 U6386 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6387) );
  INV_X1 U6387 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6398) );
  XNOR2_X1 U6388 ( .A(n4884), .B(SI_1_), .ZN(n5018) );
  NAND3_X1 U6389 ( .A1(n6357), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4883) );
  AND2_X1 U6390 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U6391 ( .A1(n6388), .A2(n4882), .ZN(n5032) );
  NAND2_X1 U6392 ( .A1(n4883), .A2(n5032), .ZN(n5017) );
  NAND2_X1 U6393 ( .A1(n5018), .A2(n5017), .ZN(n4887) );
  INV_X1 U6394 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6395 ( .A1(n4885), .A2(SI_1_), .ZN(n4886) );
  NAND2_X1 U6396 ( .A1(n4887), .A2(n4886), .ZN(n5046) );
  INV_X1 U6397 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6394) );
  INV_X1 U6398 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U6399 ( .A1(n6357), .A2(n6385), .ZN(n4888) );
  XNOR2_X1 U6400 ( .A(n4889), .B(SI_2_), .ZN(n5045) );
  NAND2_X1 U6401 ( .A1(n5046), .A2(n5045), .ZN(n4892) );
  INV_X1 U6402 ( .A(n4889), .ZN(n4890) );
  NAND2_X1 U6403 ( .A1(n4890), .A2(SI_2_), .ZN(n4891) );
  NAND2_X1 U6404 ( .A1(n4892), .A2(n4891), .ZN(n5063) );
  INV_X1 U6405 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6406 ( .A1(n4895), .A2(SI_3_), .ZN(n4896) );
  INV_X1 U6407 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6390) );
  INV_X1 U6408 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6386) );
  INV_X1 U6409 ( .A(n4897), .ZN(n4898) );
  NAND2_X1 U6410 ( .A1(n4898), .A2(SI_4_), .ZN(n4899) );
  MUX2_X1 U6411 ( .A(n6392), .B(n9027), .S(n6389), .Z(n4900) );
  INV_X1 U6412 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6413 ( .A1(n4901), .A2(SI_5_), .ZN(n4902) );
  MUX2_X1 U6414 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6389), .Z(n4905) );
  NAND2_X1 U6415 ( .A1(n5129), .A2(n4904), .ZN(n4907) );
  NAND2_X1 U6416 ( .A1(n4905), .A2(SI_7_), .ZN(n4906) );
  INV_X1 U6417 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4908) );
  INV_X1 U6418 ( .A(SI_8_), .ZN(n4909) );
  INV_X1 U6419 ( .A(n4910), .ZN(n4911) );
  NAND2_X1 U6420 ( .A1(n4911), .A2(SI_8_), .ZN(n4912) );
  MUX2_X1 U6421 ( .A(n6420), .B(n6419), .S(n6389), .Z(n4914) );
  INV_X1 U6422 ( .A(SI_9_), .ZN(n8998) );
  INV_X1 U6423 ( .A(n4914), .ZN(n4915) );
  NAND2_X1 U6424 ( .A1(n4915), .A2(SI_9_), .ZN(n4916) );
  MUX2_X1 U6425 ( .A(n6425), .B(n6423), .S(n6389), .Z(n4918) );
  INV_X1 U6426 ( .A(n4918), .ZN(n4919) );
  INV_X1 U6427 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6479) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6481) );
  MUX2_X1 U6429 ( .A(n6479), .B(n6481), .S(n6389), .Z(n4920) );
  INV_X1 U6430 ( .A(SI_11_), .ZN(n9008) );
  INV_X1 U6431 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6432 ( .A1(n4921), .A2(SI_11_), .ZN(n4922) );
  INV_X1 U6433 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6533) );
  MUX2_X1 U6434 ( .A(n8991), .B(n6533), .S(n6389), .Z(n4924) );
  INV_X1 U6435 ( .A(n4924), .ZN(n4925) );
  MUX2_X1 U6436 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6389), .Z(n4929) );
  NAND2_X1 U6437 ( .A1(n4929), .A2(SI_13_), .ZN(n4930) );
  INV_X1 U6438 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6749) );
  INV_X1 U6439 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8967) );
  MUX2_X1 U6440 ( .A(n6749), .B(n8967), .S(n6389), .Z(n4931) );
  INV_X1 U6441 ( .A(SI_14_), .ZN(n9004) );
  INV_X1 U6442 ( .A(n4931), .ZN(n4932) );
  NAND2_X1 U6443 ( .A1(n4932), .A2(SI_14_), .ZN(n4933) );
  INV_X1 U6444 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6831) );
  INV_X1 U6445 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U6446 ( .A(n6831), .B(n4935), .S(n6389), .Z(n4937) );
  XNOR2_X1 U6447 ( .A(n4937), .B(SI_15_), .ZN(n5234) );
  NAND2_X1 U6448 ( .A1(n5233), .A2(n4936), .ZN(n4940) );
  INV_X1 U6449 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6450 ( .A1(n4938), .A2(SI_15_), .ZN(n4939) );
  MUX2_X1 U6451 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6389), .Z(n4942) );
  XNOR2_X1 U6452 ( .A(n4942), .B(SI_16_), .ZN(n5248) );
  INV_X1 U6453 ( .A(n5248), .ZN(n4941) );
  NAND2_X1 U6454 ( .A1(n5249), .A2(n4941), .ZN(n4944) );
  NAND2_X1 U6455 ( .A1(n4942), .A2(SI_16_), .ZN(n4943) );
  INV_X1 U6456 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6884) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n4945) );
  MUX2_X1 U6458 ( .A(n6884), .B(n4945), .S(n6389), .Z(n4947) );
  INV_X1 U6459 ( .A(SI_17_), .ZN(n4946) );
  NAND2_X1 U6460 ( .A1(n4947), .A2(n4946), .ZN(n4950) );
  INV_X1 U6461 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6462 ( .A1(n4948), .A2(SI_17_), .ZN(n4949) );
  NAND2_X1 U6463 ( .A1(n4950), .A2(n4949), .ZN(n5264) );
  INV_X1 U6464 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6924) );
  INV_X1 U6465 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6972) );
  MUX2_X1 U6466 ( .A(n6924), .B(n6972), .S(n6389), .Z(n4951) );
  XNOR2_X1 U6467 ( .A(n4951), .B(SI_18_), .ZN(n5278) );
  INV_X1 U6468 ( .A(n5278), .ZN(n4954) );
  INV_X1 U6469 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6470 ( .A1(n4952), .A2(SI_18_), .ZN(n4953) );
  INV_X1 U6471 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7234) );
  INV_X1 U6472 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7131) );
  MUX2_X1 U6473 ( .A(n7234), .B(n7131), .S(n6389), .Z(n4956) );
  INV_X1 U6474 ( .A(SI_19_), .ZN(n4955) );
  NAND2_X1 U6475 ( .A1(n4956), .A2(n4955), .ZN(n4959) );
  INV_X1 U6476 ( .A(n4956), .ZN(n4957) );
  NAND2_X1 U6477 ( .A1(n4957), .A2(SI_19_), .ZN(n4958) );
  NAND2_X1 U6478 ( .A1(n4959), .A2(n4958), .ZN(n5296) );
  MUX2_X1 U6479 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6357), .Z(n5310) );
  INV_X1 U6480 ( .A(SI_20_), .ZN(n5312) );
  XNOR2_X1 U6481 ( .A(n5310), .B(n5312), .ZN(n4960) );
  XNOR2_X1 U6482 ( .A(n5313), .B(n4960), .ZN(n7247) );
  NOR2_X1 U6483 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4968) );
  NOR2_X1 U6484 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4967) );
  AND2_X1 U6485 ( .A1(n4968), .A2(n4967), .ZN(n4971) );
  INV_X2 U6486 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9019) );
  NOR2_X1 U6487 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4969) );
  INV_X1 U6488 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4972) );
  NOR3_X1 U6489 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5525) );
  INV_X1 U6490 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4973) );
  AND2_X1 U6491 ( .A1(n5525), .A2(n4973), .ZN(n4974) );
  INV_X1 U6492 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4999) );
  XNOR2_X2 U6493 ( .A(n4976), .B(n4999), .ZN(n7748) );
  INV_X1 U6494 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4977) );
  NAND2_X2 U6495 ( .A1(n7748), .A2(n6596), .ZN(n5034) );
  NAND2_X2 U6496 ( .A1(n5034), .A2(n6388), .ZN(n8103) );
  NAND2_X1 U6497 ( .A1(n7247), .A2(n8252), .ZN(n4979) );
  NAND2_X4 U6498 ( .A1(n5034), .A2(n6389), .ZN(n8253) );
  INV_X1 U6499 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9007) );
  OR2_X1 U6500 ( .A1(n8253), .A2(n9007), .ZN(n4978) );
  INV_X1 U6501 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n4986) );
  INV_X1 U6502 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n4988) );
  INV_X1 U6503 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n4990) );
  INV_X1 U6504 ( .A(n5240), .ZN(n4993) );
  INV_X1 U6505 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4992) );
  INV_X1 U6506 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4994) );
  INV_X1 U6507 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U6508 ( .A1(n5306), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6509 ( .A1(n5321), .A2(n4998), .ZN(n8733) );
  INV_X1 U6510 ( .A(n5003), .ZN(n5001) );
  NAND2_X1 U6511 ( .A1(n5001), .A2(n5004), .ZN(n8897) );
  INV_X1 U6512 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U6513 ( .A1(n8733), .A2(n5464), .ZN(n5011) );
  AOI22_X1 U6514 ( .A1(n5500), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7119), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5010) );
  NAND2_X2 U6515 ( .A1(n8342), .A2(n5008), .ZN(n5272) );
  INV_X1 U6516 ( .A(n7124), .ZN(n5501) );
  NAND2_X1 U6517 ( .A1(n5501), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5009) );
  INV_X1 U6518 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5012) );
  INV_X1 U6519 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6553) );
  OR2_X1 U6520 ( .A1(n7121), .A2(n6553), .ZN(n5015) );
  INV_X1 U6521 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6780) );
  OR2_X1 U6522 ( .A1(n5039), .A2(n6780), .ZN(n5014) );
  INV_X1 U6523 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U6524 ( .A(n5018), .B(n5017), .ZN(n6399) );
  OR2_X1 U6525 ( .A1(n8103), .A2(n6399), .ZN(n5023) );
  NAND2_X1 U6526 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5019) );
  MUX2_X1 U6527 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5019), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5021) );
  INV_X1 U6528 ( .A(n5047), .ZN(n5020) );
  OR2_X1 U6529 ( .A1(n5034), .A2(n6695), .ZN(n5022) );
  INV_X1 U6530 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5026) );
  INV_X1 U6531 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7769) );
  INV_X1 U6532 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7766) );
  OR2_X1 U6533 ( .A1(n5039), .A2(n7766), .ZN(n5028) );
  INV_X1 U6534 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6628) );
  OR2_X1 U6535 ( .A1(n7121), .A2(n6628), .ZN(n5027) );
  NAND2_X1 U6536 ( .A1(n6388), .A2(SI_0_), .ZN(n5031) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6538 ( .A1(n5031), .A2(n5030), .ZN(n5033) );
  AND2_X1 U6539 ( .A1(n5033), .A2(n5032), .ZN(n8908) );
  NAND2_X1 U6540 ( .A1(n6783), .A2(n7760), .ZN(n6781) );
  NAND2_X1 U6541 ( .A1(n6777), .A2(n6781), .ZN(n5036) );
  OR2_X1 U6542 ( .A1(n6625), .A2(n6648), .ZN(n5035) );
  NAND2_X1 U6543 ( .A1(n5036), .A2(n5035), .ZN(n6676) );
  INV_X1 U6544 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5037) );
  OR2_X1 U6545 ( .A1(n5038), .A2(n5037), .ZN(n5043) );
  INV_X1 U6546 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6917) );
  OR2_X1 U6547 ( .A1(n5039), .A2(n6917), .ZN(n5042) );
  INV_X1 U6548 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5040) );
  OR2_X1 U6549 ( .A1(n5272), .A2(n5040), .ZN(n5041) );
  XNOR2_X1 U6550 ( .A(n5046), .B(n5045), .ZN(n6395) );
  OR2_X1 U6551 ( .A1(n8103), .A2(n6395), .ZN(n5052) );
  OR2_X1 U6552 ( .A1(n8253), .A2(n6394), .ZN(n5051) );
  INV_X1 U6553 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5147) );
  NOR2_X1 U6554 ( .A1(n5047), .A2(n5147), .ZN(n5048) );
  OR2_X1 U6555 ( .A1(n5506), .A2(n6579), .ZN(n5050) );
  OR2_X1 U6556 ( .A1(n8476), .A2(n6916), .ZN(n8112) );
  NAND2_X1 U6557 ( .A1(n8476), .A2(n6916), .ZN(n8113) );
  INV_X1 U6558 ( .A(n6916), .ZN(n6762) );
  OR2_X1 U6559 ( .A1(n8476), .A2(n6762), .ZN(n5053) );
  INV_X1 U6560 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6561 ( .A1(n7121), .A2(n5054), .ZN(n5058) );
  OR2_X1 U6562 ( .A1(n5211), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5057) );
  INV_X1 U6563 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5055) );
  OR2_X1 U6564 ( .A1(n5272), .A2(n5055), .ZN(n5056) );
  MUX2_X1 U6565 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5060), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5061) );
  NAND2_X1 U6566 ( .A1(n5061), .A2(n5088), .ZN(n6720) );
  XNOR2_X1 U6567 ( .A(n5063), .B(n5062), .ZN(n6397) );
  OR2_X1 U6568 ( .A1(n8103), .A2(n6397), .ZN(n5065) );
  OR2_X1 U6569 ( .A1(n8253), .A2(n6396), .ZN(n5064) );
  OAI211_X1 U6570 ( .C1(n5506), .C2(n6720), .A(n5065), .B(n5064), .ZN(n7062)
         );
  NAND2_X1 U6571 ( .A1(n7119), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5070) );
  OR2_X1 U6572 ( .A1(n5272), .A2(n4708), .ZN(n5069) );
  NAND2_X1 U6573 ( .A1(n5080), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5066) );
  AND2_X1 U6574 ( .A1(n5103), .A2(n5066), .ZN(n6889) );
  OR2_X1 U6575 ( .A1(n5211), .A2(n6889), .ZN(n5068) );
  OR2_X1 U6576 ( .A1(n7121), .A2(n4569), .ZN(n5067) );
  NAND2_X1 U6577 ( .A1(n5091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5071) );
  MUX2_X1 U6578 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5071), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5073) );
  INV_X1 U6579 ( .A(n5091), .ZN(n5072) );
  INV_X1 U6580 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U6581 ( .A1(n5072), .A2(n9014), .ZN(n5124) );
  NAND2_X1 U6582 ( .A1(n5073), .A2(n5124), .ZN(n6585) );
  XNOR2_X1 U6583 ( .A(n5075), .B(n5074), .ZN(n6393) );
  OR2_X1 U6584 ( .A1(n8103), .A2(n6393), .ZN(n5077) );
  OR2_X1 U6585 ( .A1(n8253), .A2(n6392), .ZN(n5076) );
  NAND2_X1 U6586 ( .A1(n8474), .A2(n10081), .ZN(n5097) );
  NAND2_X1 U6587 ( .A1(n5500), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5085) );
  INV_X1 U6588 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5078) );
  OR2_X1 U6589 ( .A1(n5038), .A2(n5078), .ZN(n5084) );
  NAND2_X1 U6590 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5079) );
  AND2_X1 U6591 ( .A1(n5080), .A2(n5079), .ZN(n6908) );
  INV_X1 U6592 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5081) );
  OR2_X1 U6593 ( .A1(n5272), .A2(n5081), .ZN(n5082) );
  OR2_X1 U6594 ( .A1(n8103), .A2(n6391), .ZN(n5095) );
  OR2_X1 U6595 ( .A1(n8253), .A2(n6390), .ZN(n5094) );
  NAND2_X1 U6596 ( .A1(n5088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5090) );
  MUX2_X1 U6597 ( .A(n5090), .B(P2_IR_REG_31__SCAN_IN), .S(n5089), .Z(n5092)
         );
  NAND2_X1 U6598 ( .A1(n5092), .A2(n5091), .ZN(n6624) );
  OR2_X1 U6599 ( .A1(n5506), .A2(n6624), .ZN(n5093) );
  XNOR2_X1 U6600 ( .A(n5481), .B(n10076), .ZN(n8283) );
  AND2_X1 U6601 ( .A1(n5097), .A2(n8283), .ZN(n5096) );
  NAND2_X1 U6602 ( .A1(n6909), .A2(n5096), .ZN(n5102) );
  INV_X1 U6603 ( .A(n5097), .ZN(n5100) );
  OR2_X1 U6604 ( .A1(n8474), .A2(n10081), .ZN(n5098) );
  INV_X1 U6605 ( .A(n10076), .ZN(n6824) );
  OR2_X1 U6606 ( .A1(n5481), .A2(n6824), .ZN(n6976) );
  AND2_X1 U6607 ( .A1(n5098), .A2(n6976), .ZN(n5099) );
  OR2_X1 U6608 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  NAND2_X1 U6609 ( .A1(n7119), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5108) );
  INV_X1 U6610 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6588) );
  OR2_X1 U6611 ( .A1(n7121), .A2(n6588), .ZN(n5107) );
  NAND2_X1 U6612 ( .A1(n5103), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5104) );
  AND2_X1 U6613 ( .A1(n5118), .A2(n5104), .ZN(n6902) );
  OR2_X1 U6614 ( .A1(n5211), .A2(n6902), .ZN(n5106) );
  INV_X1 U6615 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6901) );
  OR2_X1 U6616 ( .A1(n7124), .A2(n6901), .ZN(n5105) );
  NAND2_X1 U6617 ( .A1(n6899), .A2(n7113), .ZN(n5114) );
  NAND2_X1 U6618 ( .A1(n5124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U6619 ( .A(n5109), .B(n5125), .ZN(n6798) );
  XNOR2_X1 U6620 ( .A(n5111), .B(n5110), .ZN(n6400) );
  OR2_X1 U6621 ( .A1(n8103), .A2(n6400), .ZN(n5113) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9005) );
  OR2_X1 U6623 ( .A1(n8253), .A2(n9005), .ZN(n5112) );
  OAI211_X1 U6624 ( .C1(n5506), .C2(n6798), .A(n5113), .B(n5112), .ZN(n6903)
         );
  NAND2_X1 U6625 ( .A1(n5114), .A2(n6903), .ZN(n5117) );
  INV_X1 U6626 ( .A(n6899), .ZN(n5115) );
  NAND2_X1 U6627 ( .A1(n5115), .A2(n8473), .ZN(n5116) );
  NAND2_X1 U6628 ( .A1(n7119), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5123) );
  OR2_X1 U6629 ( .A1(n7121), .A2(n4576), .ZN(n5122) );
  NAND2_X1 U6630 ( .A1(n5118), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5119) );
  AND2_X1 U6631 ( .A1(n5139), .A2(n5119), .ZN(n7114) );
  OR2_X1 U6632 ( .A1(n5211), .A2(n7114), .ZN(n5121) );
  INV_X1 U6633 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6792) );
  OR2_X1 U6634 ( .A1(n7124), .A2(n6792), .ZN(n5120) );
  NAND4_X1 U6635 ( .A1(n5123), .A2(n5122), .A3(n5121), .A4(n5120), .ZN(n8472)
         );
  INV_X1 U6636 ( .A(n5124), .ZN(n5126) );
  NAND2_X1 U6637 ( .A1(n5126), .A2(n5125), .ZN(n5135) );
  NAND2_X1 U6638 ( .A1(n5135), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6639 ( .A(n5127), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6927) );
  AOI22_X1 U6640 ( .A1(n5299), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6382), .B2(
        n6927), .ZN(n5131) );
  XNOR2_X1 U6641 ( .A(n5129), .B(n5128), .ZN(n6404) );
  NAND2_X1 U6642 ( .A1(n6404), .A2(n8252), .ZN(n5130) );
  OR2_X1 U6643 ( .A1(n8472), .A2(n10093), .ZN(n8145) );
  NAND2_X1 U6644 ( .A1(n8472), .A2(n10093), .ZN(n7099) );
  NAND2_X1 U6645 ( .A1(n8145), .A2(n7099), .ZN(n5483) );
  INV_X1 U6646 ( .A(n10093), .ZN(n7043) );
  NAND2_X1 U6647 ( .A1(n8472), .A2(n7043), .ZN(n5132) );
  OAI21_X1 U6648 ( .B1(n5135), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5136) );
  XNOR2_X1 U6649 ( .A(n5136), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U6650 ( .A1(n5299), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6382), .B2(
        n10048), .ZN(n5137) );
  NAND2_X1 U6651 ( .A1(n5500), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5144) );
  INV_X1 U6652 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5138) );
  OR2_X1 U6653 ( .A1(n5038), .A2(n5138), .ZN(n5143) );
  NAND2_X1 U6654 ( .A1(n5139), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5140) );
  AND2_X1 U6655 ( .A1(n5152), .A2(n5140), .ZN(n7242) );
  OR2_X1 U6656 ( .A1(n5211), .A2(n7242), .ZN(n5142) );
  INV_X1 U6657 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6943) );
  OR2_X1 U6658 ( .A1(n5272), .A2(n6943), .ZN(n5141) );
  NAND4_X1 U6659 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n8471)
         );
  AND2_X1 U6660 ( .A1(n7244), .A2(n8471), .ZN(n5145) );
  OR2_X1 U6661 ( .A1(n7244), .A2(n8471), .ZN(n5146) );
  INV_X1 U6662 ( .A(n7194), .ZN(n5158) );
  NAND2_X1 U6663 ( .A1(n6418), .A2(n8252), .ZN(n5151) );
  OR2_X1 U6664 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  XNOR2_X1 U6665 ( .A(n5149), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7134) );
  AOI22_X1 U6666 ( .A1(n5299), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6382), .B2(
        n7134), .ZN(n5150) );
  NAND2_X1 U6667 ( .A1(n5151), .A2(n5150), .ZN(n10106) );
  NAND2_X1 U6668 ( .A1(n7119), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5157) );
  INV_X1 U6669 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6932) );
  OR2_X1 U6670 ( .A1(n7124), .A2(n6932), .ZN(n5156) );
  NAND2_X1 U6671 ( .A1(n5152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5153) );
  AND2_X1 U6672 ( .A1(n5169), .A2(n5153), .ZN(n7327) );
  OR2_X1 U6673 ( .A1(n5211), .A2(n7327), .ZN(n5155) );
  INV_X1 U6674 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6931) );
  OR2_X1 U6675 ( .A1(n7121), .A2(n6931), .ZN(n5154) );
  NAND4_X1 U6676 ( .A1(n5157), .A2(n5156), .A3(n5155), .A4(n5154), .ZN(n8470)
         );
  NAND2_X1 U6677 ( .A1(n10106), .A2(n8470), .ZN(n5159) );
  XNOR2_X1 U6678 ( .A(n5162), .B(n5161), .ZN(n6422) );
  NAND2_X1 U6679 ( .A1(n6422), .A2(n8252), .ZN(n5167) );
  NAND2_X1 U6680 ( .A1(n5163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  MUX2_X1 U6681 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5164), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5165) );
  AND2_X1 U6682 ( .A1(n5165), .A2(n4310), .ZN(n7496) );
  AOI22_X1 U6683 ( .A1(n5299), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6382), .B2(
        n7496), .ZN(n5166) );
  NAND2_X1 U6684 ( .A1(n5167), .A2(n5166), .ZN(n7532) );
  NAND2_X1 U6685 ( .A1(n5500), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5174) );
  INV_X1 U6686 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6687 ( .A1(n5038), .A2(n5168), .ZN(n5173) );
  NAND2_X1 U6688 ( .A1(n5169), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5170) );
  AND2_X1 U6689 ( .A1(n5182), .A2(n5170), .ZN(n7426) );
  OR2_X1 U6690 ( .A1(n5211), .A2(n7426), .ZN(n5172) );
  INV_X1 U6691 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7489) );
  OR2_X1 U6692 ( .A1(n7124), .A2(n7489), .ZN(n5171) );
  NAND4_X1 U6693 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n8469)
         );
  AND2_X1 U6694 ( .A1(n7532), .A2(n8469), .ZN(n5176) );
  XNOR2_X1 U6695 ( .A(n5178), .B(n5177), .ZN(n6478) );
  NAND2_X1 U6696 ( .A1(n6478), .A2(n8252), .ZN(n5181) );
  NAND2_X1 U6697 ( .A1(n4310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6698 ( .A(n5179), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7508) );
  AOI22_X1 U6699 ( .A1(n5299), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6382), .B2(
        n7508), .ZN(n5180) );
  NAND2_X1 U6700 ( .A1(n5181), .A2(n5180), .ZN(n10117) );
  NAND2_X1 U6701 ( .A1(n7119), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5187) );
  INV_X1 U6702 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7505) );
  OR2_X1 U6703 ( .A1(n7121), .A2(n7505), .ZN(n5186) );
  NAND2_X1 U6704 ( .A1(n5182), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5183) );
  AND2_X1 U6705 ( .A1(n5195), .A2(n5183), .ZN(n7476) );
  OR2_X1 U6706 ( .A1(n5211), .A2(n7476), .ZN(n5185) );
  INV_X1 U6707 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7506) );
  OR2_X1 U6708 ( .A1(n7124), .A2(n7506), .ZN(n5184) );
  NAND2_X1 U6709 ( .A1(n10117), .A2(n7537), .ZN(n8157) );
  INV_X1 U6710 ( .A(n7537), .ZN(n8468) );
  NAND2_X1 U6711 ( .A1(n10117), .A2(n8468), .ZN(n5188) );
  XNOR2_X1 U6712 ( .A(n5190), .B(n5189), .ZN(n6526) );
  NAND2_X1 U6713 ( .A1(n6526), .A2(n8252), .ZN(n5194) );
  OR2_X2 U6714 ( .A1(n4310), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6715 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  INV_X1 U6716 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U6717 ( .A(n5192), .B(n5191), .ZN(n7706) );
  INV_X1 U6718 ( .A(n7706), .ZN(n7652) );
  AOI22_X1 U6719 ( .A1(n5299), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6382), .B2(
        n7652), .ZN(n5193) );
  NAND2_X1 U6720 ( .A1(n7119), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5200) );
  INV_X1 U6721 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7636) );
  OR2_X1 U6722 ( .A1(n7121), .A2(n7636), .ZN(n5199) );
  NAND2_X1 U6723 ( .A1(n5195), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5196) );
  AND2_X1 U6724 ( .A1(n5209), .A2(n5196), .ZN(n7528) );
  OR2_X1 U6725 ( .A1(n5211), .A2(n7528), .ZN(n5198) );
  INV_X1 U6726 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7637) );
  OR2_X1 U6727 ( .A1(n5272), .A2(n7637), .ZN(n5197) );
  NAND4_X1 U6728 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n8467)
         );
  OR2_X1 U6729 ( .A1(n8169), .A2(n8467), .ZN(n5202) );
  AND2_X1 U6730 ( .A1(n8169), .A2(n8467), .ZN(n5201) );
  XNOR2_X1 U6731 ( .A(n5204), .B(n5203), .ZN(n6548) );
  NAND2_X1 U6732 ( .A1(n6548), .A2(n8252), .ZN(n5208) );
  NOR2_X2 U6733 ( .A1(n5205), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5218) );
  OR2_X1 U6734 ( .A1(n5218), .A2(n5147), .ZN(n5206) );
  XNOR2_X1 U6735 ( .A(n5206), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7725) );
  AOI22_X1 U6736 ( .A1(n5299), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6382), .B2(
        n7725), .ZN(n5207) );
  NAND2_X1 U6737 ( .A1(n7119), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5215) );
  INV_X1 U6738 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7713) );
  OR2_X1 U6739 ( .A1(n7124), .A2(n7713), .ZN(n5214) );
  NAND2_X1 U6740 ( .A1(n5209), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5210) );
  AND2_X1 U6741 ( .A1(n5223), .A2(n5210), .ZN(n7588) );
  OR2_X1 U6742 ( .A1(n5211), .A2(n7588), .ZN(n5213) );
  INV_X1 U6743 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7712) );
  OR2_X1 U6744 ( .A1(n7121), .A2(n7712), .ZN(n5212) );
  NAND4_X1 U6745 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n8466)
         );
  NAND2_X1 U6746 ( .A1(n8174), .A2(n8466), .ZN(n8176) );
  NAND2_X1 U6747 ( .A1(n7456), .A2(n8177), .ZN(n7615) );
  NAND2_X1 U6748 ( .A1(n6748), .A2(n8252), .ZN(n5222) );
  NAND2_X1 U6749 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5251) );
  INV_X1 U6750 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6751 ( .A1(n5251), .A2(n5219), .ZN(n5236) );
  OR2_X1 U6752 ( .A1(n5251), .A2(n5219), .ZN(n5220) );
  NAND2_X1 U6753 ( .A1(n5236), .A2(n5220), .ZN(n8507) );
  INV_X1 U6754 ( .A(n8507), .ZN(n8505) );
  AOI22_X1 U6755 ( .A1(n5299), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6382), .B2(
        n8505), .ZN(n5221) );
  NAND2_X1 U6756 ( .A1(n7119), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5228) );
  INV_X1 U6757 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8483) );
  OR2_X1 U6758 ( .A1(n7121), .A2(n8483), .ZN(n5227) );
  NAND2_X1 U6759 ( .A1(n5223), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5224) );
  AND2_X1 U6760 ( .A1(n5240), .A2(n5224), .ZN(n7675) );
  OR2_X1 U6761 ( .A1(n5039), .A2(n7675), .ZN(n5226) );
  INV_X1 U6762 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8504) );
  OR2_X1 U6763 ( .A1(n7124), .A2(n8504), .ZN(n5225) );
  NAND4_X1 U6764 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n8465)
         );
  NAND2_X1 U6765 ( .A1(n7677), .A2(n8465), .ZN(n5229) );
  NAND2_X1 U6766 ( .A1(n7615), .A2(n5229), .ZN(n5231) );
  OR2_X1 U6767 ( .A1(n7677), .A2(n8465), .ZN(n5230) );
  NAND2_X1 U6768 ( .A1(n5231), .A2(n5230), .ZN(n7659) );
  NAND2_X1 U6769 ( .A1(n5233), .A2(n5232), .ZN(n5235) );
  XNOR2_X1 U6770 ( .A(n5235), .B(n5234), .ZN(n6808) );
  NAND2_X1 U6771 ( .A1(n6808), .A2(n8252), .ZN(n5239) );
  NAND2_X1 U6772 ( .A1(n5236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U6773 ( .A(n5237), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8524) );
  AOI22_X1 U6774 ( .A1(n5299), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6382), .B2(
        n8524), .ZN(n5238) );
  NAND2_X1 U6775 ( .A1(n7119), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5245) );
  INV_X1 U6776 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8512) );
  OR2_X1 U6777 ( .A1(n7121), .A2(n8512), .ZN(n5244) );
  NAND2_X1 U6778 ( .A1(n5240), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5241) );
  AND2_X1 U6779 ( .A1(n5256), .A2(n5241), .ZN(n7661) );
  OR2_X1 U6780 ( .A1(n5039), .A2(n7661), .ZN(n5243) );
  INV_X1 U6781 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8513) );
  OR2_X1 U6782 ( .A1(n5272), .A2(n8513), .ZN(n5242) );
  NAND2_X1 U6783 ( .A1(n7690), .A2(n8392), .ZN(n8196) );
  NAND2_X1 U6784 ( .A1(n8187), .A2(n8196), .ZN(n8186) );
  NAND2_X1 U6785 ( .A1(n7659), .A2(n8186), .ZN(n5247) );
  INV_X1 U6786 ( .A(n8392), .ZN(n8464) );
  OR2_X1 U6787 ( .A1(n7690), .A2(n8464), .ZN(n5246) );
  XNOR2_X1 U6788 ( .A(n5249), .B(n5248), .ZN(n6853) );
  NAND2_X1 U6789 ( .A1(n6853), .A2(n8252), .ZN(n5255) );
  OR2_X1 U6790 ( .A1(n5281), .A2(n5147), .ZN(n5250) );
  NAND2_X1 U6791 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  OR2_X1 U6792 ( .A1(n5252), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6793 ( .A1(n5252), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5253) );
  AND2_X1 U6794 ( .A1(n5266), .A2(n5253), .ZN(n8547) );
  AOI22_X1 U6795 ( .A1(n5299), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6382), .B2(
        n8547), .ZN(n5254) );
  NAND2_X1 U6796 ( .A1(n7119), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5261) );
  INV_X1 U6797 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9075) );
  OR2_X1 U6798 ( .A1(n7121), .A2(n9075), .ZN(n5260) );
  NAND2_X1 U6799 ( .A1(n5256), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5257) );
  AND2_X1 U6800 ( .A1(n5270), .A2(n5257), .ZN(n8393) );
  OR2_X1 U6801 ( .A1(n5039), .A2(n8393), .ZN(n5259) );
  INV_X1 U6802 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8546) );
  OR2_X1 U6803 ( .A1(n7124), .A2(n8546), .ZN(n5258) );
  NAND2_X1 U6804 ( .A1(n8829), .A2(n8774), .ZN(n8195) );
  INV_X1 U6805 ( .A(n8774), .ZN(n8463) );
  NAND2_X1 U6806 ( .A1(n8829), .A2(n8463), .ZN(n5263) );
  XNOR2_X1 U6807 ( .A(n5265), .B(n5264), .ZN(n6867) );
  NAND2_X1 U6808 ( .A1(n6867), .A2(n8252), .ZN(n5269) );
  NAND2_X1 U6809 ( .A1(n5266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5267) );
  XNOR2_X1 U6810 ( .A(n5267), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8596) );
  AOI22_X1 U6811 ( .A1(n5299), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6382), .B2(
        n8596), .ZN(n5268) );
  NAND2_X1 U6812 ( .A1(n7119), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5276) );
  INV_X1 U6813 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8824) );
  OR2_X1 U6814 ( .A1(n7121), .A2(n8824), .ZN(n5275) );
  NAND2_X1 U6815 ( .A1(n5270), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6816 ( .A1(n5287), .A2(n5271), .ZN(n8782) );
  OR2_X1 U6817 ( .A1(n5039), .A2(n8782), .ZN(n5274) );
  INV_X1 U6818 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8781) );
  OR2_X1 U6819 ( .A1(n5272), .A2(n8781), .ZN(n5273) );
  NAND2_X1 U6820 ( .A1(n8891), .A2(n8391), .ZN(n8191) );
  NAND2_X1 U6821 ( .A1(n8203), .A2(n8191), .ZN(n8771) );
  INV_X1 U6822 ( .A(n8891), .ZN(n5277) );
  XNOR2_X1 U6823 ( .A(n5279), .B(n5278), .ZN(n6923) );
  NAND2_X1 U6824 ( .A1(n6923), .A2(n8252), .ZN(n5286) );
  INV_X1 U6825 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5280) );
  NAND3_X1 U6826 ( .A1(n5281), .A2(n9019), .A3(n5280), .ZN(n5282) );
  NAND2_X1 U6827 ( .A1(n4363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5284) );
  XNOR2_X1 U6828 ( .A(n5284), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8613) );
  AOI22_X1 U6829 ( .A1(n5299), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6382), .B2(
        n8613), .ZN(n5285) );
  NAND2_X1 U6830 ( .A1(n5287), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6831 ( .A1(n5304), .A2(n5288), .ZN(n8755) );
  NAND2_X1 U6832 ( .A1(n5464), .A2(n8755), .ZN(n5293) );
  INV_X1 U6833 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5289) );
  OR2_X1 U6834 ( .A1(n5038), .A2(n5289), .ZN(n5292) );
  INV_X1 U6835 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8579) );
  OR2_X1 U6836 ( .A1(n7121), .A2(n8579), .ZN(n5291) );
  INV_X1 U6837 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8758) );
  OR2_X1 U6838 ( .A1(n7124), .A2(n8758), .ZN(n5290) );
  NAND2_X1 U6839 ( .A1(n8823), .A2(n8776), .ZN(n5295) );
  INV_X1 U6840 ( .A(n8776), .ZN(n8462) );
  XNOR2_X1 U6841 ( .A(n5297), .B(n5296), .ZN(n7130) );
  NAND2_X1 U6842 ( .A1(n7130), .A2(n8252), .ZN(n5301) );
  INV_X1 U6843 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5470) );
  AOI22_X1 U6844 ( .A1(n5299), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8622), .B2(
        n6382), .ZN(n5300) );
  INV_X1 U6845 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8884) );
  OR2_X1 U6846 ( .A1(n5038), .A2(n8884), .ZN(n5303) );
  INV_X1 U6847 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8818) );
  OR2_X1 U6848 ( .A1(n7121), .A2(n8818), .ZN(n5302) );
  AND2_X1 U6849 ( .A1(n5303), .A2(n5302), .ZN(n5309) );
  NAND2_X1 U6850 ( .A1(n5304), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6851 ( .A1(n5306), .A2(n5305), .ZN(n8744) );
  NAND2_X1 U6852 ( .A1(n8744), .A2(n5464), .ZN(n5308) );
  INV_X1 U6853 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8999) );
  OR2_X1 U6854 ( .A1(n7124), .A2(n8999), .ZN(n5307) );
  NAND2_X1 U6855 ( .A1(n8817), .A2(n8729), .ZN(n8212) );
  INV_X1 U6856 ( .A(n8817), .ZN(n8367) );
  NAND2_X1 U6857 ( .A1(n8734), .A2(n8740), .ZN(n8713) );
  INV_X1 U6858 ( .A(n5310), .ZN(n5311) );
  INV_X1 U6859 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7348) );
  INV_X1 U6860 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7347) );
  MUX2_X1 U6861 ( .A(n7348), .B(n7347), .S(n6389), .Z(n5326) );
  XNOR2_X1 U6862 ( .A(n5326), .B(SI_21_), .ZN(n5316) );
  XNOR2_X1 U6863 ( .A(n5330), .B(n5316), .ZN(n7346) );
  NAND2_X1 U6864 ( .A1(n7346), .A2(n8252), .ZN(n5318) );
  OR2_X1 U6865 ( .A1(n8253), .A2(n7348), .ZN(n5317) );
  INV_X1 U6866 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6867 ( .A1(n5321), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6868 ( .A1(n5337), .A2(n5322), .ZN(n8722) );
  NAND2_X1 U6869 ( .A1(n8722), .A2(n5464), .ZN(n5325) );
  AOI22_X1 U6870 ( .A1(n5500), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n7119), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6871 ( .A1(n5501), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6872 ( .A1(n8873), .A2(n8730), .ZN(n8220) );
  INV_X1 U6873 ( .A(n8730), .ZN(n8706) );
  INV_X1 U6874 ( .A(n5326), .ZN(n5327) );
  NOR2_X1 U6875 ( .A1(n5327), .A2(SI_21_), .ZN(n5329) );
  NAND2_X1 U6876 ( .A1(n5327), .A2(SI_21_), .ZN(n5328) );
  INV_X1 U6877 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7415) );
  INV_X1 U6878 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U6879 ( .A(n7415), .B(n7745), .S(n6389), .Z(n5332) );
  INV_X1 U6880 ( .A(SI_22_), .ZN(n5331) );
  NAND2_X1 U6881 ( .A1(n5332), .A2(n5331), .ZN(n5345) );
  INV_X1 U6882 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6883 ( .A1(n5333), .A2(SI_22_), .ZN(n5334) );
  NAND2_X1 U6884 ( .A1(n5345), .A2(n5334), .ZN(n5346) );
  XNOR2_X1 U6885 ( .A(n5347), .B(n5346), .ZN(n7414) );
  NAND2_X1 U6886 ( .A1(n7414), .A2(n8252), .ZN(n5336) );
  OR2_X1 U6887 ( .A1(n8253), .A2(n7415), .ZN(n5335) );
  NAND2_X1 U6888 ( .A1(n5337), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6889 ( .A1(n5353), .A2(n5338), .ZN(n8710) );
  NAND2_X1 U6890 ( .A1(n8710), .A2(n5464), .ZN(n5343) );
  INV_X1 U6891 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U6892 ( .A1(n5500), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6893 ( .A1(n7119), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5339) );
  OAI211_X1 U6894 ( .C1(n8709), .C2(n7124), .A(n5340), .B(n5339), .ZN(n5341)
         );
  INV_X1 U6895 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6896 ( .A1(n8867), .A2(n8692), .ZN(n8225) );
  INV_X1 U6897 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7466) );
  INV_X1 U6898 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7470) );
  MUX2_X1 U6899 ( .A(n7466), .B(n7470), .S(n6357), .Z(n5349) );
  INV_X1 U6900 ( .A(SI_23_), .ZN(n5348) );
  NAND2_X1 U6901 ( .A1(n5349), .A2(n5348), .ZN(n5365) );
  INV_X1 U6902 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6903 ( .A1(n5350), .A2(SI_23_), .ZN(n5351) );
  NOR2_X1 U6904 ( .A1(n8253), .A2(n7466), .ZN(n5352) );
  NAND2_X1 U6905 ( .A1(n5353), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6906 ( .A1(n5373), .A2(n5354), .ZN(n8696) );
  NAND2_X1 U6907 ( .A1(n8696), .A2(n5464), .ZN(n5359) );
  INV_X1 U6908 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U6909 ( .A1(n7119), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6910 ( .A1(n5500), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5355) );
  OAI211_X1 U6911 ( .C1(n8695), .C2(n7124), .A(n5356), .B(n5355), .ZN(n5357)
         );
  INV_X1 U6912 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6913 ( .A1(n5360), .A2(n8707), .ZN(n5361) );
  NAND2_X1 U6914 ( .A1(n8690), .A2(n5361), .ZN(n5362) );
  NAND2_X1 U6915 ( .A1(n5362), .A2(n4331), .ZN(n8677) );
  NAND2_X1 U6916 ( .A1(n5366), .A2(n5365), .ZN(n5381) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7773) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7554) );
  MUX2_X1 U6919 ( .A(n7773), .B(n7554), .S(n6389), .Z(n5368) );
  INV_X1 U6920 ( .A(SI_24_), .ZN(n5367) );
  NAND2_X1 U6921 ( .A1(n5368), .A2(n5367), .ZN(n5382) );
  INV_X1 U6922 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6923 ( .A1(n5369), .A2(SI_24_), .ZN(n5370) );
  AND2_X1 U6924 ( .A1(n5382), .A2(n5370), .ZN(n5380) );
  NOR2_X1 U6925 ( .A1(n8253), .A2(n7773), .ZN(n5371) );
  INV_X1 U6926 ( .A(n5373), .ZN(n5372) );
  INV_X1 U6927 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U6928 ( .A1(n5373), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6929 ( .A1(n5392), .A2(n5374), .ZN(n8685) );
  NAND2_X1 U6930 ( .A1(n8685), .A2(n5464), .ZN(n5379) );
  INV_X1 U6931 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U6932 ( .A1(n5501), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6933 ( .A1(n5500), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5375) );
  OAI211_X1 U6934 ( .C1(n5038), .C2(n8992), .A(n5376), .B(n5375), .ZN(n5377)
         );
  INV_X1 U6935 ( .A(n5377), .ZN(n5378) );
  NAND2_X1 U6936 ( .A1(n5381), .A2(n5380), .ZN(n5383) );
  NAND2_X1 U6937 ( .A1(n5383), .A2(n5382), .ZN(n5401) );
  INV_X1 U6938 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7655) );
  INV_X1 U6939 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9060) );
  MUX2_X1 U6940 ( .A(n7655), .B(n9060), .S(n6357), .Z(n5385) );
  INV_X1 U6941 ( .A(SI_25_), .ZN(n5384) );
  NAND2_X1 U6942 ( .A1(n5385), .A2(n5384), .ZN(n5402) );
  INV_X1 U6943 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6944 ( .A1(n5386), .A2(SI_25_), .ZN(n5387) );
  OR2_X1 U6945 ( .A1(n8253), .A2(n7655), .ZN(n5388) );
  INV_X1 U6946 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6947 ( .A1(n5392), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6948 ( .A1(n5410), .A2(n5393), .ZN(n8667) );
  NAND2_X1 U6949 ( .A1(n8667), .A2(n5464), .ZN(n5398) );
  INV_X1 U6950 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U6951 ( .A1(n7119), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6952 ( .A1(n5500), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5394) );
  OAI211_X1 U6953 ( .C1(n7124), .C2(n8671), .A(n5395), .B(n5394), .ZN(n5396)
         );
  INV_X1 U6954 ( .A(n5396), .ZN(n5397) );
  NAND2_X1 U6955 ( .A1(n5401), .A2(n5400), .ZN(n5403) );
  NAND2_X1 U6956 ( .A1(n5403), .A2(n5402), .ZN(n5420) );
  INV_X1 U6957 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7683) );
  INV_X1 U6958 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7681) );
  MUX2_X1 U6959 ( .A(n7683), .B(n7681), .S(n6357), .Z(n5405) );
  INV_X1 U6960 ( .A(SI_26_), .ZN(n5404) );
  NAND2_X1 U6961 ( .A1(n5405), .A2(n5404), .ZN(n5421) );
  INV_X1 U6962 ( .A(n5405), .ZN(n5406) );
  NAND2_X1 U6963 ( .A1(n5406), .A2(SI_26_), .ZN(n5407) );
  OR2_X1 U6964 ( .A1(n8253), .A2(n7683), .ZN(n5408) );
  NAND2_X1 U6965 ( .A1(n5410), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6966 ( .A1(n5431), .A2(n5411), .ZN(n8659) );
  NAND2_X1 U6967 ( .A1(n8659), .A2(n5464), .ZN(n5416) );
  INV_X1 U6968 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U6969 ( .A1(n5501), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6970 ( .A1(n7119), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5412) );
  OAI211_X1 U6971 ( .C1(n7121), .C2(n8972), .A(n5413), .B(n5412), .ZN(n5414)
         );
  INV_X1 U6972 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U6973 ( .A1(n8845), .A2(n8664), .ZN(n5418) );
  INV_X1 U6974 ( .A(n8845), .ZN(n5417) );
  NAND2_X1 U6975 ( .A1(n5420), .A2(n5419), .ZN(n5422) );
  INV_X1 U6976 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7701) );
  INV_X1 U6977 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7732) );
  MUX2_X1 U6978 ( .A(n7701), .B(n7732), .S(n6357), .Z(n5424) );
  INV_X1 U6979 ( .A(SI_27_), .ZN(n5423) );
  NAND2_X1 U6980 ( .A1(n5424), .A2(n5423), .ZN(n5444) );
  INV_X1 U6981 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6982 ( .A1(n5425), .A2(SI_27_), .ZN(n5426) );
  AND2_X1 U6983 ( .A1(n5444), .A2(n5426), .ZN(n5442) );
  NAND2_X1 U6984 ( .A1(n7700), .A2(n8252), .ZN(n5428) );
  OR2_X1 U6985 ( .A1(n8253), .A2(n7701), .ZN(n5427) );
  INV_X1 U6986 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6987 ( .A1(n5431), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6988 ( .A1(n5447), .A2(n5432), .ZN(n8347) );
  NAND2_X1 U6989 ( .A1(n8347), .A2(n5464), .ZN(n5437) );
  INV_X1 U6990 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U6991 ( .A1(n7119), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6992 ( .A1(n5500), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5433) );
  OAI211_X1 U6993 ( .C1(n9002), .C2(n7124), .A(n5434), .B(n5433), .ZN(n5435)
         );
  INV_X1 U6994 ( .A(n5435), .ZN(n5436) );
  NAND2_X1 U6995 ( .A1(n5438), .A2(n8454), .ZN(n5439) );
  NAND2_X1 U6996 ( .A1(n8642), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U6997 ( .A1(n8792), .A2(n8656), .ZN(n5440) );
  NAND2_X1 U6998 ( .A1(n5441), .A2(n5440), .ZN(n6043) );
  INV_X1 U6999 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7746) );
  INV_X1 U7000 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7730) );
  MUX2_X1 U7001 ( .A(n7746), .B(n7730), .S(n6389), .Z(n5458) );
  XNOR2_X1 U7002 ( .A(n5458), .B(SI_28_), .ZN(n5455) );
  NAND2_X1 U7003 ( .A1(n7729), .A2(n8252), .ZN(n5446) );
  OR2_X1 U7004 ( .A1(n8253), .A2(n7746), .ZN(n5445) );
  NAND2_X1 U7005 ( .A1(n5447), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7006 ( .A1(n5463), .A2(n5448), .ZN(n8635) );
  NAND2_X1 U7007 ( .A1(n8635), .A2(n5464), .ZN(n5453) );
  INV_X1 U7008 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U7009 ( .A1(n5500), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U7010 ( .A1(n5501), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U7011 ( .C1(n5038), .C2(n9022), .A(n5450), .B(n5449), .ZN(n5451)
         );
  INV_X1 U7012 ( .A(n5451), .ZN(n5452) );
  NOR2_X1 U7013 ( .A1(n8249), .A2(n8643), .ZN(n5454) );
  OAI22_X1 U7014 ( .A1(n6043), .A2(n5454), .B1(n8636), .B2(n8461), .ZN(n5469)
         );
  INV_X1 U7015 ( .A(SI_28_), .ZN(n5457) );
  NAND2_X1 U7016 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  INV_X1 U7017 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8341) );
  INV_X1 U7018 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U7019 ( .A(n8341), .B(n9798), .S(n6389), .Z(n6337) );
  NAND2_X1 U7020 ( .A1(n8340), .A2(n8252), .ZN(n5462) );
  OR2_X1 U7021 ( .A1(n8253), .A2(n8341), .ZN(n5461) );
  NAND2_X1 U7022 ( .A1(n8332), .A2(n5464), .ZN(n7128) );
  INV_X1 U7023 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U7024 ( .A1(n7119), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7025 ( .A1(n5500), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U7026 ( .C1(n7124), .C2(n8333), .A(n5466), .B(n5465), .ZN(n5467)
         );
  INV_X1 U7027 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U7028 ( .A1(n8337), .A2(n8097), .ZN(n8261) );
  XNOR2_X1 U7029 ( .A(n5469), .B(n8247), .ZN(n5509) );
  NAND2_X1 U7030 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7031 ( .A1(n5475), .A2(n5474), .ZN(n5477) );
  OR2_X1 U7032 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U7033 ( .A1(n5477), .A2(n5476), .ZN(n5511) );
  INV_X1 U7034 ( .A(n5511), .ZN(n5496) );
  NAND2_X1 U7035 ( .A1(n6643), .A2(n5496), .ZN(n8314) );
  NAND2_X1 U7036 ( .A1(n5478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U7037 ( .A(n5479), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U7038 ( .A1(n8622), .A2(n8322), .ZN(n6055) );
  INV_X1 U7039 ( .A(n7760), .ZN(n7772) );
  INV_X1 U7040 ( .A(n7062), .ZN(n10071) );
  OR2_X1 U7041 ( .A1(n8475), .A2(n10071), .ZN(n8136) );
  NAND2_X1 U7042 ( .A1(n8475), .A2(n10071), .ZN(n8121) );
  NAND2_X1 U7043 ( .A1(n7064), .A2(n8278), .ZN(n5480) );
  NAND2_X1 U7044 ( .A1(n5480), .A2(n8136), .ZN(n6906) );
  INV_X1 U7045 ( .A(n8283), .ZN(n8120) );
  NAND2_X1 U7046 ( .A1(n6906), .A2(n8120), .ZN(n6907) );
  OR2_X1 U7047 ( .A1(n5481), .A2(n10076), .ZN(n8122) );
  NAND2_X1 U7048 ( .A1(n6907), .A2(n8122), .ZN(n6974) );
  INV_X1 U7049 ( .A(n10081), .ZN(n6973) );
  NAND2_X1 U7050 ( .A1(n8474), .A2(n6973), .ZN(n8137) );
  NAND2_X1 U7051 ( .A1(n6974), .A2(n8137), .ZN(n6897) );
  OR2_X1 U7052 ( .A1(n8474), .A2(n6973), .ZN(n8123) );
  INV_X1 U7053 ( .A(n6903), .ZN(n10088) );
  OR2_X1 U7054 ( .A1(n8473), .A2(n10088), .ZN(n8127) );
  AND2_X1 U7055 ( .A1(n8123), .A2(n8127), .ZN(n8141) );
  NAND2_X1 U7056 ( .A1(n6897), .A2(n8141), .ZN(n5482) );
  NAND2_X1 U7057 ( .A1(n8473), .A2(n10088), .ZN(n8143) );
  INV_X1 U7058 ( .A(n7244), .ZN(n10098) );
  NAND2_X1 U7059 ( .A1(n10098), .A2(n8471), .ZN(n8126) );
  INV_X1 U7060 ( .A(n8471), .ZN(n7318) );
  NAND2_X1 U7061 ( .A1(n7318), .A2(n7244), .ZN(n8146) );
  INV_X1 U7062 ( .A(n7192), .ZN(n5485) );
  NAND2_X1 U7063 ( .A1(n8130), .A2(n8152), .ZN(n8285) );
  NAND2_X1 U7064 ( .A1(n5485), .A2(n5484), .ZN(n7191) );
  INV_X1 U7065 ( .A(n7532), .ZN(n10109) );
  AND2_X1 U7066 ( .A1(n10109), .A2(n8469), .ZN(n8156) );
  INV_X1 U7067 ( .A(n8469), .ZN(n7530) );
  NAND2_X1 U7068 ( .A1(n7532), .A2(n7530), .ZN(n8151) );
  AND2_X1 U7069 ( .A1(n8157), .A2(n8151), .ZN(n8161) );
  NAND2_X1 U7070 ( .A1(n5487), .A2(n8159), .ZN(n7430) );
  XNOR2_X1 U7071 ( .A(n8169), .B(n8467), .ZN(n8293) );
  NAND2_X1 U7072 ( .A1(n7430), .A2(n8293), .ZN(n7432) );
  INV_X1 U7073 ( .A(n8467), .ZN(n8168) );
  OR2_X1 U7074 ( .A1(n8169), .A2(n8168), .ZN(n8171) );
  NAND2_X1 U7075 ( .A1(n7432), .A2(n8171), .ZN(n7455) );
  INV_X1 U7076 ( .A(n8466), .ZN(n7583) );
  NAND2_X1 U7077 ( .A1(n8174), .A2(n7583), .ZN(n5488) );
  NAND2_X1 U7078 ( .A1(n7455), .A2(n5488), .ZN(n5490) );
  OR2_X1 U7079 ( .A1(n8174), .A2(n7583), .ZN(n5489) );
  NOR2_X1 U7080 ( .A1(n7677), .A2(n7694), .ZN(n8183) );
  NAND2_X1 U7081 ( .A1(n7677), .A2(n7694), .ZN(n7613) );
  NAND2_X1 U7082 ( .A1(n7610), .A2(n8275), .ZN(n7609) );
  NAND2_X1 U7083 ( .A1(n7609), .A2(n8195), .ZN(n8768) );
  NAND2_X1 U7084 ( .A1(n8760), .A2(n8776), .ZN(n8205) );
  NAND2_X1 U7085 ( .A1(n8204), .A2(n8205), .ZN(n8763) );
  AND2_X1 U7086 ( .A1(n8220), .A2(n8713), .ZN(n8215) );
  NAND2_X1 U7087 ( .A1(n5491), .A2(n8219), .ZN(n8702) );
  AND2_X1 U7088 ( .A1(n8861), .A2(n8707), .ZN(n8274) );
  NAND2_X1 U7089 ( .A1(n8856), .A2(n8693), .ZN(n8272) );
  NAND2_X1 U7090 ( .A1(n5360), .A2(n8430), .ZN(n8674) );
  AND2_X1 U7091 ( .A1(n8683), .A2(n8665), .ZN(n8271) );
  NAND2_X1 U7092 ( .A1(n5492), .A2(n8242), .ZN(n6050) );
  NAND2_X1 U7093 ( .A1(n8636), .A2(n8643), .ZN(n5493) );
  NAND2_X1 U7094 ( .A1(n6050), .A2(n5493), .ZN(n5495) );
  NAND2_X2 U7095 ( .A1(n6643), .A2(n8322), .ZN(n8256) );
  AND2_X1 U7096 ( .A1(n5511), .A2(n8609), .ZN(n5537) );
  INV_X1 U7097 ( .A(n5537), .ZN(n5497) );
  OR2_X1 U7098 ( .A1(n8256), .A2(n5497), .ZN(n6659) );
  INV_X1 U7099 ( .A(n8322), .ZN(n7416) );
  NAND2_X1 U7100 ( .A1(n6659), .A2(n10108), .ZN(n7764) );
  NAND2_X1 U7101 ( .A1(n8609), .A2(n8322), .ZN(n5514) );
  AND2_X1 U7102 ( .A1(n5497), .A2(n5514), .ZN(n5498) );
  INV_X1 U7103 ( .A(n7748), .ZN(n8319) );
  NAND2_X1 U7104 ( .A1(n8319), .A2(n8610), .ZN(n5499) );
  AND2_X1 U7105 ( .A1(n5506), .A2(n5499), .ZN(n6662) );
  INV_X1 U7106 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U7107 ( .A1(n5500), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7108 ( .A1(n5501), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5502) );
  OAI211_X1 U7109 ( .C1(n5038), .C2(n9021), .A(n5503), .B(n5502), .ZN(n5504)
         );
  INV_X1 U7110 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U7111 ( .A1(n7128), .A2(n5505), .ZN(n8460) );
  AND2_X1 U7112 ( .A1(n5506), .A2(P2_B_REG_SCAN_IN), .ZN(n5507) );
  NOR2_X1 U7113 ( .A1(n8775), .A2(n5507), .ZN(n8626) );
  AOI22_X1 U7114 ( .A1(n8750), .A2(n8461), .B1(n8460), .B2(n8626), .ZN(n5508)
         );
  INV_X1 U7115 ( .A(n6644), .ZN(n6774) );
  INV_X1 U7116 ( .A(n10082), .ZN(n10102) );
  OR2_X1 U7117 ( .A1(n5511), .A2(n5514), .ZN(n5515) );
  NAND2_X1 U7118 ( .A1(n8256), .A2(n5515), .ZN(n6769) );
  NAND2_X1 U7119 ( .A1(n5516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5552) );
  INV_X1 U7120 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7121 ( .A1(n5552), .A2(n5551), .ZN(n5517) );
  NAND2_X1 U7122 ( .A1(n5517), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5519) );
  INV_X1 U7123 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U7124 ( .A1(n5519), .A2(n5518), .ZN(n5521) );
  OR2_X1 U7125 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U7126 ( .A1(n5521), .A2(n5520), .ZN(n7775) );
  XNOR2_X1 U7127 ( .A(n7775), .B(P2_B_REG_SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7128 ( .A1(n5521), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5523) );
  INV_X1 U7129 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5522) );
  XNOR2_X1 U7130 ( .A(n5523), .B(n5522), .ZN(n7657) );
  NAND2_X1 U7131 ( .A1(n5524), .A2(n7657), .ZN(n5534) );
  NAND2_X1 U7132 ( .A1(n4975), .A2(n5525), .ZN(n5526) );
  NAND2_X1 U7133 ( .A1(n5526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5527) );
  MUX2_X1 U7134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5527), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5528) );
  AND2_X1 U7135 ( .A1(n5529), .A2(n5528), .ZN(n5531) );
  NAND2_X1 U7136 ( .A1(n5534), .A2(n5531), .ZN(n6402) );
  OR2_X1 U7137 ( .A1(n6402), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5530) );
  INV_X1 U7138 ( .A(n5531), .ZN(n7685) );
  NAND2_X1 U7139 ( .A1(n7657), .A2(n7685), .ZN(n6428) );
  NAND2_X1 U7140 ( .A1(n5530), .A2(n6428), .ZN(n6767) );
  NAND2_X1 U7141 ( .A1(n6769), .A2(n6767), .ZN(n5536) );
  INV_X1 U7142 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5532) );
  AND2_X1 U7143 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U7144 ( .A1(n5534), .A2(n5533), .ZN(n5535) );
  NAND2_X1 U7145 ( .A1(n7775), .A2(n7685), .ZN(n6431) );
  NAND2_X1 U7146 ( .A1(n5535), .A2(n6431), .ZN(n5553) );
  OR2_X1 U7147 ( .A1(n6767), .A2(n5553), .ZN(n6631) );
  AND2_X1 U7148 ( .A1(n5536), .A2(n6631), .ZN(n5557) );
  OR2_X1 U7149 ( .A1(n8256), .A2(n5537), .ZN(n6634) );
  NOR2_X1 U7150 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5541) );
  NOR4_X1 U7151 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5540) );
  NOR4_X1 U7152 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5539) );
  NOR4_X1 U7153 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5538) );
  NAND4_X1 U7154 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n5547)
         );
  NOR4_X1 U7155 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5545) );
  NOR4_X1 U7156 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5544) );
  NOR4_X1 U7157 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5543) );
  NOR4_X1 U7158 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5542) );
  NAND4_X1 U7159 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n5546)
         );
  NOR2_X1 U7160 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  OR2_X1 U7161 ( .A1(n6402), .A2(n5548), .ZN(n6054) );
  INV_X1 U7162 ( .A(n7657), .ZN(n5550) );
  NOR2_X1 U7163 ( .A1(n7775), .A2(n7685), .ZN(n5549) );
  NAND2_X1 U7164 ( .A1(n5550), .A2(n5549), .ZN(n6636) );
  XNOR2_X1 U7165 ( .A(n5552), .B(n5551), .ZN(n6642) );
  AND2_X1 U7166 ( .A1(n6054), .A2(n6403), .ZN(n6056) );
  NAND2_X1 U7167 ( .A1(n10082), .A2(n8277), .ZN(n6667) );
  INV_X1 U7168 ( .A(n5553), .ZN(n6646) );
  NAND2_X1 U7169 ( .A1(n6667), .A2(n6646), .ZN(n5555) );
  INV_X1 U7170 ( .A(n6769), .ZN(n5554) );
  NAND2_X1 U7171 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  AND3_X2 U7172 ( .A1(n5557), .A2(n6773), .A3(n5556), .ZN(n10135) );
  NAND2_X1 U7173 ( .A1(n6377), .A2(n10135), .ZN(n5560) );
  INV_X1 U7174 ( .A(n8337), .ZN(n6378) );
  NAND2_X1 U7175 ( .A1(n10135), .A2(n10118), .ZN(n8813) );
  NOR2_X1 U7176 ( .A1(n6378), .A2(n8813), .ZN(n5558) );
  NAND2_X1 U7177 ( .A1(n5560), .A2(n5559), .ZN(P2_U3488) );
  NAND3_X1 U7178 ( .A1(n5567), .A2(n5566), .A3(n5652), .ZN(n5768) );
  NOR3_X1 U7179 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n5570) );
  INV_X1 U7180 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5571) );
  NOR2_X1 U7181 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5587) );
  AND2_X1 U7182 ( .A1(n5587), .A2(n5573), .ZN(n5574) );
  NAND2_X1 U7183 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7184 ( .A1(n5578), .A2(n5577), .ZN(n5625) );
  NAND2_X1 U7185 ( .A1(n5614), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7186 ( .A1(n5645), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5582) );
  INV_X1 U7187 ( .A(n5578), .ZN(n8327) );
  NAND2_X1 U7188 ( .A1(n5635), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7189 ( .A1(n5658), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5580) );
  INV_X1 U7190 ( .A(n9286), .ZN(n6812) );
  NAND2_X1 U7191 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5584) );
  NOR2_X1 U7192 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  NAND2_X1 U7193 ( .A1(n5834), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5602) );
  OR2_X1 U7194 ( .A1(n5703), .A2(n6395), .ZN(n5600) );
  INV_X1 U7195 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9791) );
  OR2_X1 U7196 ( .A1(n5595), .A2(n9791), .ZN(n5597) );
  XNOR2_X1 U7197 ( .A(n5597), .B(n5596), .ZN(n6538) );
  NAND2_X1 U7198 ( .A1(n6812), .A2(n6842), .ZN(n5994) );
  INV_X1 U7199 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7200 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5603) );
  XNOR2_X1 U7201 ( .A(n5604), .B(n5603), .ZN(n9289) );
  OAI22_X1 U7202 ( .A1(n5605), .A2(n6387), .B1(n6416), .B2(n9289), .ZN(n5606)
         );
  INV_X1 U7203 ( .A(n5606), .ZN(n5608) );
  NAND2_X1 U7204 ( .A1(n5609), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7205 ( .A1(n5635), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7206 ( .A1(n5645), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7207 ( .A1(n5614), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7208 ( .A1(n5635), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7209 ( .A1(n5658), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5615) );
  INV_X1 U7210 ( .A(SI_0_), .ZN(n5619) );
  NOR2_X1 U7211 ( .A1(n6388), .A2(n5619), .ZN(n5621) );
  INV_X1 U7212 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U7213 ( .A(n5621), .B(n5620), .ZN(n9801) );
  INV_X1 U7214 ( .A(n7024), .ZN(n9976) );
  NAND2_X1 U7215 ( .A1(n5992), .A2(n6085), .ZN(n5622) );
  NAND2_X1 U7216 ( .A1(n9286), .A2(n5949), .ZN(n7995) );
  INV_X1 U7217 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7218 ( .A1(n5645), .A2(n5624), .ZN(n5629) );
  NAND2_X1 U7219 ( .A1(n5609), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7220 ( .A1(n5635), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7221 ( .A1(n5658), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5626) );
  OR2_X1 U7222 ( .A1(n5652), .A2(n9791), .ZN(n5631) );
  NAND2_X1 U7223 ( .A1(n5631), .A2(n5630), .ZN(n5640) );
  OAI21_X1 U7224 ( .B1(n5631), .B2(n5630), .A(n5640), .ZN(n9313) );
  OR2_X1 U7225 ( .A1(n5703), .A2(n6397), .ZN(n5632) );
  OAI211_X1 U7226 ( .C1(n6416), .C2(n9313), .A(n5633), .B(n5632), .ZN(n6814)
         );
  NAND2_X1 U7227 ( .A1(n9285), .A2(n5950), .ZN(n7854) );
  NAND2_X1 U7228 ( .A1(n5682), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7229 ( .A1(n5609), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5638) );
  INV_X1 U7230 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5634) );
  XNOR2_X1 U7231 ( .A(n5634), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U7232 ( .A1(n5645), .A2(n6963), .ZN(n5637) );
  NAND2_X1 U7233 ( .A1(n5696), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5636) );
  NAND4_X1 U7234 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(n9284)
         );
  NAND2_X1 U7235 ( .A1(n5640), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5642) );
  INV_X1 U7236 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5641) );
  XNOR2_X1 U7237 ( .A(n5642), .B(n5641), .ZN(n6518) );
  OR2_X1 U7238 ( .A1(n5703), .A2(n6391), .ZN(n5644) );
  OR2_X1 U7239 ( .A1(n5605), .A2(n6386), .ZN(n5643) );
  OAI211_X1 U7240 ( .C1(n6416), .C2(n6518), .A(n5644), .B(n5643), .ZN(n6874)
         );
  NAND2_X1 U7241 ( .A1(n9284), .A2(n6965), .ZN(n7855) );
  INV_X1 U7242 ( .A(n9284), .ZN(n6813) );
  NAND2_X1 U7243 ( .A1(n5682), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7244 ( .A1(n5614), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5649) );
  AOI21_X1 U7245 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5646) );
  NOR2_X1 U7246 ( .A1(n5646), .A2(n5693), .ZN(n9160) );
  NAND2_X1 U7247 ( .A1(n5645), .A2(n9160), .ZN(n5648) );
  NAND2_X1 U7248 ( .A1(n5696), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5647) );
  NAND4_X1 U7249 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n9283)
         );
  INV_X1 U7250 ( .A(n9283), .ZN(n6871) );
  NOR2_X1 U7251 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5651) );
  NAND2_X1 U7252 ( .A1(n5652), .A2(n5651), .ZN(n5664) );
  NAND2_X1 U7253 ( .A1(n5664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5654) );
  INV_X1 U7254 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5653) );
  XNOR2_X1 U7255 ( .A(n5654), .B(n5653), .ZN(n9866) );
  OR2_X1 U7256 ( .A1(n5703), .A2(n6393), .ZN(n5656) );
  OR2_X1 U7257 ( .A1(n5605), .A2(n9027), .ZN(n5655) );
  OAI211_X1 U7258 ( .C1(n6416), .C2(n9866), .A(n5656), .B(n5655), .ZN(n9159)
         );
  NAND2_X1 U7259 ( .A1(n6871), .A2(n9159), .ZN(n7851) );
  INV_X1 U7260 ( .A(n9159), .ZN(n10008) );
  NAND2_X1 U7261 ( .A1(n9283), .A2(n10008), .ZN(n7856) );
  NAND2_X1 U7262 ( .A1(n7851), .A2(n7856), .ZN(n7088) );
  INV_X1 U7263 ( .A(n7088), .ZN(n7807) );
  NAND2_X1 U7264 ( .A1(n7092), .A2(n7807), .ZN(n5657) );
  NAND2_X1 U7265 ( .A1(n5657), .A2(n7851), .ZN(n7050) );
  NAND2_X1 U7266 ( .A1(n5682), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7267 ( .A1(n5614), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7268 ( .A1(n5677), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5717) );
  OR2_X1 U7269 ( .A1(n5677), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5659) );
  AND2_X1 U7270 ( .A1(n5717), .A2(n5659), .ZN(n7390) );
  NAND2_X1 U7271 ( .A1(n5645), .A2(n7390), .ZN(n5661) );
  NAND2_X1 U7272 ( .A1(n5696), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5660) );
  NAND4_X1 U7273 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n9279)
         );
  INV_X1 U7274 ( .A(n9279), .ZN(n5691) );
  NAND2_X1 U7275 ( .A1(n6418), .A2(n6345), .ZN(n5668) );
  NOR2_X1 U7276 ( .A1(n5664), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5701) );
  INV_X1 U7277 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7278 ( .A1(n5701), .A2(n5665), .ZN(n5669) );
  NAND2_X1 U7279 ( .A1(n5710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U7280 ( .A(n5666), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6456) );
  AOI22_X1 U7281 ( .A1(n5834), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5833), .B2(
        n6456), .ZN(n5667) );
  NOR2_X1 U7282 ( .A1(n5691), .A2(n9959), .ZN(n7875) );
  INV_X1 U7283 ( .A(n7875), .ZN(n5706) );
  NAND2_X1 U7284 ( .A1(n5669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5688) );
  INV_X1 U7285 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U7286 ( .A1(n5688), .A2(n5670), .ZN(n5671) );
  NAND2_X1 U7287 ( .A1(n5671), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U7288 ( .A(n5672), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9819) );
  INV_X1 U7289 ( .A(n9819), .ZN(n6457) );
  NAND2_X1 U7290 ( .A1(n6408), .A2(n6345), .ZN(n5674) );
  OR2_X1 U7291 ( .A1(n5605), .A2(n6409), .ZN(n5673) );
  NAND2_X1 U7292 ( .A1(n5609), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7293 ( .A1(n5696), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5680) );
  AND2_X1 U7294 ( .A1(n5683), .A2(n5675), .ZN(n5676) );
  NOR2_X1 U7295 ( .A1(n5677), .A2(n5676), .ZN(n7254) );
  NAND2_X1 U7296 ( .A1(n5645), .A2(n7254), .ZN(n5679) );
  NAND2_X1 U7297 ( .A1(n5658), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U7298 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n9280)
         );
  NAND2_X1 U7299 ( .A1(n7257), .A2(n9280), .ZN(n9951) );
  AND2_X1 U7300 ( .A1(n5706), .A2(n9951), .ZN(n7869) );
  NAND2_X1 U7301 ( .A1(n9957), .A2(n7336), .ZN(n7865) );
  NAND2_X1 U7302 ( .A1(n5682), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7303 ( .A1(n5614), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5686) );
  OAI21_X1 U7304 ( .B1(n5695), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5683), .ZN(
        n7164) );
  INV_X1 U7305 ( .A(n7164), .ZN(n7229) );
  NAND2_X1 U7306 ( .A1(n5645), .A2(n7229), .ZN(n5685) );
  NAND2_X1 U7307 ( .A1(n5696), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U7308 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n9281)
         );
  INV_X1 U7309 ( .A(n9281), .ZN(n6001) );
  XNOR2_X1 U7310 ( .A(n5688), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9808) );
  INV_X1 U7311 ( .A(n9808), .ZN(n6470) );
  NAND2_X1 U7312 ( .A1(n6345), .A2(n6404), .ZN(n5690) );
  INV_X1 U7313 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6405) );
  OR2_X1 U7314 ( .A1(n5605), .A2(n6405), .ZN(n5689) );
  OAI211_X1 U7315 ( .C1(n6416), .C2(n6470), .A(n5690), .B(n5689), .ZN(n7167)
         );
  NAND2_X1 U7316 ( .A1(n6001), .A2(n7167), .ZN(n7209) );
  NAND2_X1 U7317 ( .A1(n7865), .A2(n7209), .ZN(n7861) );
  NAND2_X1 U7318 ( .A1(n7869), .A2(n7861), .ZN(n5692) );
  AND2_X1 U7319 ( .A1(n5691), .A2(n9959), .ZN(n7886) );
  INV_X1 U7320 ( .A(n7886), .ZN(n7876) );
  NAND2_X1 U7321 ( .A1(n5692), .A2(n7876), .ZN(n7812) );
  NAND2_X1 U7322 ( .A1(n5682), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7323 ( .A1(n5614), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5699) );
  NOR2_X1 U7324 ( .A1(n5693), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5694) );
  NOR2_X1 U7325 ( .A1(n5695), .A2(n5694), .ZN(n9630) );
  NAND2_X1 U7326 ( .A1(n5645), .A2(n9630), .ZN(n5698) );
  NAND2_X1 U7327 ( .A1(n5696), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5697) );
  NAND4_X1 U7328 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n9282)
         );
  INV_X1 U7329 ( .A(n9282), .ZN(n7163) );
  OR2_X1 U7330 ( .A1(n5701), .A2(n9791), .ZN(n5702) );
  XNOR2_X1 U7331 ( .A(n5702), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9881) );
  INV_X1 U7332 ( .A(n9881), .ZN(n6469) );
  OR2_X1 U7333 ( .A1(n5703), .A2(n6400), .ZN(n5705) );
  INV_X1 U7334 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6401) );
  OR2_X1 U7335 ( .A1(n5605), .A2(n6401), .ZN(n5704) );
  NAND2_X1 U7336 ( .A1(n7163), .A2(n9634), .ZN(n8002) );
  INV_X1 U7337 ( .A(n7167), .ZN(n10014) );
  NAND2_X1 U7338 ( .A1(n9281), .A2(n10014), .ZN(n6000) );
  NAND2_X1 U7339 ( .A1(n7866), .A2(n5706), .ZN(n7813) );
  INV_X1 U7340 ( .A(n9634), .ZN(n5999) );
  NAND2_X1 U7341 ( .A1(n9282), .A2(n5999), .ZN(n7859) );
  INV_X1 U7342 ( .A(n7859), .ZN(n5707) );
  NOR2_X1 U7343 ( .A1(n7813), .A2(n5707), .ZN(n5708) );
  NAND2_X1 U7344 ( .A1(n6422), .A2(n6345), .ZN(n5716) );
  NAND2_X1 U7345 ( .A1(n5712), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5714) );
  INV_X1 U7346 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7347 ( .A1(n5739), .A2(n5713), .ZN(n5724) );
  AOI22_X1 U7348 ( .A1(n5834), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5833), .B2(
        n6487), .ZN(n5715) );
  NAND2_X1 U7349 ( .A1(n5614), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7350 ( .A1(n5696), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7351 ( .A1(n5682), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7352 ( .A1(n5717), .A2(n9064), .ZN(n5718) );
  NAND2_X1 U7353 ( .A1(n5729), .A2(n5718), .ZN(n9855) );
  INV_X1 U7354 ( .A(n9855), .ZN(n5719) );
  NAND2_X1 U7355 ( .A1(n5645), .A2(n5719), .ZN(n5720) );
  NAND4_X1 U7356 ( .A1(n5723), .A2(n5722), .A3(n5721), .A4(n5720), .ZN(n9969)
         );
  INV_X1 U7357 ( .A(n9969), .ZN(n7389) );
  OR2_X1 U7358 ( .A1(n7379), .A2(n7389), .ZN(n7887) );
  NAND2_X1 U7359 ( .A1(n7379), .A2(n7389), .ZN(n7884) );
  NAND2_X1 U7360 ( .A1(n7887), .A2(n7884), .ZN(n7811) );
  NAND2_X1 U7361 ( .A1(n6478), .A2(n6345), .ZN(n5727) );
  NAND2_X1 U7362 ( .A1(n5724), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U7363 ( .A(n5725), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U7364 ( .A1(n5834), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5833), .B2(
        n9891), .ZN(n5726) );
  INV_X1 U7365 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7366 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  AND2_X1 U7367 ( .A1(n5745), .A2(n5730), .ZN(n9225) );
  NAND2_X1 U7368 ( .A1(n5645), .A2(n9225), .ZN(n5735) );
  NAND2_X1 U7369 ( .A1(n5609), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7370 ( .A1(n5696), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7371 ( .A1(n5682), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5732) );
  NAND4_X1 U7372 ( .A1(n5735), .A2(n5734), .A3(n5733), .A4(n5732), .ZN(n9278)
         );
  INV_X1 U7373 ( .A(n9278), .ZN(n5736) );
  NAND2_X1 U7374 ( .A1(n9224), .A2(n5736), .ZN(n7885) );
  NAND2_X1 U7375 ( .A1(n7889), .A2(n7885), .ZN(n7817) );
  INV_X1 U7376 ( .A(n7884), .ZN(n7877) );
  NOR2_X1 U7377 ( .A1(n7817), .A2(n7877), .ZN(n5737) );
  NAND2_X1 U7378 ( .A1(n6526), .A2(n6345), .ZN(n5742) );
  OAI21_X1 U7379 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U7380 ( .A1(n5739), .A2(n5738), .ZN(n5752) );
  INV_X1 U7381 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5740) );
  XNOR2_X1 U7382 ( .A(n5752), .B(n5740), .ZN(n6998) );
  AOI22_X1 U7383 ( .A1(n5834), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5833), .B2(
        n6998), .ZN(n5741) );
  NAND2_X1 U7384 ( .A1(n5682), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7385 ( .A1(n5614), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5749) );
  INV_X1 U7386 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7387 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  AND2_X1 U7388 ( .A1(n5758), .A2(n5746), .ZN(n9125) );
  NAND2_X1 U7389 ( .A1(n5645), .A2(n9125), .ZN(n5748) );
  NAND2_X1 U7390 ( .A1(n5696), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5747) );
  NAND4_X1 U7391 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n9277)
         );
  INV_X1 U7392 ( .A(n9277), .ZN(n5751) );
  NAND2_X1 U7393 ( .A1(n9130), .A2(n5751), .ZN(n8009) );
  NAND2_X1 U7394 ( .A1(n7890), .A2(n8009), .ZN(n7440) );
  INV_X1 U7395 ( .A(n7440), .ZN(n7820) );
  NAND2_X1 U7396 ( .A1(n6548), .A2(n6345), .ZN(n5755) );
  OAI21_X1 U7397 ( .B1(n5752), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5753) );
  XNOR2_X1 U7398 ( .A(n5753), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U7399 ( .A1(n5834), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5833), .B2(
        n9902), .ZN(n5754) );
  NAND2_X1 U7400 ( .A1(n5682), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7401 ( .A1(n5609), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5762) );
  INV_X1 U7402 ( .A(n5758), .ZN(n5756) );
  NAND2_X1 U7403 ( .A1(n5756), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5771) );
  INV_X1 U7404 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7405 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  AND2_X1 U7406 ( .A1(n5771), .A2(n5759), .ZN(n7571) );
  NAND2_X1 U7407 ( .A1(n5645), .A2(n7571), .ZN(n5761) );
  NAND2_X1 U7408 ( .A1(n5696), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5760) );
  NAND4_X1 U7409 ( .A1(n5763), .A2(n5762), .A3(n5761), .A4(n5760), .ZN(n9276)
         );
  INV_X1 U7410 ( .A(n9276), .ZN(n5764) );
  OR2_X1 U7411 ( .A1(n9202), .A2(n5764), .ZN(n8013) );
  NAND2_X1 U7412 ( .A1(n9202), .A2(n5764), .ZN(n8010) );
  INV_X1 U7413 ( .A(n7890), .ZN(n5765) );
  NOR2_X1 U7414 ( .A1(n7883), .A2(n5765), .ZN(n5766) );
  NAND2_X1 U7415 ( .A1(n7442), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U7416 ( .A1(n5767), .A2(n8010), .ZN(n9610) );
  INV_X1 U7417 ( .A(n9610), .ZN(n5778) );
  NAND2_X1 U7418 ( .A1(n5768), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5769) );
  XNOR2_X1 U7419 ( .A(n5769), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U7420 ( .A1(n5834), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5833), .B2(
        n9913), .ZN(n5770) );
  NAND2_X1 U7421 ( .A1(n5682), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7422 ( .A1(n5614), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5775) );
  INV_X1 U7423 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U7424 ( .A1(n5771), .A2(n8922), .ZN(n5772) );
  AND2_X1 U7425 ( .A1(n5788), .A2(n5772), .ZN(n9620) );
  NAND2_X1 U7426 ( .A1(n5645), .A2(n9620), .ZN(n5774) );
  NAND2_X1 U7427 ( .A1(n5696), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5773) );
  NAND4_X1 U7428 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n9275)
         );
  INV_X1 U7429 ( .A(n9275), .ZN(n6007) );
  NAND2_X1 U7430 ( .A1(n9723), .A2(n6007), .ZN(n7896) );
  NAND2_X1 U7431 ( .A1(n8014), .A2(n7896), .ZN(n9611) );
  NAND2_X1 U7432 ( .A1(n6808), .A2(n6345), .ZN(n5785) );
  NAND2_X1 U7433 ( .A1(n5779), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5780) );
  MUX2_X1 U7434 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5780), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5781) );
  INV_X1 U7435 ( .A(n5781), .ZN(n5783) );
  NOR2_X1 U7436 ( .A1(n5783), .A2(n5782), .ZN(n9925) );
  AOI22_X1 U7437 ( .A1(n5834), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5833), .B2(
        n9925), .ZN(n5784) );
  NAND2_X1 U7438 ( .A1(n5614), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7439 ( .A1(n5696), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5792) );
  INV_X1 U7440 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7441 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  AND2_X1 U7442 ( .A1(n5797), .A2(n5789), .ZN(n9599) );
  NAND2_X1 U7443 ( .A1(n5645), .A2(n9599), .ZN(n5791) );
  NAND2_X1 U7444 ( .A1(n5658), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5790) );
  NAND4_X1 U7445 ( .A1(n5793), .A2(n5792), .A3(n5791), .A4(n5790), .ZN(n9274)
         );
  XNOR2_X1 U7446 ( .A(n9784), .B(n9274), .ZN(n9592) );
  INV_X1 U7447 ( .A(n9274), .ZN(n7901) );
  NAND2_X1 U7448 ( .A1(n9784), .A2(n7901), .ZN(n7905) );
  NAND2_X1 U7449 ( .A1(n6853), .A2(n6345), .ZN(n5796) );
  OR2_X1 U7450 ( .A1(n5782), .A2(n9791), .ZN(n5794) );
  XNOR2_X1 U7451 ( .A(n5794), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7175) );
  AOI22_X1 U7452 ( .A1(n5834), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5833), .B2(
        n7175), .ZN(n5795) );
  NAND2_X1 U7453 ( .A1(n5614), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7454 ( .A1(n5696), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5801) );
  INV_X1 U7455 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U7456 ( .A1(n5797), .A2(n9150), .ZN(n5798) );
  AND2_X1 U7457 ( .A1(n5809), .A2(n5798), .ZN(n9584) );
  NAND2_X1 U7458 ( .A1(n5645), .A2(n9584), .ZN(n5800) );
  NAND2_X1 U7459 ( .A1(n5682), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5799) );
  NAND4_X1 U7460 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n9273)
         );
  INV_X1 U7461 ( .A(n9273), .ZN(n5803) );
  OR2_X1 U7462 ( .A1(n9583), .A2(n5803), .ZN(n8020) );
  NAND2_X1 U7463 ( .A1(n9583), .A2(n5803), .ZN(n8019) );
  NAND2_X1 U7464 ( .A1(n8020), .A2(n8019), .ZN(n6012) );
  NAND2_X1 U7465 ( .A1(n9577), .A2(n9576), .ZN(n5804) );
  NAND2_X1 U7466 ( .A1(n6867), .A2(n6345), .ZN(n5806) );
  XNOR2_X1 U7467 ( .A(n5817), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U7468 ( .A1(n5834), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5833), .B2(
        n9944), .ZN(n5805) );
  NAND2_X1 U7469 ( .A1(n5658), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7470 ( .A1(n5609), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5813) );
  INV_X1 U7471 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7472 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  AND2_X1 U7473 ( .A1(n5822), .A2(n5810), .ZN(n9568) );
  NAND2_X1 U7474 ( .A1(n5645), .A2(n9568), .ZN(n5812) );
  NAND2_X1 U7475 ( .A1(n5696), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5811) );
  NAND4_X1 U7476 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n9272)
         );
  INV_X1 U7477 ( .A(n9272), .ZN(n6013) );
  OR2_X1 U7478 ( .A1(n9775), .A2(n6013), .ZN(n9543) );
  NAND2_X1 U7479 ( .A1(n9775), .A2(n6013), .ZN(n7911) );
  NAND2_X1 U7480 ( .A1(n9543), .A2(n7911), .ZN(n9560) );
  INV_X1 U7481 ( .A(n9560), .ZN(n5815) );
  NAND2_X1 U7482 ( .A1(n6923), .A2(n6345), .ZN(n5820) );
  XNOR2_X1 U7483 ( .A(n5830), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9322) );
  AOI22_X1 U7484 ( .A1(n5834), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5833), .B2(
        n9322), .ZN(n5819) );
  NAND2_X1 U7485 ( .A1(n5682), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7486 ( .A1(n5614), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5826) );
  INV_X1 U7487 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7488 ( .A1(n5822), .A2(n5821), .ZN(n5823) );
  AND2_X1 U7489 ( .A1(n5838), .A2(n5823), .ZN(n9553) );
  NAND2_X1 U7490 ( .A1(n5645), .A2(n9553), .ZN(n5825) );
  NAND2_X1 U7491 ( .A1(n5696), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5824) );
  NAND4_X1 U7492 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n9271)
         );
  INV_X1 U7493 ( .A(n9271), .ZN(n6015) );
  OR2_X1 U7494 ( .A1(n9703), .A2(n6015), .ZN(n7916) );
  NAND2_X1 U7495 ( .A1(n9703), .A2(n6015), .ZN(n7918) );
  NAND2_X1 U7496 ( .A1(n7916), .A2(n7918), .ZN(n9544) );
  INV_X1 U7497 ( .A(n9543), .ZN(n7912) );
  NOR2_X1 U7498 ( .A1(n9544), .A2(n7912), .ZN(n5828) );
  NAND2_X1 U7499 ( .A1(n9546), .A2(n7918), .ZN(n9530) );
  NAND2_X1 U7500 ( .A1(n7130), .A2(n6345), .ZN(n5836) );
  NAND2_X1 U7501 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  AOI22_X1 U7502 ( .A1(n5834), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9330), .B2(
        n5833), .ZN(n5835) );
  NAND2_X1 U7503 ( .A1(n5609), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7504 ( .A1(n5682), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5842) );
  INV_X1 U7505 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5837) );
  INV_X1 U7506 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7507 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  AND2_X1 U7508 ( .A1(n5847), .A2(n5839), .ZN(n9533) );
  NAND2_X1 U7509 ( .A1(n5645), .A2(n9533), .ZN(n5841) );
  NAND2_X1 U7510 ( .A1(n5696), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5840) );
  NAND4_X1 U7511 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .ZN(n9270)
         );
  INV_X1 U7512 ( .A(n9270), .ZN(n6017) );
  OR2_X1 U7513 ( .A1(n9766), .A2(n6017), .ZN(n7919) );
  NAND2_X1 U7514 ( .A1(n9766), .A2(n6017), .ZN(n7989) );
  NAND2_X1 U7515 ( .A1(n7247), .A2(n6345), .ZN(n5845) );
  INV_X1 U7516 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7248) );
  OR2_X1 U7517 ( .A1(n5605), .A2(n7248), .ZN(n5844) );
  NAND2_X1 U7518 ( .A1(n5846), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5858) );
  INV_X1 U7519 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U7520 ( .A1(n5847), .A2(n9190), .ZN(n5848) );
  AND2_X1 U7521 ( .A1(n5858), .A2(n5848), .ZN(n9522) );
  NAND2_X1 U7522 ( .A1(n9522), .A2(n5645), .ZN(n5852) );
  NAND2_X1 U7523 ( .A1(n5682), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7524 ( .A1(n5609), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7525 ( .A1(n5696), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5849) );
  NAND4_X1 U7526 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n9269)
         );
  INV_X1 U7527 ( .A(n9269), .ZN(n9501) );
  NAND2_X1 U7528 ( .A1(n9521), .A2(n9501), .ZN(n7913) );
  INV_X1 U7529 ( .A(n7913), .ZN(n5853) );
  NAND2_X1 U7530 ( .A1(n7346), .A2(n6345), .ZN(n5855) );
  OR2_X1 U7531 ( .A1(n5605), .A2(n7347), .ZN(n5854) );
  INV_X1 U7532 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7533 ( .A1(n5614), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7534 ( .A1(n5682), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5856) );
  AND2_X1 U7535 ( .A1(n5857), .A2(n5856), .ZN(n5861) );
  INV_X1 U7536 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U7537 ( .A1(n5858), .A2(n9117), .ZN(n5859) );
  NAND2_X1 U7538 ( .A1(n5866), .A2(n5859), .ZN(n9505) );
  INV_X1 U7539 ( .A(n5645), .ZN(n5908) );
  OR2_X1 U7540 ( .A1(n9505), .A2(n5908), .ZN(n5860) );
  OAI211_X1 U7541 ( .C1(n5731), .C2(n5862), .A(n5861), .B(n5860), .ZN(n9268)
         );
  INV_X1 U7542 ( .A(n9268), .ZN(n9477) );
  OR2_X1 U7543 ( .A1(n9757), .A2(n9477), .ZN(n7923) );
  NAND2_X1 U7544 ( .A1(n9757), .A2(n9477), .ZN(n7925) );
  NAND2_X1 U7545 ( .A1(n7923), .A2(n7925), .ZN(n9494) );
  INV_X1 U7546 ( .A(n9492), .ZN(n7780) );
  NOR2_X1 U7547 ( .A1(n9494), .A2(n7780), .ZN(n5863) );
  NAND2_X1 U7548 ( .A1(n9496), .A2(n7925), .ZN(n9473) );
  NAND2_X1 U7549 ( .A1(n7414), .A2(n6345), .ZN(n5865) );
  OR2_X1 U7550 ( .A1(n5605), .A2(n7745), .ZN(n5864) );
  INV_X1 U7551 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U7552 ( .A1(n5866), .A2(n9208), .ZN(n5867) );
  NAND2_X1 U7553 ( .A1(n5872), .A2(n5867), .ZN(n9482) );
  AOI22_X1 U7554 ( .A1(n5614), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n5696), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7555 ( .A1(n5658), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5868) );
  OAI211_X1 U7556 ( .C1(n9482), .C2(n5908), .A(n5869), .B(n5868), .ZN(n9499)
         );
  INV_X1 U7557 ( .A(n9499), .ZN(n9118) );
  OR2_X1 U7558 ( .A1(n9752), .A2(n9118), .ZN(n7776) );
  NAND2_X1 U7559 ( .A1(n9752), .A2(n9118), .ZN(n9462) );
  NAND2_X1 U7560 ( .A1(n9472), .A2(n9462), .ZN(n5878) );
  OR2_X1 U7561 ( .A1(n5605), .A2(n7470), .ZN(n5870) );
  INV_X1 U7562 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5876) );
  INV_X1 U7563 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U7564 ( .A1(n5872), .A2(n8932), .ZN(n5873) );
  NAND2_X1 U7565 ( .A1(n5883), .A2(n5873), .ZN(n9457) );
  OR2_X1 U7566 ( .A1(n9457), .A2(n5908), .ZN(n5875) );
  AOI22_X1 U7567 ( .A1(n5682), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5614), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n5874) );
  OAI211_X1 U7568 ( .C1(n5731), .C2(n5876), .A(n5875), .B(n5874), .ZN(n9475)
         );
  INV_X1 U7569 ( .A(n6024), .ZN(n5877) );
  NAND2_X1 U7570 ( .A1(n9454), .A2(n5877), .ZN(n9461) );
  NAND2_X1 U7571 ( .A1(n5879), .A2(n6345), .ZN(n5881) );
  OR2_X1 U7572 ( .A1(n5605), .A2(n7554), .ZN(n5880) );
  INV_X1 U7573 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U7574 ( .A1(n5883), .A2(n9180), .ZN(n5884) );
  NAND2_X1 U7575 ( .A1(n5894), .A2(n5884), .ZN(n9178) );
  OR2_X1 U7576 ( .A1(n9178), .A2(n5908), .ZN(n5889) );
  INV_X1 U7577 ( .A(n5682), .ZN(n5929) );
  INV_X1 U7578 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U7579 ( .A1(n5696), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7580 ( .A1(n5614), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5885) );
  OAI211_X1 U7581 ( .C1(n5929), .C2(n9677), .A(n5886), .B(n5885), .ZN(n5887)
         );
  INV_X1 U7582 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7583 ( .A1(n5889), .A2(n5888), .ZN(n9466) );
  NAND2_X1 U7584 ( .A1(n9676), .A2(n9425), .ZN(n7785) );
  NAND2_X1 U7585 ( .A1(n7777), .A2(n7785), .ZN(n9438) );
  INV_X1 U7586 ( .A(n9475), .ZN(n9211) );
  AND2_X1 U7587 ( .A1(n9680), .A2(n9211), .ZN(n7942) );
  NOR2_X1 U7588 ( .A1(n9438), .A2(n7942), .ZN(n5890) );
  OR2_X1 U7589 ( .A1(n5605), .A2(n9060), .ZN(n5891) );
  INV_X1 U7590 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7591 ( .A1(n5894), .A2(n5893), .ZN(n5895) );
  AND2_X1 U7592 ( .A1(n5906), .A2(n5895), .ZN(n9429) );
  NAND2_X1 U7593 ( .A1(n9429), .A2(n5645), .ZN(n5900) );
  INV_X1 U7594 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U7595 ( .A1(n5696), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7596 ( .A1(n5614), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5896) );
  OAI211_X1 U7597 ( .C1(n5929), .C2(n9044), .A(n5897), .B(n5896), .ZN(n5898)
         );
  INV_X1 U7598 ( .A(n5898), .ZN(n5899) );
  INV_X1 U7599 ( .A(n9267), .ZN(n9410) );
  NAND2_X1 U7600 ( .A1(n9671), .A2(n9410), .ZN(n7956) );
  NAND2_X1 U7601 ( .A1(n7957), .A2(n7956), .ZN(n9423) );
  NAND2_X1 U7602 ( .A1(n7680), .A2(n6345), .ZN(n5903) );
  OR2_X1 U7603 ( .A1(n5605), .A2(n7681), .ZN(n5902) );
  INV_X1 U7604 ( .A(n5906), .ZN(n5904) );
  NAND2_X1 U7605 ( .A1(n5904), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5917) );
  INV_X1 U7606 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7607 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7608 ( .A1(n5917), .A2(n5907), .ZN(n9245) );
  INV_X1 U7609 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U7610 ( .A1(n5609), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U7611 ( .A1(n5696), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5909) );
  OAI211_X1 U7612 ( .C1(n9059), .C2(n5929), .A(n5910), .B(n5909), .ZN(n5911)
         );
  INV_X1 U7613 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7614 ( .A1(n5913), .A2(n5912), .ZN(n9266) );
  NAND2_X1 U7615 ( .A1(n9741), .A2(n9426), .ZN(n7962) );
  NAND2_X1 U7616 ( .A1(n9405), .A2(n7962), .ZN(n9393) );
  NAND2_X1 U7617 ( .A1(n7700), .A2(n6345), .ZN(n5915) );
  OR2_X1 U7618 ( .A1(n5605), .A2(n7732), .ZN(n5914) );
  INV_X1 U7619 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7620 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  NAND2_X1 U7621 ( .A1(n9389), .A2(n5645), .ZN(n5924) );
  INV_X1 U7622 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7623 ( .A1(n5614), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7624 ( .A1(n5696), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5919) );
  OAI211_X1 U7625 ( .C1(n5921), .C2(n5929), .A(n5920), .B(n5919), .ZN(n5922)
         );
  INV_X1 U7626 ( .A(n5922), .ZN(n5923) );
  NAND2_X1 U7627 ( .A1(n7729), .A2(n6345), .ZN(n5926) );
  OR2_X1 U7628 ( .A1(n5605), .A2(n7730), .ZN(n5925) );
  XNOR2_X1 U7629 ( .A(n9364), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9375) );
  NAND2_X1 U7630 ( .A1(n9375), .A2(n5645), .ZN(n5932) );
  INV_X1 U7631 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U7632 ( .A1(n5609), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7633 ( .A1(n5696), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5927) );
  OAI211_X1 U7634 ( .C1(n9657), .C2(n5929), .A(n5928), .B(n5927), .ZN(n5930)
         );
  INV_X1 U7635 ( .A(n5930), .ZN(n5931) );
  NAND2_X1 U7636 ( .A1(n5932), .A2(n5931), .ZN(n9359) );
  INV_X1 U7637 ( .A(n9359), .ZN(n5933) );
  NAND2_X1 U7638 ( .A1(n4340), .A2(n9352), .ZN(n5941) );
  INV_X1 U7639 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7640 ( .A1(n5937), .A2(n5935), .ZN(n5936) );
  INV_X1 U7641 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5968) );
  OR2_X1 U7642 ( .A1(n6034), .A2(n6035), .ZN(n5940) );
  NAND2_X1 U7643 ( .A1(n5938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5939) );
  XNOR2_X1 U7644 ( .A(n5939), .B(P1_IR_REG_20__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7645 ( .A1(n7993), .A2(n5962), .ZN(n7985) );
  NAND2_X1 U7646 ( .A1(n5941), .A2(n9595), .ZN(n5948) );
  INV_X1 U7647 ( .A(n7731), .ZN(n6504) );
  NAND2_X1 U7648 ( .A1(n8049), .A2(n7993), .ZN(n7797) );
  INV_X1 U7649 ( .A(n7797), .ZN(n6414) );
  NAND2_X1 U7650 ( .A1(n5645), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7651 ( .A1(n5635), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7652 ( .A1(n5614), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7653 ( .A1(n5682), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5942) );
  AND3_X1 U7654 ( .A1(n5944), .A2(n5943), .A3(n5942), .ZN(n5945) );
  OAI21_X1 U7655 ( .B1(n9364), .B2(n5946), .A(n5945), .ZN(n9265) );
  AND2_X1 U7656 ( .A1(n7731), .A2(n6414), .ZN(n9498) );
  AOI22_X1 U7657 ( .A1(n9408), .A2(n9465), .B1(n9265), .B2(n9498), .ZN(n5947)
         );
  NAND2_X1 U7658 ( .A1(n5948), .A2(n5947), .ZN(n9380) );
  NAND2_X1 U7659 ( .A1(n6859), .A2(n5950), .ZN(n6873) );
  INV_X1 U7660 ( .A(n7379), .ZN(n9850) );
  INV_X1 U7661 ( .A(n9224), .ZN(n7488) );
  NAND2_X1 U7662 ( .A1(n9455), .A2(n9460), .ZN(n9444) );
  AND2_X1 U7663 ( .A1(n6034), .A2(n7803), .ZN(n6037) );
  NAND2_X1 U7664 ( .A1(n6037), .A2(n7837), .ZN(n9617) );
  INV_X1 U7665 ( .A(n9362), .ZN(n5952) );
  AOI211_X1 U7666 ( .C1(n9655), .C2(n9388), .A(n9617), .B(n5952), .ZN(n9374)
         );
  INV_X1 U7667 ( .A(n9656), .ZN(n5988) );
  NAND2_X1 U7668 ( .A1(n4315), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5953) );
  XNOR2_X1 U7669 ( .A(n5953), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5965) );
  INV_X1 U7670 ( .A(n5965), .ZN(n7630) );
  NAND2_X1 U7671 ( .A1(n7630), .A2(P1_B_REG_SCAN_IN), .ZN(n5958) );
  INV_X1 U7672 ( .A(n5954), .ZN(n5955) );
  NAND2_X1 U7673 ( .A1(n5955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5956) );
  MUX2_X1 U7674 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5956), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5957) );
  MUX2_X1 U7675 ( .A(P1_B_REG_SCAN_IN), .B(n5958), .S(n7555), .Z(n5960) );
  INV_X1 U7676 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U7677 ( .A1(n6410), .A2(n8975), .ZN(n5961) );
  INV_X1 U7678 ( .A(n5966), .ZN(n7682) );
  NAND2_X1 U7679 ( .A1(n7682), .A2(n7630), .ZN(n6411) );
  INV_X1 U7680 ( .A(n6324), .ZN(n5963) );
  NOR2_X1 U7681 ( .A1(n6954), .A2(n5963), .ZN(n5985) );
  NAND2_X2 U7682 ( .A1(n5967), .A2(n5966), .ZN(n6074) );
  NAND2_X1 U7683 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  NAND2_X1 U7684 ( .A1(n5970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  INV_X1 U7685 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7686 ( .A(n5972), .B(n5971), .ZN(n6413) );
  NAND2_X1 U7687 ( .A1(n6074), .A2(n6384), .ZN(n8047) );
  NAND2_X1 U7688 ( .A1(n6035), .A2(n7837), .ZN(n6068) );
  INV_X1 U7689 ( .A(n6068), .ZN(n8038) );
  OR2_X1 U7690 ( .A1(n7797), .A2(n8038), .ZN(n6326) );
  INV_X1 U7691 ( .A(n6326), .ZN(n5973) );
  NOR2_X1 U7692 ( .A1(n8047), .A2(n5973), .ZN(n5984) );
  NOR2_X1 U7693 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n5977) );
  NOR4_X1 U7694 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5976) );
  NOR4_X1 U7695 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5975) );
  NOR4_X1 U7696 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U7697 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n5983)
         );
  NOR4_X1 U7698 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5981) );
  NOR4_X1 U7699 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5980) );
  NOR4_X1 U7700 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5979) );
  NOR4_X1 U7701 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7702 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n5982)
         );
  OAI21_X1 U7703 ( .B1(n5983), .B2(n5982), .A(n6410), .ZN(n6317) );
  AND2_X1 U7704 ( .A1(n5984), .A2(n6317), .ZN(n6955) );
  INV_X1 U7705 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7706 ( .A1(n6410), .A2(n5986), .ZN(n5987) );
  NAND2_X1 U7707 ( .A1(n7682), .A2(n7555), .ZN(n9790) );
  INV_X1 U7708 ( .A(n6368), .ZN(n6956) );
  AND2_X2 U7709 ( .A1(n6369), .A2(n6956), .ZN(n10030) );
  MUX2_X1 U7710 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n5988), .S(n10030), .Z(n5989) );
  NAND2_X1 U7711 ( .A1(n9288), .A2(n7024), .ZN(n7021) );
  NAND2_X1 U7712 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  NAND2_X1 U7713 ( .A1(n7020), .A2(n5993), .ZN(n6833) );
  NAND2_X1 U7714 ( .A1(n7995), .A2(n5994), .ZN(n7800) );
  NAND2_X1 U7715 ( .A1(n6833), .A2(n7800), .ZN(n6835) );
  NAND2_X1 U7716 ( .A1(n6812), .A2(n5949), .ZN(n5995) );
  NAND2_X1 U7717 ( .A1(n6835), .A2(n5995), .ZN(n6858) );
  NAND2_X1 U7718 ( .A1(n7997), .A2(n7854), .ZN(n6856) );
  NAND2_X1 U7719 ( .A1(n6858), .A2(n6856), .ZN(n6857) );
  NAND2_X1 U7720 ( .A1(n6872), .A2(n5950), .ZN(n5996) );
  NAND2_X1 U7721 ( .A1(n6857), .A2(n5996), .ZN(n6876) );
  NAND2_X1 U7722 ( .A1(n6876), .A2(n7801), .ZN(n6875) );
  NAND2_X1 U7723 ( .A1(n6813), .A2(n6965), .ZN(n5997) );
  NAND2_X1 U7724 ( .A1(n6875), .A2(n5997), .ZN(n7089) );
  NAND2_X1 U7725 ( .A1(n6871), .A2(n10008), .ZN(n5998) );
  NAND2_X1 U7726 ( .A1(n8002), .A2(n7859), .ZN(n7808) );
  NAND2_X1 U7727 ( .A1(n7209), .A2(n6000), .ZN(n7863) );
  NOR2_X1 U7728 ( .A1(n9280), .A2(n7336), .ZN(n6002) );
  NOR2_X1 U7729 ( .A1(n7875), .A2(n7886), .ZN(n9954) );
  NAND2_X1 U7730 ( .A1(n7351), .A2(n7811), .ZN(n7350) );
  OR2_X1 U7731 ( .A1(n7379), .A2(n9969), .ZN(n6003) );
  OR2_X1 U7732 ( .A1(n9224), .A2(n9278), .ZN(n6004) );
  NAND2_X1 U7733 ( .A1(n7395), .A2(n6004), .ZN(n7441) );
  NAND2_X1 U7734 ( .A1(n7439), .A2(n6005), .ZN(n7566) );
  NAND2_X1 U7735 ( .A1(n7566), .A2(n7883), .ZN(n7565) );
  NAND2_X1 U7736 ( .A1(n7565), .A2(n6006), .ZN(n9607) );
  NAND2_X1 U7737 ( .A1(n9723), .A2(n9275), .ZN(n6009) );
  NAND2_X1 U7738 ( .A1(n9590), .A2(n6010), .ZN(n6011) );
  NAND2_X1 U7739 ( .A1(n6011), .A2(n4867), .ZN(n9575) );
  AOI22_X2 U7740 ( .A1(n9575), .A2(n6012), .B1(n9273), .B2(n9583), .ZN(n9559)
         );
  INV_X1 U7741 ( .A(n9775), .ZN(n9570) );
  NAND2_X1 U7742 ( .A1(n9703), .A2(n9271), .ZN(n6016) );
  NAND2_X1 U7743 ( .A1(n9535), .A2(n6017), .ZN(n6019) );
  NAND2_X1 U7744 ( .A1(n9492), .A2(n7913), .ZN(n9515) );
  NAND2_X1 U7745 ( .A1(n9514), .A2(n9515), .ZN(n9513) );
  NAND2_X1 U7746 ( .A1(n9513), .A2(n6020), .ZN(n9491) );
  NAND2_X1 U7747 ( .A1(n9491), .A2(n4365), .ZN(n6022) );
  NOR2_X1 U7748 ( .A1(n9752), .A2(n9499), .ZN(n6023) );
  NOR2_X1 U7749 ( .A1(n9671), .A2(n9267), .ZN(n6026) );
  NAND2_X1 U7750 ( .A1(n9450), .A2(n9425), .ZN(n9418) );
  INV_X1 U7751 ( .A(n9418), .ZN(n6025) );
  NOR2_X1 U7752 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7753 ( .A1(n9417), .A2(n6027), .ZN(n6029) );
  NAND2_X1 U7754 ( .A1(n9671), .A2(n9267), .ZN(n6028) );
  NOR2_X1 U7755 ( .A1(n9404), .A2(n9426), .ZN(n9383) );
  NAND2_X1 U7756 ( .A1(n9391), .A2(n6030), .ZN(n6032) );
  INV_X1 U7757 ( .A(n6032), .ZN(n6031) );
  NAND2_X1 U7758 ( .A1(n9404), .A2(n9426), .ZN(n9384) );
  AND2_X1 U7759 ( .A1(n9384), .A2(n6032), .ZN(n6033) );
  INV_X1 U7760 ( .A(n6037), .ZN(n9975) );
  OR2_X1 U7761 ( .A1(n7797), .A2(n6068), .ZN(n8046) );
  NAND2_X1 U7762 ( .A1(n9975), .A2(n8046), .ZN(n9980) );
  AND2_X1 U7763 ( .A1(n6072), .A2(n6068), .ZN(n6036) );
  OR2_X1 U7764 ( .A1(n9980), .A2(n6036), .ZN(n6958) );
  NAND2_X1 U7765 ( .A1(n10030), .A2(n10026), .ZN(n9787) );
  NOR2_X1 U7766 ( .A1(n8097), .A2(n8775), .ZN(n6046) );
  MUX2_X1 U7767 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8633), .S(n10135), .Z(n6049) );
  INV_X1 U7768 ( .A(n6049), .ZN(n6053) );
  NAND2_X1 U7769 ( .A1(n10080), .A2(n10135), .ZN(n8828) );
  OAI22_X1 U7770 ( .A1(n8639), .A2(n8828), .B1(n8249), .B2(n8813), .ZN(n6051)
         );
  INV_X1 U7771 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7772 ( .A1(n6767), .A2(n5553), .ZN(n6772) );
  INV_X1 U7773 ( .A(n6054), .ZN(n6632) );
  NOR2_X1 U7774 ( .A1(n6639), .A2(n6666), .ZN(n6661) );
  OR2_X1 U7775 ( .A1(n5511), .A2(n6055), .ZN(n6058) );
  NAND3_X1 U7776 ( .A1(n8256), .A2(n10108), .A3(n6058), .ZN(n6653) );
  NAND2_X1 U7777 ( .A1(n6653), .A2(n8682), .ZN(n6630) );
  NAND2_X1 U7778 ( .A1(n6661), .A2(n6630), .ZN(n6062) );
  INV_X1 U7779 ( .A(n6631), .ZN(n6057) );
  AND2_X1 U7780 ( .A1(n6057), .A2(n6056), .ZN(n6665) );
  INV_X1 U7781 ( .A(n6058), .ZN(n6059) );
  NAND2_X1 U7782 ( .A1(n8277), .A2(n6059), .ZN(n6633) );
  NAND2_X1 U7783 ( .A1(n6659), .A2(n6633), .ZN(n6060) );
  NAND2_X1 U7784 ( .A1(n6665), .A2(n6060), .ZN(n6061) );
  INV_X2 U7785 ( .A(n10121), .ZN(n10119) );
  MUX2_X1 U7786 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8633), .S(n10119), .Z(n6063) );
  INV_X1 U7787 ( .A(n6063), .ZN(n6066) );
  OAI22_X1 U7788 ( .A1(n8639), .A2(n8894), .B1(n8249), .B2(n8878), .ZN(n6064)
         );
  INV_X1 U7789 ( .A(n6064), .ZN(n6065) );
  AND2_X1 U7790 ( .A1(n7993), .A2(n7837), .ZN(n6067) );
  AND2_X2 U7791 ( .A1(n6074), .A2(n6067), .ZN(n6071) );
  INV_X1 U7792 ( .A(n6071), .ZN(n6118) );
  NAND2_X2 U7793 ( .A1(n6070), .A2(n6074), .ZN(n6078) );
  OAI22_X1 U7794 ( .A1(n9485), .A2(n6118), .B1(n9118), .B2(n6078), .ZN(n9206)
         );
  NAND2_X1 U7795 ( .A1(n6072), .A2(n7803), .ZN(n6073) );
  NAND2_X4 U7796 ( .A1(n6075), .A2(n6074), .ZN(n6298) );
  NAND2_X2 U7797 ( .A1(n6078), .A2(n6298), .ZN(n6101) );
  INV_X1 U7798 ( .A(n6074), .ZN(n6076) );
  NAND2_X1 U7799 ( .A1(n6076), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7800 ( .A1(n6082), .A2(n6077), .ZN(n6501) );
  NAND2_X1 U7801 ( .A1(n9288), .A2(n6310), .ZN(n6081) );
  INV_X1 U7802 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6505) );
  NOR2_X1 U7803 ( .A1(n6074), .A2(n6505), .ZN(n6079) );
  AOI21_X1 U7804 ( .B1(n7024), .B2(n6311), .A(n6079), .ZN(n6080) );
  NAND2_X1 U7805 ( .A1(n6081), .A2(n6080), .ZN(n6500) );
  NAND2_X1 U7806 ( .A1(n6501), .A2(n6500), .ZN(n6499) );
  NAND2_X1 U7807 ( .A1(n6082), .A2(n6308), .ZN(n6083) );
  AND2_X1 U7808 ( .A1(n6499), .A2(n6083), .ZN(n9104) );
  NAND2_X1 U7809 ( .A1(n6084), .A2(n6071), .ZN(n6087) );
  NAND2_X1 U7810 ( .A1(n6085), .A2(n6101), .ZN(n6086) );
  NAND2_X1 U7811 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  INV_X2 U7812 ( .A(n6118), .ZN(n6311) );
  XNOR2_X1 U7813 ( .A(n6089), .B(n6090), .ZN(n9105) );
  NAND2_X1 U7814 ( .A1(n9104), .A2(n9105), .ZN(n9103) );
  INV_X1 U7815 ( .A(n6089), .ZN(n6091) );
  NAND2_X1 U7816 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7817 ( .A1(n9103), .A2(n6092), .ZN(n6712) );
  NAND2_X1 U7818 ( .A1(n9286), .A2(n6311), .ZN(n6094) );
  NAND2_X1 U7819 ( .A1(n6842), .A2(n6101), .ZN(n6093) );
  NAND2_X1 U7820 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  XNOR2_X1 U7821 ( .A(n6095), .B(n6298), .ZN(n6096) );
  AOI22_X1 U7822 ( .A1(n9286), .A2(n4294), .B1(n6311), .B2(n6842), .ZN(n6097)
         );
  XNOR2_X1 U7823 ( .A(n6096), .B(n6097), .ZN(n6713) );
  NAND2_X1 U7824 ( .A1(n6712), .A2(n6713), .ZN(n6100) );
  INV_X1 U7825 ( .A(n6096), .ZN(n6098) );
  NAND2_X1 U7826 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  NAND2_X1 U7827 ( .A1(n9285), .A2(n6295), .ZN(n6103) );
  NAND2_X1 U7828 ( .A1(n6814), .A2(n6305), .ZN(n6102) );
  NAND2_X1 U7829 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  XNOR2_X1 U7830 ( .A(n6104), .B(n6298), .ZN(n6105) );
  AOI22_X1 U7831 ( .A1(n9285), .A2(n4294), .B1(n6311), .B2(n6814), .ZN(n6106)
         );
  XNOR2_X1 U7832 ( .A(n6105), .B(n6106), .ZN(n6811) );
  NAND2_X1 U7833 ( .A1(n6810), .A2(n6811), .ZN(n6109) );
  INV_X1 U7834 ( .A(n6105), .ZN(n6107) );
  NAND2_X1 U7835 ( .A1(n9284), .A2(n6295), .ZN(n6111) );
  NAND2_X1 U7836 ( .A1(n6874), .A2(n6305), .ZN(n6110) );
  NAND2_X1 U7837 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  XNOR2_X1 U7838 ( .A(n6112), .B(n6308), .ZN(n6113) );
  AOI22_X1 U7839 ( .A1(n9284), .A2(n4294), .B1(n6311), .B2(n6874), .ZN(n6114)
         );
  XNOR2_X1 U7840 ( .A(n6113), .B(n6114), .ZN(n6846) );
  INV_X1 U7841 ( .A(n6113), .ZN(n6116) );
  INV_X1 U7842 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7843 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  NAND2_X1 U7844 ( .A1(n9283), .A2(n6295), .ZN(n6120) );
  NAND2_X1 U7845 ( .A1(n9159), .A2(n4295), .ZN(n6119) );
  NAND2_X1 U7846 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  XNOR2_X1 U7847 ( .A(n6121), .B(n6308), .ZN(n6122) );
  XNOR2_X2 U7848 ( .A(n6124), .B(n6122), .ZN(n9157) );
  AOI22_X1 U7849 ( .A1(n9283), .A2(n4294), .B1(n6311), .B2(n9159), .ZN(n9156)
         );
  INV_X1 U7850 ( .A(n6122), .ZN(n6123) );
  OR2_X1 U7851 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  NAND2_X1 U7852 ( .A1(n9155), .A2(n6125), .ZN(n7311) );
  NAND2_X1 U7853 ( .A1(n9282), .A2(n6295), .ZN(n6127) );
  NAND2_X1 U7854 ( .A1(n9634), .A2(n4295), .ZN(n6126) );
  NAND2_X1 U7855 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  XNOR2_X1 U7856 ( .A(n6128), .B(n6298), .ZN(n6129) );
  AOI22_X1 U7857 ( .A1(n9282), .A2(n4294), .B1(n6071), .B2(n9634), .ZN(n6130)
         );
  XNOR2_X1 U7858 ( .A(n6129), .B(n6130), .ZN(n7312) );
  NAND2_X1 U7859 ( .A1(n7311), .A2(n7312), .ZN(n6133) );
  INV_X1 U7860 ( .A(n6129), .ZN(n6131) );
  NAND2_X1 U7861 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NAND2_X1 U7862 ( .A1(n6133), .A2(n6132), .ZN(n7160) );
  NAND2_X1 U7863 ( .A1(n9281), .A2(n6295), .ZN(n6135) );
  NAND2_X1 U7864 ( .A1(n7167), .A2(n4295), .ZN(n6134) );
  NAND2_X1 U7865 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  XNOR2_X1 U7866 ( .A(n6136), .B(n6298), .ZN(n6137) );
  AOI22_X1 U7867 ( .A1(n9281), .A2(n4294), .B1(n6071), .B2(n7167), .ZN(n6138)
         );
  XNOR2_X1 U7868 ( .A(n6137), .B(n6138), .ZN(n7161) );
  NAND2_X1 U7869 ( .A1(n7160), .A2(n7161), .ZN(n6141) );
  INV_X1 U7870 ( .A(n6137), .ZN(n6139) );
  NAND2_X1 U7871 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7872 ( .A1(n9280), .A2(n6295), .ZN(n6143) );
  NAND2_X1 U7873 ( .A1(n7336), .A2(n4295), .ZN(n6142) );
  NAND2_X1 U7874 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  XNOR2_X1 U7875 ( .A(n6144), .B(n6308), .ZN(n7251) );
  NAND2_X1 U7876 ( .A1(n9280), .A2(n4294), .ZN(n6146) );
  NAND2_X1 U7877 ( .A1(n7336), .A2(n6295), .ZN(n6145) );
  AND2_X1 U7878 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  INV_X1 U7879 ( .A(n7251), .ZN(n6148) );
  INV_X1 U7880 ( .A(n6147), .ZN(n7250) );
  NAND2_X1 U7881 ( .A1(n6148), .A2(n7250), .ZN(n6149) );
  NAND2_X1 U7882 ( .A1(n9959), .A2(n4295), .ZN(n6151) );
  NAND2_X1 U7883 ( .A1(n9279), .A2(n6295), .ZN(n6150) );
  NAND2_X1 U7884 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  XNOR2_X1 U7885 ( .A(n6152), .B(n6308), .ZN(n6154) );
  AOI22_X1 U7886 ( .A1(n9959), .A2(n6311), .B1(n9279), .B2(n4294), .ZN(n6153)
         );
  NAND2_X1 U7887 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  OAI21_X1 U7888 ( .B1(n6154), .B2(n6153), .A(n6155), .ZN(n7388) );
  NAND2_X1 U7889 ( .A1(n7386), .A2(n6155), .ZN(n6162) );
  INV_X1 U7890 ( .A(n6162), .ZN(n6160) );
  NAND2_X1 U7891 ( .A1(n7379), .A2(n4295), .ZN(n6157) );
  NAND2_X1 U7892 ( .A1(n9969), .A2(n6295), .ZN(n6156) );
  NAND2_X1 U7893 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  XNOR2_X1 U7894 ( .A(n6158), .B(n6308), .ZN(n6161) );
  INV_X1 U7895 ( .A(n6161), .ZN(n6159) );
  NAND2_X1 U7896 ( .A1(n6160), .A2(n6159), .ZN(n6163) );
  AND2_X1 U7897 ( .A1(n9969), .A2(n4294), .ZN(n6164) );
  AOI21_X1 U7898 ( .B1(n7379), .B2(n6071), .A(n6164), .ZN(n9844) );
  NAND2_X1 U7899 ( .A1(n9224), .A2(n4295), .ZN(n6167) );
  NAND2_X1 U7900 ( .A1(n9278), .A2(n6295), .ZN(n6166) );
  NAND2_X1 U7901 ( .A1(n6167), .A2(n6166), .ZN(n6168) );
  XNOR2_X1 U7902 ( .A(n6168), .B(n6298), .ZN(n6171) );
  NAND2_X1 U7903 ( .A1(n9224), .A2(n6311), .ZN(n6170) );
  NAND2_X1 U7904 ( .A1(n9278), .A2(n4294), .ZN(n6169) );
  NAND2_X1 U7905 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  NAND2_X1 U7906 ( .A1(n6171), .A2(n6172), .ZN(n9220) );
  INV_X1 U7907 ( .A(n6171), .ZN(n6174) );
  INV_X1 U7908 ( .A(n6172), .ZN(n6173) );
  NAND2_X1 U7909 ( .A1(n6174), .A2(n6173), .ZN(n9219) );
  NAND2_X1 U7910 ( .A1(n9130), .A2(n4295), .ZN(n6176) );
  NAND2_X1 U7911 ( .A1(n9277), .A2(n6311), .ZN(n6175) );
  NAND2_X1 U7912 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  XNOR2_X1 U7913 ( .A(n6177), .B(n6298), .ZN(n6179) );
  AND2_X1 U7914 ( .A1(n9277), .A2(n4294), .ZN(n6178) );
  AOI21_X1 U7915 ( .B1(n9130), .B2(n6311), .A(n6178), .ZN(n6180) );
  XNOR2_X1 U7916 ( .A(n6179), .B(n6180), .ZN(n9124) );
  INV_X1 U7917 ( .A(n6179), .ZN(n6181) );
  NAND2_X1 U7918 ( .A1(n6181), .A2(n6180), .ZN(n9194) );
  NAND2_X1 U7919 ( .A1(n9202), .A2(n4295), .ZN(n6183) );
  NAND2_X1 U7920 ( .A1(n9276), .A2(n6311), .ZN(n6182) );
  NAND2_X1 U7921 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  XNOR2_X1 U7922 ( .A(n6184), .B(n6298), .ZN(n6189) );
  INV_X1 U7923 ( .A(n6189), .ZN(n6186) );
  AND2_X1 U7924 ( .A1(n9276), .A2(n4294), .ZN(n6185) );
  AOI21_X1 U7925 ( .B1(n9202), .B2(n6311), .A(n6185), .ZN(n6188) );
  NAND2_X1 U7926 ( .A1(n6186), .A2(n6188), .ZN(n6187) );
  AND2_X1 U7927 ( .A1(n9194), .A2(n6187), .ZN(n6191) );
  INV_X1 U7928 ( .A(n6187), .ZN(n6190) );
  XNOR2_X1 U7929 ( .A(n6189), .B(n6188), .ZN(n9197) );
  NAND2_X1 U7930 ( .A1(n9723), .A2(n4295), .ZN(n6193) );
  NAND2_X1 U7931 ( .A1(n9275), .A2(n6311), .ZN(n6192) );
  NAND2_X1 U7932 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  XNOR2_X1 U7933 ( .A(n6194), .B(n6298), .ZN(n6196) );
  XNOR2_X1 U7934 ( .A(n6198), .B(n6196), .ZN(n8919) );
  AND2_X1 U7935 ( .A1(n9275), .A2(n4294), .ZN(n6195) );
  AOI21_X1 U7936 ( .B1(n9723), .B2(n6311), .A(n6195), .ZN(n8920) );
  NAND2_X1 U7937 ( .A1(n8919), .A2(n8920), .ZN(n8918) );
  INV_X1 U7938 ( .A(n6196), .ZN(n6197) );
  NAND2_X1 U7939 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  NAND2_X1 U7940 ( .A1(n8918), .A2(n6199), .ZN(n9143) );
  NAND2_X1 U7941 ( .A1(n9583), .A2(n4295), .ZN(n6201) );
  NAND2_X1 U7942 ( .A1(n9273), .A2(n6311), .ZN(n6200) );
  NAND2_X1 U7943 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  XNOR2_X1 U7944 ( .A(n6202), .B(n6298), .ZN(n9142) );
  NAND2_X1 U7945 ( .A1(n9583), .A2(n6311), .ZN(n6204) );
  NAND2_X1 U7946 ( .A1(n9273), .A2(n4294), .ZN(n6203) );
  NAND2_X1 U7947 ( .A1(n6204), .A2(n6203), .ZN(n9141) );
  NAND2_X1 U7948 ( .A1(n9142), .A2(n9141), .ZN(n9140) );
  NAND2_X1 U7949 ( .A1(n9784), .A2(n4295), .ZN(n6206) );
  NAND2_X1 U7950 ( .A1(n9274), .A2(n6295), .ZN(n6205) );
  NAND2_X1 U7951 ( .A1(n6206), .A2(n6205), .ZN(n6207) );
  XNOR2_X1 U7952 ( .A(n6207), .B(n6298), .ZN(n6212) );
  NAND2_X1 U7953 ( .A1(n9784), .A2(n6295), .ZN(n6209) );
  NAND2_X1 U7954 ( .A1(n9274), .A2(n4294), .ZN(n6208) );
  NAND2_X1 U7955 ( .A1(n6209), .A2(n6208), .ZN(n9253) );
  NAND2_X1 U7956 ( .A1(n6212), .A2(n9253), .ZN(n6210) );
  AND2_X1 U7957 ( .A1(n9140), .A2(n6210), .ZN(n6211) );
  INV_X1 U7958 ( .A(n9142), .ZN(n6215) );
  OAI21_X1 U7959 ( .B1(n6212), .B2(n9253), .A(n9141), .ZN(n6214) );
  NOR2_X1 U7960 ( .A1(n9141), .A2(n9253), .ZN(n6213) );
  INV_X1 U7961 ( .A(n6212), .ZN(n9145) );
  AOI22_X1 U7962 ( .A1(n6215), .A2(n6214), .B1(n6213), .B2(n9145), .ZN(n6216)
         );
  NAND2_X1 U7963 ( .A1(n9775), .A2(n4295), .ZN(n6218) );
  NAND2_X1 U7964 ( .A1(n9272), .A2(n6295), .ZN(n6217) );
  NAND2_X1 U7965 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  XNOR2_X1 U7966 ( .A(n6219), .B(n6308), .ZN(n6221) );
  AND2_X1 U7967 ( .A1(n9272), .A2(n4294), .ZN(n6220) );
  AOI21_X1 U7968 ( .B1(n9775), .B2(n6311), .A(n6220), .ZN(n6222) );
  NAND2_X1 U7969 ( .A1(n6221), .A2(n6222), .ZN(n6226) );
  INV_X1 U7970 ( .A(n6221), .ZN(n6224) );
  INV_X1 U7971 ( .A(n6222), .ZN(n6223) );
  NAND2_X1 U7972 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AND2_X1 U7973 ( .A1(n6226), .A2(n6225), .ZN(n9167) );
  NAND2_X1 U7974 ( .A1(n9703), .A2(n6295), .ZN(n6228) );
  NAND2_X1 U7975 ( .A1(n9271), .A2(n4294), .ZN(n6227) );
  NAND2_X1 U7976 ( .A1(n6228), .A2(n6227), .ZN(n6245) );
  INV_X1 U7977 ( .A(n6245), .ZN(n9232) );
  NAND2_X1 U7978 ( .A1(n9703), .A2(n4295), .ZN(n6230) );
  NAND2_X1 U7979 ( .A1(n9271), .A2(n6295), .ZN(n6229) );
  NAND2_X1 U7980 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7981 ( .A(n6231), .B(n6298), .ZN(n9090) );
  INV_X1 U7982 ( .A(n9090), .ZN(n9093) );
  NAND2_X1 U7983 ( .A1(n9521), .A2(n4295), .ZN(n6233) );
  NAND2_X1 U7984 ( .A1(n9269), .A2(n6071), .ZN(n6232) );
  NAND2_X1 U7985 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  XNOR2_X1 U7986 ( .A(n6234), .B(n6298), .ZN(n6248) );
  NAND2_X1 U7987 ( .A1(n9521), .A2(n6071), .ZN(n6236) );
  NAND2_X1 U7988 ( .A1(n9269), .A2(n4294), .ZN(n6235) );
  NAND2_X1 U7989 ( .A1(n6236), .A2(n6235), .ZN(n6249) );
  INV_X1 U7990 ( .A(n9111), .ZN(n6243) );
  NAND2_X1 U7991 ( .A1(n9766), .A2(n4295), .ZN(n6238) );
  NAND2_X1 U7992 ( .A1(n9270), .A2(n6311), .ZN(n6237) );
  NAND2_X1 U7993 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  XNOR2_X1 U7994 ( .A(n6239), .B(n6308), .ZN(n9092) );
  INV_X1 U7995 ( .A(n9092), .ZN(n6242) );
  NAND2_X1 U7996 ( .A1(n9766), .A2(n6071), .ZN(n6241) );
  NAND2_X1 U7997 ( .A1(n9270), .A2(n4294), .ZN(n6240) );
  NAND2_X1 U7998 ( .A1(n6241), .A2(n6240), .ZN(n9091) );
  NAND2_X1 U7999 ( .A1(n6242), .A2(n9091), .ZN(n9186) );
  OAI211_X1 U8000 ( .C1(n9232), .C2(n9093), .A(n6243), .B(n9186), .ZN(n6244)
         );
  INV_X1 U8001 ( .A(n6244), .ZN(n6254) );
  OAI21_X1 U8002 ( .B1(n9090), .B2(n6245), .A(n9091), .ZN(n6247) );
  NOR2_X1 U8003 ( .A1(n9091), .A2(n6245), .ZN(n6246) );
  AOI22_X1 U8004 ( .A1(n9092), .A2(n6247), .B1(n6246), .B2(n9093), .ZN(n6252)
         );
  INV_X1 U8005 ( .A(n6248), .ZN(n6251) );
  INV_X1 U8006 ( .A(n6249), .ZN(n6250) );
  NAND2_X1 U8007 ( .A1(n6251), .A2(n6250), .ZN(n9114) );
  OAI21_X1 U8008 ( .B1(n9111), .B2(n6252), .A(n9114), .ZN(n6253) );
  NAND2_X1 U8009 ( .A1(n9757), .A2(n4295), .ZN(n6256) );
  NAND2_X1 U8010 ( .A1(n9268), .A2(n6295), .ZN(n6255) );
  NAND2_X1 U8011 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  XNOR2_X1 U8012 ( .A(n6257), .B(n6308), .ZN(n6259) );
  AND2_X1 U8013 ( .A1(n9268), .A2(n4294), .ZN(n6258) );
  AOI21_X1 U8014 ( .B1(n9757), .B2(n6071), .A(n6258), .ZN(n6260) );
  NAND2_X1 U8015 ( .A1(n6259), .A2(n6260), .ZN(n6265) );
  INV_X1 U8016 ( .A(n6259), .ZN(n6262) );
  INV_X1 U8017 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U8018 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U8019 ( .A1(n6265), .A2(n6263), .ZN(n9113) );
  AOI22_X1 U8020 ( .A1(n9752), .A2(n4295), .B1(n6071), .B2(n9499), .ZN(n6266)
         );
  XNOR2_X1 U8021 ( .A(n6266), .B(n6298), .ZN(n6267) );
  NAND2_X1 U8022 ( .A1(n9680), .A2(n4295), .ZN(n6269) );
  NAND2_X1 U8023 ( .A1(n9475), .A2(n6071), .ZN(n6268) );
  NAND2_X1 U8024 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  XNOR2_X1 U8025 ( .A(n6270), .B(n6298), .ZN(n6273) );
  NAND2_X1 U8026 ( .A1(n9680), .A2(n6071), .ZN(n6272) );
  NAND2_X1 U8027 ( .A1(n9475), .A2(n4294), .ZN(n6271) );
  NAND2_X1 U8028 ( .A1(n6272), .A2(n6271), .ZN(n6274) );
  NAND2_X1 U8029 ( .A1(n6273), .A2(n6274), .ZN(n8928) );
  INV_X1 U8030 ( .A(n6273), .ZN(n6276) );
  INV_X1 U8031 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U8032 ( .A1(n6276), .A2(n6275), .ZN(n8930) );
  NAND2_X1 U8033 ( .A1(n9676), .A2(n4295), .ZN(n6278) );
  NAND2_X1 U8034 ( .A1(n9466), .A2(n6295), .ZN(n6277) );
  NAND2_X1 U8035 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  XNOR2_X1 U8036 ( .A(n6279), .B(n6298), .ZN(n6282) );
  AOI22_X1 U8037 ( .A1(n9676), .A2(n6311), .B1(n4294), .B2(n9466), .ZN(n6280)
         );
  XNOR2_X1 U8038 ( .A(n6282), .B(n6280), .ZN(n9176) );
  INV_X1 U8039 ( .A(n6280), .ZN(n6281) );
  NAND2_X1 U8040 ( .A1(n9671), .A2(n4295), .ZN(n6285) );
  NAND2_X1 U8041 ( .A1(n9267), .A2(n6071), .ZN(n6284) );
  NAND2_X1 U8042 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  XNOR2_X1 U8043 ( .A(n6286), .B(n6298), .ZN(n6287) );
  AOI22_X1 U8044 ( .A1(n9671), .A2(n6071), .B1(n4294), .B2(n9267), .ZN(n6288)
         );
  XNOR2_X1 U8045 ( .A(n6287), .B(n6288), .ZN(n9134) );
  INV_X1 U8046 ( .A(n6287), .ZN(n6289) );
  NAND2_X1 U8047 ( .A1(n9741), .A2(n4295), .ZN(n6291) );
  NAND2_X1 U8048 ( .A1(n9266), .A2(n6295), .ZN(n6290) );
  NAND2_X1 U8049 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  XNOR2_X1 U8050 ( .A(n6292), .B(n6298), .ZN(n6300) );
  AND2_X1 U8051 ( .A1(n9266), .A2(n4294), .ZN(n6293) );
  AOI21_X1 U8052 ( .B1(n9741), .B2(n6311), .A(n6293), .ZN(n6302) );
  XNOR2_X1 U8053 ( .A(n6300), .B(n6302), .ZN(n9242) );
  AND2_X1 U8054 ( .A1(n9408), .A2(n4294), .ZN(n6294) );
  AOI21_X1 U8055 ( .B1(n9736), .B2(n6311), .A(n6294), .ZN(n6314) );
  NAND2_X1 U8056 ( .A1(n9736), .A2(n4295), .ZN(n6297) );
  NAND2_X1 U8057 ( .A1(n9408), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U8058 ( .A1(n6297), .A2(n6296), .ZN(n6299) );
  XNOR2_X1 U8059 ( .A(n6299), .B(n6298), .ZN(n6316) );
  XOR2_X1 U8060 ( .A(n6314), .B(n6316), .Z(n8912) );
  INV_X1 U8061 ( .A(n8912), .ZN(n6303) );
  INV_X1 U8062 ( .A(n6300), .ZN(n6301) );
  OR2_X1 U8063 ( .A1(n6302), .A2(n6301), .ZN(n8909) );
  AND2_X1 U8064 ( .A1(n6303), .A2(n8909), .ZN(n6304) );
  NAND2_X1 U8065 ( .A1(n9655), .A2(n4295), .ZN(n6307) );
  NAND2_X1 U8066 ( .A1(n9359), .A2(n6071), .ZN(n6306) );
  NAND2_X1 U8067 ( .A1(n6307), .A2(n6306), .ZN(n6309) );
  XNOR2_X1 U8068 ( .A(n6309), .B(n6308), .ZN(n6313) );
  AOI22_X1 U8069 ( .A1(n9655), .A2(n6311), .B1(n4294), .B2(n9359), .ZN(n6312)
         );
  XNOR2_X1 U8070 ( .A(n6313), .B(n6312), .ZN(n6333) );
  INV_X1 U8071 ( .A(n6314), .ZN(n6315) );
  NAND3_X1 U8072 ( .A1(n6368), .A2(n6954), .A3(n6317), .ZN(n6325) );
  NOR2_X1 U8073 ( .A1(n6325), .A2(n8047), .ZN(n6322) );
  INV_X1 U8074 ( .A(n9724), .ZN(n10023) );
  AND2_X1 U8075 ( .A1(n10023), .A2(n7797), .ZN(n6318) );
  NAND2_X1 U8076 ( .A1(n6322), .A2(n6318), .ZN(n9262) );
  NAND4_X1 U8077 ( .A1(n6319), .A2(n6333), .A3(n4875), .A4(n9852), .ZN(n6336)
         );
  INV_X1 U8078 ( .A(n9655), .ZN(n9378) );
  OR2_X1 U8079 ( .A1(n9975), .A2(n7837), .ZN(n9961) );
  INV_X1 U8080 ( .A(n9961), .ZN(n6962) );
  NAND2_X1 U8081 ( .A1(n6322), .A2(n6962), .ZN(n6321) );
  NAND2_X1 U8082 ( .A1(n6321), .A2(n9978), .ZN(n9260) );
  INV_X1 U8083 ( .A(n9260), .ZN(n9849) );
  NAND2_X1 U8084 ( .A1(n6322), .A2(n8038), .ZN(n9237) );
  INV_X1 U8085 ( .A(n9465), .ZN(n9956) );
  OR2_X1 U8086 ( .A1(n9237), .A2(n9956), .ZN(n9209) );
  INV_X1 U8087 ( .A(n9209), .ZN(n9246) );
  AOI22_X1 U8088 ( .A1(n9408), .A2(n9246), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6331) );
  NAND2_X1 U8089 ( .A1(n6325), .A2(n6324), .ZN(n6328) );
  AND2_X1 U8090 ( .A1(n6074), .A2(n6326), .ZN(n6327) );
  NAND2_X1 U8091 ( .A1(n6328), .A2(n6327), .ZN(n6528) );
  NAND2_X1 U8092 ( .A1(n6528), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6329) );
  OR2_X1 U8093 ( .A1(n6413), .A2(P1_U3086), .ZN(n8052) );
  INV_X1 U8094 ( .A(n9498), .ZN(n9427) );
  OR2_X1 U8095 ( .A1(n9237), .A2(n9427), .ZN(n9210) );
  INV_X1 U8096 ( .A(n9210), .ZN(n9244) );
  AOI22_X1 U8097 ( .A1(n9375), .A2(n9247), .B1(n9265), .B2(n9244), .ZN(n6330)
         );
  OAI211_X1 U8098 ( .C1(n9378), .C2(n9849), .A(n6331), .B(n6330), .ZN(n6332)
         );
  INV_X1 U8099 ( .A(n6332), .ZN(n6334) );
  NAND4_X1 U8100 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n4355), .ZN(
        P1_U3220) );
  INV_X1 U8101 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6370) );
  INV_X1 U8102 ( .A(SI_29_), .ZN(n6340) );
  INV_X1 U8103 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8328) );
  INV_X1 U8104 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8905) );
  MUX2_X1 U8105 ( .A(n8328), .B(n8905), .S(n6388), .Z(n6342) );
  NAND2_X1 U8106 ( .A1(n6342), .A2(n9066), .ZN(n6350) );
  INV_X1 U8107 ( .A(n6342), .ZN(n6343) );
  NAND2_X1 U8108 ( .A1(n6343), .A2(SI_30_), .ZN(n6344) );
  NAND2_X1 U8109 ( .A1(n6350), .A2(n6344), .ZN(n6351) );
  NAND2_X1 U8110 ( .A1(n8326), .A2(n6345), .ZN(n6347) );
  OR2_X1 U8111 ( .A1(n5605), .A2(n8328), .ZN(n6346) );
  NAND2_X1 U8112 ( .A1(n8340), .A2(n6345), .ZN(n6349) );
  OR2_X1 U8113 ( .A1(n5605), .A2(n9798), .ZN(n6348) );
  OAI21_X1 U8114 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6356) );
  INV_X1 U8115 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6353) );
  INV_X1 U8116 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U8117 ( .A(n6353), .B(n8900), .S(n6388), .Z(n6354) );
  XNOR2_X1 U8118 ( .A(n6354), .B(SI_31_), .ZN(n6355) );
  XNOR2_X1 U8119 ( .A(n6356), .B(n6355), .ZN(n8102) );
  MUX2_X1 U8120 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8102), .S(n6357), .Z(n6358) );
  XNOR2_X1 U8121 ( .A(n9341), .B(n6359), .ZN(n6360) );
  NAND2_X1 U8122 ( .A1(n5682), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8123 ( .A1(n5614), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8124 ( .A1(n5696), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6361) );
  NAND3_X1 U8125 ( .A1(n6363), .A2(n6362), .A3(n6361), .ZN(n9264) );
  INV_X1 U8126 ( .A(n9427), .ZN(n9968) );
  INV_X1 U8127 ( .A(P1_B_REG_SCAN_IN), .ZN(n6365) );
  OR2_X1 U8128 ( .A1(n4296), .A2(n6365), .ZN(n6366) );
  NAND2_X1 U8129 ( .A1(n9968), .A2(n6366), .ZN(n9356) );
  INV_X1 U8130 ( .A(n9356), .ZN(n6367) );
  AND2_X1 U8131 ( .A1(n9264), .A2(n6367), .ZN(n9337) );
  NOR2_X1 U8132 ( .A1(n9336), .A2(n9337), .ZN(n6373) );
  AND2_X2 U8133 ( .A1(n6369), .A2(n6368), .ZN(n10042) );
  INV_X1 U8134 ( .A(n9719), .ZN(n9715) );
  NAND2_X1 U8135 ( .A1(n6372), .A2(n6371), .ZN(P1_U3553) );
  INV_X1 U8136 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U8137 ( .A1(n6376), .A2(n6375), .ZN(P1_U3521) );
  NAND2_X1 U8138 ( .A1(n6379), .A2(n4357), .ZN(P2_U3456) );
  INV_X1 U8139 ( .A(n6642), .ZN(n6380) );
  OR2_X1 U8140 ( .A1(n8256), .A2(n6380), .ZN(n6381) );
  NAND2_X1 U8141 ( .A1(n6381), .A2(n6591), .ZN(n6575) );
  OR2_X1 U8142 ( .A1(n6575), .A2(n6382), .ZN(n6383) );
  NAND2_X1 U8143 ( .A1(n6383), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8144 ( .A(n8588), .ZN(P2_U3893) );
  INV_X1 U8145 ( .A(n6384), .ZN(n6527) );
  OR2_X2 U8146 ( .A1(n6074), .A2(n6527), .ZN(n9287) );
  INV_X1 U8147 ( .A(n9287), .ZN(P1_U3973) );
  NAND2_X1 U8148 ( .A1(n6388), .A2(P1_U3086), .ZN(n8329) );
  AND2_X1 U8149 ( .A1(n6389), .A2(P1_U3086), .ZN(n7467) );
  INV_X2 U8150 ( .A(n7467), .ZN(n9800) );
  OAI222_X1 U8151 ( .A1(n8329), .A2(n6385), .B1(n9800), .B2(n6395), .C1(
        P1_U3086), .C2(n6538), .ZN(P1_U3353) );
  OAI222_X1 U8152 ( .A1(n8329), .A2(n9028), .B1(n9800), .B2(n6397), .C1(
        P1_U3086), .C2(n9313), .ZN(P1_U3352) );
  OAI222_X1 U8153 ( .A1(n8329), .A2(n6386), .B1(n9800), .B2(n6391), .C1(
        P1_U3086), .C2(n6518), .ZN(P1_U3351) );
  INV_X1 U8154 ( .A(n8329), .ZN(n9794) );
  INV_X1 U8155 ( .A(n9794), .ZN(n9797) );
  OAI222_X1 U8156 ( .A1(n9797), .A2(n6387), .B1(n9800), .B2(n6399), .C1(
        P1_U3086), .C2(n9289), .ZN(P1_U3354) );
  OAI222_X1 U8157 ( .A1(n8329), .A2(n9027), .B1(n9800), .B2(n6393), .C1(
        P1_U3086), .C2(n9866), .ZN(P1_U3350) );
  NAND2_X1 U8158 ( .A1(n6388), .A2(P2_U3151), .ZN(n8907) );
  INV_X1 U8159 ( .A(n8907), .ZN(n7464) );
  INV_X1 U8160 ( .A(n7464), .ZN(n8331) );
  NAND2_X1 U8161 ( .A1(n6389), .A2(P2_U3151), .ZN(n8904) );
  OAI222_X1 U8162 ( .A1(n6624), .A2(P2_U3151), .B1(n8331), .B2(n6391), .C1(
        n6390), .C2(n8904), .ZN(P2_U3291) );
  OAI222_X1 U8163 ( .A1(n6585), .A2(P2_U3151), .B1(n8331), .B2(n6393), .C1(
        n6392), .C2(n8904), .ZN(P2_U3290) );
  OAI222_X1 U8164 ( .A1(n6579), .A2(P2_U3151), .B1(n8331), .B2(n6395), .C1(
        n6394), .C2(n8904), .ZN(P2_U3293) );
  OAI222_X1 U8165 ( .A1(n6720), .A2(P2_U3151), .B1(n8331), .B2(n6397), .C1(
        n6396), .C2(n8904), .ZN(P2_U3292) );
  OAI222_X1 U8166 ( .A1(n6695), .A2(P2_U3151), .B1(n8331), .B2(n6399), .C1(
        n6398), .C2(n8904), .ZN(P2_U3294) );
  OAI222_X1 U8167 ( .A1(n6798), .A2(P2_U3151), .B1(n8331), .B2(n6400), .C1(
        n9005), .C2(n8904), .ZN(P2_U3289) );
  OAI222_X1 U8168 ( .A1(n8329), .A2(n6401), .B1(n9800), .B2(n6400), .C1(
        P1_U3086), .C2(n6469), .ZN(P1_U3349) );
  NAND2_X1 U8169 ( .A1(n6403), .A2(n6402), .ZN(n6427) );
  AND2_X1 U8170 ( .A1(n6427), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8171 ( .A1(n6427), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8172 ( .A1(n6427), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8173 ( .A1(n6427), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8174 ( .A1(n6427), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8175 ( .A1(n6427), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8176 ( .A1(n6427), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8177 ( .A1(n6427), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8178 ( .A1(n6427), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8179 ( .A1(n6427), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8180 ( .A1(n6427), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8181 ( .A1(n6427), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8182 ( .A1(n6427), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  INV_X1 U8183 ( .A(n6404), .ZN(n6407) );
  OAI222_X1 U8184 ( .A1(n8329), .A2(n6405), .B1(n9800), .B2(n6407), .C1(
        P1_U3086), .C2(n6470), .ZN(P1_U3348) );
  INV_X1 U8185 ( .A(n6927), .ZN(n6939) );
  INV_X1 U8186 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6406) );
  INV_X1 U8187 ( .A(n8904), .ZN(n7749) );
  INV_X1 U8188 ( .A(n7749), .ZN(n8899) );
  OAI222_X1 U8189 ( .A1(n6939), .A2(P2_U3151), .B1(n8331), .B2(n6407), .C1(
        n6406), .C2(n8899), .ZN(P2_U3288) );
  INV_X1 U8190 ( .A(n6408), .ZN(n7751) );
  OAI222_X1 U8191 ( .A1(n8329), .A2(n6409), .B1(n9800), .B2(n7751), .C1(
        P1_U3086), .C2(n6457), .ZN(P1_U3347) );
  NOR2_X1 U8192 ( .A1(n8047), .A2(n6410), .ZN(n9992) );
  NAND2_X1 U8193 ( .A1(n9992), .A2(n6411), .ZN(n6412) );
  OAI21_X1 U8194 ( .B1(n9992), .B2(n8975), .A(n6412), .ZN(P1_U3440) );
  NAND2_X1 U8195 ( .A1(n8047), .A2(n8052), .ZN(n6437) );
  INV_X1 U8196 ( .A(n6437), .ZN(n6417) );
  NAND2_X1 U8197 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  AND2_X1 U8198 ( .A1(n6416), .A2(n6415), .ZN(n6438) );
  OR2_X1 U8199 ( .A1(n6417), .A2(n6438), .ZN(n9950) );
  INV_X1 U8200 ( .A(n9950), .ZN(n9924) );
  NOR2_X1 U8201 ( .A1(n9924), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8202 ( .A(n6418), .ZN(n6421) );
  INV_X1 U8203 ( .A(n6456), .ZN(n9836) );
  OAI222_X1 U8204 ( .A1(n9800), .A2(n6421), .B1(n9836), .B2(P1_U3086), .C1(
        n6419), .C2(n9797), .ZN(P1_U3346) );
  INV_X1 U8205 ( .A(n7134), .ZN(n7145) );
  OAI222_X1 U8206 ( .A1(P2_U3151), .A2(n7145), .B1(n8331), .B2(n6421), .C1(
        n6420), .C2(n8899), .ZN(P2_U3286) );
  INV_X1 U8207 ( .A(n6422), .ZN(n6426) );
  INV_X1 U8208 ( .A(n6487), .ZN(n6477) );
  OAI222_X1 U8209 ( .A1(n9800), .A2(n6426), .B1(n6477), .B2(P1_U3086), .C1(
        n6423), .C2(n9797), .ZN(P1_U3345) );
  NAND2_X1 U8210 ( .A1(n6783), .A2(P2_U3893), .ZN(n6424) );
  OAI21_X1 U8211 ( .B1(P2_U3893), .B2(n5620), .A(n6424), .ZN(P2_U3491) );
  INV_X1 U8212 ( .A(n7496), .ZN(n7149) );
  OAI222_X1 U8213 ( .A1(P2_U3151), .A2(n7149), .B1(n8331), .B2(n6426), .C1(
        n6425), .C2(n8899), .ZN(P2_U3285) );
  INV_X1 U8214 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6430) );
  INV_X1 U8215 ( .A(n6428), .ZN(n6429) );
  AOI22_X1 U8216 ( .A1(n6427), .A2(n6430), .B1(n6753), .B2(n6429), .ZN(
        P2_U3377) );
  INV_X1 U8217 ( .A(n6431), .ZN(n6432) );
  AOI22_X1 U8218 ( .A1(n6427), .A2(n5532), .B1(n6753), .B2(n6432), .ZN(
        P2_U3376) );
  AND2_X1 U8219 ( .A1(n6427), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8220 ( .A1(n6427), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8221 ( .A1(n6427), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8222 ( .A1(n6427), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8223 ( .A1(n6427), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8224 ( .A1(n6427), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8225 ( .A1(n6427), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8226 ( .A1(n6427), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8227 ( .A1(n6427), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8228 ( .A1(n6427), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8229 ( .A1(n6427), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8230 ( .A1(n6427), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8231 ( .A1(n6427), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8232 ( .A1(n6427), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8233 ( .A1(n6427), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8234 ( .A1(n6427), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8235 ( .A1(n6427), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  NAND2_X1 U8236 ( .A1(n5682), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8237 ( .A1(n5609), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8238 ( .A1(n5696), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6433) );
  AND3_X1 U8239 ( .A1(n6435), .A2(n6434), .A3(n6433), .ZN(n9357) );
  NAND2_X1 U8240 ( .A1(n9287), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6436) );
  OAI21_X1 U8241 ( .B1(n9357), .B2(n9287), .A(n6436), .ZN(P1_U3584) );
  NAND2_X1 U8242 ( .A1(n6438), .A2(n6437), .ZN(n9865) );
  OR2_X1 U8243 ( .A1(n9865), .A2(n6504), .ZN(n9837) );
  NOR2_X1 U8244 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9064), .ZN(n9845) );
  INV_X1 U8245 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7285) );
  INV_X1 U8246 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U8247 ( .A1(n6456), .A2(n10040), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n9836), .ZN(n9831) );
  NAND2_X1 U8248 ( .A1(n9819), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6449) );
  INV_X1 U8249 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U8250 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6439), .S(n9819), .Z(n9814)
         );
  INV_X1 U8251 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10037) );
  MUX2_X1 U8252 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10037), .S(n9808), .Z(n9806)
         );
  INV_X1 U8253 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6448) );
  MUX2_X1 U8254 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6448), .S(n9881), .Z(n9886)
         );
  INV_X1 U8255 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10035) );
  INV_X1 U8256 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6877) );
  INV_X1 U8257 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6445) );
  MUX2_X1 U8258 ( .A(n6445), .B(P1_REG1_REG_3__SCAN_IN), .S(n9313), .Z(n6444)
         );
  INV_X1 U8259 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6440) );
  MUX2_X1 U8260 ( .A(n6440), .B(P1_REG1_REG_2__SCAN_IN), .S(n6538), .Z(n6442)
         );
  MUX2_X1 U8261 ( .A(n10033), .B(P1_REG1_REG_1__SCAN_IN), .S(n9289), .Z(n9295)
         );
  AND2_X1 U8262 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9296) );
  NAND2_X1 U8263 ( .A1(n9295), .A2(n9296), .ZN(n9294) );
  INV_X1 U8264 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10033) );
  OR2_X1 U8265 ( .A1(n9289), .A2(n10033), .ZN(n6539) );
  NAND2_X1 U8266 ( .A1(n9294), .A2(n6539), .ZN(n6441) );
  NAND2_X1 U8267 ( .A1(n6442), .A2(n6441), .ZN(n9309) );
  NAND2_X1 U8268 ( .A1(n5598), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U8269 ( .A1(n9309), .A2(n9308), .ZN(n6443) );
  NAND2_X1 U8270 ( .A1(n6444), .A2(n6443), .ZN(n9312) );
  OR2_X1 U8271 ( .A1(n9313), .A2(n6445), .ZN(n6514) );
  NAND2_X1 U8272 ( .A1(n9312), .A2(n6514), .ZN(n6447) );
  MUX2_X1 U8273 ( .A(n6877), .B(P1_REG1_REG_4__SCAN_IN), .S(n6518), .Z(n6446)
         );
  NAND2_X1 U8274 ( .A1(n6447), .A2(n6446), .ZN(n6516) );
  OAI21_X1 U8275 ( .B1(n6877), .B2(n6518), .A(n6516), .ZN(n9870) );
  MUX2_X1 U8276 ( .A(n10035), .B(P1_REG1_REG_5__SCAN_IN), .S(n9866), .Z(n9869)
         );
  NAND2_X1 U8277 ( .A1(n9870), .A2(n9869), .ZN(n9868) );
  OAI21_X1 U8278 ( .B1(n10035), .B2(n9866), .A(n9868), .ZN(n9887) );
  NAND2_X1 U8279 ( .A1(n9886), .A2(n9887), .ZN(n9885) );
  OAI21_X1 U8280 ( .B1(n6469), .B2(n6448), .A(n9885), .ZN(n9807) );
  NAND2_X1 U8281 ( .A1(n9806), .A2(n9807), .ZN(n9805) );
  OAI21_X1 U8282 ( .B1(n6470), .B2(n10037), .A(n9805), .ZN(n9815) );
  NAND2_X1 U8283 ( .A1(n9814), .A2(n9815), .ZN(n9813) );
  NAND2_X1 U8284 ( .A1(n6449), .A2(n9813), .ZN(n9830) );
  NOR2_X1 U8285 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  NOR2_X1 U8286 ( .A1(n6456), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6450) );
  NOR2_X1 U8287 ( .A1(n9829), .A2(n6450), .ZN(n6453) );
  INV_X1 U8288 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6451) );
  MUX2_X1 U8289 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6451), .S(n6487), .Z(n6452)
         );
  INV_X1 U8290 ( .A(n4296), .ZN(n6502) );
  OR2_X1 U8291 ( .A1(n9865), .A2(n6502), .ZN(n9832) );
  INV_X1 U8292 ( .A(n9832), .ZN(n9941) );
  NAND2_X1 U8293 ( .A1(n6452), .A2(n6453), .ZN(n6482) );
  OAI211_X1 U8294 ( .C1(n6453), .C2(n6452), .A(n9941), .B(n6482), .ZN(n6454)
         );
  OAI21_X1 U8295 ( .B1(n9950), .B2(n7285), .A(n6454), .ZN(n6455) );
  NOR2_X1 U8296 ( .A1(n9845), .A2(n6455), .ZN(n6476) );
  INV_X1 U8297 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U8298 ( .A1(n6456), .A2(n9974), .B1(P1_REG2_REG_9__SCAN_IN), .B2(
        n9836), .ZN(n9826) );
  NAND2_X1 U8299 ( .A1(n9819), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6472) );
  INV_X1 U8300 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6458) );
  AOI22_X1 U8301 ( .A1(n9819), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6458), .B2(
        n6457), .ZN(n9818) );
  INV_X1 U8302 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6471) );
  AOI22_X1 U8303 ( .A1(n9808), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6471), .B2(
        n6470), .ZN(n9804) );
  INV_X1 U8304 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9632) );
  AOI22_X1 U8305 ( .A1(n9881), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9632), .B2(
        n6469), .ZN(n9884) );
  INV_X1 U8306 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6468) );
  INV_X1 U8307 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6509) );
  INV_X1 U8308 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6465) );
  MUX2_X1 U8309 ( .A(n6465), .B(P1_REG2_REG_3__SCAN_IN), .S(n9313), .Z(n6464)
         );
  INV_X1 U8310 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6459) );
  MUX2_X1 U8311 ( .A(n6459), .B(P1_REG2_REG_2__SCAN_IN), .S(n6538), .Z(n6462)
         );
  INV_X1 U8312 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6460) );
  MUX2_X1 U8313 ( .A(n6460), .B(P1_REG2_REG_1__SCAN_IN), .S(n9289), .Z(n9298)
         );
  AND2_X1 U8314 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9299) );
  NAND2_X1 U8315 ( .A1(n9298), .A2(n9299), .ZN(n9297) );
  OR2_X1 U8316 ( .A1(n9289), .A2(n6460), .ZN(n6535) );
  NAND2_X1 U8317 ( .A1(n9297), .A2(n6535), .ZN(n6461) );
  NAND2_X1 U8318 ( .A1(n6462), .A2(n6461), .ZN(n9304) );
  NAND2_X1 U8319 ( .A1(n5598), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U8320 ( .A1(n9304), .A2(n9303), .ZN(n6463) );
  NAND2_X1 U8321 ( .A1(n6464), .A2(n6463), .ZN(n9307) );
  OR2_X1 U8322 ( .A1(n9313), .A2(n6465), .ZN(n6510) );
  NAND2_X1 U8323 ( .A1(n9307), .A2(n6510), .ZN(n6467) );
  MUX2_X1 U8324 ( .A(n6509), .B(P1_REG2_REG_4__SCAN_IN), .S(n6518), .Z(n6466)
         );
  NAND2_X1 U8325 ( .A1(n6467), .A2(n6466), .ZN(n6512) );
  OAI21_X1 U8326 ( .B1(n6509), .B2(n6518), .A(n6512), .ZN(n9873) );
  MUX2_X1 U8327 ( .A(n6468), .B(P1_REG2_REG_5__SCAN_IN), .S(n9866), .Z(n9872)
         );
  NAND2_X1 U8328 ( .A1(n9873), .A2(n9872), .ZN(n9871) );
  OAI21_X1 U8329 ( .B1(n6468), .B2(n9866), .A(n9871), .ZN(n9883) );
  NAND2_X1 U8330 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U8331 ( .B1(n9632), .B2(n6469), .A(n9882), .ZN(n9803) );
  NAND2_X1 U8332 ( .A1(n9804), .A2(n9803), .ZN(n9802) );
  OAI21_X1 U8333 ( .B1(n6471), .B2(n6470), .A(n9802), .ZN(n9817) );
  NAND2_X1 U8334 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  NAND2_X1 U8335 ( .A1(n6472), .A2(n9816), .ZN(n9825) );
  NOR2_X1 U8336 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  AOI21_X1 U8337 ( .B1(n9836), .B2(n9974), .A(n9824), .ZN(n6474) );
  INV_X1 U8338 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7354) );
  AOI22_X1 U8339 ( .A1(n6487), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7354), .B2(
        n6477), .ZN(n6473) );
  OR2_X1 U8340 ( .A1(n7731), .A2(n4296), .ZN(n8048) );
  OR2_X1 U8341 ( .A1(n9865), .A2(n8048), .ZN(n9827) );
  INV_X1 U8342 ( .A(n9827), .ZN(n9945) );
  NAND2_X1 U8343 ( .A1(n6473), .A2(n6474), .ZN(n6488) );
  OAI211_X1 U8344 ( .C1(n6474), .C2(n6473), .A(n9945), .B(n6488), .ZN(n6475)
         );
  OAI211_X1 U8345 ( .C1(n9837), .C2(n6477), .A(n6476), .B(n6475), .ZN(P1_U3253) );
  INV_X1 U8346 ( .A(n7508), .ZN(n7519) );
  INV_X1 U8347 ( .A(n6478), .ZN(n6480) );
  OAI222_X1 U8348 ( .A1(n7519), .A2(P2_U3151), .B1(n8331), .B2(n6480), .C1(
        n6479), .C2(n8899), .ZN(P2_U3284) );
  INV_X1 U8349 ( .A(n9891), .ZN(n6486) );
  OAI222_X1 U8350 ( .A1(n8329), .A2(n6481), .B1(n9800), .B2(n6480), .C1(
        P1_U3086), .C2(n6486), .ZN(P1_U3344) );
  INV_X1 U8351 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7486) );
  MUX2_X1 U8352 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7486), .S(n9891), .Z(n9893)
         );
  NAND2_X1 U8353 ( .A1(n6487), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8354 ( .A1(n6483), .A2(n6482), .ZN(n9894) );
  NAND2_X1 U8355 ( .A1(n9893), .A2(n9894), .ZN(n9892) );
  OAI21_X1 U8356 ( .B1(n7486), .B2(n6486), .A(n9892), .ZN(n6485) );
  INV_X1 U8357 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7559) );
  INV_X1 U8358 ( .A(n6998), .ZN(n6990) );
  AOI22_X1 U8359 ( .A1(n6998), .A2(n7559), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n6990), .ZN(n6484) );
  NOR2_X1 U8360 ( .A1(n6485), .A2(n6484), .ZN(n7000) );
  AOI21_X1 U8361 ( .B1(n6485), .B2(n6484), .A(n7000), .ZN(n6498) );
  INV_X1 U8362 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U8363 ( .A1(n6998), .A2(n6989), .B1(P1_REG2_REG_12__SCAN_IN), .B2(
        n6990), .ZN(n6492) );
  NAND2_X1 U8364 ( .A1(n9891), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6490) );
  INV_X1 U8365 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U8366 ( .A1(n9891), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7400), .B2(
        n6486), .ZN(n9897) );
  NAND2_X1 U8367 ( .A1(n6487), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8368 ( .A1(n6489), .A2(n6488), .ZN(n9896) );
  NAND2_X1 U8369 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  NAND2_X1 U8370 ( .A1(n6490), .A2(n9895), .ZN(n6491) );
  NOR2_X1 U8371 ( .A1(n6492), .A2(n6491), .ZN(n6988) );
  AOI21_X1 U8372 ( .B1(n6492), .B2(n6491), .A(n6988), .ZN(n6493) );
  OR2_X1 U8373 ( .A1(n6493), .A2(n9827), .ZN(n6497) );
  AND2_X1 U8374 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6495) );
  NOR2_X1 U8375 ( .A1(n9837), .A2(n6990), .ZN(n6494) );
  AOI211_X1 U8376 ( .C1(n9924), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6495), .B(
        n6494), .ZN(n6496) );
  OAI211_X1 U8377 ( .C1(n6498), .C2(n9832), .A(n6497), .B(n6496), .ZN(P1_U3255) );
  OAI21_X1 U8378 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(n6531) );
  NOR2_X1 U8379 ( .A1(n6502), .A2(n7731), .ZN(n6508) );
  INV_X1 U8380 ( .A(n9299), .ZN(n6506) );
  OR2_X1 U8381 ( .A1(n4296), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8382 ( .A1(n6504), .A2(n6503), .ZN(n9857) );
  NAND2_X1 U8383 ( .A1(n9857), .A2(n6505), .ZN(n9860) );
  OAI211_X1 U8384 ( .C1(n6506), .C2(n8048), .A(n9860), .B(P1_U3973), .ZN(n6507) );
  AOI21_X1 U8385 ( .B1(n6531), .B2(n6508), .A(n6507), .ZN(n6547) );
  MUX2_X1 U8386 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6509), .S(n6518), .Z(n6511)
         );
  NAND3_X1 U8387 ( .A1(n6511), .A2(n9307), .A3(n6510), .ZN(n6513) );
  NAND3_X1 U8388 ( .A1(n9945), .A2(n6513), .A3(n6512), .ZN(n6524) );
  MUX2_X1 U8389 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6877), .S(n6518), .Z(n6515)
         );
  NAND3_X1 U8390 ( .A1(n6515), .A2(n9312), .A3(n6514), .ZN(n6517) );
  NAND3_X1 U8391 ( .A1(n9941), .A2(n6517), .A3(n6516), .ZN(n6523) );
  INV_X1 U8392 ( .A(n6518), .ZN(n6519) );
  NAND2_X1 U8393 ( .A1(n9943), .A2(n6519), .ZN(n6522) );
  NOR2_X1 U8394 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5634), .ZN(n6520) );
  AOI21_X1 U8395 ( .B1(n9924), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6520), .ZN(
        n6521) );
  NAND4_X1 U8396 ( .A1(n6524), .A2(n6523), .A3(n6522), .A4(n6521), .ZN(n6525)
         );
  OR2_X1 U8397 ( .A1(n6547), .A2(n6525), .ZN(P1_U3247) );
  INV_X1 U8398 ( .A(n6526), .ZN(n6532) );
  OAI222_X1 U8399 ( .A1(P2_U3151), .A2(n7706), .B1(n8331), .B2(n6532), .C1(
        n8991), .C2(n8904), .ZN(P2_U3283) );
  INV_X1 U8400 ( .A(n9237), .ZN(n9847) );
  AND2_X1 U8401 ( .A1(n6084), .A2(n9968), .ZN(n9998) );
  OR2_X1 U8402 ( .A1(n6528), .A2(n6527), .ZN(n9107) );
  AOI22_X1 U8403 ( .A1(n9847), .A2(n9998), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9107), .ZN(n6530) );
  NAND2_X1 U8404 ( .A1(n9260), .A2(n7024), .ZN(n6529) );
  OAI211_X1 U8405 ( .C1(n6531), .C2(n9262), .A(n6530), .B(n6529), .ZN(P1_U3232) );
  OAI222_X1 U8406 ( .A1(n8329), .A2(n6533), .B1(P1_U3086), .B2(n6990), .C1(
        n6532), .C2(n9800), .ZN(P1_U3343) );
  NOR2_X1 U8407 ( .A1(n9837), .A2(n6538), .ZN(n6546) );
  INV_X1 U8408 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6534) );
  INV_X1 U8409 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7737) );
  OAI22_X1 U8410 ( .A1(n9950), .A2(n6534), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7737), .ZN(n6545) );
  MUX2_X1 U8411 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6459), .S(n6538), .Z(n6536)
         );
  NAND3_X1 U8412 ( .A1(n6536), .A2(n9297), .A3(n6535), .ZN(n6537) );
  NAND2_X1 U8413 ( .A1(n6537), .A2(n9304), .ZN(n6543) );
  MUX2_X1 U8414 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6440), .S(n6538), .Z(n6540)
         );
  NAND3_X1 U8415 ( .A1(n6540), .A2(n9294), .A3(n6539), .ZN(n6541) );
  NAND2_X1 U8416 ( .A1(n6541), .A2(n9309), .ZN(n6542) );
  OAI22_X1 U8417 ( .A1(n9827), .A2(n6543), .B1(n9832), .B2(n6542), .ZN(n6544)
         );
  OR4_X1 U8418 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(P1_U3245)
         );
  INV_X1 U8419 ( .A(n7725), .ZN(n7709) );
  INV_X1 U8420 ( .A(n6548), .ZN(n6550) );
  INV_X1 U8421 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6549) );
  OAI222_X1 U8422 ( .A1(n7709), .A2(P2_U3151), .B1(n8331), .B2(n6550), .C1(
        n6549), .C2(n8904), .ZN(P2_U3282) );
  INV_X1 U8423 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6551) );
  INV_X1 U8424 ( .A(n9902), .ZN(n7002) );
  OAI222_X1 U8425 ( .A1(n8329), .A2(n6551), .B1(n9800), .B2(n6550), .C1(
        P1_U3086), .C2(n7002), .ZN(P1_U3342) );
  MUX2_X1 U8426 ( .A(n6901), .B(n6588), .S(n8318), .Z(n6552) );
  INV_X1 U8427 ( .A(n6798), .ZN(n6599) );
  NAND2_X1 U8428 ( .A1(n6552), .A2(n6599), .ZN(n6789) );
  OAI21_X1 U8429 ( .B1(n6552), .B2(n6599), .A(n6789), .ZN(n6564) );
  MUX2_X1 U8430 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8318), .Z(n6560) );
  MUX2_X1 U8431 ( .A(n6554), .B(n6553), .S(n8318), .Z(n6555) );
  MUX2_X1 U8432 ( .A(n7769), .B(n6628), .S(n8318), .Z(n7753) );
  NAND2_X1 U8433 ( .A1(n7753), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7752) );
  INV_X1 U8434 ( .A(n6555), .ZN(n6556) );
  AOI22_X1 U8435 ( .A1(n6689), .A2(n7752), .B1(n6556), .B2(n6695), .ZN(n6697)
         );
  MUX2_X1 U8436 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8318), .Z(n6557) );
  XNOR2_X1 U8437 ( .A(n6557), .B(n6579), .ZN(n6696) );
  INV_X1 U8438 ( .A(n6579), .ZN(n6709) );
  INV_X1 U8439 ( .A(n6557), .ZN(n6558) );
  MUX2_X1 U8440 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8318), .Z(n6559) );
  XNOR2_X1 U8441 ( .A(n6559), .B(n6720), .ZN(n6719) );
  NOR2_X1 U8442 ( .A1(n6718), .A2(n6719), .ZN(n6717) );
  NOR2_X1 U8443 ( .A1(n6559), .A2(n6720), .ZN(n6605) );
  XNOR2_X1 U8444 ( .A(n6560), .B(n6624), .ZN(n6604) );
  MUX2_X1 U8445 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8318), .Z(n6561) );
  XNOR2_X1 U8446 ( .A(n6561), .B(n6585), .ZN(n6733) );
  INV_X1 U8447 ( .A(n6561), .ZN(n6562) );
  AOI21_X1 U8448 ( .B1(n6564), .B2(n6563), .A(n6791), .ZN(n6602) );
  NAND2_X1 U8449 ( .A1(P2_U3893), .A2(n7748), .ZN(n10055) );
  NOR2_X1 U8450 ( .A1(n7769), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8451 ( .A1(n5047), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6566) );
  OAI21_X1 U8452 ( .B1(n6695), .B2(n6565), .A(n6566), .ZN(n6681) );
  OR2_X1 U8453 ( .A1(n6681), .A2(n6554), .ZN(n6683) );
  NAND2_X1 U8454 ( .A1(n6683), .A2(n6566), .ZN(n6702) );
  NAND2_X1 U8455 ( .A1(n6579), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8456 ( .A1(n6701), .A2(n6567), .ZN(n6568) );
  NAND2_X1 U8457 ( .A1(n6568), .A2(n6720), .ZN(n6609) );
  NAND2_X1 U8458 ( .A1(n6723), .A2(n6609), .ZN(n6570) );
  MUX2_X1 U8459 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5081), .S(n6624), .Z(n6608)
         );
  NAND2_X1 U8460 ( .A1(n6570), .A2(n6608), .ZN(n6612) );
  NAND2_X1 U8461 ( .A1(n6624), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8462 ( .A1(n6572), .A2(n6585), .ZN(n6574) );
  NAND3_X1 U8463 ( .A1(n6737), .A2(n4383), .A3(n6574), .ZN(n6576) );
  OR2_X1 U8464 ( .A1(n6575), .A2(P2_U3151), .ZN(n6597) );
  NOR2_X1 U8465 ( .A1(n6597), .A2(n7748), .ZN(n7755) );
  NAND2_X1 U8466 ( .A1(n7755), .A2(n8610), .ZN(n8620) );
  AOI21_X1 U8467 ( .B1(n6800), .B2(n6576), .A(n8620), .ZN(n6595) );
  INV_X1 U8468 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6678) );
  NOR2_X1 U8469 ( .A1(n6628), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U8470 ( .A1(n5047), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6578) );
  OAI21_X1 U8471 ( .B1(n6695), .B2(n6577), .A(n6578), .ZN(n6684) );
  OR2_X1 U8472 ( .A1(n6684), .A2(n6553), .ZN(n6686) );
  NAND2_X1 U8473 ( .A1(n6686), .A2(n6578), .ZN(n6699) );
  NAND2_X1 U8474 ( .A1(n6579), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8475 ( .A1(n6581), .A2(n6720), .ZN(n6614) );
  AND2_X1 U8476 ( .A1(n6614), .A2(n6582), .ZN(n6722) );
  NAND2_X1 U8477 ( .A1(n6721), .A2(n6614), .ZN(n6583) );
  INV_X1 U8478 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10124) );
  MUX2_X1 U8479 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10124), .S(n6624), .Z(n6613)
         );
  NAND2_X1 U8480 ( .A1(n6583), .A2(n6613), .ZN(n6617) );
  NAND2_X1 U8481 ( .A1(n6624), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6584) );
  NAND2_X1 U8482 ( .A1(n6617), .A2(n6584), .ZN(n6586) );
  NAND2_X1 U8483 ( .A1(n6586), .A2(n6585), .ZN(n6589) );
  AND2_X1 U8484 ( .A1(n6587), .A2(n6589), .ZN(n6736) );
  NAND3_X1 U8485 ( .A1(n6735), .A2(n4380), .A3(n6589), .ZN(n6590) );
  NAND2_X1 U8486 ( .A1(n7755), .A2(n8318), .ZN(n8624) );
  AOI21_X1 U8487 ( .B1(n6795), .B2(n6590), .A(n8624), .ZN(n6594) );
  AND2_X1 U8488 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7076) );
  INV_X1 U8489 ( .A(n6591), .ZN(n6592) );
  INV_X1 U8490 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7272) );
  NOR2_X1 U8491 ( .A1(n8594), .A2(n7272), .ZN(n6593) );
  NOR4_X1 U8492 ( .A1(n6595), .A2(n6594), .A3(n7076), .A4(n6593), .ZN(n6601)
         );
  NOR2_X1 U8493 ( .A1(n6597), .A2(n8318), .ZN(n6598) );
  MUX2_X1 U8494 ( .A(P2_U3893), .B(n6598), .S(n7748), .Z(n10047) );
  NAND2_X1 U8495 ( .A1(n10047), .A2(n6599), .ZN(n6600) );
  OAI211_X1 U8496 ( .C1(n6602), .C2(n10055), .A(n6601), .B(n6600), .ZN(
        P2_U3188) );
  INV_X1 U8497 ( .A(n10047), .ZN(n8587) );
  INV_X1 U8498 ( .A(n6603), .ZN(n6607) );
  INV_X1 U8499 ( .A(n10055), .ZN(n8589) );
  OAI21_X1 U8500 ( .B1(n6717), .B2(n6605), .A(n6604), .ZN(n6606) );
  NAND3_X1 U8501 ( .A1(n6607), .A2(n8589), .A3(n6606), .ZN(n6623) );
  INV_X1 U8502 ( .A(n6608), .ZN(n6610) );
  NAND3_X1 U8503 ( .A1(n6723), .A2(n6610), .A3(n6609), .ZN(n6611) );
  AOI21_X1 U8504 ( .B1(n6612), .B2(n6611), .A(n8620), .ZN(n6621) );
  INV_X1 U8505 ( .A(n6613), .ZN(n6615) );
  NAND3_X1 U8506 ( .A1(n6721), .A2(n6615), .A3(n6614), .ZN(n6616) );
  AOI21_X1 U8507 ( .B1(n6617), .B2(n6616), .A(n8624), .ZN(n6620) );
  INV_X1 U8508 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8509 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6822) );
  OAI21_X1 U8510 ( .B1(n8594), .B2(n6618), .A(n6822), .ZN(n6619) );
  NOR3_X1 U8511 ( .A1(n6621), .A2(n6620), .A3(n6619), .ZN(n6622) );
  OAI211_X1 U8512 ( .C1(n8587), .C2(n6624), .A(n6623), .B(n6622), .ZN(P2_U3186) );
  NAND2_X1 U8513 ( .A1(n10113), .A2(n8738), .ZN(n6627) );
  NAND2_X1 U8514 ( .A1(n6783), .A2(n7772), .ZN(n8106) );
  NAND2_X1 U8515 ( .A1(n6778), .A2(n8106), .ZN(n8276) );
  NAND2_X1 U8516 ( .A1(n8477), .A2(n8752), .ZN(n7765) );
  OAI21_X1 U8517 ( .B1(n10108), .B2(n7772), .A(n7765), .ZN(n6626) );
  AOI21_X1 U8518 ( .B1(n6627), .B2(n8276), .A(n6626), .ZN(n10066) );
  MUX2_X1 U8519 ( .A(n6628), .B(n10066), .S(n10135), .Z(n6629) );
  INV_X1 U8520 ( .A(n6629), .ZN(P2_U3459) );
  OAI21_X1 U8521 ( .B1(n6632), .B2(n6631), .A(n6630), .ZN(n6637) );
  INV_X1 U8522 ( .A(n6633), .ZN(n6652) );
  NAND2_X1 U8523 ( .A1(n6652), .A2(n6639), .ZN(n6635) );
  NAND4_X1 U8524 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6638)
         );
  NAND2_X1 U8525 ( .A1(n6638), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6641) );
  NOR2_X1 U8526 ( .A1(n6659), .A2(n6666), .ZN(n8320) );
  NAND2_X1 U8527 ( .A1(n8320), .A2(n6639), .ZN(n6640) );
  AND2_X1 U8528 ( .A1(n6641), .A2(n6640), .ZN(n6754) );
  OR2_X1 U8529 ( .A1(n6642), .A2(P2_U3151), .ZN(n8324) );
  OR2_X1 U8530 ( .A1(n6644), .A2(n6643), .ZN(n6645) );
  NAND3_X2 U8531 ( .A1(n6646), .A2(n6645), .A3(n8314), .ZN(n6650) );
  INV_X1 U8532 ( .A(n6778), .ZN(n6647) );
  AOI21_X1 U8533 ( .B1(n7772), .B2(n6650), .A(n6647), .ZN(n6751) );
  XNOR2_X1 U8534 ( .A(n6650), .B(n6648), .ZN(n6649) );
  XNOR2_X1 U8535 ( .A(n6649), .B(n8477), .ZN(n6752) );
  OAI22_X1 U8536 ( .A1(n6751), .A2(n6752), .B1(n8477), .B2(n6649), .ZN(n6760)
         );
  XNOR2_X1 U8537 ( .A(n6650), .B(n6916), .ZN(n6651) );
  XNOR2_X1 U8538 ( .A(n6651), .B(n8476), .ZN(n6761) );
  INV_X1 U8539 ( .A(n8476), .ZN(n6756) );
  XNOR2_X1 U8540 ( .A(n8090), .B(n10071), .ZN(n6819) );
  XNOR2_X1 U8541 ( .A(n6819), .B(n8475), .ZN(n6657) );
  NAND2_X1 U8542 ( .A1(n6658), .A2(n6657), .ZN(n6818) );
  NAND2_X1 U8543 ( .A1(n6661), .A2(n6652), .ZN(n6656) );
  INV_X1 U8544 ( .A(n6653), .ZN(n6654) );
  NAND2_X1 U8545 ( .A1(n6665), .A2(n6654), .ZN(n6655) );
  OAI211_X1 U8546 ( .C1(n6658), .C2(n6657), .A(n6818), .B(n8439), .ZN(n6673)
         );
  INV_X1 U8547 ( .A(n6659), .ZN(n6660) );
  NAND2_X1 U8548 ( .A1(n6661), .A2(n6660), .ZN(n6664) );
  INV_X1 U8549 ( .A(n6662), .ZN(n6663) );
  NAND2_X1 U8550 ( .A1(n6665), .A2(n10118), .ZN(n6668) );
  NAND2_X1 U8551 ( .A1(n6668), .A2(n8756), .ZN(n8456) );
  NAND2_X1 U8552 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6727) );
  INV_X1 U8553 ( .A(n6727), .ZN(n6669) );
  AOI21_X1 U8554 ( .B1(n8456), .B2(n7062), .A(n6669), .ZN(n6670) );
  OAI21_X1 U8555 ( .B1(n8429), .B2(n6756), .A(n6670), .ZN(n6671) );
  AOI21_X1 U8556 ( .B1(n8420), .B2(n5481), .A(n6671), .ZN(n6672) );
  OAI211_X1 U8557 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8404), .A(n6673), .B(
        n6672), .ZN(P2_U3158) );
  OAI21_X1 U8558 ( .B1(n6675), .B2(n8279), .A(n6674), .ZN(n6920) );
  INV_X1 U8559 ( .A(n8475), .ZN(n6826) );
  XNOR2_X1 U8560 ( .A(n8279), .B(n6676), .ZN(n6677) );
  OAI222_X1 U8561 ( .A1(n8775), .A2(n6826), .B1(n8773), .B2(n5025), .C1(n8738), 
        .C2(n6677), .ZN(n6919) );
  AOI21_X1 U8562 ( .B1(n10080), .B2(n6920), .A(n6919), .ZN(n6747) );
  OAI22_X1 U8563 ( .A1(n8813), .A2(n6916), .B1(n10135), .B2(n6678), .ZN(n6679)
         );
  INV_X1 U8564 ( .A(n6679), .ZN(n6680) );
  OAI21_X1 U8565 ( .B1(n6747), .B2(n10133), .A(n6680), .ZN(P2_U3461) );
  INV_X1 U8566 ( .A(n8594), .ZN(n10049) );
  NAND2_X1 U8567 ( .A1(n6681), .A2(n6554), .ZN(n6682) );
  AOI21_X1 U8568 ( .B1(n6683), .B2(n6682), .A(n8620), .ZN(n6688) );
  NAND2_X1 U8569 ( .A1(n6684), .A2(n6553), .ZN(n6685) );
  AOI21_X1 U8570 ( .B1(n6686), .B2(n6685), .A(n8624), .ZN(n6687) );
  AOI211_X1 U8571 ( .C1(n10049), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6688), .B(
        n6687), .ZN(n6694) );
  XOR2_X1 U8572 ( .A(n7752), .B(n6689), .Z(n6690) );
  NAND2_X1 U8573 ( .A1(n6690), .A2(n8589), .ZN(n6691) );
  OAI21_X1 U8574 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6780), .A(n6691), .ZN(n6692) );
  INV_X1 U8575 ( .A(n6692), .ZN(n6693) );
  OAI211_X1 U8576 ( .C1(n8587), .C2(n6695), .A(n6694), .B(n6693), .ZN(P2_U3183) );
  XNOR2_X1 U8577 ( .A(n6697), .B(n6696), .ZN(n6711) );
  INV_X1 U8578 ( .A(n8624), .ZN(n10050) );
  OAI21_X1 U8579 ( .B1(n6700), .B2(n6699), .A(n6698), .ZN(n6705) );
  INV_X1 U8580 ( .A(n8620), .ZN(n10060) );
  OAI21_X1 U8581 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n6704) );
  AOI22_X1 U8582 ( .A1(n10050), .A2(n6705), .B1(n10060), .B2(n6704), .ZN(n6707) );
  NAND2_X1 U8583 ( .A1(n10049), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n6706) );
  OAI211_X1 U8584 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6917), .A(n6707), .B(n6706), .ZN(n6708) );
  AOI21_X1 U8585 ( .B1(n6709), .B2(n10047), .A(n6708), .ZN(n6710) );
  OAI21_X1 U8586 ( .B1(n10055), .B2(n6711), .A(n6710), .ZN(P2_U3184) );
  XOR2_X1 U8587 ( .A(n6712), .B(n6713), .Z(n6716) );
  AOI22_X1 U8588 ( .A1(n9260), .A2(n6842), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9107), .ZN(n6715) );
  AOI22_X1 U8589 ( .A1(n9246), .A2(n6084), .B1(n9244), .B2(n9285), .ZN(n6714)
         );
  OAI211_X1 U8590 ( .C1(n6716), .C2(n9262), .A(n6715), .B(n6714), .ZN(P1_U3237) );
  AOI21_X1 U8591 ( .B1(n6719), .B2(n6718), .A(n6717), .ZN(n6732) );
  INV_X1 U8592 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6729) );
  OAI21_X1 U8593 ( .B1(n6722), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6721), .ZN(
        n6726) );
  OAI21_X1 U8594 ( .B1(n6724), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6723), .ZN(
        n6725) );
  AOI22_X1 U8595 ( .A1(n10050), .A2(n6726), .B1(n10060), .B2(n6725), .ZN(n6728) );
  OAI211_X1 U8596 ( .C1(n8594), .C2(n6729), .A(n6728), .B(n6727), .ZN(n6730)
         );
  AOI21_X1 U8597 ( .B1(n4391), .B2(n10047), .A(n6730), .ZN(n6731) );
  OAI21_X1 U8598 ( .B1(n6732), .B2(n10055), .A(n6731), .ZN(P2_U3185) );
  XNOR2_X1 U8599 ( .A(n6734), .B(n6733), .ZN(n6744) );
  INV_X1 U8600 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7269) );
  OAI21_X1 U8601 ( .B1(n6736), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6735), .ZN(
        n6739) );
  OAI21_X1 U8602 ( .B1(n4381), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6737), .ZN(
        n6738) );
  AOI22_X1 U8603 ( .A1(n10050), .A2(n6739), .B1(n10060), .B2(n6738), .ZN(n6741) );
  AND2_X1 U8604 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6890) );
  INV_X1 U8605 ( .A(n6890), .ZN(n6740) );
  OAI211_X1 U8606 ( .C1(n7269), .C2(n8594), .A(n6741), .B(n6740), .ZN(n6742)
         );
  AOI21_X1 U8607 ( .B1(n4393), .B2(n10047), .A(n6742), .ZN(n6743) );
  OAI21_X1 U8608 ( .B1(n6744), .B2(n10055), .A(n6743), .ZN(P2_U3187) );
  OAI22_X1 U8609 ( .A1(n6916), .A2(n8878), .B1(n10119), .B2(n5037), .ZN(n6745)
         );
  INV_X1 U8610 ( .A(n6745), .ZN(n6746) );
  OAI21_X1 U8611 ( .B1(n6747), .B2(n10121), .A(n6746), .ZN(P2_U3396) );
  INV_X1 U8612 ( .A(n6748), .ZN(n6750) );
  OAI222_X1 U8613 ( .A1(n8507), .A2(P2_U3151), .B1(n8331), .B2(n6750), .C1(
        n6749), .C2(n8904), .ZN(P2_U3281) );
  INV_X1 U8614 ( .A(n9913), .ZN(n7003) );
  OAI222_X1 U8615 ( .A1(n9797), .A2(n8967), .B1(n9800), .B2(n6750), .C1(
        P1_U3086), .C2(n7003), .ZN(P1_U3341) );
  XOR2_X1 U8616 ( .A(n6752), .B(n6751), .Z(n6759) );
  NAND2_X1 U8617 ( .A1(n6754), .A2(n6753), .ZN(n7761) );
  INV_X1 U8618 ( .A(n8429), .ZN(n8449) );
  AOI22_X1 U8619 ( .A1(n8449), .A2(n6783), .B1(n6648), .B2(n8456), .ZN(n6755)
         );
  OAI21_X1 U8620 ( .B1(n6756), .B2(n8453), .A(n6755), .ZN(n6757) );
  AOI21_X1 U8621 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7761), .A(n6757), .ZN(
        n6758) );
  OAI21_X1 U8622 ( .B1(n8458), .B2(n6759), .A(n6758), .ZN(P2_U3162) );
  XOR2_X1 U8623 ( .A(n6761), .B(n6760), .Z(n6766) );
  AOI22_X1 U8624 ( .A1(n8449), .A2(n8477), .B1(n6762), .B2(n8456), .ZN(n6763)
         );
  OAI21_X1 U8625 ( .B1(n6826), .B2(n8453), .A(n6763), .ZN(n6764) );
  AOI21_X1 U8626 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7761), .A(n6764), .ZN(
        n6765) );
  OAI21_X1 U8627 ( .B1(n6766), .B2(n8458), .A(n6765), .ZN(P2_U3177) );
  INV_X1 U8628 ( .A(n6767), .ZN(n6768) );
  NAND2_X1 U8629 ( .A1(n6769), .A2(n6768), .ZN(n6771) );
  OR2_X1 U8630 ( .A1(n6769), .A2(n5553), .ZN(n6770) );
  NAND4_X1 U8631 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6779)
         );
  AND2_X1 U8632 ( .A1(n6643), .A2(n6774), .ZN(n6975) );
  INV_X1 U8633 ( .A(n6975), .ZN(n6775) );
  AND2_X1 U8634 ( .A1(n7198), .A2(n6775), .ZN(n6776) );
  INV_X1 U8635 ( .A(n8788), .ZN(n8764) );
  XNOR2_X1 U8636 ( .A(n6778), .B(n6777), .ZN(n10070) );
  OR2_X1 U8637 ( .A1(n6779), .A2(n8682), .ZN(n8698) );
  OAI22_X1 U8638 ( .A1(n8698), .A2(n10067), .B1(n8756), .B2(n6780), .ZN(n6787)
         );
  XNOR2_X1 U8639 ( .A(n6777), .B(n6781), .ZN(n6782) );
  NAND2_X1 U8640 ( .A1(n6782), .A2(n8769), .ZN(n6785) );
  AOI22_X1 U8641 ( .A1(n8750), .A2(n6783), .B1(n8476), .B2(n8752), .ZN(n6784)
         );
  NAND2_X1 U8642 ( .A1(n6785), .A2(n6784), .ZN(n10068) );
  MUX2_X1 U8643 ( .A(n10068), .B(P2_REG2_REG_1__SCAN_IN), .S(n8767), .Z(n6786)
         );
  AOI211_X1 U8644 ( .C1(n8764), .C2(n10070), .A(n6787), .B(n6786), .ZN(n6788)
         );
  INV_X1 U8645 ( .A(n6788), .ZN(P2_U3232) );
  INV_X1 U8646 ( .A(n6789), .ZN(n6790) );
  MUX2_X1 U8647 ( .A(n6792), .B(n4576), .S(n8318), .Z(n6926) );
  XNOR2_X1 U8648 ( .A(n6926), .B(n6927), .ZN(n6793) );
  NOR2_X1 U8649 ( .A1(n6794), .A2(n6793), .ZN(n6925) );
  AOI21_X1 U8650 ( .B1(n6794), .B2(n6793), .A(n6925), .ZN(n6807) );
  NAND2_X1 U8651 ( .A1(n6796), .A2(n6939), .ZN(n10043) );
  OAI21_X1 U8652 ( .B1(n4377), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10044), .ZN(
        n6805) );
  NAND2_X1 U8653 ( .A1(n6798), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8654 ( .A1(n6800), .A2(n6799), .ZN(n6940) );
  XNOR2_X1 U8655 ( .A(n6938), .B(n6792), .ZN(n6801) );
  NOR2_X1 U8656 ( .A1(n8620), .A2(n6801), .ZN(n6804) );
  INV_X1 U8657 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8658 ( .A1(n10047), .A2(n6927), .ZN(n6802) );
  NAND2_X1 U8659 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7112) );
  OAI211_X1 U8660 ( .C1(n7275), .C2(n8594), .A(n6802), .B(n7112), .ZN(n6803)
         );
  AOI211_X1 U8661 ( .C1(n10050), .C2(n6805), .A(n6804), .B(n6803), .ZN(n6806)
         );
  OAI21_X1 U8662 ( .B1(n6807), .B2(n10055), .A(n6806), .ZN(P2_U3189) );
  INV_X1 U8663 ( .A(n6808), .ZN(n6832) );
  AOI22_X1 U8664 ( .A1(n9925), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9794), .ZN(n6809) );
  OAI21_X1 U8665 ( .B1(n6832), .B2(n9800), .A(n6809), .ZN(P1_U3340) );
  XOR2_X1 U8666 ( .A(n6810), .B(n6811), .Z(n6817) );
  OAI22_X1 U8667 ( .A1(n6813), .A2(n9427), .B1(n6812), .B2(n9956), .ZN(n6861)
         );
  AOI22_X1 U8668 ( .A1(n6861), .A2(n9847), .B1(n6814), .B2(n9260), .ZN(n6816)
         );
  MUX2_X1 U8669 ( .A(n9856), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6815) );
  OAI211_X1 U8670 ( .C1(n6817), .C2(n9262), .A(n6816), .B(n6815), .ZN(P1_U3218) );
  INV_X2 U8671 ( .A(n7534), .ZN(n8090) );
  XNOR2_X1 U8672 ( .A(n6824), .B(n8090), .ZN(n6886) );
  XNOR2_X1 U8673 ( .A(n6886), .B(n5481), .ZN(n6821) );
  OAI21_X1 U8674 ( .B1(n6826), .B2(n6819), .A(n6818), .ZN(n6820) );
  AOI21_X1 U8675 ( .B1(n6821), .B2(n6820), .A(n6887), .ZN(n6830) );
  INV_X1 U8676 ( .A(n6822), .ZN(n6823) );
  AOI21_X1 U8677 ( .B1(n8456), .B2(n6824), .A(n6823), .ZN(n6825) );
  OAI21_X1 U8678 ( .B1(n8429), .B2(n6826), .A(n6825), .ZN(n6828) );
  NOR2_X1 U8679 ( .A1(n8404), .A2(n6908), .ZN(n6827) );
  AOI211_X1 U8680 ( .C1(n8420), .C2(n8474), .A(n6828), .B(n6827), .ZN(n6829)
         );
  OAI21_X1 U8681 ( .B1(n6830), .B2(n8458), .A(n6829), .ZN(P2_U3170) );
  INV_X1 U8682 ( .A(n8524), .ZN(n8534) );
  OAI222_X1 U8683 ( .A1(P2_U3151), .A2(n8534), .B1(n8331), .B2(n6832), .C1(
        n6831), .C2(n8904), .ZN(P2_U3280) );
  INV_X1 U8684 ( .A(n9727), .ZN(n10016) );
  OR2_X1 U8685 ( .A1(n6833), .A2(n7800), .ZN(n6834) );
  NAND2_X1 U8686 ( .A1(n6835), .A2(n6834), .ZN(n7736) );
  OAI21_X1 U8687 ( .B1(n7027), .B2(n5949), .A(n9966), .ZN(n6836) );
  NOR2_X1 U8688 ( .A1(n6836), .A2(n6859), .ZN(n7739) );
  XNOR2_X1 U8689 ( .A(n7800), .B(n6837), .ZN(n6840) );
  AOI22_X1 U8690 ( .A1(n9465), .A2(n6084), .B1(n9285), .B2(n9498), .ZN(n6839)
         );
  INV_X1 U8691 ( .A(n6958), .ZN(n9615) );
  NAND2_X1 U8692 ( .A1(n7736), .A2(n9615), .ZN(n6838) );
  OAI211_X1 U8693 ( .C1(n6840), .C2(n9995), .A(n6839), .B(n6838), .ZN(n7734)
         );
  AOI211_X1 U8694 ( .C1(n10016), .C2(n7736), .A(n7739), .B(n7734), .ZN(n6844)
         );
  AOI22_X1 U8695 ( .A1(n9785), .A2(n6842), .B1(n10028), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n6841) );
  OAI21_X1 U8696 ( .B1(n6844), .B2(n10028), .A(n6841), .ZN(P1_U3459) );
  AOI22_X1 U8697 ( .A1(n9719), .A2(n6842), .B1(n10039), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6843) );
  OAI21_X1 U8698 ( .B1(n6844), .B2(n10039), .A(n6843), .ZN(P1_U3524) );
  AOI21_X1 U8699 ( .B1(n6845), .B2(n6846), .A(n9262), .ZN(n6848) );
  NAND2_X1 U8700 ( .A1(n6848), .A2(n6847), .ZN(n6852) );
  OAI22_X1 U8701 ( .A1(n9849), .A2(n6965), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5634), .ZN(n6850) );
  OAI22_X1 U8702 ( .A1(n6871), .A2(n9210), .B1(n9209), .B2(n6872), .ZN(n6849)
         );
  AOI211_X1 U8703 ( .C1(n6963), .C2(n9247), .A(n6850), .B(n6849), .ZN(n6851)
         );
  NAND2_X1 U8704 ( .A1(n6852), .A2(n6851), .ZN(P1_U3230) );
  INV_X1 U8705 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6854) );
  INV_X1 U8706 ( .A(n6853), .ZN(n6855) );
  INV_X1 U8707 ( .A(n7175), .ZN(n7171) );
  OAI222_X1 U8708 ( .A1(n9797), .A2(n6854), .B1(n9800), .B2(n6855), .C1(
        P1_U3086), .C2(n7171), .ZN(P1_U3339) );
  INV_X1 U8709 ( .A(n8547), .ZN(n8561) );
  INV_X1 U8710 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9073) );
  OAI222_X1 U8711 ( .A1(n8561), .A2(P2_U3151), .B1(n8331), .B2(n6855), .C1(
        n9073), .C2(n8904), .ZN(P2_U3279) );
  OAI21_X1 U8712 ( .B1(n6858), .B2(n6856), .A(n6857), .ZN(n7074) );
  INV_X1 U8713 ( .A(n6859), .ZN(n6860) );
  AOI211_X1 U8714 ( .C1(n6814), .C2(n6860), .A(n9617), .B(n4487), .ZN(n7068)
         );
  XNOR2_X1 U8715 ( .A(n6856), .B(n8001), .ZN(n6863) );
  INV_X1 U8716 ( .A(n6861), .ZN(n6862) );
  OAI21_X1 U8717 ( .B1(n6863), .B2(n9995), .A(n6862), .ZN(n7071) );
  AOI211_X1 U8718 ( .C1(n10026), .C2(n7074), .A(n7068), .B(n7071), .ZN(n6866)
         );
  AOI22_X1 U8719 ( .A1(n9785), .A2(n6814), .B1(n10028), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8720 ( .B1(n6866), .B2(n10028), .A(n6864), .ZN(P1_U3462) );
  AOI22_X1 U8721 ( .A1(n9719), .A2(n6814), .B1(n10039), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6865) );
  OAI21_X1 U8722 ( .B1(n6866), .B2(n10039), .A(n6865), .ZN(P1_U3525) );
  INV_X1 U8723 ( .A(n6867), .ZN(n6885) );
  AOI22_X1 U8724 ( .A1(n9944), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9794), .ZN(n6868) );
  OAI21_X1 U8725 ( .B1(n6885), .B2(n9800), .A(n6868), .ZN(P1_U3338) );
  XNOR2_X1 U8726 ( .A(n6869), .B(n7801), .ZN(n6870) );
  OAI222_X1 U8727 ( .A1(n9956), .A2(n6872), .B1(n9427), .B2(n6871), .C1(n6870), 
        .C2(n9995), .ZN(n6960) );
  AOI211_X1 U8728 ( .C1(n6874), .C2(n6873), .A(n9617), .B(n4369), .ZN(n6967)
         );
  NOR2_X1 U8729 ( .A1(n6960), .A2(n6967), .ZN(n6883) );
  OAI21_X1 U8730 ( .B1(n6876), .B2(n7801), .A(n6875), .ZN(n6953) );
  NAND2_X1 U8731 ( .A1(n10042), .A2(n10026), .ZN(n9721) );
  INV_X1 U8732 ( .A(n9721), .ZN(n7599) );
  OAI22_X1 U8733 ( .A1(n9715), .A2(n6965), .B1(n10042), .B2(n6877), .ZN(n6878)
         );
  AOI21_X1 U8734 ( .B1(n6953), .B2(n7599), .A(n6878), .ZN(n6879) );
  OAI21_X1 U8735 ( .B1(n6883), .B2(n10039), .A(n6879), .ZN(P1_U3526) );
  INV_X1 U8736 ( .A(n9787), .ZN(n7596) );
  INV_X1 U8737 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6880) );
  OAI22_X1 U8738 ( .A1(n9781), .A2(n6965), .B1(n10030), .B2(n6880), .ZN(n6881)
         );
  AOI21_X1 U8739 ( .B1(n6953), .B2(n7596), .A(n6881), .ZN(n6882) );
  OAI21_X1 U8740 ( .B1(n6883), .B2(n10028), .A(n6882), .ZN(P1_U3465) );
  INV_X1 U8741 ( .A(n8596), .ZN(n8569) );
  OAI222_X1 U8742 ( .A1(n8569), .A2(P2_U3151), .B1(n8331), .B2(n6885), .C1(
        n6884), .C2(n8904), .ZN(P2_U3278) );
  XNOR2_X1 U8743 ( .A(n8090), .B(n10081), .ZN(n7079) );
  XNOR2_X1 U8744 ( .A(n7079), .B(n8474), .ZN(n7080) );
  INV_X1 U8745 ( .A(n6886), .ZN(n6888) );
  INV_X1 U8746 ( .A(n5481), .ZN(n6893) );
  XOR2_X1 U8747 ( .A(n7080), .B(n4373), .Z(n6896) );
  INV_X1 U8748 ( .A(n6889), .ZN(n6983) );
  OR2_X1 U8749 ( .A1(n8453), .A2(n7113), .ZN(n6892) );
  AOI21_X1 U8750 ( .B1(n8456), .B2(n10081), .A(n6890), .ZN(n6891) );
  OAI211_X1 U8751 ( .C1(n6893), .C2(n8429), .A(n6892), .B(n6891), .ZN(n6894)
         );
  AOI21_X1 U8752 ( .B1(n8450), .B2(n6983), .A(n6894), .ZN(n6895) );
  OAI21_X1 U8753 ( .B1(n6896), .B2(n8458), .A(n6895), .ZN(P2_U3167) );
  NAND2_X1 U8754 ( .A1(n6897), .A2(n8123), .ZN(n6898) );
  NAND2_X1 U8755 ( .A1(n8127), .A2(n8143), .ZN(n8281) );
  XNOR2_X1 U8756 ( .A(n6898), .B(n8281), .ZN(n10089) );
  XNOR2_X1 U8757 ( .A(n6899), .B(n8281), .ZN(n6900) );
  AOI222_X1 U8758 ( .A1(n8769), .A2(n6900), .B1(n8474), .B2(n8750), .C1(n8472), 
        .C2(n8752), .ZN(n10087) );
  MUX2_X1 U8759 ( .A(n6901), .B(n10087), .S(n8780), .Z(n6905) );
  INV_X1 U8760 ( .A(n8756), .ZN(n8784) );
  INV_X1 U8761 ( .A(n6902), .ZN(n7085) );
  AOI22_X1 U8762 ( .A1(n8785), .A2(n6903), .B1(n8784), .B2(n7085), .ZN(n6904)
         );
  OAI211_X1 U8763 ( .C1(n8788), .C2(n10089), .A(n6905), .B(n6904), .ZN(
        P2_U3227) );
  OAI21_X1 U8764 ( .B1(n6906), .B2(n8120), .A(n6907), .ZN(n10079) );
  OAI22_X1 U8765 ( .A1(n8698), .A2(n10076), .B1(n6908), .B2(n8756), .ZN(n6914)
         );
  NAND2_X1 U8766 ( .A1(n6909), .A2(n8283), .ZN(n6977) );
  OAI21_X1 U8767 ( .B1(n8283), .B2(n6909), .A(n6977), .ZN(n6910) );
  NAND2_X1 U8768 ( .A1(n6910), .A2(n8769), .ZN(n6912) );
  AOI22_X1 U8769 ( .A1(n8752), .A2(n8474), .B1(n8475), .B2(n8750), .ZN(n6911)
         );
  NAND2_X1 U8770 ( .A1(n6912), .A2(n6911), .ZN(n10077) );
  MUX2_X1 U8771 ( .A(n10077), .B(P2_REG2_REG_4__SCAN_IN), .S(n8767), .Z(n6913)
         );
  AOI211_X1 U8772 ( .C1(n8764), .C2(n10079), .A(n6914), .B(n6913), .ZN(n6915)
         );
  INV_X1 U8773 ( .A(n6915), .ZN(P2_U3229) );
  OAI22_X1 U8774 ( .A1(n8756), .A2(n6917), .B1(n6916), .B2(n8682), .ZN(n6918)
         );
  OAI21_X1 U8775 ( .B1(n6919), .B2(n6918), .A(n8780), .ZN(n6922) );
  NAND2_X1 U8776 ( .A1(n8764), .A2(n6920), .ZN(n6921) );
  OAI211_X1 U8777 ( .C1(n5040), .C2(n8780), .A(n6922), .B(n6921), .ZN(P2_U3231) );
  INV_X1 U8778 ( .A(n8613), .ZN(n8618) );
  INV_X1 U8779 ( .A(n6923), .ZN(n6971) );
  OAI222_X1 U8780 ( .A1(P2_U3151), .A2(n8618), .B1(n8331), .B2(n6971), .C1(
        n6924), .C2(n8904), .ZN(P2_U3277) );
  INV_X1 U8781 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10129) );
  MUX2_X1 U8782 ( .A(n6943), .B(n10129), .S(n8318), .Z(n6928) );
  NAND2_X1 U8783 ( .A1(n6928), .A2(n10048), .ZN(n6929) );
  OAI21_X1 U8784 ( .B1(n6928), .B2(n10048), .A(n6929), .ZN(n10053) );
  INV_X1 U8785 ( .A(n6929), .ZN(n6930) );
  MUX2_X1 U8786 ( .A(n6932), .B(n6931), .S(n8318), .Z(n7133) );
  XNOR2_X1 U8787 ( .A(n7133), .B(n7134), .ZN(n6933) );
  AOI21_X1 U8788 ( .B1(n6934), .B2(n6933), .A(n7132), .ZN(n6952) );
  OR2_X1 U8789 ( .A1(n10048), .A2(n10129), .ZN(n6935) );
  NAND2_X1 U8790 ( .A1(n10046), .A2(n6935), .ZN(n7139) );
  OAI21_X1 U8791 ( .B1(n6936), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7141), .ZN(
        n6950) );
  AND2_X1 U8792 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7324) );
  AOI21_X1 U8793 ( .B1(n10049), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7324), .ZN(
        n6937) );
  OAI21_X1 U8794 ( .B1(n8587), .B2(n7145), .A(n6937), .ZN(n6949) );
  NAND2_X1 U8795 ( .A1(n6938), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6942) );
  NAND2_X1 U8796 ( .A1(n6940), .A2(n6939), .ZN(n6941) );
  NAND2_X1 U8797 ( .A1(n6942), .A2(n6941), .ZN(n10058) );
  XNOR2_X1 U8798 ( .A(n10048), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U8799 ( .A1(n10058), .A2(n10059), .ZN(n10057) );
  OR2_X1 U8800 ( .A1(n10048), .A2(n6943), .ZN(n6944) );
  NAND2_X1 U8801 ( .A1(n10057), .A2(n6944), .ZN(n7146) );
  XNOR2_X1 U8802 ( .A(n7146), .B(n7134), .ZN(n6946) );
  INV_X1 U8803 ( .A(n6946), .ZN(n6945) );
  NAND2_X1 U8804 ( .A1(n6945), .A2(n6932), .ZN(n6947) );
  AOI21_X1 U8805 ( .B1(n6947), .B2(n7148), .A(n8620), .ZN(n6948) );
  AOI211_X1 U8806 ( .C1(n10050), .C2(n6950), .A(n6949), .B(n6948), .ZN(n6951)
         );
  OAI21_X1 U8807 ( .B1(n6952), .B2(n10055), .A(n6951), .ZN(P2_U3191) );
  INV_X1 U8808 ( .A(n6953), .ZN(n6970) );
  NAND3_X1 U8809 ( .A1(n6956), .A2(n6955), .A3(n6954), .ZN(n6957) );
  NAND2_X1 U8810 ( .A1(n6958), .A2(n7030), .ZN(n6959) );
  INV_X1 U8811 ( .A(n6960), .ZN(n6961) );
  MUX2_X1 U8812 ( .A(n6509), .B(n6961), .S(n9984), .Z(n6969) );
  NAND2_X2 U8813 ( .A1(n9984), .A2(n6962), .ZN(n9622) );
  INV_X1 U8814 ( .A(n6963), .ZN(n6964) );
  OAI22_X1 U8815 ( .A1(n9622), .A2(n6965), .B1(n9978), .B2(n6964), .ZN(n6966)
         );
  AOI21_X1 U8816 ( .B1(n6967), .B2(n9637), .A(n6966), .ZN(n6968) );
  OAI211_X1 U8817 ( .C1(n6970), .C2(n9606), .A(n6969), .B(n6968), .ZN(P1_U3289) );
  INV_X1 U8818 ( .A(n9322), .ZN(n7183) );
  OAI222_X1 U8819 ( .A1(n8329), .A2(n6972), .B1(n7183), .B2(P1_U3086), .C1(
        n9800), .C2(n6971), .ZN(P1_U3337) );
  XNOR2_X1 U8820 ( .A(n8474), .B(n6973), .ZN(n8282) );
  XOR2_X1 U8821 ( .A(n6974), .B(n8282), .Z(n10083) );
  INV_X1 U8822 ( .A(n10083), .ZN(n6986) );
  NAND2_X1 U8823 ( .A1(n8780), .A2(n6975), .ZN(n8334) );
  INV_X1 U8824 ( .A(n7198), .ZN(n6982) );
  NAND2_X1 U8825 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  XOR2_X1 U8826 ( .A(n6978), .B(n8282), .Z(n6980) );
  AOI22_X1 U8827 ( .A1(n8473), .A2(n8752), .B1(n8750), .B2(n5481), .ZN(n6979)
         );
  OAI21_X1 U8828 ( .B1(n6980), .B2(n8738), .A(n6979), .ZN(n6981) );
  AOI21_X1 U8829 ( .B1(n6982), .B2(n10083), .A(n6981), .ZN(n10085) );
  MUX2_X1 U8830 ( .A(n4708), .B(n10085), .S(n8780), .Z(n6985) );
  AOI22_X1 U8831 ( .A1(n8785), .A2(n10081), .B1(n8784), .B2(n6983), .ZN(n6984)
         );
  OAI211_X1 U8832 ( .C1(n6986), .C2(n8334), .A(n6985), .B(n6984), .ZN(P2_U3228) );
  INV_X1 U8833 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U8834 ( .A1(n7175), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n6987), .B2(
        n7171), .ZN(n6995) );
  INV_X1 U8835 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U8836 ( .A1(n9913), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n6991), .B2(
        n7003), .ZN(n9916) );
  INV_X1 U8837 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7572) );
  AOI22_X1 U8838 ( .A1(n9902), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7572), .B2(
        n7002), .ZN(n9908) );
  AOI21_X1 U8839 ( .B1(n6990), .B2(n6989), .A(n6988), .ZN(n9907) );
  NAND2_X1 U8840 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  OAI21_X1 U8841 ( .B1(n7572), .B2(n7002), .A(n9906), .ZN(n9915) );
  NAND2_X1 U8842 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  OAI21_X1 U8843 ( .B1(n6991), .B2(n7003), .A(n9914), .ZN(n6992) );
  NAND2_X1 U8844 ( .A1(n9925), .A2(n6992), .ZN(n6993) );
  XOR2_X1 U8845 ( .A(n9925), .B(n6992), .Z(n9929) );
  NAND2_X1 U8846 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9929), .ZN(n9928) );
  NAND2_X1 U8847 ( .A1(n6993), .A2(n9928), .ZN(n6994) );
  NAND2_X1 U8848 ( .A1(n6995), .A2(n6994), .ZN(n7176) );
  OAI21_X1 U8849 ( .B1(n6995), .B2(n6994), .A(n7176), .ZN(n7012) );
  NOR2_X1 U8850 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9150), .ZN(n6997) );
  NOR2_X1 U8851 ( .A1(n9837), .A2(n7171), .ZN(n6996) );
  AOI211_X1 U8852 ( .C1(n9924), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n6997), .B(
        n6996), .ZN(n7011) );
  INV_X1 U8853 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U8854 ( .A1(n7175), .A2(n9713), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n7171), .ZN(n7008) );
  INV_X1 U8855 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7004) );
  XNOR2_X1 U8856 ( .A(n7003), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9919) );
  INV_X1 U8857 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7001) );
  XNOR2_X1 U8858 ( .A(n9902), .B(n7001), .ZN(n9904) );
  NOR2_X1 U8859 ( .A1(n6998), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8860 ( .A1(n7000), .A2(n6999), .ZN(n9905) );
  NAND2_X1 U8861 ( .A1(n9904), .A2(n9905), .ZN(n9903) );
  OAI21_X1 U8862 ( .B1(n7002), .B2(n7001), .A(n9903), .ZN(n9918) );
  NAND2_X1 U8863 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  OAI21_X1 U8864 ( .B1(n7004), .B2(n7003), .A(n9917), .ZN(n7005) );
  NAND2_X1 U8865 ( .A1(n9925), .A2(n7005), .ZN(n7006) );
  XOR2_X1 U8866 ( .A(n7005), .B(n9925), .Z(n9927) );
  NAND2_X1 U8867 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9927), .ZN(n9926) );
  NAND2_X1 U8868 ( .A1(n7006), .A2(n9926), .ZN(n7007) );
  NOR2_X1 U8869 ( .A1(n7008), .A2(n7007), .ZN(n7170) );
  AOI21_X1 U8870 ( .B1(n7008), .B2(n7007), .A(n7170), .ZN(n7009) );
  OR2_X1 U8871 ( .A1(n7009), .A2(n9832), .ZN(n7010) );
  OAI211_X1 U8872 ( .C1(n7012), .C2(n9827), .A(n7011), .B(n7010), .ZN(P1_U3259) );
  INV_X1 U8873 ( .A(n7802), .ZN(n7013) );
  NAND2_X1 U8874 ( .A1(n7013), .A2(n5990), .ZN(n7015) );
  NAND2_X1 U8875 ( .A1(n7015), .A2(n7014), .ZN(n7019) );
  NAND2_X1 U8876 ( .A1(n9288), .A2(n9465), .ZN(n7017) );
  NAND2_X1 U8877 ( .A1(n9286), .A2(n9498), .ZN(n7016) );
  NAND2_X1 U8878 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  AOI21_X1 U8879 ( .B1(n7019), .B2(n9595), .A(n7018), .ZN(n7023) );
  OAI21_X1 U8880 ( .B1(n5990), .B2(n7021), .A(n7020), .ZN(n10003) );
  NAND2_X1 U8881 ( .A1(n10003), .A2(n9615), .ZN(n7022) );
  AND2_X1 U8882 ( .A1(n7023), .A2(n7022), .ZN(n10005) );
  INV_X1 U8883 ( .A(n9622), .ZN(n9635) );
  INV_X1 U8884 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9290) );
  OAI22_X1 U8885 ( .A1(n9978), .A2(n9290), .B1(n6460), .B2(n9984), .ZN(n7029)
         );
  NAND2_X1 U8886 ( .A1(n6085), .A2(n7024), .ZN(n7025) );
  NAND2_X1 U8887 ( .A1(n7025), .A2(n9966), .ZN(n7026) );
  OR2_X1 U8888 ( .A1(n7027), .A2(n7026), .ZN(n10001) );
  NOR2_X1 U8889 ( .A1(n9970), .A2(n10001), .ZN(n7028) );
  AOI211_X1 U8890 ( .C1(n9635), .C2(n6085), .A(n7029), .B(n7028), .ZN(n7033)
         );
  INV_X1 U8891 ( .A(n7030), .ZN(n7031) );
  NAND2_X1 U8892 ( .A1(n9984), .A2(n7031), .ZN(n9625) );
  INV_X1 U8893 ( .A(n9625), .ZN(n7735) );
  NAND2_X1 U8894 ( .A1(n10003), .A2(n7735), .ZN(n7032) );
  OAI211_X1 U8895 ( .C1(n10005), .C2(n9987), .A(n7033), .B(n7032), .ZN(
        P1_U3292) );
  NAND2_X1 U8896 ( .A1(n8588), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7034) );
  OAI21_X1 U8897 ( .B1(n8097), .B2(n8588), .A(n7034), .ZN(P2_U3520) );
  OR2_X1 U8898 ( .A1(n7036), .A2(n8287), .ZN(n7037) );
  NAND2_X1 U8899 ( .A1(n7035), .A2(n7037), .ZN(n10094) );
  XNOR2_X1 U8900 ( .A(n7038), .B(n8287), .ZN(n7039) );
  NAND2_X1 U8901 ( .A1(n7039), .A2(n8769), .ZN(n7041) );
  AOI22_X1 U8902 ( .A1(n8473), .A2(n8750), .B1(n8752), .B2(n8471), .ZN(n7040)
         );
  OAI211_X1 U8903 ( .C1(n7198), .C2(n10094), .A(n7041), .B(n7040), .ZN(n10096)
         );
  NAND2_X1 U8904 ( .A1(n10096), .A2(n8780), .ZN(n7045) );
  OAI22_X1 U8905 ( .A1(n8780), .A2(n6792), .B1(n7114), .B2(n8756), .ZN(n7042)
         );
  AOI21_X1 U8906 ( .B1(n8785), .B2(n7043), .A(n7042), .ZN(n7044) );
  OAI211_X1 U8907 ( .C1(n10094), .C2(n8334), .A(n7045), .B(n7044), .ZN(
        P2_U3226) );
  OAI21_X1 U8908 ( .B1(n7047), .B2(n7808), .A(n7046), .ZN(n9636) );
  NAND2_X1 U8909 ( .A1(n7090), .A2(n9634), .ZN(n7048) );
  NAND2_X1 U8910 ( .A1(n7048), .A2(n9966), .ZN(n7049) );
  NOR2_X1 U8911 ( .A1(n7228), .A2(n7049), .ZN(n9638) );
  XNOR2_X1 U8912 ( .A(n7050), .B(n7808), .ZN(n7053) );
  NAND2_X1 U8913 ( .A1(n9283), .A2(n9465), .ZN(n7052) );
  NAND2_X1 U8914 ( .A1(n9281), .A2(n9498), .ZN(n7051) );
  AND2_X1 U8915 ( .A1(n7052), .A2(n7051), .ZN(n7310) );
  OAI21_X1 U8916 ( .B1(n7053), .B2(n9995), .A(n7310), .ZN(n9629) );
  AOI211_X1 U8917 ( .C1(n10026), .C2(n9636), .A(n9638), .B(n9629), .ZN(n7056)
         );
  AOI22_X1 U8918 ( .A1(n9719), .A2(n9634), .B1(n10039), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7054) );
  OAI21_X1 U8919 ( .B1(n7056), .B2(n10039), .A(n7054), .ZN(P1_U3528) );
  AOI22_X1 U8920 ( .A1(n9785), .A2(n9634), .B1(n10028), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n7055) );
  OAI21_X1 U8921 ( .B1(n7056), .B2(n10028), .A(n7055), .ZN(P1_U3471) );
  INV_X1 U8922 ( .A(n8278), .ZN(n7058) );
  XNOR2_X1 U8923 ( .A(n7057), .B(n7058), .ZN(n7059) );
  NAND2_X1 U8924 ( .A1(n7059), .A2(n8769), .ZN(n7061) );
  AOI22_X1 U8925 ( .A1(n8750), .A2(n8476), .B1(n5481), .B2(n8752), .ZN(n7060)
         );
  NAND2_X1 U8926 ( .A1(n7061), .A2(n7060), .ZN(n10073) );
  AOI22_X1 U8927 ( .A1(n8785), .A2(n7062), .B1(n4981), .B2(n8784), .ZN(n7063)
         );
  OAI21_X1 U8928 ( .B1(n5055), .B2(n8780), .A(n7063), .ZN(n7066) );
  XOR2_X1 U8929 ( .A(n7064), .B(n8278), .Z(n10072) );
  NOR2_X1 U8930 ( .A1(n10072), .A2(n8788), .ZN(n7065) );
  AOI211_X1 U8931 ( .C1(n8780), .C2(n10073), .A(n7066), .B(n7065), .ZN(n7067)
         );
  INV_X1 U8932 ( .A(n7067), .ZN(P2_U3230) );
  INV_X1 U8933 ( .A(n9606), .ZN(n9964) );
  INV_X1 U8934 ( .A(n7068), .ZN(n7070) );
  INV_X1 U8935 ( .A(n9978), .ZN(n9619) );
  AOI22_X1 U8936 ( .A1(n9635), .A2(n6814), .B1(n5624), .B2(n9619), .ZN(n7069)
         );
  OAI21_X1 U8937 ( .B1(n7070), .B2(n9970), .A(n7069), .ZN(n7073) );
  MUX2_X1 U8938 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7071), .S(n9984), .Z(n7072)
         );
  AOI211_X1 U8939 ( .C1(n9964), .C2(n7074), .A(n7073), .B(n7072), .ZN(n7075)
         );
  INV_X1 U8940 ( .A(n7075), .ZN(P1_U3290) );
  INV_X1 U8941 ( .A(n8456), .ZN(n8446) );
  AOI21_X1 U8942 ( .B1(n8449), .B2(n8474), .A(n7076), .ZN(n7078) );
  NAND2_X1 U8943 ( .A1(n8420), .A2(n8472), .ZN(n7077) );
  OAI211_X1 U8944 ( .C1(n10088), .C2(n8446), .A(n7078), .B(n7077), .ZN(n7084)
         );
  XNOR2_X1 U8945 ( .A(n8090), .B(n10088), .ZN(n7106) );
  XNOR2_X1 U8946 ( .A(n7106), .B(n7113), .ZN(n7082) );
  AOI211_X1 U8947 ( .C1(n7082), .C2(n7081), .A(n8458), .B(n7108), .ZN(n7083)
         );
  AOI211_X1 U8948 ( .C1(n7085), .C2(n8450), .A(n7084), .B(n7083), .ZN(n7086)
         );
  INV_X1 U8949 ( .A(n7086), .ZN(P2_U3179) );
  OAI21_X1 U8950 ( .B1(n7089), .B2(n7088), .A(n7087), .ZN(n10011) );
  OAI211_X1 U8951 ( .C1(n4369), .C2(n10008), .A(n9966), .B(n7090), .ZN(n10007)
         );
  AOI22_X1 U8952 ( .A1(n9635), .A2(n9159), .B1(n9160), .B2(n9619), .ZN(n7091)
         );
  OAI21_X1 U8953 ( .B1(n10007), .B2(n9970), .A(n7091), .ZN(n7097) );
  XNOR2_X1 U8954 ( .A(n7092), .B(n7807), .ZN(n7093) );
  NAND2_X1 U8955 ( .A1(n7093), .A2(n9595), .ZN(n7095) );
  AOI22_X1 U8956 ( .A1(n9465), .A2(n9284), .B1(n9282), .B2(n9498), .ZN(n7094)
         );
  NAND2_X1 U8957 ( .A1(n7095), .A2(n7094), .ZN(n10009) );
  MUX2_X1 U8958 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10009), .S(n9984), .Z(n7096)
         );
  AOI211_X1 U8959 ( .C1(n9964), .C2(n10011), .A(n7097), .B(n7096), .ZN(n7098)
         );
  INV_X1 U8960 ( .A(n7098), .ZN(P1_U3288) );
  NAND2_X1 U8961 ( .A1(n7035), .A2(n7099), .ZN(n7100) );
  AND2_X1 U8962 ( .A1(n8126), .A2(n8146), .ZN(n8286) );
  XNOR2_X1 U8963 ( .A(n7100), .B(n8286), .ZN(n10099) );
  XOR2_X1 U8964 ( .A(n7101), .B(n8286), .Z(n7102) );
  OAI222_X1 U8965 ( .A1(n8775), .A2(n7418), .B1(n8773), .B2(n7237), .C1(n7102), 
        .C2(n8738), .ZN(n10101) );
  NAND2_X1 U8966 ( .A1(n10101), .A2(n8780), .ZN(n7105) );
  OAI22_X1 U8967 ( .A1(n8780), .A2(n6943), .B1(n7242), .B2(n8756), .ZN(n7103)
         );
  AOI21_X1 U8968 ( .B1(n8785), .B2(n7244), .A(n7103), .ZN(n7104) );
  OAI211_X1 U8969 ( .C1(n10099), .C2(n8788), .A(n7105), .B(n7104), .ZN(
        P2_U3225) );
  XNOR2_X1 U8970 ( .A(n10093), .B(n8090), .ZN(n7236) );
  XNOR2_X1 U8971 ( .A(n7236), .B(n8472), .ZN(n7110) );
  INV_X1 U8972 ( .A(n7106), .ZN(n7107) );
  NOR2_X1 U8973 ( .A1(n7108), .A2(n4333), .ZN(n7109) );
  NAND2_X1 U8974 ( .A1(n7109), .A2(n7110), .ZN(n7239) );
  OAI21_X1 U8975 ( .B1(n7110), .B2(n7109), .A(n7239), .ZN(n7111) );
  NAND2_X1 U8976 ( .A1(n7111), .A2(n8439), .ZN(n7118) );
  OAI21_X1 U8977 ( .B1(n8429), .B2(n7113), .A(n7112), .ZN(n7116) );
  NOR2_X1 U8978 ( .A1(n8404), .A2(n7114), .ZN(n7115) );
  AOI211_X1 U8979 ( .C1(n8420), .C2(n8471), .A(n7116), .B(n7115), .ZN(n7117)
         );
  OAI211_X1 U8980 ( .C1(n10093), .C2(n8446), .A(n7118), .B(n7117), .ZN(
        P2_U3153) );
  INV_X1 U8981 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7125) );
  NAND2_X1 U8982 ( .A1(n7119), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7123) );
  INV_X1 U8983 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7120) );
  OR2_X1 U8984 ( .A1(n7121), .A2(n7120), .ZN(n7122) );
  OAI211_X1 U8985 ( .C1(n7125), .C2(n7124), .A(n7123), .B(n7122), .ZN(n7126)
         );
  INV_X1 U8986 ( .A(n7126), .ZN(n7127) );
  INV_X1 U8987 ( .A(n8628), .ZN(n8313) );
  NAND2_X1 U8988 ( .A1(n8313), .A2(P2_U3893), .ZN(n7129) );
  OAI21_X1 U8989 ( .B1(P2_U3893), .B2(n6353), .A(n7129), .ZN(P2_U3522) );
  INV_X1 U8990 ( .A(n7130), .ZN(n7235) );
  OAI222_X1 U8991 ( .A1(n8329), .A2(n7131), .B1(n9800), .B2(n7235), .C1(
        P1_U3086), .C2(n6035), .ZN(P1_U3336) );
  AOI21_X1 U8992 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7138) );
  INV_X1 U8993 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7495) );
  MUX2_X1 U8994 ( .A(n7489), .B(n7495), .S(n8318), .Z(n7136) );
  AND2_X1 U8995 ( .A1(n7136), .A2(n7496), .ZN(n7510) );
  INV_X1 U8996 ( .A(n7510), .ZN(n7135) );
  OAI21_X1 U8997 ( .B1(n7496), .B2(n7136), .A(n7135), .ZN(n7137) );
  AOI21_X1 U8998 ( .B1(n7138), .B2(n7137), .A(n7509), .ZN(n7159) );
  NAND2_X1 U8999 ( .A1(n7139), .A2(n7145), .ZN(n7140) );
  AOI22_X1 U9000 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7496), .B1(n7149), .B2(
        n7495), .ZN(n7142) );
  AOI21_X1 U9001 ( .B1(n4376), .B2(n7142), .A(n7497), .ZN(n7156) );
  INV_X1 U9002 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7284) );
  INV_X1 U9003 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U9004 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9077), .ZN(n7423) );
  INV_X1 U9005 ( .A(n7423), .ZN(n7143) );
  OAI21_X1 U9006 ( .B1(n8594), .B2(n7284), .A(n7143), .ZN(n7144) );
  AOI21_X1 U9007 ( .B1(n7496), .B2(n10047), .A(n7144), .ZN(n7155) );
  NAND2_X1 U9008 ( .A1(n7146), .A2(n7145), .ZN(n7147) );
  AOI22_X1 U9009 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7496), .B1(n7149), .B2(
        n7489), .ZN(n7151) );
  AOI21_X1 U9010 ( .B1(n7152), .B2(n7151), .A(n7150), .ZN(n7153) );
  OR2_X1 U9011 ( .A1(n7153), .A2(n8620), .ZN(n7154) );
  OAI211_X1 U9012 ( .C1(n7156), .C2(n8624), .A(n7155), .B(n7154), .ZN(n7157)
         );
  INV_X1 U9013 ( .A(n7157), .ZN(n7158) );
  OAI21_X1 U9014 ( .B1(n7159), .B2(n10055), .A(n7158), .ZN(P2_U3192) );
  XOR2_X1 U9015 ( .A(n7160), .B(n7161), .Z(n7169) );
  INV_X1 U9016 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7162) );
  OAI22_X1 U9017 ( .A1(n9209), .A2(n7163), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7162), .ZN(n7166) );
  OAI22_X1 U9018 ( .A1(n9957), .A2(n9210), .B1(n9856), .B2(n7164), .ZN(n7165)
         );
  AOI211_X1 U9019 ( .C1(n7167), .C2(n9260), .A(n7166), .B(n7165), .ZN(n7168)
         );
  OAI21_X1 U9020 ( .B1(n7169), .B2(n9262), .A(n7168), .ZN(P1_U3213) );
  AOI21_X1 U9021 ( .B1(n7171), .B2(n9713), .A(n7170), .ZN(n9938) );
  XNOR2_X1 U9022 ( .A(n9944), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9937) );
  OR2_X1 U9023 ( .A1(n9938), .A2(n9937), .ZN(n9940) );
  OR2_X1 U9024 ( .A1(n9944), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7172) );
  INV_X1 U9025 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9704) );
  XNOR2_X1 U9026 ( .A(n9322), .B(n9704), .ZN(n7173) );
  AOI21_X1 U9027 ( .B1(n9940), .B2(n7172), .A(n7173), .ZN(n7190) );
  AND2_X1 U9028 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  NAND2_X1 U9029 ( .A1(n9940), .A2(n7174), .ZN(n9324) );
  NAND2_X1 U9030 ( .A1(n9324), .A2(n9941), .ZN(n7189) );
  NAND2_X1 U9031 ( .A1(n7175), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7177) );
  AND2_X1 U9032 ( .A1(n7177), .A2(n7176), .ZN(n9935) );
  OR2_X1 U9033 ( .A1(n9944), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U9034 ( .A1(n9944), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7178) );
  AND2_X1 U9035 ( .A1(n7179), .A2(n7178), .ZN(n9936) );
  NAND2_X1 U9036 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  NAND2_X1 U9037 ( .A1(n9934), .A2(n7179), .ZN(n7182) );
  NAND2_X1 U9038 ( .A1(n9322), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9319) );
  OAI21_X1 U9039 ( .B1(n9322), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9319), .ZN(
        n7180) );
  OR2_X1 U9040 ( .A1(n7182), .A2(n7180), .ZN(n9320) );
  NAND2_X1 U9041 ( .A1(n7183), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7181) );
  OAI211_X1 U9042 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n7183), .A(n7182), .B(
        n7181), .ZN(n7184) );
  NAND3_X1 U9043 ( .A1(n9320), .A2(n7184), .A3(n9945), .ZN(n7188) );
  INV_X1 U9044 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U9045 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9236) );
  OAI21_X1 U9046 ( .B1(n9950), .B2(n7185), .A(n9236), .ZN(n7186) );
  AOI21_X1 U9047 ( .B1(n9322), .B2(n9943), .A(n7186), .ZN(n7187) );
  OAI211_X1 U9048 ( .C1(n7190), .C2(n7189), .A(n7188), .B(n7187), .ZN(P1_U3261) );
  NAND2_X1 U9049 ( .A1(n7192), .A2(n8285), .ZN(n7193) );
  NAND2_X1 U9050 ( .A1(n7191), .A2(n7193), .ZN(n10103) );
  XNOR2_X1 U9051 ( .A(n7194), .B(n8285), .ZN(n7195) );
  NAND2_X1 U9052 ( .A1(n7195), .A2(n8769), .ZN(n7197) );
  AOI22_X1 U9053 ( .A1(n8752), .A2(n8469), .B1(n8471), .B2(n8750), .ZN(n7196)
         );
  OAI211_X1 U9054 ( .C1(n7198), .C2(n10103), .A(n7197), .B(n7196), .ZN(n10104)
         );
  NAND2_X1 U9055 ( .A1(n10104), .A2(n8780), .ZN(n7201) );
  OAI22_X1 U9056 ( .A1(n8780), .A2(n6932), .B1(n7327), .B2(n8756), .ZN(n7199)
         );
  AOI21_X1 U9057 ( .B1(n8785), .B2(n10106), .A(n7199), .ZN(n7200) );
  OAI211_X1 U9058 ( .C1(n10103), .C2(n8334), .A(n7201), .B(n7200), .ZN(
        P2_U3224) );
  AOI21_X1 U9059 ( .B1(n7203), .B2(n7210), .A(n7202), .ZN(n7331) );
  AOI21_X1 U9060 ( .B1(n7227), .B2(n7336), .A(n9617), .ZN(n7204) );
  AND2_X1 U9061 ( .A1(n7204), .A2(n9965), .ZN(n7333) );
  INV_X2 U9062 ( .A(n9984), .ZN(n9987) );
  NAND2_X1 U9063 ( .A1(n9987), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U9064 ( .A1(n9619), .A2(n7254), .ZN(n7205) );
  OAI211_X1 U9065 ( .C1(n9622), .C2(n7257), .A(n7206), .B(n7205), .ZN(n7207)
         );
  AOI21_X1 U9066 ( .B1(n7333), .B2(n9637), .A(n7207), .ZN(n7216) );
  NAND2_X1 U9067 ( .A1(n7050), .A2(n7859), .ZN(n7220) );
  NAND2_X1 U9068 ( .A1(n7220), .A2(n8002), .ZN(n7208) );
  INV_X1 U9069 ( .A(n7863), .ZN(n7848) );
  NAND2_X1 U9070 ( .A1(n7208), .A2(n7848), .ZN(n7222) );
  NAND2_X1 U9071 ( .A1(n7222), .A2(n7209), .ZN(n9953) );
  XOR2_X1 U9072 ( .A(n7210), .B(n9953), .Z(n7214) );
  NAND2_X1 U9073 ( .A1(n9281), .A2(n9465), .ZN(n7212) );
  NAND2_X1 U9074 ( .A1(n9279), .A2(n9498), .ZN(n7211) );
  NAND2_X1 U9075 ( .A1(n7212), .A2(n7211), .ZN(n7253) );
  INV_X1 U9076 ( .A(n7253), .ZN(n7213) );
  OAI21_X1 U9077 ( .B1(n7214), .B2(n9995), .A(n7213), .ZN(n7332) );
  NAND2_X1 U9078 ( .A1(n7332), .A2(n9984), .ZN(n7215) );
  OAI211_X1 U9079 ( .C1(n7331), .C2(n9606), .A(n7216), .B(n7215), .ZN(P1_U3285) );
  NOR2_X1 U9080 ( .A1(n7217), .A2(n7863), .ZN(n7218) );
  OR2_X1 U9081 ( .A1(n7219), .A2(n7218), .ZN(n10017) );
  NAND3_X1 U9082 ( .A1(n7220), .A2(n8002), .A3(n7863), .ZN(n7221) );
  NAND2_X1 U9083 ( .A1(n7222), .A2(n7221), .ZN(n7223) );
  NAND2_X1 U9084 ( .A1(n7223), .A2(n9595), .ZN(n7225) );
  AOI22_X1 U9085 ( .A1(n9465), .A2(n9282), .B1(n9280), .B2(n9498), .ZN(n7224)
         );
  NAND2_X1 U9086 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  AOI21_X1 U9087 ( .B1(n10017), .B2(n9615), .A(n7226), .ZN(n10019) );
  OAI211_X1 U9088 ( .C1(n7228), .C2(n10014), .A(n9966), .B(n7227), .ZN(n10013)
         );
  NOR2_X1 U9089 ( .A1(n10013), .A2(n9970), .ZN(n7232) );
  AOI22_X1 U9090 ( .A1(n9987), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7229), .B2(
        n9619), .ZN(n7230) );
  OAI21_X1 U9091 ( .B1(n10014), .B2(n9622), .A(n7230), .ZN(n7231) );
  AOI211_X1 U9092 ( .C1(n10017), .C2(n7735), .A(n7232), .B(n7231), .ZN(n7233)
         );
  OAI21_X1 U9093 ( .B1(n10019), .B2(n9987), .A(n7233), .ZN(P1_U3286) );
  OAI222_X1 U9094 ( .A1(P2_U3151), .A2(n8609), .B1(n8331), .B2(n7235), .C1(
        n7234), .C2(n8899), .ZN(P2_U3276) );
  XNOR2_X1 U9095 ( .A(n7244), .B(n8090), .ZN(n7317) );
  XNOR2_X1 U9096 ( .A(n7317), .B(n7318), .ZN(n7320) );
  NAND2_X1 U9097 ( .A1(n7239), .A2(n7238), .ZN(n7321) );
  XOR2_X1 U9098 ( .A(n7320), .B(n7321), .Z(n7246) );
  NAND2_X1 U9099 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n10064) );
  OAI21_X1 U9100 ( .B1(n8429), .B2(n7237), .A(n10064), .ZN(n7240) );
  AOI21_X1 U9101 ( .B1(n8420), .B2(n8470), .A(n7240), .ZN(n7241) );
  OAI21_X1 U9102 ( .B1(n7242), .B2(n8404), .A(n7241), .ZN(n7243) );
  AOI21_X1 U9103 ( .B1(n7244), .B2(n8456), .A(n7243), .ZN(n7245) );
  OAI21_X1 U9104 ( .B1(n7246), .B2(n8458), .A(n7245), .ZN(P2_U3161) );
  INV_X1 U9105 ( .A(n7247), .ZN(n8330) );
  OAI222_X1 U9106 ( .A1(n9800), .A2(n8330), .B1(n7837), .B2(P1_U3086), .C1(
        n7248), .C2(n9797), .ZN(P1_U3335) );
  XNOR2_X1 U9107 ( .A(n7251), .B(n7250), .ZN(n7252) );
  XNOR2_X1 U9108 ( .A(n7249), .B(n7252), .ZN(n7259) );
  AOI22_X1 U9109 ( .A1(n9847), .A2(n7253), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7256) );
  NAND2_X1 U9110 ( .A1(n9247), .A2(n7254), .ZN(n7255) );
  OAI211_X1 U9111 ( .C1(n7257), .C2(n9849), .A(n7256), .B(n7255), .ZN(n7258)
         );
  AOI21_X1 U9112 ( .B1(n7259), .B2(n9852), .A(n7258), .ZN(n7260) );
  INV_X1 U9113 ( .A(n7260), .ZN(P1_U3221) );
  INV_X1 U9114 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8559) );
  INV_X1 U9115 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U9116 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7303) );
  NOR2_X1 U9117 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7300) );
  NOR2_X1 U9118 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7297) );
  NOR2_X1 U9119 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7295) );
  NOR2_X1 U9120 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7292) );
  NOR2_X1 U9121 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7290) );
  NOR2_X1 U9122 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7287) );
  NOR2_X1 U9123 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7283) );
  NOR2_X1 U9124 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7280) );
  NOR2_X1 U9125 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7278) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7274) );
  NOR2_X1 U9127 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7271) );
  NOR2_X1 U9128 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7268) );
  NAND2_X1 U9129 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7266) );
  XOR2_X1 U9130 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10171) );
  NAND2_X1 U9131 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7264) );
  AOI21_X1 U9132 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10137) );
  INV_X1 U9133 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U9134 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7261) );
  NOR2_X1 U9135 ( .A1(n9291), .A2(n7261), .ZN(n10136) );
  NOR2_X1 U9136 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10136), .ZN(n7262) );
  NOR2_X1 U9137 ( .A1(n10137), .A2(n7262), .ZN(n10169) );
  XOR2_X1 U9138 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10168) );
  NAND2_X1 U9139 ( .A1(n10169), .A2(n10168), .ZN(n7263) );
  NAND2_X1 U9140 ( .A1(n7264), .A2(n7263), .ZN(n10170) );
  NAND2_X1 U9141 ( .A1(n10171), .A2(n10170), .ZN(n7265) );
  NAND2_X1 U9142 ( .A1(n7266), .A2(n7265), .ZN(n10173) );
  XNOR2_X1 U9143 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10172) );
  NOR2_X1 U9144 ( .A1(n10173), .A2(n10172), .ZN(n7267) );
  NOR2_X1 U9145 ( .A1(n7268), .A2(n7267), .ZN(n10161) );
  XOR2_X1 U9146 ( .A(n7269), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10160) );
  NOR2_X1 U9147 ( .A1(n10161), .A2(n10160), .ZN(n7270) );
  NOR2_X1 U9148 ( .A1(n7271), .A2(n7270), .ZN(n10159) );
  INV_X1 U9149 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U9150 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n9879), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(n7272), .ZN(n10158) );
  NOR2_X1 U9151 ( .A1(n10159), .A2(n10158), .ZN(n7273) );
  NOR2_X1 U9152 ( .A1(n7274), .A2(n7273), .ZN(n10165) );
  INV_X1 U9153 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7276) );
  AOI22_X1 U9154 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n7276), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n7275), .ZN(n10164) );
  NOR2_X1 U9155 ( .A1(n10165), .A2(n10164), .ZN(n7277) );
  NOR2_X1 U9156 ( .A1(n7278), .A2(n7277), .ZN(n10167) );
  XNOR2_X1 U9157 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10166) );
  NOR2_X1 U9158 ( .A1(n10167), .A2(n10166), .ZN(n7279) );
  NOR2_X1 U9159 ( .A1(n7280), .A2(n7279), .ZN(n10163) );
  INV_X1 U9160 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9841) );
  INV_X1 U9161 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7281) );
  AOI22_X1 U9162 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9841), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7281), .ZN(n10162) );
  NOR2_X1 U9163 ( .A1(n10163), .A2(n10162), .ZN(n7282) );
  NOR2_X1 U9164 ( .A1(n7283), .A2(n7282), .ZN(n10157) );
  AOI22_X1 U9165 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n7285), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7284), .ZN(n10156) );
  NOR2_X1 U9166 ( .A1(n10157), .A2(n10156), .ZN(n7286) );
  NOR2_X1 U9167 ( .A1(n7287), .A2(n7286), .ZN(n10155) );
  INV_X1 U9168 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7288) );
  INV_X1 U9169 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7504) );
  AOI22_X1 U9170 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n7288), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7504), .ZN(n10154) );
  NOR2_X1 U9171 ( .A1(n10155), .A2(n10154), .ZN(n7289) );
  NOR2_X1 U9172 ( .A1(n7290), .A2(n7289), .ZN(n10153) );
  XNOR2_X1 U9173 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10152) );
  NOR2_X1 U9174 ( .A1(n10153), .A2(n10152), .ZN(n7291) );
  NOR2_X1 U9175 ( .A1(n7292), .A2(n7291), .ZN(n10151) );
  INV_X1 U9176 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7722) );
  INV_X1 U9177 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7293) );
  AOI22_X1 U9178 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n7722), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(n7293), .ZN(n10150) );
  NOR2_X1 U9179 ( .A1(n10151), .A2(n10150), .ZN(n7294) );
  NOR2_X1 U9180 ( .A1(n7295), .A2(n7294), .ZN(n10149) );
  XNOR2_X1 U9181 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10148) );
  NOR2_X1 U9182 ( .A1(n10149), .A2(n10148), .ZN(n7296) );
  NOR2_X1 U9183 ( .A1(n7297), .A2(n7296), .ZN(n10147) );
  INV_X1 U9184 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7298) );
  INV_X1 U9185 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8521) );
  AOI22_X1 U9186 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7298), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8521), .ZN(n10146) );
  NOR2_X1 U9187 ( .A1(n10147), .A2(n10146), .ZN(n7299) );
  NOR2_X1 U9188 ( .A1(n7300), .A2(n7299), .ZN(n10145) );
  INV_X1 U9189 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7301) );
  INV_X1 U9190 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8533) );
  AOI22_X1 U9191 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7301), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8533), .ZN(n10144) );
  NOR2_X1 U9192 ( .A1(n10145), .A2(n10144), .ZN(n7302) );
  NOR2_X1 U9193 ( .A1(n7303), .A2(n7302), .ZN(n10143) );
  AOI22_X1 U9194 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9949), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8559), .ZN(n10142) );
  NOR2_X1 U9195 ( .A1(n10143), .A2(n10142), .ZN(n7304) );
  AOI21_X1 U9196 ( .B1(n8559), .B2(n9949), .A(n7304), .ZN(n7305) );
  AND2_X1 U9197 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7305), .ZN(n10140) );
  NOR2_X1 U9198 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10140), .ZN(n7306) );
  NOR2_X1 U9199 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7305), .ZN(n10139) );
  NOR2_X1 U9200 ( .A1(n7306), .A2(n10139), .ZN(n7308) );
  XNOR2_X1 U9201 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7307) );
  XNOR2_X1 U9202 ( .A(n7308), .B(n7307), .ZN(ADD_1068_U4) );
  NAND2_X1 U9203 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U9204 ( .A1(n9260), .A2(n9634), .ZN(n7309) );
  OAI211_X1 U9205 ( .C1(n7310), .C2(n9237), .A(n9878), .B(n7309), .ZN(n7315)
         );
  XOR2_X1 U9206 ( .A(n7311), .B(n7312), .Z(n7313) );
  NOR2_X1 U9207 ( .A1(n7313), .A2(n9262), .ZN(n7314) );
  AOI211_X1 U9208 ( .C1(n9630), .C2(n9247), .A(n7315), .B(n7314), .ZN(n7316)
         );
  INV_X1 U9209 ( .A(n7316), .ZN(P1_U3239) );
  INV_X1 U9210 ( .A(n7317), .ZN(n7319) );
  XNOR2_X1 U9211 ( .A(n10106), .B(n8090), .ZN(n7417) );
  XNOR2_X1 U9212 ( .A(n7417), .B(n7418), .ZN(n7322) );
  NAND2_X1 U9213 ( .A1(n7323), .A2(n7322), .ZN(n7422) );
  OAI211_X1 U9214 ( .C1(n7323), .C2(n7322), .A(n7422), .B(n8439), .ZN(n7330)
         );
  AOI21_X1 U9215 ( .B1(n8449), .B2(n8471), .A(n7324), .ZN(n7326) );
  NAND2_X1 U9216 ( .A1(n8420), .A2(n8469), .ZN(n7325) );
  OAI211_X1 U9217 ( .C1(n8404), .C2(n7327), .A(n7326), .B(n7325), .ZN(n7328)
         );
  AOI21_X1 U9218 ( .B1(n10106), .B2(n8456), .A(n7328), .ZN(n7329) );
  NAND2_X1 U9219 ( .A1(n7330), .A2(n7329), .ZN(P2_U3171) );
  INV_X1 U9220 ( .A(n7331), .ZN(n7334) );
  AOI211_X1 U9221 ( .C1(n7334), .C2(n10026), .A(n7333), .B(n7332), .ZN(n7338)
         );
  AOI22_X1 U9222 ( .A1(n9719), .A2(n7336), .B1(n10039), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U9223 ( .B1(n7338), .B2(n10039), .A(n7335), .ZN(P1_U3530) );
  AOI22_X1 U9224 ( .A1(n9785), .A2(n7336), .B1(n10028), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n7337) );
  OAI21_X1 U9225 ( .B1(n7338), .B2(n10028), .A(n7337), .ZN(P1_U3477) );
  INV_X1 U9226 ( .A(n8151), .ZN(n7339) );
  OR2_X1 U9227 ( .A1(n8156), .A2(n7339), .ZN(n8290) );
  XOR2_X1 U9228 ( .A(n7340), .B(n8290), .Z(n10110) );
  XNOR2_X1 U9229 ( .A(n7341), .B(n8290), .ZN(n7342) );
  OAI222_X1 U9230 ( .A1(n8775), .A2(n7537), .B1(n8773), .B2(n7418), .C1(n7342), 
        .C2(n8738), .ZN(n10112) );
  NAND2_X1 U9231 ( .A1(n10112), .A2(n8780), .ZN(n7345) );
  OAI22_X1 U9232 ( .A1(n8780), .A2(n7489), .B1(n7426), .B2(n8756), .ZN(n7343)
         );
  AOI21_X1 U9233 ( .B1(n8785), .B2(n7532), .A(n7343), .ZN(n7344) );
  OAI211_X1 U9234 ( .C1(n8788), .C2(n10110), .A(n7345), .B(n7344), .ZN(
        P2_U3223) );
  INV_X1 U9235 ( .A(n7346), .ZN(n7349) );
  OAI222_X1 U9236 ( .A1(n9800), .A2(n7349), .B1(n7803), .B2(P1_U3086), .C1(
        n7347), .C2(n9797), .ZN(P1_U3334) );
  OAI222_X1 U9237 ( .A1(n8277), .A2(P2_U3151), .B1(n8331), .B2(n7349), .C1(
        n7348), .C2(n8899), .ZN(P2_U3274) );
  OAI21_X1 U9238 ( .B1(n7351), .B2(n7811), .A(n7350), .ZN(n7378) );
  INV_X1 U9239 ( .A(n7378), .ZN(n7365) );
  INV_X1 U9240 ( .A(n7352), .ZN(n9967) );
  AOI211_X1 U9241 ( .C1(n7379), .C2(n9967), .A(n9617), .B(n7353), .ZN(n7377)
         );
  NOR2_X1 U9242 ( .A1(n9850), .A2(n9622), .ZN(n7356) );
  OAI22_X1 U9243 ( .A1(n9984), .A2(n7354), .B1(n9855), .B2(n9978), .ZN(n7355)
         );
  AOI211_X1 U9244 ( .C1(n7377), .C2(n9637), .A(n7356), .B(n7355), .ZN(n7364)
         );
  INV_X1 U9245 ( .A(n7403), .ZN(n7357) );
  AOI21_X1 U9246 ( .B1(n7811), .B2(n7358), .A(n7357), .ZN(n7362) );
  NAND2_X1 U9247 ( .A1(n9279), .A2(n9465), .ZN(n7360) );
  NAND2_X1 U9248 ( .A1(n9278), .A2(n9498), .ZN(n7359) );
  NAND2_X1 U9249 ( .A1(n7360), .A2(n7359), .ZN(n9846) );
  INV_X1 U9250 ( .A(n9846), .ZN(n7361) );
  OAI21_X1 U9251 ( .B1(n7362), .B2(n9995), .A(n7361), .ZN(n7376) );
  NAND2_X1 U9252 ( .A1(n7376), .A2(n9984), .ZN(n7363) );
  OAI211_X1 U9253 ( .C1(n7365), .C2(n9606), .A(n7364), .B(n7363), .ZN(P1_U3283) );
  NAND2_X1 U9254 ( .A1(n7366), .A2(n8151), .ZN(n7367) );
  XNOR2_X1 U9255 ( .A(n7367), .B(n8291), .ZN(n10114) );
  INV_X1 U9256 ( .A(n7368), .ZN(n7370) );
  OAI211_X1 U9257 ( .C1(n7370), .C2(n8291), .A(n8769), .B(n7369), .ZN(n7372)
         );
  AOI22_X1 U9258 ( .A1(n8750), .A2(n8469), .B1(n8467), .B2(n8752), .ZN(n7371)
         );
  NAND2_X1 U9259 ( .A1(n7372), .A2(n7371), .ZN(n10115) );
  NAND2_X1 U9260 ( .A1(n10115), .A2(n8780), .ZN(n7375) );
  OAI22_X1 U9261 ( .A1(n8780), .A2(n7506), .B1(n7476), .B2(n8756), .ZN(n7373)
         );
  AOI21_X1 U9262 ( .B1(n8785), .B2(n10117), .A(n7373), .ZN(n7374) );
  OAI211_X1 U9263 ( .C1(n8788), .C2(n10114), .A(n7375), .B(n7374), .ZN(
        P2_U3222) );
  AOI211_X1 U9264 ( .C1(n7378), .C2(n10026), .A(n7377), .B(n7376), .ZN(n7384)
         );
  AOI22_X1 U9265 ( .A1(n9719), .A2(n7379), .B1(n10039), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7380) );
  OAI21_X1 U9266 ( .B1(n7384), .B2(n10039), .A(n7380), .ZN(P1_U3532) );
  INV_X1 U9267 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7381) );
  OAI22_X1 U9268 ( .A1(n9781), .A2(n9850), .B1(n10030), .B2(n7381), .ZN(n7382)
         );
  INV_X1 U9269 ( .A(n7382), .ZN(n7383) );
  OAI21_X1 U9270 ( .B1(n7384), .B2(n10028), .A(n7383), .ZN(P1_U3483) );
  INV_X1 U9271 ( .A(n7386), .ZN(n7387) );
  AOI21_X1 U9272 ( .B1(n7388), .B2(n7385), .A(n7387), .ZN(n7394) );
  NAND2_X1 U9273 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9839) );
  OAI21_X1 U9274 ( .B1(n9210), .B2(n7389), .A(n9839), .ZN(n7392) );
  INV_X1 U9275 ( .A(n7390), .ZN(n9960) );
  OAI22_X1 U9276 ( .A1(n9957), .A2(n9209), .B1(n9856), .B2(n9960), .ZN(n7391)
         );
  AOI211_X1 U9277 ( .C1(n9959), .C2(n9260), .A(n7392), .B(n7391), .ZN(n7393)
         );
  OAI21_X1 U9278 ( .B1(n7394), .B2(n9262), .A(n7393), .ZN(P1_U3231) );
  OAI21_X1 U9279 ( .B1(n7396), .B2(n7817), .A(n7395), .ZN(n7482) );
  INV_X1 U9280 ( .A(n7482), .ZN(n7413) );
  INV_X1 U9281 ( .A(n7353), .ZN(n7398) );
  INV_X1 U9282 ( .A(n7449), .ZN(n7397) );
  AOI211_X1 U9283 ( .C1(n9224), .C2(n7398), .A(n9617), .B(n7397), .ZN(n7481)
         );
  NOR2_X1 U9284 ( .A1(n7488), .A2(n9622), .ZN(n7402) );
  INV_X1 U9285 ( .A(n9225), .ZN(n7399) );
  OAI22_X1 U9286 ( .A1(n9984), .A2(n7400), .B1(n7399), .B2(n9978), .ZN(n7401)
         );
  AOI211_X1 U9287 ( .C1(n7481), .C2(n9637), .A(n7402), .B(n7401), .ZN(n7412)
         );
  NAND2_X1 U9288 ( .A1(n7403), .A2(n7884), .ZN(n7404) );
  NAND2_X1 U9289 ( .A1(n7404), .A2(n7817), .ZN(n7406) );
  NAND3_X1 U9290 ( .A1(n7406), .A2(n7405), .A3(n9595), .ZN(n7410) );
  NAND2_X1 U9291 ( .A1(n9277), .A2(n9498), .ZN(n7408) );
  NAND2_X1 U9292 ( .A1(n9969), .A2(n9465), .ZN(n7407) );
  NAND2_X1 U9293 ( .A1(n7408), .A2(n7407), .ZN(n9223) );
  INV_X1 U9294 ( .A(n9223), .ZN(n7409) );
  NAND2_X1 U9295 ( .A1(n7410), .A2(n7409), .ZN(n7480) );
  NAND2_X1 U9296 ( .A1(n7480), .A2(n9984), .ZN(n7411) );
  OAI211_X1 U9297 ( .C1(n7413), .C2(n9606), .A(n7412), .B(n7411), .ZN(P1_U3282) );
  INV_X1 U9298 ( .A(n7414), .ZN(n7744) );
  OAI222_X1 U9299 ( .A1(P2_U3151), .A2(n7416), .B1(n8331), .B2(n7744), .C1(
        n7415), .C2(n8899), .ZN(P2_U3273) );
  INV_X1 U9300 ( .A(n7417), .ZN(n7419) );
  INV_X1 U9301 ( .A(n7420), .ZN(n7421) );
  XNOR2_X1 U9302 ( .A(n7542), .B(n8469), .ZN(n7472) );
  XNOR2_X1 U9303 ( .A(n10109), .B(n6650), .ZN(n7531) );
  XNOR2_X1 U9304 ( .A(n7472), .B(n7531), .ZN(n7429) );
  AOI21_X1 U9305 ( .B1(n8449), .B2(n8470), .A(n7423), .ZN(n7425) );
  NAND2_X1 U9306 ( .A1(n8420), .A2(n8468), .ZN(n7424) );
  OAI211_X1 U9307 ( .C1(n8404), .C2(n7426), .A(n7425), .B(n7424), .ZN(n7427)
         );
  AOI21_X1 U9308 ( .B1(n7532), .B2(n8456), .A(n7427), .ZN(n7428) );
  OAI21_X1 U9309 ( .B1(n7429), .B2(n8458), .A(n7428), .ZN(P2_U3157) );
  OR2_X1 U9310 ( .A1(n7430), .A2(n8293), .ZN(n7431) );
  NAND2_X1 U9311 ( .A1(n7432), .A2(n7431), .ZN(n7553) );
  XOR2_X1 U9312 ( .A(n7433), .B(n8293), .Z(n7434) );
  OAI222_X1 U9313 ( .A1(n8775), .A2(n7583), .B1(n8773), .B2(n7537), .C1(n8738), 
        .C2(n7434), .ZN(n7548) );
  NAND2_X1 U9314 ( .A1(n7548), .A2(n8780), .ZN(n7438) );
  NAND2_X1 U9315 ( .A1(n8767), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7435) );
  OAI21_X1 U9316 ( .B1(n7528), .B2(n8756), .A(n7435), .ZN(n7436) );
  AOI21_X1 U9317 ( .B1(n8169), .B2(n8785), .A(n7436), .ZN(n7437) );
  OAI211_X1 U9318 ( .C1(n7553), .C2(n8788), .A(n7438), .B(n7437), .ZN(P2_U3221) );
  OAI21_X1 U9319 ( .B1(n7441), .B2(n7440), .A(n7439), .ZN(n7558) );
  INV_X1 U9320 ( .A(n7558), .ZN(n7454) );
  OAI211_X1 U9321 ( .C1(n7820), .C2(n7443), .A(n7442), .B(n9595), .ZN(n7447)
         );
  NAND2_X1 U9322 ( .A1(n9276), .A2(n9968), .ZN(n7445) );
  NAND2_X1 U9323 ( .A1(n9278), .A2(n9465), .ZN(n7444) );
  NAND2_X1 U9324 ( .A1(n7445), .A2(n7444), .ZN(n9126) );
  INV_X1 U9325 ( .A(n9126), .ZN(n7446) );
  NAND2_X1 U9326 ( .A1(n7447), .A2(n7446), .ZN(n7556) );
  INV_X1 U9327 ( .A(n9130), .ZN(n7564) );
  INV_X1 U9328 ( .A(n7567), .ZN(n7448) );
  AOI211_X1 U9329 ( .C1(n9130), .C2(n7449), .A(n9617), .B(n7448), .ZN(n7557)
         );
  NAND2_X1 U9330 ( .A1(n7557), .A2(n9637), .ZN(n7451) );
  AOI22_X1 U9331 ( .A1(n9987), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9125), .B2(
        n9619), .ZN(n7450) );
  OAI211_X1 U9332 ( .C1(n7564), .C2(n9622), .A(n7451), .B(n7450), .ZN(n7452)
         );
  AOI21_X1 U9333 ( .B1(n9984), .B2(n7556), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9334 ( .B1(n7454), .B2(n9606), .A(n7453), .ZN(P1_U3281) );
  XOR2_X1 U9335 ( .A(n7455), .B(n8292), .Z(n7523) );
  OAI21_X1 U9336 ( .B1(n8292), .B2(n7457), .A(n7456), .ZN(n7458) );
  NAND2_X1 U9337 ( .A1(n7458), .A2(n8769), .ZN(n7460) );
  AOI22_X1 U9338 ( .A1(n8752), .A2(n8465), .B1(n8467), .B2(n8750), .ZN(n7459)
         );
  NAND2_X1 U9339 ( .A1(n7460), .A2(n7459), .ZN(n7522) );
  INV_X1 U9340 ( .A(n8174), .ZN(n7593) );
  OAI22_X1 U9341 ( .A1(n7593), .A2(n8682), .B1(n7588), .B2(n8756), .ZN(n7461)
         );
  OAI21_X1 U9342 ( .B1(n7522), .B2(n7461), .A(n8780), .ZN(n7463) );
  NAND2_X1 U9343 ( .A1(n8767), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7462) );
  OAI211_X1 U9344 ( .C1(n7523), .C2(n8788), .A(n7463), .B(n7462), .ZN(P2_U3220) );
  NAND2_X1 U9345 ( .A1(n7468), .A2(n7464), .ZN(n7465) );
  OAI211_X1 U9346 ( .C1(n7466), .C2(n8899), .A(n7465), .B(n8324), .ZN(P2_U3272) );
  NAND2_X1 U9347 ( .A1(n7468), .A2(n7467), .ZN(n7469) );
  OAI211_X1 U9348 ( .C1(n7470), .C2(n8329), .A(n7469), .B(n8052), .ZN(P1_U3332) );
  INV_X1 U9349 ( .A(n7531), .ZN(n7471) );
  OAI22_X1 U9350 ( .A1(n7472), .A2(n7471), .B1(n8469), .B2(n7542), .ZN(n7473)
         );
  XNOR2_X1 U9351 ( .A(n7536), .B(n8090), .ZN(n7529) );
  XNOR2_X1 U9352 ( .A(n7473), .B(n7529), .ZN(n7479) );
  AND2_X1 U9353 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7515) );
  AOI21_X1 U9354 ( .B1(n8449), .B2(n8469), .A(n7515), .ZN(n7475) );
  NAND2_X1 U9355 ( .A1(n8420), .A2(n8467), .ZN(n7474) );
  OAI211_X1 U9356 ( .C1(n8404), .C2(n7476), .A(n7475), .B(n7474), .ZN(n7477)
         );
  AOI21_X1 U9357 ( .B1(n10117), .B2(n8456), .A(n7477), .ZN(n7478) );
  OAI21_X1 U9358 ( .B1(n7479), .B2(n8458), .A(n7478), .ZN(P2_U3176) );
  INV_X1 U9359 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7483) );
  AOI211_X1 U9360 ( .C1(n7482), .C2(n10026), .A(n7481), .B(n7480), .ZN(n7485)
         );
  MUX2_X1 U9361 ( .A(n7483), .B(n7485), .S(n10030), .Z(n7484) );
  OAI21_X1 U9362 ( .B1(n7488), .B2(n9781), .A(n7484), .ZN(P1_U3486) );
  MUX2_X1 U9363 ( .A(n7486), .B(n7485), .S(n10042), .Z(n7487) );
  OAI21_X1 U9364 ( .B1(n7488), .B2(n9715), .A(n7487), .ZN(P1_U3533) );
  OR2_X1 U9365 ( .A1(n7496), .A2(n7489), .ZN(n7491) );
  NAND2_X1 U9366 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  AOI21_X1 U9367 ( .B1(n7494), .B2(n7506), .A(n7631), .ZN(n7503) );
  OR2_X1 U9368 ( .A1(n7496), .A2(n7495), .ZN(n7499) );
  INV_X1 U9369 ( .A(n7497), .ZN(n7498) );
  NAND2_X1 U9370 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  AOI21_X1 U9371 ( .B1(n7501), .B2(n7505), .A(n4372), .ZN(n7502) );
  OAI22_X1 U9372 ( .A1(n7503), .A2(n8620), .B1(n8624), .B2(n7502), .ZN(n7517)
         );
  NOR2_X1 U9373 ( .A1(n8594), .A2(n7504), .ZN(n7516) );
  MUX2_X1 U9374 ( .A(n7506), .B(n7505), .S(n8318), .Z(n7507) );
  OAI21_X1 U9375 ( .B1(n7508), .B2(n7507), .A(n4374), .ZN(n7512) );
  AOI21_X1 U9376 ( .B1(n7512), .B2(n7511), .A(n7640), .ZN(n7513) );
  NOR2_X1 U9377 ( .A1(n7513), .A2(n10055), .ZN(n7514) );
  NOR4_X1 U9378 ( .A1(n7517), .A2(n7516), .A3(n7515), .A4(n7514), .ZN(n7518)
         );
  OAI21_X1 U9379 ( .B1(n7519), .B2(n8587), .A(n7518), .ZN(P2_U3193) );
  MUX2_X1 U9380 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7522), .S(n10135), .Z(n7521) );
  OAI22_X1 U9381 ( .A1(n7523), .A2(n8828), .B1(n7593), .B2(n8813), .ZN(n7520)
         );
  OR2_X1 U9382 ( .A1(n7521), .A2(n7520), .ZN(P2_U3472) );
  MUX2_X1 U9383 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n7522), .S(n10119), .Z(n7525) );
  OAI22_X1 U9384 ( .A1(n7523), .A2(n8894), .B1(n7593), .B2(n8878), .ZN(n7524)
         );
  OR2_X1 U9385 ( .A1(n7525), .A2(n7524), .ZN(P2_U3429) );
  NAND2_X1 U9386 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .ZN(n7643) );
  OAI21_X1 U9387 ( .B1(n8453), .B2(n7583), .A(n7643), .ZN(n7526) );
  AOI21_X1 U9388 ( .B1(n8449), .B2(n8468), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9389 ( .B1(n7528), .B2(n8404), .A(n7527), .ZN(n7546) );
  AOI21_X1 U9390 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7541) );
  NAND3_X1 U9391 ( .A1(n7532), .A2(n8469), .A3(n6650), .ZN(n7533) );
  OAI211_X1 U9392 ( .C1(n7537), .C2(n6650), .A(n8291), .B(n7533), .ZN(n7539)
         );
  INV_X1 U9393 ( .A(n8090), .ZN(n8074) );
  NAND3_X1 U9394 ( .A1(n10109), .A2(n7534), .A3(n8469), .ZN(n7535) );
  OAI211_X1 U9395 ( .C1(n7537), .C2(n8074), .A(n7536), .B(n7535), .ZN(n7538)
         );
  XNOR2_X1 U9396 ( .A(n8169), .B(n8090), .ZN(n7584) );
  XNOR2_X1 U9397 ( .A(n7584), .B(n8467), .ZN(n7543) );
  AOI211_X1 U9398 ( .C1(n7544), .C2(n7543), .A(n8458), .B(n4368), .ZN(n7545)
         );
  AOI211_X1 U9399 ( .C1(n8169), .C2(n8456), .A(n7546), .B(n7545), .ZN(n7547)
         );
  INV_X1 U9400 ( .A(n7547), .ZN(P2_U3164) );
  INV_X1 U9401 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7549) );
  AOI21_X1 U9402 ( .B1(n10118), .B2(n8169), .A(n7548), .ZN(n7551) );
  MUX2_X1 U9403 ( .A(n7549), .B(n7551), .S(n10119), .Z(n7550) );
  OAI21_X1 U9404 ( .B1(n7553), .B2(n8894), .A(n7550), .ZN(P2_U3426) );
  MUX2_X1 U9405 ( .A(n7636), .B(n7551), .S(n10135), .Z(n7552) );
  OAI21_X1 U9406 ( .B1(n8828), .B2(n7553), .A(n7552), .ZN(P2_U3471) );
  INV_X1 U9407 ( .A(n5879), .ZN(n7774) );
  OAI222_X1 U9408 ( .A1(n9800), .A2(n7774), .B1(P1_U3086), .B2(n7555), .C1(
        n7554), .C2(n9797), .ZN(P1_U3331) );
  AOI211_X1 U9409 ( .C1(n7558), .C2(n10026), .A(n7557), .B(n7556), .ZN(n7561)
         );
  MUX2_X1 U9410 ( .A(n7559), .B(n7561), .S(n10042), .Z(n7560) );
  OAI21_X1 U9411 ( .B1(n7564), .B2(n9715), .A(n7560), .ZN(P1_U3534) );
  INV_X1 U9412 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7562) );
  MUX2_X1 U9413 ( .A(n7562), .B(n7561), .S(n10030), .Z(n7563) );
  OAI21_X1 U9414 ( .B1(n7564), .B2(n9781), .A(n7563), .ZN(P1_U3489) );
  OAI21_X1 U9415 ( .B1(n7566), .B2(n7883), .A(n7565), .ZN(n7600) );
  INV_X1 U9416 ( .A(n7600), .ZN(n7582) );
  NAND2_X1 U9417 ( .A1(n7567), .A2(n9202), .ZN(n7568) );
  NAND2_X1 U9418 ( .A1(n7568), .A2(n9966), .ZN(n7569) );
  NOR2_X1 U9419 ( .A1(n9616), .A2(n7569), .ZN(n7594) );
  INV_X1 U9420 ( .A(n9202), .ZN(n7570) );
  NOR2_X1 U9421 ( .A1(n7570), .A2(n9622), .ZN(n7574) );
  INV_X1 U9422 ( .A(n7571), .ZN(n9200) );
  OAI22_X1 U9423 ( .A1(n9984), .A2(n7572), .B1(n9200), .B2(n9978), .ZN(n7573)
         );
  AOI211_X1 U9424 ( .C1(n7594), .C2(n9637), .A(n7574), .B(n7573), .ZN(n7581)
         );
  NAND2_X1 U9425 ( .A1(n7442), .A2(n7890), .ZN(n7575) );
  XOR2_X1 U9426 ( .A(n7883), .B(n7575), .Z(n7579) );
  NAND2_X1 U9427 ( .A1(n9277), .A2(n9465), .ZN(n7577) );
  NAND2_X1 U9428 ( .A1(n9275), .A2(n9498), .ZN(n7576) );
  NAND2_X1 U9429 ( .A1(n7577), .A2(n7576), .ZN(n9198) );
  INV_X1 U9430 ( .A(n9198), .ZN(n7578) );
  OAI21_X1 U9431 ( .B1(n7579), .B2(n9995), .A(n7578), .ZN(n7595) );
  NAND2_X1 U9432 ( .A1(n7595), .A2(n9984), .ZN(n7580) );
  OAI211_X1 U9433 ( .C1(n7582), .C2(n9606), .A(n7581), .B(n7580), .ZN(P1_U3280) );
  XNOR2_X1 U9434 ( .A(n8174), .B(n8090), .ZN(n7672) );
  XNOR2_X1 U9435 ( .A(n7672), .B(n7583), .ZN(n7586) );
  NAND2_X1 U9436 ( .A1(n7585), .A2(n7586), .ZN(n7671) );
  OAI21_X1 U9437 ( .B1(n7586), .B2(n7585), .A(n7671), .ZN(n7587) );
  NAND2_X1 U9438 ( .A1(n7587), .A2(n8439), .ZN(n7592) );
  NAND2_X1 U9439 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7720) );
  OAI21_X1 U9440 ( .B1(n8429), .B2(n8168), .A(n7720), .ZN(n7590) );
  NOR2_X1 U9441 ( .A1(n8404), .A2(n7588), .ZN(n7589) );
  AOI211_X1 U9442 ( .C1(n8420), .C2(n8465), .A(n7590), .B(n7589), .ZN(n7591)
         );
  OAI211_X1 U9443 ( .C1(n7593), .C2(n8446), .A(n7592), .B(n7591), .ZN(P2_U3174) );
  NOR2_X1 U9444 ( .A1(n7595), .A2(n7594), .ZN(n7603) );
  NAND2_X1 U9445 ( .A1(n7600), .A2(n7596), .ZN(n7598) );
  AOI22_X1 U9446 ( .A1(n9202), .A2(n9785), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10028), .ZN(n7597) );
  OAI211_X1 U9447 ( .C1(n7603), .C2(n10028), .A(n7598), .B(n7597), .ZN(
        P1_U3492) );
  NAND2_X1 U9448 ( .A1(n7600), .A2(n7599), .ZN(n7602) );
  AOI22_X1 U9449 ( .A1(n9202), .A2(n9719), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10039), .ZN(n7601) );
  OAI211_X1 U9450 ( .C1(n7603), .C2(n10039), .A(n7602), .B(n7601), .ZN(
        P1_U3535) );
  AOI21_X1 U9451 ( .B1(n7604), .B2(n8275), .A(n8738), .ZN(n7607) );
  OAI22_X1 U9452 ( .A1(n8391), .A2(n8775), .B1(n8392), .B2(n8773), .ZN(n7605)
         );
  AOI21_X1 U9453 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n8832) );
  OAI22_X1 U9454 ( .A1(n8780), .A2(n8546), .B1(n8393), .B2(n8756), .ZN(n7608)
         );
  AOI21_X1 U9455 ( .B1(n8829), .B2(n8785), .A(n7608), .ZN(n7612) );
  OAI21_X1 U9456 ( .B1(n7610), .B2(n8275), .A(n7609), .ZN(n8830) );
  NAND2_X1 U9457 ( .A1(n8830), .A2(n8764), .ZN(n7611) );
  OAI211_X1 U9458 ( .C1(n8832), .C2(n8767), .A(n7612), .B(n7611), .ZN(P2_U3217) );
  INV_X1 U9459 ( .A(n7613), .ZN(n8184) );
  OR2_X1 U9460 ( .A1(n8183), .A2(n8184), .ZN(n8180) );
  XNOR2_X1 U9461 ( .A(n7614), .B(n4539), .ZN(n7628) );
  XNOR2_X1 U9462 ( .A(n7615), .B(n8180), .ZN(n7616) );
  AOI222_X1 U9463 ( .A1(n8769), .A2(n7616), .B1(n8464), .B2(n8752), .C1(n8466), 
        .C2(n8750), .ZN(n7622) );
  MUX2_X1 U9464 ( .A(n8483), .B(n7622), .S(n10135), .Z(n7618) );
  INV_X1 U9465 ( .A(n8813), .ZN(n8825) );
  NAND2_X1 U9466 ( .A1(n7677), .A2(n8825), .ZN(n7617) );
  OAI211_X1 U9467 ( .C1(n7628), .C2(n8828), .A(n7618), .B(n7617), .ZN(P2_U3473) );
  INV_X1 U9468 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7619) );
  MUX2_X1 U9469 ( .A(n7619), .B(n7622), .S(n10119), .Z(n7621) );
  NAND2_X1 U9470 ( .A1(n7677), .A2(n8890), .ZN(n7620) );
  OAI211_X1 U9471 ( .C1(n7628), .C2(n8894), .A(n7621), .B(n7620), .ZN(P2_U3432) );
  INV_X1 U9472 ( .A(n7622), .ZN(n7625) );
  INV_X1 U9473 ( .A(n7677), .ZN(n7623) );
  OAI22_X1 U9474 ( .A1(n7623), .A2(n8682), .B1(n7675), .B2(n8756), .ZN(n7624)
         );
  OAI21_X1 U9475 ( .B1(n7625), .B2(n7624), .A(n8780), .ZN(n7627) );
  NAND2_X1 U9476 ( .A1(n8767), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7626) );
  OAI211_X1 U9477 ( .C1(n7628), .C2(n8788), .A(n7627), .B(n7626), .ZN(P2_U3219) );
  INV_X1 U9478 ( .A(n7629), .ZN(n7656) );
  OAI222_X1 U9479 ( .A1(n9800), .A2(n7656), .B1(P1_U3086), .B2(n7630), .C1(
        n9060), .C2(n9797), .ZN(P1_U3330) );
  NAND2_X1 U9480 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7706), .ZN(n7633) );
  OAI21_X1 U9481 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7706), .A(n7633), .ZN(
        n7634) );
  AOI21_X1 U9482 ( .B1(n7635), .B2(n7634), .A(n7702), .ZN(n7654) );
  MUX2_X1 U9483 ( .A(n7637), .B(n7636), .S(n8318), .Z(n7639) );
  AND2_X1 U9484 ( .A1(n7639), .A2(n7652), .ZN(n7717) );
  INV_X1 U9485 ( .A(n7717), .ZN(n7638) );
  OAI21_X1 U9486 ( .B1(n7652), .B2(n7639), .A(n7638), .ZN(n7642) );
  AOI21_X1 U9487 ( .B1(n7642), .B2(n7641), .A(n7716), .ZN(n7645) );
  NAND2_X1 U9488 ( .A1(n10049), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7644) );
  OAI211_X1 U9489 ( .C1(n7645), .C2(n10055), .A(n7644), .B(n7643), .ZN(n7651)
         );
  NAND2_X1 U9490 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7706), .ZN(n7646) );
  OAI21_X1 U9491 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7706), .A(n7646), .ZN(
        n7647) );
  NOR2_X1 U9492 ( .A1(n7648), .A2(n7647), .ZN(n7708) );
  AOI21_X1 U9493 ( .B1(n7648), .B2(n7647), .A(n7708), .ZN(n7649) );
  NOR2_X1 U9494 ( .A1(n7649), .A2(n8624), .ZN(n7650) );
  AOI211_X1 U9495 ( .C1(n10047), .C2(n7652), .A(n7651), .B(n7650), .ZN(n7653)
         );
  OAI21_X1 U9496 ( .B1(n7654), .B2(n8620), .A(n7653), .ZN(P2_U3194) );
  OAI222_X1 U9497 ( .A1(n7657), .A2(P2_U3151), .B1(n8331), .B2(n7656), .C1(
        n7655), .C2(n8899), .ZN(P2_U3270) );
  XNOR2_X1 U9498 ( .A(n7658), .B(n8186), .ZN(n7670) );
  XNOR2_X1 U9499 ( .A(n7659), .B(n8186), .ZN(n7660) );
  AOI222_X1 U9500 ( .A1(n8769), .A2(n7660), .B1(n8465), .B2(n8750), .C1(n8463), 
        .C2(n8752), .ZN(n7667) );
  MUX2_X1 U9501 ( .A(n8513), .B(n7667), .S(n8780), .Z(n7663) );
  INV_X1 U9502 ( .A(n7661), .ZN(n7696) );
  AOI22_X1 U9503 ( .A1(n7690), .A2(n8785), .B1(n8784), .B2(n7696), .ZN(n7662)
         );
  OAI211_X1 U9504 ( .C1(n7670), .C2(n8788), .A(n7663), .B(n7662), .ZN(P2_U3218) );
  INV_X1 U9505 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7664) );
  MUX2_X1 U9506 ( .A(n7664), .B(n7667), .S(n10119), .Z(n7666) );
  NAND2_X1 U9507 ( .A1(n7690), .A2(n8890), .ZN(n7665) );
  OAI211_X1 U9508 ( .C1(n7670), .C2(n8894), .A(n7666), .B(n7665), .ZN(P2_U3435) );
  MUX2_X1 U9509 ( .A(n8512), .B(n7667), .S(n10135), .Z(n7669) );
  NAND2_X1 U9510 ( .A1(n7690), .A2(n8825), .ZN(n7668) );
  OAI211_X1 U9511 ( .C1(n8828), .C2(n7670), .A(n7669), .B(n7668), .ZN(P2_U3474) );
  XNOR2_X1 U9512 ( .A(n7677), .B(n8090), .ZN(n7686) );
  XNOR2_X1 U9513 ( .A(n7686), .B(n7694), .ZN(n7688) );
  OAI21_X2 U9514 ( .B1(n7672), .B2(n8466), .A(n7671), .ZN(n7689) );
  XOR2_X1 U9515 ( .A(n7688), .B(n7689), .Z(n7679) );
  AOI22_X1 U9516 ( .A1(n8420), .A2(n8464), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7674) );
  NAND2_X1 U9517 ( .A1(n8449), .A2(n8466), .ZN(n7673) );
  OAI211_X1 U9518 ( .C1(n8404), .C2(n7675), .A(n7674), .B(n7673), .ZN(n7676)
         );
  AOI21_X1 U9519 ( .B1(n7677), .B2(n8456), .A(n7676), .ZN(n7678) );
  OAI21_X1 U9520 ( .B1(n7679), .B2(n8458), .A(n7678), .ZN(P2_U3155) );
  INV_X1 U9521 ( .A(n7680), .ZN(n7684) );
  OAI222_X1 U9522 ( .A1(n9800), .A2(n7684), .B1(P1_U3086), .B2(n7682), .C1(
        n7681), .C2(n9797), .ZN(P1_U3329) );
  OAI222_X1 U9523 ( .A1(n7685), .A2(P2_U3151), .B1(n8907), .B2(n7684), .C1(
        n7683), .C2(n8899), .ZN(P2_U3269) );
  INV_X1 U9524 ( .A(n7690), .ZN(n7699) );
  INV_X1 U9525 ( .A(n7686), .ZN(n7687) );
  XNOR2_X1 U9526 ( .A(n7690), .B(n6650), .ZN(n8054) );
  XNOR2_X1 U9527 ( .A(n8054), .B(n8392), .ZN(n7691) );
  OAI211_X1 U9528 ( .C1(n7692), .C2(n7691), .A(n8056), .B(n8439), .ZN(n7698)
         );
  NAND2_X1 U9529 ( .A1(n8420), .A2(n8463), .ZN(n7693) );
  NAND2_X1 U9530 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8519) );
  OAI211_X1 U9531 ( .C1(n7694), .C2(n8429), .A(n7693), .B(n8519), .ZN(n7695)
         );
  AOI21_X1 U9532 ( .B1(n8450), .B2(n7696), .A(n7695), .ZN(n7697) );
  OAI211_X1 U9533 ( .C1(n7699), .C2(n8446), .A(n7698), .B(n7697), .ZN(P2_U3181) );
  INV_X1 U9534 ( .A(n7700), .ZN(n7733) );
  OAI222_X1 U9535 ( .A1(P2_U3151), .A2(n8318), .B1(n8907), .B2(n7733), .C1(
        n7701), .C2(n8899), .ZN(P2_U3268) );
  AOI21_X1 U9536 ( .B1(n7705), .B2(n7713), .A(n8479), .ZN(n7728) );
  AND2_X1 U9537 ( .A1(n7706), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9538 ( .A1(n7710), .A2(n7709), .ZN(n8492) );
  NOR2_X1 U9539 ( .A1(n4358), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7711) );
  OAI21_X1 U9540 ( .B1(n7711), .B2(n8493), .A(n10050), .ZN(n7727) );
  MUX2_X1 U9541 ( .A(n7713), .B(n7712), .S(n8318), .Z(n7715) );
  AND2_X1 U9542 ( .A1(n7715), .A2(n7725), .ZN(n8486) );
  INV_X1 U9543 ( .A(n8486), .ZN(n7714) );
  OAI21_X1 U9544 ( .B1(n7725), .B2(n7715), .A(n7714), .ZN(n7719) );
  NOR2_X1 U9545 ( .A1(n7717), .A2(n7716), .ZN(n7718) );
  AOI21_X1 U9546 ( .B1(n7719), .B2(n7718), .A(n8485), .ZN(n7721) );
  OAI21_X1 U9547 ( .B1(n7721), .B2(n10055), .A(n7720), .ZN(n7724) );
  NOR2_X1 U9548 ( .A1(n8594), .A2(n7722), .ZN(n7723) );
  AOI211_X1 U9549 ( .C1(n10047), .C2(n7725), .A(n7724), .B(n7723), .ZN(n7726)
         );
  OAI211_X1 U9550 ( .C1(n7728), .C2(n8620), .A(n7727), .B(n7726), .ZN(P2_U3195) );
  INV_X1 U9551 ( .A(n7729), .ZN(n7747) );
  OAI222_X1 U9552 ( .A1(n9800), .A2(n7747), .B1(n7731), .B2(P1_U3086), .C1(
        n7730), .C2(n9797), .ZN(P1_U3327) );
  OAI222_X1 U9553 ( .A1(n9800), .A2(n7733), .B1(P1_U3086), .B2(n4296), .C1(
        n7732), .C2(n9797), .ZN(P1_U3328) );
  MUX2_X1 U9554 ( .A(n7734), .B(P1_REG2_REG_2__SCAN_IN), .S(n9987), .Z(n7743)
         );
  NAND2_X1 U9555 ( .A1(n7736), .A2(n7735), .ZN(n7741) );
  OAI22_X1 U9556 ( .A1(n9622), .A2(n5949), .B1(n9978), .B2(n7737), .ZN(n7738)
         );
  AOI21_X1 U9557 ( .B1(n7739), .B2(n9637), .A(n7738), .ZN(n7740) );
  NAND2_X1 U9558 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  OR2_X1 U9559 ( .A1(n7743), .A2(n7742), .ZN(P1_U3291) );
  OAI222_X1 U9560 ( .A1(n9797), .A2(n7745), .B1(n9800), .B2(n7744), .C1(
        P1_U3086), .C2(n6034), .ZN(P1_U3333) );
  OAI222_X1 U9561 ( .A1(P2_U3151), .A2(n7748), .B1(n8907), .B2(n7747), .C1(
        n7746), .C2(n8899), .ZN(P2_U3267) );
  AOI22_X1 U9562 ( .A1(n10048), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n7749), .ZN(n7750) );
  OAI21_X1 U9563 ( .B1(n7751), .B2(n8907), .A(n7750), .ZN(P2_U3287) );
  INV_X1 U9564 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7759) );
  OAI21_X1 U9565 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7753), .A(n7752), .ZN(n7754) );
  OAI21_X1 U9566 ( .B1(n7755), .B2(n8589), .A(n7754), .ZN(n7756) );
  OAI21_X1 U9567 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7766), .A(n7756), .ZN(n7757) );
  AOI21_X1 U9568 ( .B1(n10049), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7757), .ZN(
        n7758) );
  OAI21_X1 U9569 ( .B1(n7759), .B2(n8587), .A(n7758), .ZN(P2_U3182) );
  AOI22_X1 U9570 ( .A1(n8439), .A2(n8276), .B1(n7760), .B2(n8456), .ZN(n7763)
         );
  NAND2_X1 U9571 ( .A1(n7761), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7762) );
  OAI211_X1 U9572 ( .C1(n5025), .C2(n8453), .A(n7763), .B(n7762), .ZN(P2_U3172) );
  INV_X1 U9573 ( .A(n7764), .ZN(n7768) );
  OAI21_X1 U9574 ( .B1(n8756), .B2(n7766), .A(n7765), .ZN(n7767) );
  AOI21_X1 U9575 ( .B1(n7768), .B2(n8276), .A(n7767), .ZN(n7770) );
  MUX2_X1 U9576 ( .A(n7770), .B(n7769), .S(n8767), .Z(n7771) );
  OAI21_X1 U9577 ( .B1(n8698), .B2(n7772), .A(n7771), .ZN(P2_U3233) );
  OAI222_X1 U9578 ( .A1(n7775), .A2(P2_U3151), .B1(n8331), .B2(n7774), .C1(
        n7773), .C2(n8899), .ZN(P2_U3271) );
  NAND2_X1 U9579 ( .A1(n7952), .A2(n7958), .ZN(n7789) );
  INV_X1 U9580 ( .A(n7942), .ZN(n9440) );
  AND2_X1 U9581 ( .A1(n7940), .A2(n7776), .ZN(n7841) );
  INV_X1 U9582 ( .A(n7841), .ZN(n7778) );
  INV_X1 U9583 ( .A(n7777), .ZN(n7947) );
  AOI21_X1 U9584 ( .B1(n9440), .B2(n7778), .A(n7947), .ZN(n7779) );
  INV_X1 U9585 ( .A(n7785), .ZN(n7946) );
  OAI21_X1 U9586 ( .B1(n7779), .B2(n7946), .A(n7957), .ZN(n7784) );
  INV_X1 U9587 ( .A(n7923), .ZN(n7782) );
  NOR4_X1 U9588 ( .A1(n7789), .A2(n7784), .A3(n7782), .A4(n7780), .ZN(n8027)
         );
  OAI211_X1 U9589 ( .C1(n7782), .C2(n7913), .A(n9462), .B(n7925), .ZN(n7783)
         );
  NOR2_X1 U9590 ( .A1(n7942), .A2(n7783), .ZN(n7786) );
  AOI21_X1 U9591 ( .B1(n7786), .B2(n7785), .A(n7784), .ZN(n7787) );
  NAND2_X1 U9592 ( .A1(n7962), .A2(n7956), .ZN(n7950) );
  NOR2_X1 U9593 ( .A1(n7787), .A2(n7950), .ZN(n7790) );
  NAND2_X1 U9594 ( .A1(n9351), .A2(n7954), .ZN(n7964) );
  INV_X1 U9595 ( .A(n7964), .ZN(n7788) );
  OAI21_X1 U9596 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n7988) );
  AOI21_X1 U9597 ( .B1(n8027), .B2(n7781), .A(n7988), .ZN(n7792) );
  INV_X1 U9598 ( .A(n9265), .ZN(n7791) );
  OAI21_X1 U9599 ( .B1(n9363), .B2(n7791), .A(n7963), .ZN(n8029) );
  OAI22_X1 U9600 ( .A1(n7792), .A2(n8029), .B1(n9732), .B2(n9264), .ZN(n7795)
         );
  INV_X1 U9601 ( .A(n9363), .ZN(n9649) );
  NAND2_X1 U9602 ( .A1(n7973), .A2(n9357), .ZN(n7833) );
  OAI21_X1 U9603 ( .B1(n9649), .B2(n9265), .A(n7833), .ZN(n8032) );
  INV_X1 U9604 ( .A(n9264), .ZN(n7793) );
  NOR2_X1 U9605 ( .A1(n7793), .A2(n9357), .ZN(n7971) );
  INV_X1 U9606 ( .A(n7971), .ZN(n7794) );
  OAI22_X1 U9607 ( .A1(n7795), .A2(n8032), .B1(n7973), .B2(n7794), .ZN(n7798)
         );
  INV_X1 U9608 ( .A(n7986), .ZN(n8034) );
  INV_X1 U9609 ( .A(n7983), .ZN(n7796) );
  AOI211_X1 U9610 ( .C1(n7798), .C2(n8034), .A(n7797), .B(n7796), .ZN(n7836)
         );
  OR2_X1 U9611 ( .A1(n7973), .A2(n9357), .ZN(n7799) );
  NAND2_X1 U9612 ( .A1(n7983), .A2(n7799), .ZN(n8036) );
  INV_X1 U9613 ( .A(n9494), .ZN(n9490) );
  INV_X1 U9614 ( .A(n9544), .ZN(n9540) );
  NOR2_X1 U9615 ( .A1(n6856), .A2(n7800), .ZN(n7805) );
  INV_X1 U9616 ( .A(n7801), .ZN(n7804) );
  AND2_X1 U9617 ( .A1(n9288), .A2(n9976), .ZN(n7991) );
  NOR2_X1 U9618 ( .A1(n7802), .A2(n7991), .ZN(n9994) );
  NAND4_X1 U9619 ( .A1(n7805), .A2(n7804), .A3(n9994), .A4(n7803), .ZN(n7810)
         );
  NAND2_X1 U9620 ( .A1(n7807), .A2(n7806), .ZN(n7809) );
  NOR3_X1 U9621 ( .A1(n7810), .A2(n7809), .A3(n7808), .ZN(n7816) );
  INV_X1 U9622 ( .A(n7811), .ZN(n7815) );
  INV_X1 U9623 ( .A(n7812), .ZN(n8003) );
  INV_X1 U9624 ( .A(n7813), .ZN(n7814) );
  AND4_X1 U9625 ( .A1(n7816), .A2(n7815), .A3(n8003), .A4(n7814), .ZN(n7819)
         );
  INV_X1 U9626 ( .A(n7817), .ZN(n7818) );
  NAND3_X1 U9627 ( .A1(n7820), .A2(n7819), .A3(n7818), .ZN(n7821) );
  NOR2_X1 U9628 ( .A1(n7883), .A2(n7821), .ZN(n7822) );
  NAND4_X1 U9629 ( .A1(n9576), .A2(n5777), .A3(n7822), .A4(n9592), .ZN(n7823)
         );
  NOR2_X1 U9630 ( .A1(n7823), .A2(n9560), .ZN(n7824) );
  NAND3_X1 U9631 ( .A1(n9529), .A2(n9540), .A3(n7824), .ZN(n7825) );
  NOR2_X1 U9632 ( .A1(n9515), .A2(n7825), .ZN(n7826) );
  NAND4_X1 U9633 ( .A1(n9461), .A2(n9474), .A3(n9490), .A4(n7826), .ZN(n7827)
         );
  NOR2_X1 U9634 ( .A1(n9438), .A2(n7827), .ZN(n7828) );
  NAND3_X1 U9635 ( .A1(n9407), .A2(n5901), .A3(n7828), .ZN(n7829) );
  NOR2_X1 U9636 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND4_X1 U9637 ( .A1(n7833), .A2(n9353), .A3(n7832), .A4(n7831), .ZN(n7834)
         );
  INV_X1 U9638 ( .A(n7979), .ZN(n7835) );
  NOR2_X1 U9639 ( .A1(n7836), .A2(n7835), .ZN(n7838) );
  INV_X1 U9640 ( .A(n9462), .ZN(n7839) );
  NOR2_X1 U9641 ( .A1(n7942), .A2(n7839), .ZN(n7840) );
  MUX2_X1 U9642 ( .A(n7841), .B(n7840), .S(n7984), .Z(n7945) );
  INV_X1 U9643 ( .A(n7997), .ZN(n7845) );
  NOR2_X1 U9644 ( .A1(n8001), .A2(n7845), .ZN(n7844) );
  NAND2_X1 U9645 ( .A1(n7842), .A2(n7852), .ZN(n7843) );
  INV_X1 U9646 ( .A(n7984), .ZN(n7975) );
  MUX2_X1 U9647 ( .A(n7844), .B(n7843), .S(n7975), .Z(n7853) );
  OAI21_X1 U9648 ( .B1(n7853), .B2(n7845), .A(n7855), .ZN(n7847) );
  NAND2_X1 U9649 ( .A1(n7859), .A2(n7856), .ZN(n7846) );
  AOI21_X1 U9650 ( .B1(n7847), .B2(n7851), .A(n7846), .ZN(n7850) );
  NAND4_X1 U9651 ( .A1(n7848), .A2(n7975), .A3(n7865), .A4(n8002), .ZN(n7849)
         );
  AND2_X1 U9652 ( .A1(n7852), .A2(n7851), .ZN(n7998) );
  NAND2_X1 U9653 ( .A1(n7853), .A2(n7998), .ZN(n7860) );
  NAND2_X1 U9654 ( .A1(n7855), .A2(n7854), .ZN(n7858) );
  INV_X1 U9655 ( .A(n7856), .ZN(n7857) );
  AOI21_X1 U9656 ( .B1(n7998), .B2(n7858), .A(n7857), .ZN(n7999) );
  NAND3_X1 U9657 ( .A1(n7860), .A2(n7999), .A3(n7859), .ZN(n7862) );
  INV_X1 U9658 ( .A(n7861), .ZN(n7864) );
  NAND4_X1 U9659 ( .A1(n7862), .A2(n7864), .A3(n7984), .A4(n8002), .ZN(n7872)
         );
  NAND3_X1 U9660 ( .A1(n7864), .A2(n7984), .A3(n7863), .ZN(n7868) );
  INV_X1 U9661 ( .A(n7865), .ZN(n9952) );
  OAI21_X1 U9662 ( .B1(n9952), .B2(n7866), .A(n7975), .ZN(n7867) );
  OAI211_X1 U9663 ( .C1(n7869), .C2(n7975), .A(n7868), .B(n7867), .ZN(n7870)
         );
  INV_X1 U9664 ( .A(n7870), .ZN(n7871) );
  NAND2_X1 U9665 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  NAND2_X1 U9666 ( .A1(n7874), .A2(n7873), .ZN(n7892) );
  AOI21_X1 U9667 ( .B1(n7892), .B2(n7876), .A(n7875), .ZN(n7878) );
  OAI211_X1 U9668 ( .C1(n7878), .C2(n7877), .A(n7889), .B(n7887), .ZN(n7881)
         );
  NAND3_X1 U9669 ( .A1(n8009), .A2(n7975), .A3(n7885), .ZN(n7879) );
  NOR2_X1 U9670 ( .A1(n7883), .A2(n7879), .ZN(n7880) );
  NAND2_X1 U9671 ( .A1(n7881), .A2(n7880), .ZN(n7898) );
  AND2_X1 U9672 ( .A1(n7890), .A2(n7975), .ZN(n7882) );
  NOR2_X1 U9673 ( .A1(n7883), .A2(n7882), .ZN(n7895) );
  NAND2_X1 U9674 ( .A1(n7885), .A2(n7884), .ZN(n8005) );
  OR2_X1 U9675 ( .A1(n8005), .A2(n7886), .ZN(n7891) );
  OR2_X1 U9676 ( .A1(n8005), .A2(n7887), .ZN(n7888) );
  AND3_X1 U9677 ( .A1(n7890), .A2(n7889), .A3(n7888), .ZN(n8008) );
  OAI21_X1 U9678 ( .B1(n7892), .B2(n7891), .A(n8008), .ZN(n7893) );
  NAND4_X1 U9679 ( .A1(n7893), .A2(n5777), .A3(n7984), .A4(n8009), .ZN(n7894)
         );
  OAI21_X1 U9680 ( .B1(n7895), .B2(n9611), .A(n7894), .ZN(n7897) );
  NAND2_X1 U9681 ( .A1(n7905), .A2(n7896), .ZN(n7990) );
  INV_X1 U9682 ( .A(n8010), .ZN(n7900) );
  NOR2_X1 U9683 ( .A1(n7990), .A2(n8013), .ZN(n7899) );
  MUX2_X1 U9684 ( .A(n7900), .B(n7899), .S(n7975), .Z(n7902) );
  NOR2_X1 U9685 ( .A1(n9784), .A2(n7901), .ZN(n8016) );
  INV_X1 U9686 ( .A(n8016), .ZN(n7903) );
  NAND2_X1 U9687 ( .A1(n7903), .A2(n8014), .ZN(n7904) );
  NAND2_X1 U9688 ( .A1(n7904), .A2(n7984), .ZN(n7907) );
  OAI21_X1 U9689 ( .B1(n7975), .B2(n7905), .A(n9576), .ZN(n7906) );
  INV_X1 U9690 ( .A(n8020), .ZN(n7909) );
  NAND2_X1 U9691 ( .A1(n7911), .A2(n8019), .ZN(n7908) );
  MUX2_X1 U9692 ( .A(n7909), .B(n7908), .S(n7975), .Z(n7910) );
  AND2_X1 U9693 ( .A1(n7918), .A2(n7911), .ZN(n8026) );
  OAI21_X1 U9694 ( .B1(n7917), .B2(n7912), .A(n8026), .ZN(n7915) );
  AND2_X1 U9695 ( .A1(n7919), .A2(n7916), .ZN(n8023) );
  NAND3_X1 U9696 ( .A1(n7913), .A2(n7989), .A3(n7984), .ZN(n7914) );
  AOI21_X1 U9697 ( .B1(n7915), .B2(n8023), .A(n7914), .ZN(n7926) );
  NAND3_X1 U9698 ( .A1(n7917), .A2(n7916), .A3(n9543), .ZN(n7922) );
  AND2_X1 U9699 ( .A1(n7989), .A2(n7918), .ZN(n7921) );
  NAND3_X1 U9700 ( .A1(n9492), .A2(n7975), .A3(n7919), .ZN(n7920) );
  AOI21_X1 U9701 ( .B1(n7922), .B2(n7921), .A(n7920), .ZN(n7924) );
  AOI22_X1 U9702 ( .A1(n7926), .A2(n7925), .B1(n7924), .B2(n7923), .ZN(n7939)
         );
  NAND2_X1 U9703 ( .A1(n9269), .A2(n7984), .ZN(n7927) );
  OAI22_X1 U9704 ( .A1(n9521), .A2(n7927), .B1(n9477), .B2(n7975), .ZN(n7932)
         );
  NAND2_X1 U9705 ( .A1(n9501), .A2(n7975), .ZN(n7933) );
  OAI21_X1 U9706 ( .B1(n9268), .B2(n7933), .A(n9521), .ZN(n7931) );
  INV_X1 U9707 ( .A(n7927), .ZN(n7928) );
  AND2_X1 U9708 ( .A1(n7928), .A2(n9268), .ZN(n7929) );
  OR2_X1 U9709 ( .A1(n9521), .A2(n7929), .ZN(n7930) );
  AOI22_X1 U9710 ( .A1(n9508), .A2(n7932), .B1(n7931), .B2(n7930), .ZN(n7938)
         );
  INV_X1 U9711 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U9712 ( .A1(n9521), .A2(n7934), .ZN(n7935) );
  OAI21_X1 U9713 ( .B1(n7984), .B2(n9268), .A(n7935), .ZN(n7936) );
  NAND2_X1 U9714 ( .A1(n9757), .A2(n7936), .ZN(n7937) );
  NAND4_X1 U9715 ( .A1(n7939), .A2(n9474), .A3(n7938), .A4(n7937), .ZN(n7944)
         );
  INV_X1 U9716 ( .A(n7940), .ZN(n7941) );
  MUX2_X1 U9717 ( .A(n7942), .B(n7941), .S(n7984), .Z(n7943) );
  MUX2_X1 U9718 ( .A(n7947), .B(n7946), .S(n7984), .Z(n7948) );
  INV_X1 U9719 ( .A(n7957), .ZN(n7949) );
  NOR2_X1 U9720 ( .A1(n7960), .A2(n7949), .ZN(n7951) );
  OAI21_X1 U9721 ( .B1(n7951), .B2(n7950), .A(n7958), .ZN(n7955) );
  INV_X1 U9722 ( .A(n7963), .ZN(n7953) );
  INV_X1 U9723 ( .A(n7952), .ZN(n7961) );
  AOI211_X1 U9724 ( .C1(n7955), .C2(n7954), .A(n7953), .B(n7961), .ZN(n7968)
         );
  INV_X1 U9725 ( .A(n7956), .ZN(n7959) );
  OAI21_X1 U9726 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(n7966) );
  INV_X1 U9727 ( .A(n9351), .ZN(n7967) );
  NAND2_X1 U9728 ( .A1(n9363), .A2(n9265), .ZN(n7970) );
  MUX2_X1 U9729 ( .A(n9363), .B(n9265), .S(n7984), .Z(n7969) );
  MUX2_X1 U9730 ( .A(n7974), .B(n7984), .S(n7973), .Z(n7972) );
  MUX2_X1 U9731 ( .A(n7975), .B(n7974), .S(n7973), .Z(n7976) );
  NOR3_X1 U9732 ( .A1(n7976), .A2(n9357), .A3(n9340), .ZN(n7977) );
  OAI21_X1 U9733 ( .B1(n7982), .B2(n6034), .A(n7993), .ZN(n7980) );
  NAND2_X1 U9734 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  AOI211_X1 U9735 ( .C1(n7986), .C2(n9330), .A(n8049), .B(n7985), .ZN(n7987)
         );
  INV_X1 U9736 ( .A(n9983), .ZN(n8039) );
  INV_X1 U9737 ( .A(n7988), .ZN(n8031) );
  INV_X1 U9738 ( .A(n7990), .ZN(n8018) );
  INV_X1 U9739 ( .A(n7991), .ZN(n7994) );
  NAND2_X1 U9740 ( .A1(n6084), .A2(n5991), .ZN(n7992) );
  NAND4_X1 U9741 ( .A1(n7995), .A2(n7994), .A3(n7993), .A4(n7992), .ZN(n7996)
         );
  NAND3_X1 U9742 ( .A1(n7998), .A2(n7997), .A3(n7996), .ZN(n8000) );
  OAI21_X1 U9743 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(n8004) );
  NAND3_X1 U9744 ( .A1(n8004), .A2(n8003), .A3(n8002), .ZN(n8007) );
  AOI21_X1 U9745 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8012) );
  INV_X1 U9746 ( .A(n8008), .ZN(n8011) );
  OAI211_X1 U9747 ( .C1(n8012), .C2(n8011), .A(n8010), .B(n8009), .ZN(n8015)
         );
  NAND3_X1 U9748 ( .A1(n8015), .A2(n8014), .A3(n8013), .ZN(n8017) );
  AOI21_X1 U9749 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8022) );
  INV_X1 U9750 ( .A(n8019), .ZN(n8021) );
  OAI211_X1 U9751 ( .C1(n8022), .C2(n8021), .A(n9543), .B(n8020), .ZN(n8025)
         );
  INV_X1 U9752 ( .A(n8023), .ZN(n8024) );
  AOI21_X1 U9753 ( .B1(n8026), .B2(n8025), .A(n8024), .ZN(n8028) );
  OAI21_X1 U9754 ( .B1(n4632), .B2(n8028), .A(n8027), .ZN(n8030) );
  AOI21_X1 U9755 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n8033) );
  NOR2_X1 U9756 ( .A1(n8033), .A2(n8032), .ZN(n8035) );
  OAI21_X1 U9757 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8037) );
  MUX2_X1 U9758 ( .A(n8039), .B(n8038), .S(n8037), .Z(n8040) );
  NAND2_X1 U9759 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NOR3_X1 U9760 ( .A1(n8048), .A2(n8047), .A3(n8046), .ZN(n8051) );
  OAI21_X1 U9761 ( .B1(n8052), .B2(n8049), .A(P1_B_REG_SCAN_IN), .ZN(n8050) );
  OAI22_X1 U9762 ( .A1(n8053), .A2(n8052), .B1(n8051), .B2(n8050), .ZN(
        P1_U3242) );
  INV_X1 U9763 ( .A(n8054), .ZN(n8055) );
  XNOR2_X1 U9764 ( .A(n8829), .B(n8090), .ZN(n8388) );
  XNOR2_X1 U9765 ( .A(n8891), .B(n8074), .ZN(n8057) );
  NAND2_X1 U9766 ( .A1(n8057), .A2(n8391), .ZN(n8436) );
  OAI21_X1 U9767 ( .B1(n8057), .B2(n8391), .A(n8436), .ZN(n8401) );
  XNOR2_X1 U9768 ( .A(n8823), .B(n8090), .ZN(n8058) );
  NAND2_X1 U9769 ( .A1(n8058), .A2(n8776), .ZN(n8359) );
  INV_X1 U9770 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U9771 ( .A1(n8059), .A2(n8462), .ZN(n8060) );
  AND2_X1 U9772 ( .A1(n8359), .A2(n8060), .ZN(n8437) );
  XNOR2_X1 U9773 ( .A(n8817), .B(n8074), .ZN(n8061) );
  NAND2_X1 U9774 ( .A1(n8061), .A2(n8729), .ZN(n8415) );
  INV_X1 U9775 ( .A(n8061), .ZN(n8062) );
  INV_X1 U9776 ( .A(n8729), .ZN(n8753) );
  NAND2_X1 U9777 ( .A1(n8062), .A2(n8753), .ZN(n8063) );
  INV_X1 U9778 ( .A(n8360), .ZN(n8064) );
  OR2_X1 U9779 ( .A1(n8064), .A2(n8359), .ZN(n8065) );
  INV_X1 U9780 ( .A(n8065), .ZN(n8066) );
  XNOR2_X1 U9781 ( .A(n8734), .B(n8074), .ZN(n8067) );
  NAND2_X1 U9782 ( .A1(n8067), .A2(n8740), .ZN(n8070) );
  INV_X1 U9783 ( .A(n8067), .ZN(n8068) );
  INV_X1 U9784 ( .A(n8740), .ZN(n8719) );
  NAND2_X1 U9785 ( .A1(n8068), .A2(n8719), .ZN(n8069) );
  AND2_X1 U9786 ( .A1(n8070), .A2(n8069), .ZN(n8416) );
  NAND2_X1 U9787 ( .A1(n8417), .A2(n8070), .ZN(n8369) );
  XNOR2_X1 U9788 ( .A(n8873), .B(n6650), .ZN(n8071) );
  XNOR2_X1 U9789 ( .A(n8071), .B(n8730), .ZN(n8370) );
  NAND2_X1 U9790 ( .A1(n8369), .A2(n8370), .ZN(n8368) );
  XNOR2_X1 U9791 ( .A(n8867), .B(n8074), .ZN(n8425) );
  XNOR2_X1 U9792 ( .A(n8861), .B(n8074), .ZN(n8075) );
  NAND2_X1 U9793 ( .A1(n8352), .A2(n8430), .ZN(n8378) );
  INV_X1 U9794 ( .A(n8075), .ZN(n8076) );
  NAND2_X1 U9795 ( .A1(n8077), .A2(n8076), .ZN(n8377) );
  XNOR2_X1 U9796 ( .A(n8683), .B(n8090), .ZN(n8084) );
  NAND2_X1 U9797 ( .A1(n8084), .A2(n8693), .ZN(n8379) );
  XNOR2_X1 U9798 ( .A(n8851), .B(n8090), .ZN(n8081) );
  INV_X1 U9799 ( .A(n8081), .ZN(n8078) );
  NAND2_X1 U9800 ( .A1(n8078), .A2(n8080), .ZN(n8079) );
  AND2_X1 U9801 ( .A1(n8379), .A2(n8079), .ZN(n8083) );
  AND2_X1 U9802 ( .A1(n8377), .A2(n8083), .ZN(n8086) );
  INV_X1 U9803 ( .A(n8079), .ZN(n8082) );
  XNOR2_X1 U9804 ( .A(n8081), .B(n8080), .ZN(n8382) );
  INV_X1 U9805 ( .A(n8083), .ZN(n8085) );
  XNOR2_X1 U9806 ( .A(n8084), .B(n8665), .ZN(n8409) );
  XNOR2_X1 U9807 ( .A(n8845), .B(n8090), .ZN(n8087) );
  XNOR2_X1 U9808 ( .A(n8087), .B(n8644), .ZN(n8448) );
  INV_X1 U9809 ( .A(n8087), .ZN(n8088) );
  NAND2_X1 U9810 ( .A1(n8088), .A2(n8644), .ZN(n8089) );
  XNOR2_X1 U9811 ( .A(n8792), .B(n8090), .ZN(n8091) );
  NAND2_X1 U9812 ( .A1(n8091), .A2(n8656), .ZN(n8092) );
  OAI21_X1 U9813 ( .B1(n8091), .B2(n8656), .A(n8092), .ZN(n8343) );
  XNOR2_X1 U9814 ( .A(n8302), .B(n8090), .ZN(n8093) );
  XNOR2_X1 U9815 ( .A(n8094), .B(n8093), .ZN(n8101) );
  INV_X1 U9816 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8095) );
  OAI22_X1 U9817 ( .A1(n8454), .A2(n8429), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8095), .ZN(n8099) );
  INV_X1 U9818 ( .A(n8635), .ZN(n8096) );
  OAI22_X1 U9819 ( .A1(n8097), .A2(n8453), .B1(n8096), .B2(n8404), .ZN(n8098)
         );
  AOI211_X1 U9820 ( .C1(n8636), .C2(n8456), .A(n8099), .B(n8098), .ZN(n8100)
         );
  OAI21_X1 U9821 ( .B1(n8101), .B2(n8458), .A(n8100), .ZN(P2_U3160) );
  INV_X1 U9822 ( .A(n8102), .ZN(n9796) );
  OAI22_X1 U9823 ( .A1(n9796), .A2(n8103), .B1(n8253), .B2(n8900), .ZN(n8307)
         );
  MUX2_X1 U9824 ( .A(n8461), .B(n8636), .S(n8256), .Z(n8250) );
  INV_X1 U9825 ( .A(n8106), .ZN(n8105) );
  AND2_X1 U9826 ( .A1(n8106), .A2(n6643), .ZN(n8109) );
  OAI21_X1 U9827 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n8110) );
  NAND2_X1 U9828 ( .A1(n8136), .A2(n8112), .ZN(n8115) );
  NAND2_X1 U9829 ( .A1(n8121), .A2(n8113), .ZN(n8114) );
  MUX2_X1 U9830 ( .A(n8115), .B(n8114), .S(n8264), .Z(n8116) );
  INV_X1 U9831 ( .A(n8116), .ZN(n8117) );
  INV_X1 U9832 ( .A(n8121), .ZN(n8124) );
  OAI211_X1 U9833 ( .C1(n8140), .C2(n8124), .A(n8123), .B(n8122), .ZN(n8125)
         );
  NAND3_X1 U9834 ( .A1(n8125), .A2(n8143), .A3(n8137), .ZN(n8128) );
  NAND4_X1 U9835 ( .A1(n8128), .A2(n8149), .A3(n8287), .A4(n8127), .ZN(n8135)
         );
  INV_X1 U9836 ( .A(n8129), .ZN(n8132) );
  OAI21_X1 U9837 ( .B1(n8132), .B2(n8131), .A(n8130), .ZN(n8133) );
  NOR2_X1 U9838 ( .A1(n8156), .A2(n8133), .ZN(n8134) );
  NAND2_X1 U9839 ( .A1(n8135), .A2(n8134), .ZN(n8155) );
  INV_X1 U9840 ( .A(n8136), .ZN(n8139) );
  NAND2_X1 U9841 ( .A1(n5481), .A2(n10076), .ZN(n8138) );
  OAI211_X1 U9842 ( .C1(n8140), .C2(n8139), .A(n8138), .B(n8137), .ZN(n8142)
         );
  NAND2_X1 U9843 ( .A1(n8142), .A2(n8141), .ZN(n8144) );
  NAND3_X1 U9844 ( .A1(n8144), .A2(n8287), .A3(n8143), .ZN(n8148) );
  NAND2_X1 U9845 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  NAND3_X1 U9846 ( .A1(n8153), .A2(n8152), .A3(n8151), .ZN(n8154) );
  NAND2_X1 U9847 ( .A1(n5486), .A2(n8159), .ZN(n8158) );
  AND2_X1 U9848 ( .A1(n8158), .A2(n8157), .ZN(n8163) );
  INV_X1 U9849 ( .A(n8159), .ZN(n8160) );
  NOR2_X1 U9850 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  MUX2_X1 U9851 ( .A(n8163), .B(n8162), .S(n8256), .Z(n8164) );
  INV_X1 U9852 ( .A(n8164), .ZN(n8165) );
  NAND2_X1 U9853 ( .A1(n8167), .A2(n8293), .ZN(n8173) );
  NAND2_X1 U9854 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  MUX2_X1 U9855 ( .A(n8171), .B(n8170), .S(n8256), .Z(n8172) );
  NAND2_X1 U9856 ( .A1(n8173), .A2(n8172), .ZN(n8179) );
  MUX2_X1 U9857 ( .A(n8466), .B(n8174), .S(n8256), .Z(n8175) );
  OAI21_X1 U9858 ( .B1(n8179), .B2(n8176), .A(n8175), .ZN(n8182) );
  INV_X1 U9859 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U9860 ( .A1(n8179), .A2(n8178), .ZN(n8181) );
  MUX2_X1 U9861 ( .A(n8184), .B(n8183), .S(n8264), .Z(n8185) );
  INV_X1 U9862 ( .A(n8186), .ZN(n8295) );
  NAND3_X1 U9863 ( .A1(n8188), .A2(n8264), .A3(n8195), .ZN(n8190) );
  INV_X1 U9864 ( .A(n8771), .ZN(n8189) );
  NAND2_X1 U9865 ( .A1(n8190), .A2(n8189), .ZN(n8194) );
  NAND2_X1 U9866 ( .A1(n8205), .A2(n8191), .ZN(n8192) );
  NAND2_X1 U9867 ( .A1(n8192), .A2(n8264), .ZN(n8193) );
  NAND2_X1 U9868 ( .A1(n8194), .A2(n8193), .ZN(n8201) );
  NAND3_X1 U9869 ( .A1(n8197), .A2(n8196), .A3(n8195), .ZN(n8199) );
  NAND3_X1 U9870 ( .A1(n8199), .A2(n8256), .A3(n8198), .ZN(n8200) );
  NAND2_X1 U9871 ( .A1(n8201), .A2(n8200), .ZN(n8208) );
  NAND2_X1 U9872 ( .A1(n8742), .A2(n8204), .ZN(n8202) );
  NOR2_X1 U9873 ( .A1(n8208), .A2(n8202), .ZN(n8210) );
  AND2_X1 U9874 ( .A1(n8204), .A2(n8203), .ZN(n8207) );
  NAND2_X1 U9875 ( .A1(n8212), .A2(n8205), .ZN(n8206) );
  AOI21_X1 U9876 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8209) );
  NAND2_X1 U9877 ( .A1(n8727), .A2(n8211), .ZN(n8214) );
  NAND2_X1 U9878 ( .A1(n8713), .A2(n8212), .ZN(n8213) );
  MUX2_X1 U9879 ( .A(n8214), .B(n8213), .S(n8264), .Z(n8216) );
  AOI21_X1 U9880 ( .B1(n8219), .B2(n8217), .A(n8256), .ZN(n8218) );
  NOR2_X1 U9881 ( .A1(n8220), .A2(n8256), .ZN(n8221) );
  INV_X1 U9882 ( .A(n8222), .ZN(n8223) );
  NOR2_X1 U9883 ( .A1(n8274), .A2(n8223), .ZN(n8224) );
  MUX2_X1 U9884 ( .A(n8225), .B(n8224), .S(n8264), .Z(n8226) );
  NAND2_X1 U9885 ( .A1(n8227), .A2(n8226), .ZN(n8232) );
  INV_X1 U9886 ( .A(n8674), .ZN(n8273) );
  OR2_X1 U9887 ( .A1(n8232), .A2(n8273), .ZN(n8230) );
  NOR2_X1 U9888 ( .A1(n8271), .A2(n8274), .ZN(n8229) );
  INV_X1 U9889 ( .A(n8272), .ZN(n8228) );
  AOI21_X1 U9890 ( .B1(n8232), .B2(n8231), .A(n8271), .ZN(n8233) );
  MUX2_X1 U9891 ( .A(n8235), .B(n8234), .S(n8264), .Z(n8236) );
  MUX2_X1 U9892 ( .A(n8238), .B(n4433), .S(n8264), .Z(n8239) );
  NOR2_X1 U9893 ( .A1(n8641), .A2(n8239), .ZN(n8240) );
  NAND2_X1 U9894 ( .A1(n8241), .A2(n8240), .ZN(n8245) );
  MUX2_X1 U9895 ( .A(n8243), .B(n8242), .S(n8256), .Z(n8244) );
  NAND2_X1 U9896 ( .A1(n8251), .A2(n8250), .ZN(n8265) );
  NAND2_X1 U9897 ( .A1(n8326), .A2(n8252), .ZN(n8255) );
  OR2_X1 U9898 ( .A1(n8253), .A2(n8905), .ZN(n8254) );
  INV_X1 U9899 ( .A(n8460), .ZN(n8263) );
  OAI21_X1 U9900 ( .B1(n8263), .B2(n8256), .A(n8311), .ZN(n8257) );
  INV_X1 U9901 ( .A(n8257), .ZN(n8259) );
  INV_X1 U9902 ( .A(n8261), .ZN(n8262) );
  AOI21_X1 U9903 ( .B1(n8263), .B2(n8311), .A(n8262), .ZN(n8308) );
  NOR2_X1 U9904 ( .A1(n4799), .A2(n8264), .ZN(n8266) );
  OAI211_X1 U9905 ( .C1(n8267), .C2(n8461), .A(n8266), .B(n8265), .ZN(n8268)
         );
  NOR2_X1 U9906 ( .A1(n8307), .A2(n8628), .ZN(n8316) );
  INV_X1 U9907 ( .A(n8316), .ZN(n8304) );
  INV_X1 U9908 ( .A(n8270), .ZN(n8309) );
  INV_X1 U9909 ( .A(n8670), .ZN(n8300) );
  NAND2_X1 U9910 ( .A1(n4441), .A2(n8272), .ZN(n8679) );
  NOR2_X1 U9911 ( .A1(n6777), .A2(n8276), .ZN(n8280) );
  NAND4_X1 U9912 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), .ZN(n8284)
         );
  NOR4_X1 U9913 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n8288)
         );
  NAND4_X1 U9914 ( .A1(n8288), .A2(n8287), .A3(n5484), .A4(n8286), .ZN(n8289)
         );
  NOR4_X1 U9915 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n8294)
         );
  NAND4_X1 U9916 ( .A1(n8295), .A2(n4539), .A3(n8294), .A4(n8293), .ZN(n8296)
         );
  NOR4_X1 U9917 ( .A1(n8763), .A2(n8771), .A3(n5262), .A4(n8296), .ZN(n8297)
         );
  NAND4_X1 U9918 ( .A1(n8727), .A2(n8716), .A3(n8742), .A4(n8297), .ZN(n8298)
         );
  NOR4_X1 U9919 ( .A1(n8679), .A2(n8704), .A3(n8689), .A4(n8298), .ZN(n8299)
         );
  NAND3_X1 U9920 ( .A1(n8655), .A2(n8300), .A3(n8299), .ZN(n8301) );
  NOR4_X1 U9921 ( .A1(n8309), .A2(n8302), .A3(n8641), .A4(n8301), .ZN(n8303)
         );
  NAND4_X1 U9922 ( .A1(n8304), .A2(n8308), .A3(n8303), .A4(n8312), .ZN(n8305)
         );
  INV_X1 U9923 ( .A(n8307), .ZN(n8835) );
  AOI21_X1 U9924 ( .B1(n8313), .B2(n8312), .A(n8835), .ZN(n8315) );
  XNOR2_X1 U9925 ( .A(n8317), .B(n8609), .ZN(n8325) );
  NAND3_X1 U9926 ( .A1(n8320), .A2(n8319), .A3(n8318), .ZN(n8321) );
  OAI211_X1 U9927 ( .C1(n8322), .C2(n8324), .A(n8321), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8323) );
  OAI21_X1 U9928 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(P2_U3296) );
  INV_X1 U9929 ( .A(n8326), .ZN(n8906) );
  OAI222_X1 U9930 ( .A1(n8329), .A2(n8328), .B1(n9800), .B2(n8906), .C1(
        P1_U3086), .C2(n8327), .ZN(P1_U3325) );
  OAI222_X1 U9931 ( .A1(n5511), .A2(P2_U3151), .B1(n8331), .B2(n8330), .C1(
        n9007), .C2(n8899), .ZN(P2_U3275) );
  NAND2_X1 U9932 ( .A1(n8332), .A2(n8784), .ZN(n8629) );
  OAI21_X1 U9933 ( .B1(n8780), .B2(n8333), .A(n8629), .ZN(n8336) );
  NOR2_X1 U9934 ( .A1(n5510), .A2(n8334), .ZN(n8335) );
  OAI21_X1 U9935 ( .B1(n8339), .B2(n8767), .A(n8338), .ZN(P2_U3204) );
  INV_X1 U9936 ( .A(n8340), .ZN(n9799) );
  OAI222_X1 U9937 ( .A1(P2_U3151), .A2(n8342), .B1(n8907), .B2(n9799), .C1(
        n8341), .C2(n8899), .ZN(P2_U3266) );
  AOI21_X1 U9938 ( .B1(n8344), .B2(n8343), .A(n8458), .ZN(n8346) );
  NAND2_X1 U9939 ( .A1(n8346), .A2(n8345), .ZN(n8351) );
  INV_X1 U9940 ( .A(n8347), .ZN(n8649) );
  AOI22_X1 U9941 ( .A1(n8664), .A2(n8449), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8348) );
  OAI21_X1 U9942 ( .B1(n8649), .B2(n8404), .A(n8348), .ZN(n8349) );
  AOI21_X1 U9943 ( .B1(n8461), .B2(n8420), .A(n8349), .ZN(n8350) );
  OAI211_X1 U9944 ( .C1(n5438), .C2(n8446), .A(n8351), .B(n8350), .ZN(P2_U3154) );
  XNOR2_X1 U9945 ( .A(n8352), .B(n8707), .ZN(n8357) );
  AOI22_X1 U9946 ( .A1(n8665), .A2(n8420), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8354) );
  NAND2_X1 U9947 ( .A1(n8450), .A2(n8696), .ZN(n8353) );
  OAI211_X1 U9948 ( .C1(n8692), .C2(n8429), .A(n8354), .B(n8353), .ZN(n8355)
         );
  AOI21_X1 U9949 ( .B1(n5360), .B2(n8456), .A(n8355), .ZN(n8356) );
  OAI21_X1 U9950 ( .B1(n8357), .B2(n8458), .A(n8356), .ZN(P2_U3156) );
  AND2_X1 U9951 ( .A1(n8358), .A2(n8437), .ZN(n8440) );
  INV_X1 U9952 ( .A(n8359), .ZN(n8361) );
  NOR3_X1 U9953 ( .A1(n8440), .A2(n8361), .A3(n8360), .ZN(n8362) );
  OAI21_X1 U9954 ( .B1(n8362), .B2(n4314), .A(n8439), .ZN(n8366) );
  NAND2_X1 U9955 ( .A1(n8449), .A2(n8462), .ZN(n8363) );
  NAND2_X1 U9956 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8617) );
  OAI211_X1 U9957 ( .C1(n8740), .C2(n8453), .A(n8363), .B(n8617), .ZN(n8364)
         );
  AOI21_X1 U9958 ( .B1(n8450), .B2(n8744), .A(n8364), .ZN(n8365) );
  OAI211_X1 U9959 ( .C1(n8367), .C2(n8446), .A(n8366), .B(n8365), .ZN(P2_U3159) );
  INV_X1 U9960 ( .A(n8873), .ZN(n8376) );
  OAI21_X1 U9961 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8371) );
  NAND2_X1 U9962 ( .A1(n8371), .A2(n8439), .ZN(n8375) );
  AOI22_X1 U9963 ( .A1(n8718), .A2(n8420), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8372) );
  OAI21_X1 U9964 ( .B1(n8740), .B2(n8429), .A(n8372), .ZN(n8373) );
  AOI21_X1 U9965 ( .B1(n8722), .B2(n8450), .A(n8373), .ZN(n8374) );
  OAI211_X1 U9966 ( .C1(n8376), .C2(n8446), .A(n8375), .B(n8374), .ZN(P2_U3163) );
  NAND2_X1 U9967 ( .A1(n8378), .A2(n8377), .ZN(n8408) );
  NAND2_X1 U9968 ( .A1(n8408), .A2(n8409), .ZN(n8380) );
  NAND2_X1 U9969 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  XOR2_X1 U9970 ( .A(n8382), .B(n8381), .Z(n8387) );
  AOI22_X1 U9971 ( .A1(n8665), .A2(n8449), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8384) );
  NAND2_X1 U9972 ( .A1(n8667), .A2(n8450), .ZN(n8383) );
  OAI211_X1 U9973 ( .C1(n8644), .C2(n8453), .A(n8384), .B(n8383), .ZN(n8385)
         );
  AOI21_X1 U9974 ( .B1(n8851), .B2(n8456), .A(n8385), .ZN(n8386) );
  OAI21_X1 U9975 ( .B1(n8387), .B2(n8458), .A(n8386), .ZN(P2_U3165) );
  XNOR2_X1 U9976 ( .A(n8388), .B(n8774), .ZN(n8389) );
  XNOR2_X1 U9977 ( .A(n8390), .B(n8389), .ZN(n8398) );
  INV_X1 U9978 ( .A(n8391), .ZN(n8751) );
  NAND2_X1 U9979 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8532) );
  OAI21_X1 U9980 ( .B1(n8429), .B2(n8392), .A(n8532), .ZN(n8395) );
  NOR2_X1 U9981 ( .A1(n8404), .A2(n8393), .ZN(n8394) );
  AOI211_X1 U9982 ( .C1(n8420), .C2(n8751), .A(n8395), .B(n8394), .ZN(n8397)
         );
  NAND2_X1 U9983 ( .A1(n8829), .A2(n8456), .ZN(n8396) );
  OAI211_X1 U9984 ( .C1(n8398), .C2(n8458), .A(n8397), .B(n8396), .ZN(P2_U3166) );
  INV_X1 U9985 ( .A(n8399), .ZN(n8438) );
  AOI21_X1 U9986 ( .B1(n8401), .B2(n8400), .A(n8438), .ZN(n8407) );
  NAND2_X1 U9987 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8558) );
  OAI21_X1 U9988 ( .B1(n8453), .B2(n8776), .A(n8558), .ZN(n8402) );
  AOI21_X1 U9989 ( .B1(n8449), .B2(n8463), .A(n8402), .ZN(n8403) );
  OAI21_X1 U9990 ( .B1(n8782), .B2(n8404), .A(n8403), .ZN(n8405) );
  AOI21_X1 U9991 ( .B1(n8891), .B2(n8456), .A(n8405), .ZN(n8406) );
  OAI21_X1 U9992 ( .B1(n8407), .B2(n8458), .A(n8406), .ZN(P2_U3168) );
  XOR2_X1 U9993 ( .A(n8409), .B(n8408), .Z(n8414) );
  AOI22_X1 U9994 ( .A1(n8680), .A2(n8420), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8411) );
  NAND2_X1 U9995 ( .A1(n8450), .A2(n8685), .ZN(n8410) );
  OAI211_X1 U9996 ( .C1(n8430), .C2(n8429), .A(n8411), .B(n8410), .ZN(n8412)
         );
  AOI21_X1 U9997 ( .B1(n8856), .B2(n8456), .A(n8412), .ZN(n8413) );
  OAI21_X1 U9998 ( .B1(n8414), .B2(n8458), .A(n8413), .ZN(P2_U3169) );
  NOR3_X1 U9999 ( .A1(n4314), .A2(n4657), .A3(n8416), .ZN(n8419) );
  INV_X1 U10000 ( .A(n8417), .ZN(n8418) );
  OAI21_X1 U10001 ( .B1(n8419), .B2(n8418), .A(n8439), .ZN(n8424) );
  AOI22_X1 U10002 ( .A1(n8706), .A2(n8420), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8421) );
  OAI21_X1 U10003 ( .B1(n8729), .B2(n8429), .A(n8421), .ZN(n8422) );
  AOI21_X1 U10004 ( .B1(n8733), .B2(n8450), .A(n8422), .ZN(n8423) );
  OAI211_X1 U10005 ( .C1(n8879), .C2(n8446), .A(n8424), .B(n8423), .ZN(
        P2_U3173) );
  XNOR2_X1 U10006 ( .A(n8425), .B(n8692), .ZN(n8426) );
  XNOR2_X1 U10007 ( .A(n8427), .B(n8426), .ZN(n8435) );
  INV_X1 U10008 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8428) );
  OAI22_X1 U10009 ( .A1(n8730), .A2(n8429), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8428), .ZN(n8432) );
  NOR2_X1 U10010 ( .A1(n8430), .A2(n8453), .ZN(n8431) );
  AOI211_X1 U10011 ( .C1(n8710), .C2(n8450), .A(n8432), .B(n8431), .ZN(n8434)
         );
  NAND2_X1 U10012 ( .A1(n8867), .A2(n8456), .ZN(n8433) );
  OAI211_X1 U10013 ( .C1(n8435), .C2(n8458), .A(n8434), .B(n8433), .ZN(
        P2_U3175) );
  NOR3_X1 U10014 ( .A1(n8438), .A2(n4662), .A3(n8437), .ZN(n8441) );
  OAI21_X1 U10015 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8445) );
  NAND2_X1 U10016 ( .A1(n8449), .A2(n8751), .ZN(n8442) );
  NAND2_X1 U10017 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8592) );
  OAI211_X1 U10018 ( .C1(n8729), .C2(n8453), .A(n8442), .B(n8592), .ZN(n8443)
         );
  AOI21_X1 U10019 ( .B1(n8450), .B2(n8755), .A(n8443), .ZN(n8444) );
  OAI211_X1 U10020 ( .C1(n8823), .C2(n8446), .A(n8445), .B(n8444), .ZN(
        P2_U3178) );
  XOR2_X1 U10021 ( .A(n8448), .B(n8447), .Z(n8459) );
  AOI22_X1 U10022 ( .A1(n8680), .A2(n8449), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8452) );
  NAND2_X1 U10023 ( .A1(n8659), .A2(n8450), .ZN(n8451) );
  OAI211_X1 U10024 ( .C1(n8454), .C2(n8453), .A(n8452), .B(n8451), .ZN(n8455)
         );
  AOI21_X1 U10025 ( .B1(n8845), .B2(n8456), .A(n8455), .ZN(n8457) );
  OAI21_X1 U10026 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(P2_U3180) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8460), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8461), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8656), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10030 ( .A(n8664), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8588), .Z(
        P2_U3517) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8680), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8665), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10033 ( .A(n8707), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8588), .Z(
        P2_U3514) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8718), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8706), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8719), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8753), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8462), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8751), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8463), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8464), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8465), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10043 ( .A(n8466), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8588), .Z(
        P2_U3504) );
  MUX2_X1 U10044 ( .A(n8467), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8588), .Z(
        P2_U3503) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8468), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10046 ( .A(n8469), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8588), .Z(
        P2_U3501) );
  MUX2_X1 U10047 ( .A(n8470), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8588), .Z(
        P2_U3500) );
  MUX2_X1 U10048 ( .A(n8471), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8588), .Z(
        P2_U3499) );
  MUX2_X1 U10049 ( .A(n8472), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8588), .Z(
        P2_U3498) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8473), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10051 ( .A(n8474), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8588), .Z(
        P2_U3496) );
  MUX2_X1 U10052 ( .A(n5481), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8588), .Z(
        P2_U3495) );
  MUX2_X1 U10053 ( .A(n8475), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8588), .Z(
        P2_U3494) );
  MUX2_X1 U10054 ( .A(n8476), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8588), .Z(
        P2_U3493) );
  MUX2_X1 U10055 ( .A(n8477), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8588), .Z(
        P2_U3492) );
  NAND2_X1 U10056 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8507), .ZN(n8480) );
  OAI21_X1 U10057 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8507), .A(n8480), .ZN(
        n8481) );
  AOI21_X1 U10058 ( .B1(n8482), .B2(n8481), .A(n8502), .ZN(n8501) );
  MUX2_X1 U10059 ( .A(n8504), .B(n8483), .S(n8318), .Z(n8484) );
  OAI21_X1 U10060 ( .B1(n8505), .B2(n8484), .A(n4371), .ZN(n8487) );
  AOI21_X1 U10061 ( .B1(n8487), .B2(n4366), .A(n8516), .ZN(n8491) );
  NAND2_X1 U10062 ( .A1(n10049), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10063 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8489) );
  OAI211_X1 U10064 ( .C1(n8491), .C2(n10055), .A(n8490), .B(n8489), .ZN(n8499)
         );
  INV_X1 U10065 ( .A(n8492), .ZN(n8494) );
  NAND2_X1 U10066 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8507), .ZN(n8495) );
  OAI21_X1 U10067 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8507), .A(n8495), .ZN(
        n8496) );
  AOI21_X1 U10068 ( .B1(n4361), .B2(n8496), .A(n8509), .ZN(n8497) );
  NOR2_X1 U10069 ( .A1(n8497), .A2(n8624), .ZN(n8498) );
  AOI211_X1 U10070 ( .C1(n10047), .C2(n8505), .A(n8499), .B(n8498), .ZN(n8500)
         );
  OAI21_X1 U10071 ( .B1(n8501), .B2(n8620), .A(n8500), .ZN(P2_U3196) );
  INV_X1 U10072 ( .A(n8502), .ZN(n8503) );
  OAI21_X1 U10073 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8535) );
  XNOR2_X1 U10074 ( .A(n8535), .B(n8534), .ZN(n8506) );
  AOI21_X1 U10075 ( .B1(n8506), .B2(n8513), .A(n8537), .ZN(n8527) );
  AND2_X1 U10076 ( .A1(n8507), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8508) );
  NOR2_X1 U10077 ( .A1(n4359), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8511) );
  OAI21_X1 U10078 ( .B1(n8511), .B2(n8529), .A(n10050), .ZN(n8526) );
  MUX2_X1 U10079 ( .A(n8513), .B(n8512), .S(n8318), .Z(n8515) );
  AND2_X1 U10080 ( .A1(n8515), .A2(n8524), .ZN(n8545) );
  INV_X1 U10081 ( .A(n8545), .ZN(n8514) );
  OAI21_X1 U10082 ( .B1(n8524), .B2(n8515), .A(n8514), .ZN(n8518) );
  AOI21_X1 U10083 ( .B1(n8518), .B2(n8517), .A(n8544), .ZN(n8520) );
  OAI21_X1 U10084 ( .B1(n8520), .B2(n10055), .A(n8519), .ZN(n8523) );
  NOR2_X1 U10085 ( .A1(n8594), .A2(n8521), .ZN(n8522) );
  AOI211_X1 U10086 ( .C1(n10047), .C2(n8524), .A(n8523), .B(n8522), .ZN(n8525)
         );
  OAI211_X1 U10087 ( .C1(n8527), .C2(n8620), .A(n8526), .B(n8525), .ZN(
        P2_U3197) );
  AOI22_X1 U10088 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8547), .B1(n8561), .B2(
        n9075), .ZN(n8530) );
  NOR2_X1 U10089 ( .A1(n8531), .A2(n8530), .ZN(n8556) );
  AOI21_X1 U10090 ( .B1(n8531), .B2(n8530), .A(n8556), .ZN(n8555) );
  OAI21_X1 U10091 ( .B1(n8594), .B2(n8533), .A(n8532), .ZN(n8543) );
  AND2_X1 U10092 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  MUX2_X1 U10093 ( .A(n8546), .B(P2_REG2_REG_16__SCAN_IN), .S(n8547), .Z(n8538) );
  INV_X1 U10094 ( .A(n8538), .ZN(n8539) );
  AOI21_X1 U10095 ( .B1(n8540), .B2(n8539), .A(n8560), .ZN(n8541) );
  NOR2_X1 U10096 ( .A1(n8541), .A2(n8620), .ZN(n8542) );
  AOI211_X1 U10097 ( .C1(n10047), .C2(n8547), .A(n8543), .B(n8542), .ZN(n8554)
         );
  MUX2_X1 U10098 ( .A(n8546), .B(n9075), .S(n8318), .Z(n8548) );
  NAND2_X1 U10099 ( .A1(n8548), .A2(n8547), .ZN(n8566) );
  MUX2_X1 U10100 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8318), .Z(n8549) );
  AND2_X1 U10101 ( .A1(n8549), .A2(n8561), .ZN(n8568) );
  INV_X1 U10102 ( .A(n8568), .ZN(n8550) );
  NAND2_X1 U10103 ( .A1(n8566), .A2(n8550), .ZN(n8551) );
  XNOR2_X1 U10104 ( .A(n8567), .B(n8551), .ZN(n8552) );
  NAND2_X1 U10105 ( .A1(n8552), .A2(n8589), .ZN(n8553) );
  OAI211_X1 U10106 ( .C1(n8555), .C2(n8624), .A(n8554), .B(n8553), .ZN(
        P2_U3198) );
  AOI21_X1 U10107 ( .B1(n8824), .B2(n8557), .A(n8577), .ZN(n8575) );
  OAI21_X1 U10108 ( .B1(n8594), .B2(n8559), .A(n8558), .ZN(n8565) );
  NOR2_X1 U10109 ( .A1(n8781), .A2(n8562), .ZN(n8597) );
  AOI21_X1 U10110 ( .B1(n8562), .B2(n8781), .A(n8597), .ZN(n8563) );
  NOR2_X1 U10111 ( .A1(n8620), .A2(n8563), .ZN(n8564) );
  AOI211_X1 U10112 ( .C1(n10047), .C2(n8596), .A(n8565), .B(n8564), .ZN(n8574)
         );
  MUX2_X1 U10113 ( .A(n8781), .B(n8824), .S(n8318), .Z(n8583) );
  XNOR2_X1 U10114 ( .A(n8583), .B(n8569), .ZN(n8570) );
  OAI21_X1 U10115 ( .B1(n8571), .B2(n8570), .A(n8582), .ZN(n8572) );
  NAND2_X1 U10116 ( .A1(n8572), .A2(n8589), .ZN(n8573) );
  OAI211_X1 U10117 ( .C1(n8575), .C2(n8624), .A(n8574), .B(n8573), .ZN(
        P2_U3199) );
  NOR2_X1 U10118 ( .A1(n8596), .A2(n8576), .ZN(n8578) );
  AOI22_X1 U10119 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8613), .B1(n8618), .B2(
        n8579), .ZN(n8580) );
  AOI21_X1 U10120 ( .B1(n8581), .B2(n8580), .A(n4326), .ZN(n8606) );
  MUX2_X1 U10121 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8318), .Z(n8584) );
  INV_X1 U10122 ( .A(n8614), .ZN(n8586) );
  NAND2_X1 U10123 ( .A1(n8585), .A2(n8584), .ZN(n8612) );
  NAND2_X1 U10124 ( .A1(n8586), .A2(n8612), .ZN(n8590) );
  OAI21_X1 U10125 ( .B1(n8588), .B2(n8590), .A(n8587), .ZN(n8605) );
  INV_X1 U10126 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8593) );
  NAND3_X1 U10127 ( .A1(n8590), .A2(n8589), .A3(n8618), .ZN(n8591) );
  OAI211_X1 U10128 ( .C1(n8594), .C2(n8593), .A(n8592), .B(n8591), .ZN(n8604)
         );
  NOR2_X1 U10129 ( .A1(n8596), .A2(n8595), .ZN(n8598) );
  NAND2_X1 U10130 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8618), .ZN(n8599) );
  OAI21_X1 U10131 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8618), .A(n8599), .ZN(
        n8600) );
  NOR2_X1 U10132 ( .A1(n8602), .A2(n8620), .ZN(n8603) );
  AOI21_X1 U10133 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8618), .A(n4326), .ZN(
        n8608) );
  XNOR2_X1 U10134 ( .A(n8609), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8611) );
  INV_X1 U10135 ( .A(n8611), .ZN(n8607) );
  XNOR2_X1 U10136 ( .A(n8608), .B(n8607), .ZN(n8625) );
  XNOR2_X1 U10137 ( .A(n8609), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8619) );
  MUX2_X1 U10138 ( .A(n8611), .B(n8619), .S(n8610), .Z(n8615) );
  NAND2_X1 U10139 ( .A1(n10049), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8616) );
  OAI21_X1 U10140 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(P2_U3201) );
  INV_X1 U10141 ( .A(n8626), .ZN(n8627) );
  AOI21_X1 U10142 ( .B1(n8629), .B2(n8833), .A(n8767), .ZN(n8631) );
  AOI21_X1 U10143 ( .B1(n8767), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8631), .ZN(
        n8630) );
  OAI21_X1 U10144 ( .B1(n8835), .B2(n8698), .A(n8630), .ZN(P2_U3202) );
  AOI21_X1 U10145 ( .B1(n8767), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8631), .ZN(
        n8632) );
  OAI21_X1 U10146 ( .B1(n8838), .B2(n8698), .A(n8632), .ZN(P2_U3203) );
  MUX2_X1 U10147 ( .A(P2_REG2_REG_28__SCAN_IN), .B(n8633), .S(n8780), .Z(n8634) );
  INV_X1 U10148 ( .A(n8634), .ZN(n8638) );
  AOI22_X1 U10149 ( .A1(n8636), .A2(n8785), .B1(n8784), .B2(n8635), .ZN(n8637)
         );
  OAI211_X1 U10150 ( .C1(n8639), .C2(n8788), .A(n8638), .B(n8637), .ZN(
        P2_U3205) );
  XNOR2_X1 U10151 ( .A(n8642), .B(n8641), .ZN(n8648) );
  NAND2_X1 U10152 ( .A1(n8794), .A2(n8780), .ZN(n8652) );
  OAI22_X1 U10153 ( .A1(n8649), .A2(n8756), .B1(n8780), .B2(n9002), .ZN(n8650)
         );
  AOI21_X1 U10154 ( .B1(n8792), .B2(n8785), .A(n8650), .ZN(n8651) );
  OAI211_X1 U10155 ( .C1(n8842), .C2(n8788), .A(n8652), .B(n8651), .ZN(
        P2_U3206) );
  INV_X1 U10156 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8658) );
  XOR2_X1 U10157 ( .A(n8655), .B(n8654), .Z(n8657) );
  AOI222_X1 U10158 ( .A1(n8769), .A2(n8657), .B1(n8680), .B2(n8750), .C1(n8656), .C2(n8752), .ZN(n8843) );
  MUX2_X1 U10159 ( .A(n8658), .B(n8843), .S(n8780), .Z(n8661) );
  AOI22_X1 U10160 ( .A1(n8845), .A2(n8785), .B1(n8784), .B2(n8659), .ZN(n8660)
         );
  OAI211_X1 U10161 ( .C1(n8848), .C2(n8788), .A(n8661), .B(n8660), .ZN(
        P2_U3207) );
  OAI21_X1 U10162 ( .B1(n8663), .B2(n8670), .A(n8662), .ZN(n8666) );
  AOI222_X1 U10163 ( .A1(n8769), .A2(n8666), .B1(n8665), .B2(n8750), .C1(n8664), .C2(n8752), .ZN(n8849) );
  INV_X1 U10164 ( .A(n8682), .ZN(n8668) );
  AOI22_X1 U10165 ( .A1(n8851), .A2(n8668), .B1(n8784), .B2(n8667), .ZN(n8669)
         );
  AOI21_X1 U10166 ( .B1(n8849), .B2(n8669), .A(n8767), .ZN(n8673) );
  XNOR2_X1 U10167 ( .A(n4436), .B(n8670), .ZN(n8854) );
  OAI22_X1 U10168 ( .A1(n8854), .A2(n8788), .B1(n8671), .B2(n8780), .ZN(n8672)
         );
  OR2_X1 U10169 ( .A1(n8673), .A2(n8672), .ZN(P2_U3208) );
  NAND2_X1 U10170 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  XNOR2_X1 U10171 ( .A(n8676), .B(n8679), .ZN(n8859) );
  XNOR2_X1 U10172 ( .A(n8678), .B(n8679), .ZN(n8681) );
  AOI222_X1 U10173 ( .A1(n8769), .A2(n8681), .B1(n8680), .B2(n8752), .C1(n8707), .C2(n8750), .ZN(n8855) );
  OAI21_X1 U10174 ( .B1(n8683), .B2(n8682), .A(n8855), .ZN(n8684) );
  NAND2_X1 U10175 ( .A1(n8684), .A2(n8780), .ZN(n8687) );
  AOI22_X1 U10176 ( .A1(n8685), .A2(n8784), .B1(n8767), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8686) );
  OAI211_X1 U10177 ( .C1(n8859), .C2(n8788), .A(n8687), .B(n8686), .ZN(
        P2_U3209) );
  XOR2_X1 U10178 ( .A(n8688), .B(n8689), .Z(n8862) );
  XOR2_X1 U10179 ( .A(n8690), .B(n8689), .Z(n8691) );
  OAI222_X1 U10180 ( .A1(n8775), .A2(n8693), .B1(n8773), .B2(n8692), .C1(n8738), .C2(n8691), .ZN(n8860) );
  INV_X1 U10181 ( .A(n8860), .ZN(n8694) );
  MUX2_X1 U10182 ( .A(n8695), .B(n8694), .S(n8780), .Z(n8701) );
  INV_X1 U10183 ( .A(n8696), .ZN(n8697) );
  OAI22_X1 U10184 ( .A1(n8861), .A2(n8698), .B1(n8697), .B2(n8756), .ZN(n8699)
         );
  INV_X1 U10185 ( .A(n8699), .ZN(n8700) );
  OAI211_X1 U10186 ( .C1(n8862), .C2(n8788), .A(n8701), .B(n8700), .ZN(
        P2_U3210) );
  XOR2_X1 U10187 ( .A(n8702), .B(n8704), .Z(n8870) );
  OAI21_X1 U10188 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8708) );
  AOI222_X1 U10189 ( .A1(n8769), .A2(n8708), .B1(n8707), .B2(n8752), .C1(n8706), .C2(n8750), .ZN(n8865) );
  MUX2_X1 U10190 ( .A(n8709), .B(n8865), .S(n8780), .Z(n8712) );
  AOI22_X1 U10191 ( .A1(n8867), .A2(n8785), .B1(n8784), .B2(n8710), .ZN(n8711)
         );
  OAI211_X1 U10192 ( .C1(n8870), .C2(n8788), .A(n8712), .B(n8711), .ZN(
        P2_U3211) );
  NAND2_X1 U10193 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  XOR2_X1 U10194 ( .A(n8716), .B(n8715), .Z(n8876) );
  INV_X1 U10195 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8721) );
  XNOR2_X1 U10196 ( .A(n8717), .B(n8716), .ZN(n8720) );
  AOI222_X1 U10197 ( .A1(n8769), .A2(n8720), .B1(n8719), .B2(n8750), .C1(n8718), .C2(n8752), .ZN(n8871) );
  MUX2_X1 U10198 ( .A(n8721), .B(n8871), .S(n8780), .Z(n8724) );
  AOI22_X1 U10199 ( .A1(n8873), .A2(n8785), .B1(n8784), .B2(n8722), .ZN(n8723)
         );
  OAI211_X1 U10200 ( .C1(n8876), .C2(n8788), .A(n8724), .B(n8723), .ZN(
        P2_U3212) );
  XNOR2_X1 U10201 ( .A(n8725), .B(n8727), .ZN(n8880) );
  INV_X1 U10202 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8732) );
  AOI21_X1 U10203 ( .B1(n8727), .B2(n8726), .A(n4335), .ZN(n8728) );
  OAI222_X1 U10204 ( .A1(n8775), .A2(n8730), .B1(n8773), .B2(n8729), .C1(n8738), .C2(n8728), .ZN(n8877) );
  INV_X1 U10205 ( .A(n8877), .ZN(n8731) );
  MUX2_X1 U10206 ( .A(n8732), .B(n8731), .S(n8780), .Z(n8736) );
  AOI22_X1 U10207 ( .A1(n8734), .A2(n8785), .B1(n8784), .B2(n8733), .ZN(n8735)
         );
  OAI211_X1 U10208 ( .C1(n8880), .C2(n8788), .A(n8736), .B(n8735), .ZN(
        P2_U3213) );
  XNOR2_X1 U10209 ( .A(n8737), .B(n8742), .ZN(n8739) );
  OAI222_X1 U10210 ( .A1(n8775), .A2(n8740), .B1(n8773), .B2(n8776), .C1(n8739), .C2(n8738), .ZN(n8816) );
  OAI21_X1 U10211 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8886) );
  AOI22_X1 U10212 ( .A1(n8767), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8784), .B2(
        n8744), .ZN(n8746) );
  NAND2_X1 U10213 ( .A1(n8817), .A2(n8785), .ZN(n8745) );
  OAI211_X1 U10214 ( .C1(n8886), .C2(n8788), .A(n8746), .B(n8745), .ZN(n8747)
         );
  AOI21_X1 U10215 ( .B1(n8816), .B2(n8780), .A(n8747), .ZN(n8748) );
  INV_X1 U10216 ( .A(n8748), .ZN(P2_U3214) );
  XOR2_X1 U10217 ( .A(n8749), .B(n8763), .Z(n8754) );
  AOI222_X1 U10218 ( .A1(n8769), .A2(n8754), .B1(n8753), .B2(n8752), .C1(n8751), .C2(n8750), .ZN(n8822) );
  INV_X1 U10219 ( .A(n8755), .ZN(n8757) );
  OAI22_X1 U10220 ( .A1(n8780), .A2(n8758), .B1(n8757), .B2(n8756), .ZN(n8759)
         );
  AOI21_X1 U10221 ( .B1(n8760), .B2(n8785), .A(n8759), .ZN(n8766) );
  NAND2_X1 U10222 ( .A1(n8762), .A2(n8763), .ZN(n8820) );
  NAND3_X1 U10223 ( .A1(n8761), .A2(n8820), .A3(n8764), .ZN(n8765) );
  OAI211_X1 U10224 ( .C1(n8822), .C2(n8767), .A(n8766), .B(n8765), .ZN(
        P2_U3215) );
  XNOR2_X1 U10225 ( .A(n8768), .B(n8771), .ZN(n8895) );
  OAI211_X1 U10226 ( .C1(n8772), .C2(n8771), .A(n8770), .B(n8769), .ZN(n8779)
         );
  OAI22_X1 U10227 ( .A1(n8776), .A2(n8775), .B1(n8774), .B2(n8773), .ZN(n8777)
         );
  INV_X1 U10228 ( .A(n8777), .ZN(n8778) );
  MUX2_X1 U10229 ( .A(n8781), .B(n8888), .S(n8780), .Z(n8787) );
  INV_X1 U10230 ( .A(n8782), .ZN(n8783) );
  AOI22_X1 U10231 ( .A1(n8891), .A2(n8785), .B1(n8784), .B2(n8783), .ZN(n8786)
         );
  OAI211_X1 U10232 ( .C1(n8895), .C2(n8788), .A(n8787), .B(n8786), .ZN(
        P2_U3216) );
  NOR2_X1 U10233 ( .A1(n8833), .A2(n10133), .ZN(n8790) );
  AOI21_X1 U10234 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10133), .A(n8790), .ZN(
        n8789) );
  OAI21_X1 U10235 ( .B1(n8835), .B2(n8813), .A(n8789), .ZN(P2_U3490) );
  AOI21_X1 U10236 ( .B1(n10133), .B2(P2_REG1_REG_30__SCAN_IN), .A(n8790), .ZN(
        n8791) );
  OAI21_X1 U10237 ( .B1(n8838), .B2(n8813), .A(n8791), .ZN(P2_U3489) );
  INV_X1 U10238 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8795) );
  MUX2_X1 U10239 ( .A(n8795), .B(n8839), .S(n10135), .Z(n8796) );
  OAI21_X1 U10240 ( .B1(n8842), .B2(n8828), .A(n8796), .ZN(P2_U3486) );
  MUX2_X1 U10241 ( .A(n8972), .B(n8843), .S(n10135), .Z(n8798) );
  NAND2_X1 U10242 ( .A1(n8845), .A2(n8825), .ZN(n8797) );
  OAI211_X1 U10243 ( .C1(n8828), .C2(n8848), .A(n8798), .B(n8797), .ZN(
        P2_U3485) );
  INV_X1 U10244 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8799) );
  MUX2_X1 U10245 ( .A(n8799), .B(n8849), .S(n10135), .Z(n8801) );
  NAND2_X1 U10246 ( .A1(n8851), .A2(n8825), .ZN(n8800) );
  OAI211_X1 U10247 ( .C1(n8854), .C2(n8828), .A(n8801), .B(n8800), .ZN(
        P2_U3484) );
  INV_X1 U10248 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10249 ( .A(n8802), .B(n8855), .S(n10135), .Z(n8804) );
  NAND2_X1 U10250 ( .A1(n8856), .A2(n8825), .ZN(n8803) );
  OAI211_X1 U10251 ( .C1(n8828), .C2(n8859), .A(n8804), .B(n8803), .ZN(
        P2_U3483) );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8860), .S(n10135), .Z(
        n8806) );
  OAI22_X1 U10253 ( .A1(n8862), .A2(n8828), .B1(n8861), .B2(n8813), .ZN(n8805)
         );
  OR2_X1 U10254 ( .A1(n8806), .A2(n8805), .ZN(P2_U3482) );
  INV_X1 U10255 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8807) );
  MUX2_X1 U10256 ( .A(n8807), .B(n8865), .S(n10135), .Z(n8809) );
  NAND2_X1 U10257 ( .A1(n8867), .A2(n8825), .ZN(n8808) );
  OAI211_X1 U10258 ( .C1(n8870), .C2(n8828), .A(n8809), .B(n8808), .ZN(
        P2_U3481) );
  INV_X1 U10259 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8810) );
  MUX2_X1 U10260 ( .A(n8810), .B(n8871), .S(n10135), .Z(n8812) );
  NAND2_X1 U10261 ( .A1(n8873), .A2(n8825), .ZN(n8811) );
  OAI211_X1 U10262 ( .C1(n8828), .C2(n8876), .A(n8812), .B(n8811), .ZN(
        P2_U3480) );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8877), .S(n10135), .Z(
        n8815) );
  OAI22_X1 U10264 ( .A1(n8880), .A2(n8828), .B1(n8879), .B2(n8813), .ZN(n8814)
         );
  OR2_X1 U10265 ( .A1(n8815), .A2(n8814), .ZN(P2_U3479) );
  AOI21_X1 U10266 ( .B1(n10118), .B2(n8817), .A(n8816), .ZN(n8883) );
  MUX2_X1 U10267 ( .A(n8818), .B(n8883), .S(n10135), .Z(n8819) );
  OAI21_X1 U10268 ( .B1(n8828), .B2(n8886), .A(n8819), .ZN(P2_U3478) );
  NAND3_X1 U10269 ( .A1(n8761), .A2(n10080), .A3(n8820), .ZN(n8821) );
  OAI211_X1 U10270 ( .C1(n8823), .C2(n10108), .A(n8822), .B(n8821), .ZN(n8887)
         );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8887), .S(n10135), .Z(
        P2_U3477) );
  MUX2_X1 U10272 ( .A(n8824), .B(n8888), .S(n10135), .Z(n8827) );
  NAND2_X1 U10273 ( .A1(n8891), .A2(n8825), .ZN(n8826) );
  OAI211_X1 U10274 ( .C1(n8828), .C2(n8895), .A(n8827), .B(n8826), .ZN(
        P2_U3476) );
  AOI22_X1 U10275 ( .A1(n8830), .A2(n10080), .B1(n10118), .B2(n8829), .ZN(
        n8831) );
  NAND2_X1 U10276 ( .A1(n8832), .A2(n8831), .ZN(n8896) );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8896), .S(n10135), .Z(
        P2_U3475) );
  NOR2_X1 U10278 ( .A1(n8833), .A2(n10121), .ZN(n8836) );
  AOI21_X1 U10279 ( .B1(n10121), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8836), .ZN(
        n8834) );
  OAI21_X1 U10280 ( .B1(n8835), .B2(n8878), .A(n8834), .ZN(P2_U3458) );
  AOI21_X1 U10281 ( .B1(n10121), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8836), .ZN(
        n8837) );
  OAI21_X1 U10282 ( .B1(n8838), .B2(n8878), .A(n8837), .ZN(P2_U3457) );
  INV_X1 U10283 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U10284 ( .A(n8840), .B(n8839), .S(n10119), .Z(n8841) );
  OAI21_X1 U10285 ( .B1(n8842), .B2(n8894), .A(n8841), .ZN(P2_U3454) );
  INV_X1 U10286 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U10287 ( .A(n8844), .B(n8843), .S(n10119), .Z(n8847) );
  NAND2_X1 U10288 ( .A1(n8845), .A2(n8890), .ZN(n8846) );
  OAI211_X1 U10289 ( .C1(n8848), .C2(n8894), .A(n8847), .B(n8846), .ZN(
        P2_U3453) );
  INV_X1 U10290 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8850) );
  MUX2_X1 U10291 ( .A(n8850), .B(n8849), .S(n10119), .Z(n8853) );
  NAND2_X1 U10292 ( .A1(n8851), .A2(n8890), .ZN(n8852) );
  OAI211_X1 U10293 ( .C1(n8854), .C2(n8894), .A(n8853), .B(n8852), .ZN(
        P2_U3452) );
  MUX2_X1 U10294 ( .A(n8992), .B(n8855), .S(n10119), .Z(n8858) );
  NAND2_X1 U10295 ( .A1(n8856), .A2(n8890), .ZN(n8857) );
  OAI211_X1 U10296 ( .C1(n8859), .C2(n8894), .A(n8858), .B(n8857), .ZN(
        P2_U3451) );
  MUX2_X1 U10297 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8860), .S(n10119), .Z(
        n8864) );
  OAI22_X1 U10298 ( .A1(n8862), .A2(n8894), .B1(n8861), .B2(n8878), .ZN(n8863)
         );
  OR2_X1 U10299 ( .A1(n8864), .A2(n8863), .ZN(P2_U3450) );
  INV_X1 U10300 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U10301 ( .A(n8866), .B(n8865), .S(n10119), .Z(n8869) );
  NAND2_X1 U10302 ( .A1(n8867), .A2(n8890), .ZN(n8868) );
  OAI211_X1 U10303 ( .C1(n8870), .C2(n8894), .A(n8869), .B(n8868), .ZN(
        P2_U3449) );
  INV_X1 U10304 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8872) );
  MUX2_X1 U10305 ( .A(n8872), .B(n8871), .S(n10119), .Z(n8875) );
  NAND2_X1 U10306 ( .A1(n8873), .A2(n8890), .ZN(n8874) );
  OAI211_X1 U10307 ( .C1(n8876), .C2(n8894), .A(n8875), .B(n8874), .ZN(
        P2_U3448) );
  MUX2_X1 U10308 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8877), .S(n10119), .Z(
        n8882) );
  OAI22_X1 U10309 ( .A1(n8880), .A2(n8894), .B1(n8879), .B2(n8878), .ZN(n8881)
         );
  OR2_X1 U10310 ( .A1(n8882), .A2(n8881), .ZN(P2_U3447) );
  MUX2_X1 U10311 ( .A(n8884), .B(n8883), .S(n10119), .Z(n8885) );
  OAI21_X1 U10312 ( .B1(n8886), .B2(n8894), .A(n8885), .ZN(P2_U3446) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8887), .S(n10119), .Z(
        P2_U3444) );
  INV_X1 U10314 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U10315 ( .A(n8889), .B(n8888), .S(n10119), .Z(n8893) );
  NAND2_X1 U10316 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  OAI211_X1 U10317 ( .C1(n8895), .C2(n8894), .A(n8893), .B(n8892), .ZN(
        P2_U3441) );
  MUX2_X1 U10318 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8896), .S(n10119), .Z(
        P2_U3438) );
  NAND3_X1 U10319 ( .A1(n8898), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8901) );
  OAI22_X1 U10320 ( .A1(n8897), .A2(n8901), .B1(n8900), .B2(n8899), .ZN(n8902)
         );
  INV_X1 U10321 ( .A(n8902), .ZN(n8903) );
  OAI21_X1 U10322 ( .B1(n9796), .B2(n8907), .A(n8903), .ZN(P2_U3264) );
  MUX2_X1 U10323 ( .A(n8908), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10324 ( .A1(n8909), .A2(n9241), .ZN(n8911) );
  AOI21_X1 U10325 ( .B1(n8912), .B2(n8911), .A(n8910), .ZN(n8917) );
  AND2_X1 U10326 ( .A1(n9266), .A2(n9465), .ZN(n8913) );
  AOI21_X1 U10327 ( .B1(n9359), .B2(n9968), .A(n8913), .ZN(n9394) );
  AOI22_X1 U10328 ( .A1(n9389), .A2(n9247), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8914) );
  OAI21_X1 U10329 ( .B1(n9394), .B2(n9237), .A(n8914), .ZN(n8915) );
  AOI21_X1 U10330 ( .B1(n9736), .B2(n9260), .A(n8915), .ZN(n8916) );
  OAI21_X1 U10331 ( .B1(n8917), .B2(n9262), .A(n8916), .ZN(P1_U3214) );
  OAI21_X1 U10332 ( .B1(n8920), .B2(n8919), .A(n8918), .ZN(n8921) );
  NAND2_X1 U10333 ( .A1(n8921), .A2(n9852), .ZN(n8925) );
  AOI22_X1 U10334 ( .A1(n9465), .A2(n9276), .B1(n9274), .B2(n9498), .ZN(n9612)
         );
  OAI22_X1 U10335 ( .A1(n9612), .A2(n9237), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8922), .ZN(n8923) );
  AOI21_X1 U10336 ( .B1(n9620), .B2(n9247), .A(n8923), .ZN(n8924) );
  OAI211_X1 U10337 ( .C1(n9623), .C2(n9849), .A(n8925), .B(n8924), .ZN(
        P1_U3215) );
  INV_X1 U10338 ( .A(n8926), .ZN(n8931) );
  AOI21_X1 U10339 ( .B1(n8928), .B2(n8930), .A(n8927), .ZN(n8929) );
  AOI21_X1 U10340 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n8936) );
  OAI22_X1 U10341 ( .A1(n9425), .A2(n9210), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8932), .ZN(n8934) );
  OAI22_X1 U10342 ( .A1(n9118), .A2(n9209), .B1(n9856), .B2(n9457), .ZN(n8933)
         );
  AOI211_X1 U10343 ( .C1(n9680), .C2(n9260), .A(n8934), .B(n8933), .ZN(n8935)
         );
  OAI21_X1 U10344 ( .B1(n8936), .B2(n9262), .A(n8935), .ZN(P1_U3216) );
  NAND2_X1 U10345 ( .A1(keyinput13), .A2(keyinput33), .ZN(n8937) );
  NOR3_X1 U10346 ( .A1(keyinput38), .A2(keyinput46), .A3(n8937), .ZN(n8942) );
  NOR3_X1 U10347 ( .A1(keyinput23), .A2(keyinput60), .A3(keyinput58), .ZN(
        n8941) );
  NAND3_X1 U10348 ( .A1(keyinput47), .A2(keyinput61), .A3(keyinput30), .ZN(
        n8939) );
  NAND3_X1 U10349 ( .A1(keyinput12), .A2(keyinput55), .A3(keyinput32), .ZN(
        n8938) );
  NOR4_X1 U10350 ( .A1(keyinput22), .A2(keyinput2), .A3(n8939), .A4(n8938), 
        .ZN(n8940) );
  NAND4_X1 U10351 ( .A1(n8942), .A2(keyinput11), .A3(n8941), .A4(n8940), .ZN(
        n8957) );
  NOR4_X1 U10352 ( .A1(keyinput37), .A2(keyinput45), .A3(keyinput5), .A4(
        keyinput20), .ZN(n8944) );
  NOR2_X1 U10353 ( .A1(keyinput29), .A2(keyinput10), .ZN(n8943) );
  NAND4_X1 U10354 ( .A1(n8944), .A2(keyinput6), .A3(keyinput43), .A4(n8943), 
        .ZN(n8956) );
  NOR3_X1 U10355 ( .A1(keyinput15), .A2(keyinput18), .A3(keyinput0), .ZN(n8947) );
  INV_X1 U10356 ( .A(keyinput26), .ZN(n8945) );
  NOR3_X1 U10357 ( .A1(keyinput19), .A2(keyinput4), .A3(n8945), .ZN(n8946) );
  NAND4_X1 U10358 ( .A1(keyinput51), .A2(n8947), .A3(keyinput63), .A4(n8946), 
        .ZN(n8955) );
  NOR3_X1 U10359 ( .A1(keyinput36), .A2(keyinput39), .A3(keyinput40), .ZN(
        n8949) );
  NOR3_X1 U10360 ( .A1(keyinput44), .A2(keyinput7), .A3(keyinput16), .ZN(n8948) );
  NAND4_X1 U10361 ( .A1(keyinput34), .A2(n8949), .A3(keyinput1), .A4(n8948), 
        .ZN(n8953) );
  NOR2_X1 U10362 ( .A1(keyinput14), .A2(keyinput31), .ZN(n8950) );
  NAND3_X1 U10363 ( .A1(keyinput25), .A2(keyinput53), .A3(n8950), .ZN(n8952)
         );
  NAND3_X1 U10364 ( .A1(keyinput56), .A2(keyinput41), .A3(keyinput28), .ZN(
        n8951) );
  OR4_X1 U10365 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(keyinput21), .ZN(
        n8954) );
  NOR4_X1 U10366 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n9057)
         );
  NOR2_X1 U10367 ( .A1(keyinput59), .A2(keyinput49), .ZN(n8964) );
  NAND2_X1 U10368 ( .A1(keyinput48), .A2(keyinput9), .ZN(n8962) );
  NOR3_X1 U10369 ( .A1(keyinput57), .A2(keyinput35), .A3(keyinput62), .ZN(
        n8960) );
  INV_X1 U10370 ( .A(keyinput8), .ZN(n8958) );
  NOR3_X1 U10371 ( .A1(keyinput42), .A2(keyinput50), .A3(n8958), .ZN(n8959) );
  NAND4_X1 U10372 ( .A1(keyinput54), .A2(n8960), .A3(keyinput17), .A4(n8959), 
        .ZN(n8961) );
  NOR4_X1 U10373 ( .A1(keyinput3), .A2(keyinput24), .A3(n8962), .A4(n8961), 
        .ZN(n8963) );
  AND4_X1 U10374 ( .A1(keyinput27), .A2(keyinput52), .A3(n8964), .A4(n8963), 
        .ZN(n9056) );
  INV_X1 U10375 ( .A(keyinput36), .ZN(n8966) );
  AOI22_X1 U10376 ( .A1(n8967), .A2(keyinput34), .B1(P2_ADDR_REG_9__SCAN_IN), 
        .B2(n8966), .ZN(n8965) );
  OAI221_X1 U10377 ( .B1(n8967), .B2(keyinput34), .C1(n8966), .C2(
        P2_ADDR_REG_9__SCAN_IN), .A(n8965), .ZN(n8979) );
  INV_X1 U10378 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9990) );
  INV_X1 U10379 ( .A(keyinput40), .ZN(n8969) );
  AOI22_X1 U10380 ( .A1(n9990), .A2(keyinput39), .B1(P2_ADDR_REG_11__SCAN_IN), 
        .B2(n8969), .ZN(n8968) );
  OAI221_X1 U10381 ( .B1(n9990), .B2(keyinput39), .C1(n8969), .C2(
        P2_ADDR_REG_11__SCAN_IN), .A(n8968), .ZN(n8978) );
  INV_X1 U10382 ( .A(keyinput14), .ZN(n8971) );
  AOI22_X1 U10383 ( .A1(n8972), .A2(keyinput31), .B1(P2_ADDR_REG_12__SCAN_IN), 
        .B2(n8971), .ZN(n8970) );
  OAI221_X1 U10384 ( .B1(n8972), .B2(keyinput31), .C1(n8971), .C2(
        P2_ADDR_REG_12__SCAN_IN), .A(n8970), .ZN(n8977) );
  INV_X1 U10385 ( .A(keyinput37), .ZN(n8974) );
  AOI22_X1 U10386 ( .A1(n8975), .A2(keyinput45), .B1(P2_WR_REG_SCAN_IN), .B2(
        n8974), .ZN(n8973) );
  OAI221_X1 U10387 ( .B1(n8975), .B2(keyinput45), .C1(n8974), .C2(
        P2_WR_REG_SCAN_IN), .A(n8973), .ZN(n8976) );
  OR4_X1 U10388 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(n8987)
         );
  INV_X1 U10389 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8982) );
  INV_X1 U10390 ( .A(SI_15_), .ZN(n8981) );
  AOI22_X1 U10391 ( .A1(n8982), .A2(keyinput30), .B1(n8981), .B2(keyinput22), 
        .ZN(n8980) );
  OAI221_X1 U10392 ( .B1(n8982), .B2(keyinput30), .C1(n8981), .C2(keyinput22), 
        .A(n8980), .ZN(n8986) );
  AOI22_X1 U10393 ( .A1(n9208), .A2(keyinput21), .B1(n5168), .B2(keyinput56), 
        .ZN(n8983) );
  OAI221_X1 U10394 ( .B1(n9208), .B2(keyinput21), .C1(n5168), .C2(keyinput56), 
        .A(n8983), .ZN(n8985) );
  INV_X1 U10395 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9989) );
  XNOR2_X1 U10396 ( .A(n9989), .B(keyinput53), .ZN(n8984) );
  NOR4_X1 U10397 ( .A1(n8987), .A2(n8986), .A3(n8985), .A4(n8984), .ZN(n9054)
         );
  INV_X1 U10398 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8989) );
  AOI22_X1 U10399 ( .A1(n8989), .A2(keyinput27), .B1(n5624), .B2(keyinput59), 
        .ZN(n8988) );
  OAI221_X1 U10400 ( .B1(n8989), .B2(keyinput27), .C1(n5624), .C2(keyinput59), 
        .A(n8988), .ZN(n8996) );
  AOI22_X1 U10401 ( .A1(n8992), .A2(keyinput7), .B1(n8991), .B2(keyinput16), 
        .ZN(n8990) );
  OAI221_X1 U10402 ( .B1(n8992), .B2(keyinput7), .C1(n8991), .C2(keyinput16), 
        .A(n8990), .ZN(n8995) );
  INV_X1 U10403 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10031) );
  XNOR2_X1 U10404 ( .A(keyinput32), .B(n10031), .ZN(n8994) );
  XNOR2_X1 U10405 ( .A(keyinput3), .B(n5054), .ZN(n8993) );
  NOR4_X1 U10406 ( .A1(n8996), .A2(n8995), .A3(n8994), .A4(n8993), .ZN(n9053)
         );
  AOI22_X1 U10407 ( .A1(n8999), .A2(keyinput57), .B1(n8998), .B2(keyinput35), 
        .ZN(n8997) );
  OAI221_X1 U10408 ( .B1(n8999), .B2(keyinput57), .C1(n8998), .C2(keyinput35), 
        .A(n8997), .ZN(n9012) );
  AOI22_X1 U10409 ( .A1(n9002), .A2(keyinput42), .B1(n9001), .B2(keyinput17), 
        .ZN(n9000) );
  OAI221_X1 U10410 ( .B1(n9002), .B2(keyinput42), .C1(n9001), .C2(keyinput17), 
        .A(n9000), .ZN(n9011) );
  AOI22_X1 U10411 ( .A1(n9005), .A2(keyinput47), .B1(n9004), .B2(keyinput61), 
        .ZN(n9003) );
  OAI221_X1 U10412 ( .B1(n9005), .B2(keyinput47), .C1(n9004), .C2(keyinput61), 
        .A(n9003), .ZN(n9010) );
  AOI22_X1 U10413 ( .A1(n9008), .A2(keyinput51), .B1(n9007), .B2(keyinput0), 
        .ZN(n9006) );
  OAI221_X1 U10414 ( .B1(n9008), .B2(keyinput51), .C1(n9007), .C2(keyinput0), 
        .A(n9006), .ZN(n9009) );
  NOR4_X1 U10415 ( .A1(n9012), .A2(n9011), .A3(n9010), .A4(n9009), .ZN(n9052)
         );
  XNOR2_X1 U10416 ( .A(n5630), .B(keyinput28), .ZN(n9018) );
  XNOR2_X1 U10417 ( .A(n9013), .B(keyinput48), .ZN(n9017) );
  XNOR2_X1 U10418 ( .A(n9014), .B(keyinput25), .ZN(n9016) );
  XNOR2_X1 U10419 ( .A(n9180), .B(keyinput8), .ZN(n9015) );
  NOR4_X1 U10420 ( .A1(n9018), .A2(n9017), .A3(n9016), .A4(n9015), .ZN(n9041)
         );
  XNOR2_X1 U10421 ( .A(n9019), .B(keyinput62), .ZN(n9026) );
  XNOR2_X1 U10422 ( .A(n9020), .B(keyinput24), .ZN(n9025) );
  XNOR2_X1 U10423 ( .A(n9021), .B(keyinput41), .ZN(n9024) );
  XNOR2_X1 U10424 ( .A(n9022), .B(keyinput9), .ZN(n9023) );
  NOR4_X1 U10425 ( .A1(n9026), .A2(n9025), .A3(n9024), .A4(n9023), .ZN(n9040)
         );
  XOR2_X1 U10426 ( .A(SI_16_), .B(keyinput18), .Z(n9032) );
  XOR2_X1 U10427 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput15), .Z(n9031) );
  XNOR2_X1 U10428 ( .A(n9027), .B(keyinput50), .ZN(n9030) );
  XNOR2_X1 U10429 ( .A(n9028), .B(keyinput54), .ZN(n9029) );
  NOR4_X1 U10430 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(n9039)
         );
  XOR2_X1 U10431 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput2), .Z(n9037) );
  XOR2_X1 U10432 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput55), .Z(n9036) );
  XNOR2_X1 U10433 ( .A(n9033), .B(keyinput5), .ZN(n9035) );
  INV_X1 U10434 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10075) );
  XNOR2_X1 U10435 ( .A(keyinput20), .B(n10075), .ZN(n9034) );
  NOR4_X1 U10436 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n9038)
         );
  NAND4_X1 U10437 ( .A1(n9041), .A2(n9040), .A3(n9039), .A4(n9038), .ZN(n9050)
         );
  AOI22_X1 U10438 ( .A1(n6353), .A2(keyinput49), .B1(n4569), .B2(keyinput52), 
        .ZN(n9042) );
  OAI221_X1 U10439 ( .B1(n6353), .B2(keyinput49), .C1(n4569), .C2(keyinput52), 
        .A(n9042), .ZN(n9049) );
  INV_X1 U10440 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9045) );
  AOI22_X1 U10441 ( .A1(n9045), .A2(keyinput1), .B1(keyinput44), .B2(n9044), 
        .ZN(n9043) );
  OAI221_X1 U10442 ( .B1(n9045), .B2(keyinput1), .C1(n9044), .C2(keyinput44), 
        .A(n9043), .ZN(n9048) );
  INV_X1 U10443 ( .A(keyinput12), .ZN(n9046) );
  XNOR2_X1 U10444 ( .A(n9046), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(n9047) );
  NOR4_X1 U10445 ( .A1(n9050), .A2(n9049), .A3(n9048), .A4(n9047), .ZN(n9051)
         );
  NAND4_X1 U10446 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n9055)
         );
  AOI21_X1 U10447 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9085) );
  AOI22_X1 U10448 ( .A1(n9060), .A2(keyinput13), .B1(keyinput33), .B2(n9059), 
        .ZN(n9058) );
  OAI221_X1 U10449 ( .B1(n9060), .B2(keyinput13), .C1(n9059), .C2(keyinput33), 
        .A(n9058), .ZN(n9070) );
  INV_X1 U10450 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U10451 ( .A1(n9988), .A2(keyinput38), .B1(n6780), .B2(keyinput46), 
        .ZN(n9061) );
  OAI221_X1 U10452 ( .B1(n9988), .B2(keyinput38), .C1(n6780), .C2(keyinput46), 
        .A(n9061), .ZN(n9069) );
  INV_X1 U10453 ( .A(keyinput60), .ZN(n9063) );
  AOI22_X1 U10454 ( .A1(n9064), .A2(keyinput23), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n9063), .ZN(n9062) );
  OAI221_X1 U10455 ( .B1(n9064), .B2(keyinput23), .C1(n9063), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n9062), .ZN(n9068) );
  INV_X1 U10456 ( .A(SI_30_), .ZN(n9066) );
  AOI22_X1 U10457 ( .A1(n9677), .A2(keyinput58), .B1(keyinput11), .B2(n9066), 
        .ZN(n9065) );
  OAI221_X1 U10458 ( .B1(n9677), .B2(keyinput58), .C1(n9066), .C2(keyinput11), 
        .A(n9065), .ZN(n9067) );
  NOR4_X1 U10459 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n9084)
         );
  INV_X1 U10460 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9645) );
  INV_X1 U10461 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U10462 ( .A1(n9645), .A2(keyinput6), .B1(n9991), .B2(keyinput29), 
        .ZN(n9071) );
  OAI221_X1 U10463 ( .B1(n9645), .B2(keyinput6), .C1(n9991), .C2(keyinput29), 
        .A(n9071), .ZN(n9082) );
  AOI22_X1 U10464 ( .A1(n5620), .A2(keyinput10), .B1(n9073), .B2(keyinput43), 
        .ZN(n9072) );
  OAI221_X1 U10465 ( .B1(n5620), .B2(keyinput10), .C1(n9073), .C2(keyinput43), 
        .A(n9072), .ZN(n9081) );
  AOI22_X1 U10466 ( .A1(n9075), .A2(keyinput63), .B1(keyinput19), .B2(n5081), 
        .ZN(n9074) );
  OAI221_X1 U10467 ( .B1(n9075), .B2(keyinput63), .C1(n5081), .C2(keyinput19), 
        .A(n9074), .ZN(n9080) );
  INV_X1 U10468 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9078) );
  AOI22_X1 U10469 ( .A1(n9078), .A2(keyinput4), .B1(n9077), .B2(keyinput26), 
        .ZN(n9076) );
  OAI221_X1 U10470 ( .B1(n9078), .B2(keyinput4), .C1(n9077), .C2(keyinput26), 
        .A(n9076), .ZN(n9079) );
  NOR4_X1 U10471 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n9083)
         );
  NAND3_X1 U10472 ( .A1(n9085), .A2(n9084), .A3(n9083), .ZN(n9102) );
  INV_X1 U10473 ( .A(n9533), .ZN(n9089) );
  NAND2_X1 U10474 ( .A1(n9271), .A2(n9465), .ZN(n9087) );
  NAND2_X1 U10475 ( .A1(n9269), .A2(n9968), .ZN(n9086) );
  NAND2_X1 U10476 ( .A1(n9087), .A2(n9086), .ZN(n9531) );
  AOI22_X1 U10477 ( .A1(n9847), .A2(n9531), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9088) );
  OAI21_X1 U10478 ( .B1(n9856), .B2(n9089), .A(n9088), .ZN(n9100) );
  NAND2_X1 U10479 ( .A1(n9231), .A2(n9232), .ZN(n9230) );
  XNOR2_X1 U10480 ( .A(n9092), .B(n9091), .ZN(n9095) );
  NAND2_X1 U10481 ( .A1(n9094), .A2(n9093), .ZN(n9096) );
  NAND3_X1 U10482 ( .A1(n9230), .A2(n9095), .A3(n9096), .ZN(n9187) );
  INV_X1 U10483 ( .A(n9187), .ZN(n9098) );
  AOI21_X1 U10484 ( .B1(n9230), .B2(n9096), .A(n9095), .ZN(n9097) );
  NOR3_X1 U10485 ( .A1(n9098), .A2(n9097), .A3(n9262), .ZN(n9099) );
  XOR2_X1 U10486 ( .A(n9102), .B(n9101), .Z(P1_U3219) );
  OAI21_X1 U10487 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9106) );
  NAND2_X1 U10488 ( .A1(n9106), .A2(n9852), .ZN(n9110) );
  AOI22_X1 U10489 ( .A1(n9260), .A2(n6085), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9107), .ZN(n9109) );
  AOI22_X1 U10490 ( .A1(n9246), .A2(n9288), .B1(n9244), .B2(n9286), .ZN(n9108)
         );
  NAND3_X1 U10491 ( .A1(n9110), .A2(n9109), .A3(n9108), .ZN(P1_U3222) );
  INV_X1 U10492 ( .A(n9114), .ZN(n9112) );
  NOR2_X1 U10493 ( .A1(n9112), .A2(n9111), .ZN(n9185) );
  NAND3_X1 U10494 ( .A1(n9187), .A2(n9185), .A3(n9186), .ZN(n9184) );
  NAND3_X1 U10495 ( .A1(n9184), .A2(n9114), .A3(n9113), .ZN(n9115) );
  AND2_X1 U10496 ( .A1(n9116), .A2(n9115), .ZN(n9122) );
  OAI22_X1 U10497 ( .A1(n9118), .A2(n9210), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9117), .ZN(n9120) );
  OAI22_X1 U10498 ( .A1(n9501), .A2(n9209), .B1(n9856), .B2(n9505), .ZN(n9119)
         );
  AOI211_X1 U10499 ( .C1(n9757), .C2(n9260), .A(n9120), .B(n9119), .ZN(n9121)
         );
  OAI21_X1 U10500 ( .B1(n9122), .B2(n9262), .A(n9121), .ZN(P1_U3223) );
  XOR2_X1 U10501 ( .A(n9123), .B(n9124), .Z(n9132) );
  INV_X1 U10502 ( .A(n9125), .ZN(n9128) );
  AOI22_X1 U10503 ( .A1(n9847), .A2(n9126), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3086), .ZN(n9127) );
  OAI21_X1 U10504 ( .B1(n9856), .B2(n9128), .A(n9127), .ZN(n9129) );
  AOI21_X1 U10505 ( .B1(n9130), .B2(n9260), .A(n9129), .ZN(n9131) );
  OAI21_X1 U10506 ( .B1(n9132), .B2(n9262), .A(n9131), .ZN(P1_U3224) );
  XOR2_X1 U10507 ( .A(n9134), .B(n9133), .Z(n9139) );
  AOI22_X1 U10508 ( .A1(n9266), .A2(n9244), .B1(n9429), .B2(n9247), .ZN(n9136)
         );
  AOI22_X1 U10509 ( .A1(n9466), .A2(n9246), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9135) );
  NAND2_X1 U10510 ( .A1(n9136), .A2(n9135), .ZN(n9137) );
  AOI21_X1 U10511 ( .B1(n9671), .B2(n9260), .A(n9137), .ZN(n9138) );
  OAI21_X1 U10512 ( .B1(n9139), .B2(n9262), .A(n9138), .ZN(P1_U3225) );
  OAI21_X1 U10513 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n9147) );
  XNOR2_X1 U10514 ( .A(n9144), .B(n9145), .ZN(n9254) );
  NOR2_X1 U10515 ( .A1(n9254), .A2(n9253), .ZN(n9252) );
  AOI21_X1 U10516 ( .B1(n9145), .B2(n9144), .A(n9252), .ZN(n9146) );
  XOR2_X1 U10517 ( .A(n9147), .B(n9146), .Z(n9154) );
  NAND2_X1 U10518 ( .A1(n9274), .A2(n9465), .ZN(n9149) );
  NAND2_X1 U10519 ( .A1(n9272), .A2(n9498), .ZN(n9148) );
  AND2_X1 U10520 ( .A1(n9149), .A2(n9148), .ZN(n9579) );
  OAI22_X1 U10521 ( .A1(n9579), .A2(n9237), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9150), .ZN(n9151) );
  AOI21_X1 U10522 ( .B1(n9584), .B2(n9247), .A(n9151), .ZN(n9153) );
  NAND2_X1 U10523 ( .A1(n9583), .A2(n9260), .ZN(n9152) );
  OAI211_X1 U10524 ( .C1(n9154), .C2(n9262), .A(n9153), .B(n9152), .ZN(
        P1_U3226) );
  OAI21_X1 U10525 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9158) );
  NAND2_X1 U10526 ( .A1(n9158), .A2(n9852), .ZN(n9164) );
  AOI22_X1 U10527 ( .A1(n9246), .A2(n9284), .B1(n9244), .B2(n9282), .ZN(n9163)
         );
  AOI22_X1 U10528 ( .A1(n9260), .A2(n9159), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n9162) );
  NAND2_X1 U10529 ( .A1(n9247), .A2(n9160), .ZN(n9161) );
  NAND4_X1 U10530 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(
        P1_U3227) );
  OAI21_X1 U10531 ( .B1(n9167), .B2(n9165), .A(n9166), .ZN(n9168) );
  NAND2_X1 U10532 ( .A1(n9168), .A2(n9852), .ZN(n9173) );
  NAND2_X1 U10533 ( .A1(n9271), .A2(n9498), .ZN(n9170) );
  NAND2_X1 U10534 ( .A1(n9273), .A2(n9465), .ZN(n9169) );
  AND2_X1 U10535 ( .A1(n9170), .A2(n9169), .ZN(n9562) );
  NAND2_X1 U10536 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9947) );
  OAI21_X1 U10537 ( .B1(n9562), .B2(n9237), .A(n9947), .ZN(n9171) );
  AOI21_X1 U10538 ( .B1(n9568), .B2(n9247), .A(n9171), .ZN(n9172) );
  OAI211_X1 U10539 ( .C1(n9570), .C2(n9849), .A(n9173), .B(n9172), .ZN(
        P1_U3228) );
  OAI21_X1 U10540 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9177) );
  NAND2_X1 U10541 ( .A1(n9177), .A2(n9852), .ZN(n9183) );
  INV_X1 U10542 ( .A(n9178), .ZN(n9447) );
  AND2_X1 U10543 ( .A1(n9475), .A2(n9465), .ZN(n9179) );
  AOI21_X1 U10544 ( .B1(n9267), .B2(n9968), .A(n9179), .ZN(n9441) );
  OAI22_X1 U10545 ( .A1(n9441), .A2(n9237), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9180), .ZN(n9181) );
  AOI21_X1 U10546 ( .B1(n9447), .B2(n9247), .A(n9181), .ZN(n9182) );
  OAI211_X1 U10547 ( .C1(n9450), .C2(n9849), .A(n9183), .B(n9182), .ZN(
        P1_U3229) );
  INV_X1 U10548 ( .A(n9521), .ZN(n9763) );
  INV_X1 U10549 ( .A(n9184), .ZN(n9189) );
  AOI21_X1 U10550 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9188) );
  OAI21_X1 U10551 ( .B1(n9189), .B2(n9188), .A(n9852), .ZN(n9193) );
  AOI22_X1 U10552 ( .A1(n9268), .A2(n9968), .B1(n9270), .B2(n9465), .ZN(n9518)
         );
  OAI22_X1 U10553 ( .A1(n9518), .A2(n9237), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9190), .ZN(n9191) );
  AOI21_X1 U10554 ( .B1(n9522), .B2(n9247), .A(n9191), .ZN(n9192) );
  OAI211_X1 U10555 ( .C1(n9763), .C2(n9849), .A(n9193), .B(n9192), .ZN(
        P1_U3233) );
  NAND2_X1 U10556 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  XOR2_X1 U10557 ( .A(n9197), .B(n9196), .Z(n9204) );
  AOI22_X1 U10558 ( .A1(n9847), .A2(n9198), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9199) );
  OAI21_X1 U10559 ( .B1(n9856), .B2(n9200), .A(n9199), .ZN(n9201) );
  AOI21_X1 U10560 ( .B1(n9202), .B2(n9260), .A(n9201), .ZN(n9203) );
  OAI21_X1 U10561 ( .B1(n9204), .B2(n9262), .A(n9203), .ZN(P1_U3234) );
  NOR2_X1 U10562 ( .A1(n9205), .A2(n4325), .ZN(n9207) );
  XNOR2_X1 U10563 ( .A(n9207), .B(n9206), .ZN(n9215) );
  OAI22_X1 U10564 ( .A1(n9209), .A2(n9477), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9208), .ZN(n9213) );
  OAI22_X1 U10565 ( .A1(n9211), .A2(n9210), .B1(n9856), .B2(n9482), .ZN(n9212)
         );
  AOI211_X1 U10566 ( .C1(n9752), .C2(n9260), .A(n9213), .B(n9212), .ZN(n9214)
         );
  OAI21_X1 U10567 ( .B1(n9215), .B2(n9262), .A(n9214), .ZN(P1_U3235) );
  INV_X1 U10568 ( .A(n9219), .ZN(n9216) );
  NOR2_X1 U10569 ( .A1(n9217), .A2(n9216), .ZN(n9222) );
  AOI21_X1 U10570 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9221) );
  OAI21_X1 U10571 ( .B1(n9222), .B2(n9221), .A(n9852), .ZN(n9229) );
  AOI22_X1 U10572 ( .A1(n9847), .A2(n9223), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9228) );
  NAND2_X1 U10573 ( .A1(n9224), .A2(n9260), .ZN(n9227) );
  NAND2_X1 U10574 ( .A1(n9247), .A2(n9225), .ZN(n9226) );
  NAND4_X1 U10575 ( .A1(n9229), .A2(n9228), .A3(n9227), .A4(n9226), .ZN(
        P1_U3236) );
  OAI21_X1 U10576 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9233) );
  NAND2_X1 U10577 ( .A1(n9233), .A2(n9852), .ZN(n9240) );
  NAND2_X1 U10578 ( .A1(n9272), .A2(n9465), .ZN(n9235) );
  NAND2_X1 U10579 ( .A1(n9270), .A2(n9498), .ZN(n9234) );
  AND2_X1 U10580 ( .A1(n9235), .A2(n9234), .ZN(n9549) );
  OAI21_X1 U10581 ( .B1(n9549), .B2(n9237), .A(n9236), .ZN(n9238) );
  AOI21_X1 U10582 ( .B1(n9553), .B2(n9247), .A(n9238), .ZN(n9239) );
  OAI211_X1 U10583 ( .C1(n9556), .C2(n9849), .A(n9240), .B(n9239), .ZN(
        P1_U3238) );
  OAI211_X1 U10584 ( .C1(n9243), .C2(n9242), .A(n9241), .B(n9852), .ZN(n9251)
         );
  AOI22_X1 U10585 ( .A1(n9408), .A2(n9244), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9250) );
  INV_X1 U10586 ( .A(n9245), .ZN(n9402) );
  AOI22_X1 U10587 ( .A1(n9402), .A2(n9247), .B1(n9267), .B2(n9246), .ZN(n9249)
         );
  NAND2_X1 U10588 ( .A1(n9741), .A2(n9260), .ZN(n9248) );
  NAND4_X1 U10589 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(
        P1_U3240) );
  AOI21_X1 U10590 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9263) );
  INV_X1 U10591 ( .A(n9599), .ZN(n9258) );
  NAND2_X1 U10592 ( .A1(n9275), .A2(n9465), .ZN(n9256) );
  NAND2_X1 U10593 ( .A1(n9273), .A2(n9498), .ZN(n9255) );
  NAND2_X1 U10594 ( .A1(n9256), .A2(n9255), .ZN(n9594) );
  AOI22_X1 U10595 ( .A1(n9847), .A2(n9594), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9257) );
  OAI21_X1 U10596 ( .B1(n9856), .B2(n9258), .A(n9257), .ZN(n9259) );
  AOI21_X1 U10597 ( .B1(n9784), .B2(n9260), .A(n9259), .ZN(n9261) );
  OAI21_X1 U10598 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(P1_U3241) );
  MUX2_X1 U10599 ( .A(n9264), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9287), .Z(
        P1_U3585) );
  MUX2_X1 U10600 ( .A(n9265), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9287), .Z(
        P1_U3583) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9359), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10602 ( .A(n9408), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9287), .Z(
        P1_U3581) );
  MUX2_X1 U10603 ( .A(n9266), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9287), .Z(
        P1_U3580) );
  MUX2_X1 U10604 ( .A(n9267), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9287), .Z(
        P1_U3579) );
  MUX2_X1 U10605 ( .A(n9466), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9287), .Z(
        P1_U3578) );
  MUX2_X1 U10606 ( .A(n9475), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9287), .Z(
        P1_U3577) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9499), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10608 ( .A(n9268), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9287), .Z(
        P1_U3575) );
  MUX2_X1 U10609 ( .A(n9269), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9287), .Z(
        P1_U3574) );
  MUX2_X1 U10610 ( .A(n9270), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9287), .Z(
        P1_U3573) );
  MUX2_X1 U10611 ( .A(n9271), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9287), .Z(
        P1_U3572) );
  MUX2_X1 U10612 ( .A(n9272), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9287), .Z(
        P1_U3571) );
  MUX2_X1 U10613 ( .A(n9273), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9287), .Z(
        P1_U3570) );
  MUX2_X1 U10614 ( .A(n9274), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9287), .Z(
        P1_U3569) );
  MUX2_X1 U10615 ( .A(n9275), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9287), .Z(
        P1_U3568) );
  MUX2_X1 U10616 ( .A(n9276), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9287), .Z(
        P1_U3567) );
  MUX2_X1 U10617 ( .A(n9277), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9287), .Z(
        P1_U3566) );
  MUX2_X1 U10618 ( .A(n9278), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9287), .Z(
        P1_U3565) );
  MUX2_X1 U10619 ( .A(n9969), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9287), .Z(
        P1_U3564) );
  MUX2_X1 U10620 ( .A(n9279), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9287), .Z(
        P1_U3563) );
  MUX2_X1 U10621 ( .A(n9280), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9287), .Z(
        P1_U3562) );
  MUX2_X1 U10622 ( .A(n9281), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9287), .Z(
        P1_U3561) );
  MUX2_X1 U10623 ( .A(n9282), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9287), .Z(
        P1_U3560) );
  MUX2_X1 U10624 ( .A(n9283), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9287), .Z(
        P1_U3559) );
  MUX2_X1 U10625 ( .A(n9284), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9287), .Z(
        P1_U3558) );
  MUX2_X1 U10626 ( .A(n9285), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9287), .Z(
        P1_U3557) );
  MUX2_X1 U10627 ( .A(n9286), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9287), .Z(
        P1_U3556) );
  MUX2_X1 U10628 ( .A(n6084), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9287), .Z(
        P1_U3555) );
  MUX2_X1 U10629 ( .A(n9288), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9287), .Z(
        P1_U3554) );
  INV_X1 U10630 ( .A(n9289), .ZN(n9293) );
  OAI22_X1 U10631 ( .A1(n9950), .A2(n9291), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9290), .ZN(n9292) );
  AOI21_X1 U10632 ( .B1(n9293), .B2(n9943), .A(n9292), .ZN(n9302) );
  OAI211_X1 U10633 ( .C1(n9296), .C2(n9295), .A(n9941), .B(n9294), .ZN(n9301)
         );
  OAI211_X1 U10634 ( .C1(n9299), .C2(n9298), .A(n9945), .B(n9297), .ZN(n9300)
         );
  NAND3_X1 U10635 ( .A1(n9302), .A2(n9301), .A3(n9300), .ZN(P1_U3244) );
  MUX2_X1 U10636 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6465), .S(n9313), .Z(n9305)
         );
  NAND3_X1 U10637 ( .A1(n9305), .A2(n9304), .A3(n9303), .ZN(n9306) );
  NAND3_X1 U10638 ( .A1(n9945), .A2(n9307), .A3(n9306), .ZN(n9318) );
  AOI22_X1 U10639 ( .A1(n9924), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n9317) );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6445), .S(n9313), .Z(n9310)
         );
  NAND3_X1 U10641 ( .A1(n9310), .A2(n9309), .A3(n9308), .ZN(n9311) );
  NAND3_X1 U10642 ( .A1(n9941), .A2(n9312), .A3(n9311), .ZN(n9316) );
  INV_X1 U10643 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U10644 ( .A1(n9943), .A2(n9314), .ZN(n9315) );
  NAND4_X1 U10645 ( .A1(n9318), .A2(n9317), .A3(n9316), .A4(n9315), .ZN(
        P1_U3246) );
  NAND2_X1 U10646 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  XNOR2_X1 U10647 ( .A(n9321), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U10648 ( .A1(n9322), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U10649 ( .A1(n9324), .A2(n9323), .ZN(n9325) );
  XNOR2_X1 U10650 ( .A(n9325), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9327) );
  OAI22_X1 U10651 ( .A1(n9326), .A2(n9827), .B1(n9327), .B2(n9832), .ZN(n9332)
         );
  INV_X1 U10652 ( .A(n9326), .ZN(n9329) );
  AOI21_X1 U10653 ( .B1(n9327), .B2(n9941), .A(n9943), .ZN(n9328) );
  OAI21_X1 U10654 ( .B1(n9329), .B2(n9827), .A(n9328), .ZN(n9331) );
  MUX2_X1 U10655 ( .A(n9332), .B(n9331), .S(n9330), .Z(n9333) );
  INV_X1 U10656 ( .A(n9333), .ZN(n9335) );
  NAND2_X1 U10657 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9334) );
  OAI211_X1 U10658 ( .C1(n4498), .C2(n9950), .A(n9335), .B(n9334), .ZN(
        P1_U3262) );
  NAND2_X1 U10659 ( .A1(n9336), .A2(n9637), .ZN(n9339) );
  INV_X1 U10660 ( .A(n9337), .ZN(n9643) );
  NOR2_X1 U10661 ( .A1(n9643), .A2(n9987), .ZN(n9343) );
  AOI21_X1 U10662 ( .B1(n9987), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9343), .ZN(
        n9338) );
  OAI211_X1 U10663 ( .C1(n9622), .C2(n9340), .A(n9339), .B(n9338), .ZN(
        P1_U3263) );
  OAI211_X1 U10664 ( .C1(n9732), .C2(n9361), .A(n9966), .B(n9341), .ZN(n9644)
         );
  NOR2_X1 U10665 ( .A1(n9732), .A2(n9622), .ZN(n9342) );
  AOI211_X1 U10666 ( .C1(n9987), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9343), .B(
        n9342), .ZN(n9344) );
  OAI21_X1 U10667 ( .B1(n9970), .B2(n9644), .A(n9344), .ZN(P1_U3264) );
  NOR2_X1 U10668 ( .A1(n9655), .A2(n9359), .ZN(n9347) );
  XNOR2_X1 U10669 ( .A(n9350), .B(n9353), .ZN(n9647) );
  INV_X1 U10670 ( .A(n9647), .ZN(n9373) );
  OAI22_X1 U10671 ( .A1(n9358), .A2(n9995), .B1(n9357), .B2(n9356), .ZN(n9652)
         );
  INV_X1 U10672 ( .A(n9652), .ZN(n9360) );
  NAND2_X1 U10673 ( .A1(n9359), .A2(n9465), .ZN(n9648) );
  AOI211_X1 U10674 ( .C1(n9363), .C2(n9362), .A(n9617), .B(n9361), .ZN(n9651)
         );
  INV_X1 U10675 ( .A(n9364), .ZN(n9365) );
  NAND3_X1 U10676 ( .A1(n9365), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n9619), .ZN(
        n9367) );
  NAND2_X1 U10677 ( .A1(n9987), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9366) );
  OAI211_X1 U10678 ( .C1(n9649), .C2(n9622), .A(n9367), .B(n9366), .ZN(n9368)
         );
  OAI21_X1 U10679 ( .B1(n9373), .B2(n9606), .A(n9372), .ZN(P1_U3356) );
  NAND2_X1 U10680 ( .A1(n9374), .A2(n9637), .ZN(n9377) );
  AOI22_X1 U10681 ( .A1(n9375), .A2(n9619), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9987), .ZN(n9376) );
  OAI211_X1 U10682 ( .C1(n9378), .C2(n9622), .A(n9377), .B(n9376), .ZN(n9379)
         );
  AOI21_X1 U10683 ( .B1(n9380), .B2(n9984), .A(n9379), .ZN(n9381) );
  OAI21_X1 U10684 ( .B1(n9660), .B2(n9606), .A(n9381), .ZN(P1_U3265) );
  OAI211_X1 U10685 ( .C1(n9387), .C2(n9391), .A(n9966), .B(n9388), .ZN(n9661)
         );
  INV_X1 U10686 ( .A(n9661), .ZN(n9399) );
  AOI22_X1 U10687 ( .A1(n9389), .A2(n9619), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9987), .ZN(n9390) );
  OAI21_X1 U10688 ( .B1(n9391), .B2(n9622), .A(n9390), .ZN(n9398) );
  XNOR2_X1 U10689 ( .A(n9393), .B(n9392), .ZN(n9396) );
  INV_X1 U10690 ( .A(n9394), .ZN(n9395) );
  AOI21_X1 U10691 ( .B1(n9396), .B2(n9595), .A(n9395), .ZN(n9662) );
  NOR2_X1 U10692 ( .A1(n9662), .A2(n9987), .ZN(n9397) );
  AOI211_X1 U10693 ( .C1(n9399), .C2(n9637), .A(n9398), .B(n9397), .ZN(n9400)
         );
  OAI21_X1 U10694 ( .B1(n9738), .B2(n9606), .A(n9400), .ZN(P1_U3266) );
  INV_X1 U10695 ( .A(n9387), .ZN(n9401) );
  OAI211_X1 U10696 ( .C1(n9404), .C2(n9428), .A(n9401), .B(n9966), .ZN(n9665)
         );
  INV_X1 U10697 ( .A(n9665), .ZN(n9415) );
  AOI22_X1 U10698 ( .A1(n9402), .A2(n9619), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9987), .ZN(n9403) );
  OAI21_X1 U10699 ( .B1(n9404), .B2(n9622), .A(n9403), .ZN(n9414) );
  OAI21_X1 U10700 ( .B1(n9407), .B2(n9406), .A(n9405), .ZN(n9412) );
  NAND2_X1 U10701 ( .A1(n9408), .A2(n9968), .ZN(n9409) );
  OAI21_X1 U10702 ( .B1(n9410), .B2(n9956), .A(n9409), .ZN(n9411) );
  AOI21_X1 U10703 ( .B1(n9412), .B2(n9595), .A(n9411), .ZN(n9666) );
  NOR2_X1 U10704 ( .A1(n9666), .A2(n9987), .ZN(n9413) );
  AOI211_X1 U10705 ( .C1(n9415), .C2(n9637), .A(n9414), .B(n9413), .ZN(n9416)
         );
  OAI21_X1 U10706 ( .B1(n9743), .B2(n9606), .A(n9416), .ZN(P1_U3267) );
  NAND2_X1 U10707 ( .A1(n9417), .A2(n9418), .ZN(n9419) );
  INV_X1 U10708 ( .A(n9420), .ZN(n9421) );
  AOI21_X1 U10709 ( .B1(n9423), .B2(n9422), .A(n9421), .ZN(n9424) );
  OAI222_X1 U10710 ( .A1(n9427), .A2(n9426), .B1(n9956), .B2(n9425), .C1(n9995), .C2(n9424), .ZN(n9669) );
  INV_X1 U10711 ( .A(n9671), .ZN(n9432) );
  AOI211_X1 U10712 ( .C1(n9671), .C2(n9445), .A(n9617), .B(n9428), .ZN(n9670)
         );
  NAND2_X1 U10713 ( .A1(n9670), .A2(n9637), .ZN(n9431) );
  AOI22_X1 U10714 ( .A1(n9429), .A2(n9619), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9987), .ZN(n9430) );
  OAI211_X1 U10715 ( .C1(n9432), .C2(n9622), .A(n9431), .B(n9430), .ZN(n9433)
         );
  AOI21_X1 U10716 ( .B1(n9669), .B2(n9984), .A(n9433), .ZN(n9434) );
  OAI21_X1 U10717 ( .B1(n9673), .B2(n9606), .A(n9434), .ZN(P1_U3268) );
  XOR2_X1 U10718 ( .A(n9435), .B(n9438), .Z(n9748) );
  NAND2_X1 U10719 ( .A1(n9436), .A2(n9595), .ZN(n9443) );
  INV_X1 U10720 ( .A(n9438), .ZN(n9439) );
  AOI21_X1 U10721 ( .B1(n9437), .B2(n9440), .A(n9439), .ZN(n9442) );
  OAI21_X1 U10722 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9674) );
  INV_X1 U10723 ( .A(n9445), .ZN(n9446) );
  AOI211_X1 U10724 ( .C1(n9676), .C2(n9444), .A(n9617), .B(n9446), .ZN(n9675)
         );
  NAND2_X1 U10725 ( .A1(n9675), .A2(n9637), .ZN(n9449) );
  AOI22_X1 U10726 ( .A1(n9447), .A2(n9619), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9987), .ZN(n9448) );
  OAI211_X1 U10727 ( .C1(n9450), .C2(n9622), .A(n9449), .B(n9448), .ZN(n9451)
         );
  AOI21_X1 U10728 ( .B1(n9984), .B2(n9674), .A(n9451), .ZN(n9452) );
  OAI21_X1 U10729 ( .B1(n9748), .B2(n9606), .A(n9452), .ZN(P1_U3269) );
  AOI22_X1 U10730 ( .A1(n4327), .A2(n9454), .B1(n9461), .B2(n9453), .ZN(n9683)
         );
  INV_X1 U10731 ( .A(n9455), .ZN(n9480) );
  INV_X1 U10732 ( .A(n9444), .ZN(n9456) );
  AOI211_X1 U10733 ( .C1(n9680), .C2(n9480), .A(n9617), .B(n9456), .ZN(n9679)
         );
  INV_X1 U10734 ( .A(n9457), .ZN(n9458) );
  AOI22_X1 U10735 ( .A1(n9458), .A2(n9619), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9987), .ZN(n9459) );
  OAI21_X1 U10736 ( .B1(n9460), .B2(n9622), .A(n9459), .ZN(n9469) );
  INV_X1 U10737 ( .A(n9461), .ZN(n9463) );
  NAND3_X1 U10738 ( .A1(n9472), .A2(n9463), .A3(n9462), .ZN(n9464) );
  NAND2_X1 U10739 ( .A1(n9437), .A2(n9464), .ZN(n9467) );
  AOI222_X1 U10740 ( .A1(n9595), .A2(n9467), .B1(n9466), .B2(n9968), .C1(n9499), .C2(n9465), .ZN(n9682) );
  NOR2_X1 U10741 ( .A1(n9682), .A2(n9987), .ZN(n9468) );
  AOI211_X1 U10742 ( .C1(n9679), .C2(n9637), .A(n9469), .B(n9468), .ZN(n9470)
         );
  OAI21_X1 U10743 ( .B1(n9683), .B2(n9606), .A(n9470), .ZN(P1_U3270) );
  XNOR2_X1 U10744 ( .A(n9471), .B(n9474), .ZN(n9754) );
  OAI21_X1 U10745 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n9479) );
  NAND2_X1 U10746 ( .A1(n9475), .A2(n9968), .ZN(n9476) );
  OAI21_X1 U10747 ( .B1(n9477), .B2(n9956), .A(n9476), .ZN(n9478) );
  AOI21_X1 U10748 ( .B1(n9479), .B2(n9595), .A(n9478), .ZN(n9685) );
  INV_X1 U10749 ( .A(n9685), .ZN(n9488) );
  INV_X1 U10750 ( .A(n9504), .ZN(n9481) );
  OAI211_X1 U10751 ( .C1(n9485), .C2(n9481), .A(n9480), .B(n9966), .ZN(n9684)
         );
  NOR2_X1 U10752 ( .A1(n9684), .A2(n9970), .ZN(n9487) );
  INV_X1 U10753 ( .A(n9482), .ZN(n9483) );
  AOI22_X1 U10754 ( .A1(n9987), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9483), .B2(
        n9619), .ZN(n9484) );
  OAI21_X1 U10755 ( .B1(n9485), .B2(n9622), .A(n9484), .ZN(n9486) );
  AOI211_X1 U10756 ( .C1(n9488), .C2(n9984), .A(n9487), .B(n9486), .ZN(n9489)
         );
  OAI21_X1 U10757 ( .B1(n9754), .B2(n9606), .A(n9489), .ZN(P1_U3271) );
  XNOR2_X1 U10758 ( .A(n9491), .B(n9490), .ZN(n9759) );
  NAND2_X1 U10759 ( .A1(n9493), .A2(n9492), .ZN(n9495) );
  NAND2_X1 U10760 ( .A1(n9495), .A2(n9494), .ZN(n9497) );
  NAND2_X1 U10761 ( .A1(n9497), .A2(n9496), .ZN(n9503) );
  NAND2_X1 U10762 ( .A1(n9499), .A2(n9498), .ZN(n9500) );
  OAI21_X1 U10763 ( .B1(n9501), .B2(n9956), .A(n9500), .ZN(n9502) );
  AOI21_X1 U10764 ( .B1(n9503), .B2(n9595), .A(n9502), .ZN(n9689) );
  INV_X1 U10765 ( .A(n9689), .ZN(n9511) );
  OAI211_X1 U10766 ( .C1(n9508), .C2(n4307), .A(n9504), .B(n9966), .ZN(n9688)
         );
  NOR2_X1 U10767 ( .A1(n9688), .A2(n9970), .ZN(n9510) );
  INV_X1 U10768 ( .A(n9505), .ZN(n9506) );
  AOI22_X1 U10769 ( .A1(n9987), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9506), .B2(
        n9619), .ZN(n9507) );
  OAI21_X1 U10770 ( .B1(n9508), .B2(n9622), .A(n9507), .ZN(n9509) );
  AOI211_X1 U10771 ( .C1(n9511), .C2(n9984), .A(n9510), .B(n9509), .ZN(n9512)
         );
  OAI21_X1 U10772 ( .B1(n9759), .B2(n9606), .A(n9512), .ZN(P1_U3272) );
  OAI21_X1 U10773 ( .B1(n9514), .B2(n9515), .A(n9513), .ZN(n9694) );
  INV_X1 U10774 ( .A(n9694), .ZN(n9527) );
  INV_X1 U10775 ( .A(n9515), .ZN(n9516) );
  XNOR2_X1 U10776 ( .A(n7781), .B(n9516), .ZN(n9517) );
  NAND2_X1 U10777 ( .A1(n9517), .A2(n9595), .ZN(n9519) );
  NAND2_X1 U10778 ( .A1(n9519), .A2(n9518), .ZN(n9692) );
  AOI211_X1 U10779 ( .C1(n9521), .C2(n9520), .A(n9617), .B(n4307), .ZN(n9693)
         );
  NAND2_X1 U10780 ( .A1(n9693), .A2(n9637), .ZN(n9524) );
  AOI22_X1 U10781 ( .A1(n9987), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9522), .B2(
        n9619), .ZN(n9523) );
  OAI211_X1 U10782 ( .C1(n9763), .C2(n9622), .A(n9524), .B(n9523), .ZN(n9525)
         );
  AOI21_X1 U10783 ( .B1(n9984), .B2(n9692), .A(n9525), .ZN(n9526) );
  OAI21_X1 U10784 ( .B1(n9527), .B2(n9606), .A(n9526), .ZN(P1_U3273) );
  XOR2_X1 U10785 ( .A(n9528), .B(n9529), .Z(n9768) );
  XNOR2_X1 U10786 ( .A(n9530), .B(n9529), .ZN(n9532) );
  AOI21_X1 U10787 ( .B1(n9532), .B2(n9595), .A(n9531), .ZN(n9698) );
  INV_X1 U10788 ( .A(n9698), .ZN(n9538) );
  OAI211_X1 U10789 ( .C1(n9535), .C2(n9551), .A(n9520), .B(n9966), .ZN(n9697)
         );
  NOR2_X1 U10790 ( .A1(n9697), .A2(n9970), .ZN(n9537) );
  AOI22_X1 U10791 ( .A1(n9987), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9533), .B2(
        n9619), .ZN(n9534) );
  OAI21_X1 U10792 ( .B1(n9535), .B2(n9622), .A(n9534), .ZN(n9536) );
  AOI211_X1 U10793 ( .C1(n9538), .C2(n9984), .A(n9537), .B(n9536), .ZN(n9539)
         );
  OAI21_X1 U10794 ( .B1(n9768), .B2(n9606), .A(n9539), .ZN(P1_U3274) );
  XNOR2_X1 U10795 ( .A(n9541), .B(n9540), .ZN(n9772) );
  NAND2_X1 U10796 ( .A1(n9542), .A2(n9543), .ZN(n9545) );
  NAND2_X1 U10797 ( .A1(n9545), .A2(n9544), .ZN(n9547) );
  NAND2_X1 U10798 ( .A1(n9547), .A2(n9546), .ZN(n9548) );
  NAND2_X1 U10799 ( .A1(n9548), .A2(n9595), .ZN(n9550) );
  NAND2_X1 U10800 ( .A1(n9550), .A2(n9549), .ZN(n9701) );
  OAI21_X1 U10801 ( .B1(n9567), .B2(n9556), .A(n9966), .ZN(n9552) );
  NOR2_X1 U10802 ( .A1(n9552), .A2(n9551), .ZN(n9702) );
  NAND2_X1 U10803 ( .A1(n9702), .A2(n9637), .ZN(n9555) );
  AOI22_X1 U10804 ( .A1(n9987), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9553), .B2(
        n9619), .ZN(n9554) );
  OAI211_X1 U10805 ( .C1(n9556), .C2(n9622), .A(n9555), .B(n9554), .ZN(n9557)
         );
  AOI21_X1 U10806 ( .B1(n9701), .B2(n9984), .A(n9557), .ZN(n9558) );
  OAI21_X1 U10807 ( .B1(n9772), .B2(n9606), .A(n9558), .ZN(P1_U3275) );
  XOR2_X1 U10808 ( .A(n9560), .B(n9559), .Z(n9777) );
  AOI21_X1 U10809 ( .B1(n9561), .B2(n9560), .A(n9995), .ZN(n9564) );
  INV_X1 U10810 ( .A(n9562), .ZN(n9563) );
  AOI21_X1 U10811 ( .B1(n9564), .B2(n9542), .A(n9563), .ZN(n9707) );
  INV_X1 U10812 ( .A(n9707), .ZN(n9573) );
  NAND2_X1 U10813 ( .A1(n9581), .A2(n9775), .ZN(n9565) );
  NAND2_X1 U10814 ( .A1(n9565), .A2(n9966), .ZN(n9566) );
  OR2_X1 U10815 ( .A1(n9567), .A2(n9566), .ZN(n9706) );
  NOR2_X1 U10816 ( .A1(n9706), .A2(n9970), .ZN(n9572) );
  AOI22_X1 U10817 ( .A1(n9987), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9568), .B2(
        n9619), .ZN(n9569) );
  OAI21_X1 U10818 ( .B1(n9570), .B2(n9622), .A(n9569), .ZN(n9571) );
  AOI211_X1 U10819 ( .C1(n9573), .C2(n9984), .A(n9572), .B(n9571), .ZN(n9574)
         );
  OAI21_X1 U10820 ( .B1(n9777), .B2(n9606), .A(n9574), .ZN(P1_U3276) );
  XNOR2_X1 U10821 ( .A(n9575), .B(n9576), .ZN(n9712) );
  INV_X1 U10822 ( .A(n9712), .ZN(n9589) );
  XNOR2_X1 U10823 ( .A(n9577), .B(n9576), .ZN(n9578) );
  NAND2_X1 U10824 ( .A1(n9578), .A2(n9595), .ZN(n9580) );
  NAND2_X1 U10825 ( .A1(n9580), .A2(n9579), .ZN(n9710) );
  INV_X1 U10826 ( .A(n9581), .ZN(n9582) );
  AOI211_X1 U10827 ( .C1(n9583), .C2(n9598), .A(n9617), .B(n9582), .ZN(n9711)
         );
  NAND2_X1 U10828 ( .A1(n9711), .A2(n9637), .ZN(n9586) );
  AOI22_X1 U10829 ( .A1(n9987), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9584), .B2(
        n9619), .ZN(n9585) );
  OAI211_X1 U10830 ( .C1(n4479), .C2(n9622), .A(n9586), .B(n9585), .ZN(n9587)
         );
  AOI21_X1 U10831 ( .B1(n9984), .B2(n9710), .A(n9587), .ZN(n9588) );
  OAI21_X1 U10832 ( .B1(n9589), .B2(n9606), .A(n9588), .ZN(P1_U3277) );
  XOR2_X1 U10833 ( .A(n9590), .B(n9592), .Z(n9788) );
  OAI21_X1 U10834 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9596) );
  AOI21_X1 U10835 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9717) );
  INV_X1 U10836 ( .A(n9717), .ZN(n9604) );
  OAI211_X1 U10837 ( .C1(n9597), .C2(n9601), .A(n9966), .B(n9598), .ZN(n9716)
         );
  NOR2_X1 U10838 ( .A1(n9716), .A2(n9970), .ZN(n9603) );
  AOI22_X1 U10839 ( .A1(n9987), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9599), .B2(
        n9619), .ZN(n9600) );
  OAI21_X1 U10840 ( .B1(n9601), .B2(n9622), .A(n9600), .ZN(n9602) );
  AOI211_X1 U10841 ( .C1(n9604), .C2(n9984), .A(n9603), .B(n9602), .ZN(n9605)
         );
  OAI21_X1 U10842 ( .B1(n9788), .B2(n9606), .A(n9605), .ZN(P1_U3278) );
  XNOR2_X1 U10843 ( .A(n9607), .B(n9611), .ZN(n9624) );
  INV_X1 U10844 ( .A(n9608), .ZN(n9609) );
  AOI211_X1 U10845 ( .C1(n9611), .C2(n9610), .A(n9995), .B(n9609), .ZN(n9614)
         );
  INV_X1 U10846 ( .A(n9612), .ZN(n9613) );
  AOI211_X1 U10847 ( .C1(n9624), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9726)
         );
  INV_X1 U10848 ( .A(n9616), .ZN(n9618) );
  AOI211_X1 U10849 ( .C1(n9723), .C2(n9618), .A(n9617), .B(n9597), .ZN(n9722)
         );
  AOI22_X1 U10850 ( .A1(n9987), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9620), .B2(
        n9619), .ZN(n9621) );
  OAI21_X1 U10851 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9627) );
  INV_X1 U10852 ( .A(n9624), .ZN(n9728) );
  NOR2_X1 U10853 ( .A1(n9728), .A2(n9625), .ZN(n9626) );
  AOI211_X1 U10854 ( .C1(n9722), .C2(n9637), .A(n9627), .B(n9626), .ZN(n9628)
         );
  OAI21_X1 U10855 ( .B1(n9987), .B2(n9726), .A(n9628), .ZN(P1_U3279) );
  NAND2_X1 U10856 ( .A1(n9629), .A2(n9984), .ZN(n9642) );
  INV_X1 U10857 ( .A(n9630), .ZN(n9631) );
  OAI22_X1 U10858 ( .A1(n9984), .A2(n9632), .B1(n9631), .B2(n9978), .ZN(n9633)
         );
  AOI21_X1 U10859 ( .B1(n9635), .B2(n9634), .A(n9633), .ZN(n9641) );
  NAND2_X1 U10860 ( .A1(n9636), .A2(n9964), .ZN(n9640) );
  NAND2_X1 U10861 ( .A1(n9638), .A2(n9637), .ZN(n9639) );
  NAND4_X1 U10862 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(
        P1_U3287) );
  AND2_X1 U10863 ( .A1(n9644), .A2(n9643), .ZN(n9729) );
  MUX2_X1 U10864 ( .A(n9645), .B(n9729), .S(n10042), .Z(n9646) );
  OAI21_X1 U10865 ( .B1(n9732), .B2(n9715), .A(n9646), .ZN(P1_U3552) );
  NAND2_X1 U10866 ( .A1(n9647), .A2(n10026), .ZN(n9654) );
  OAI21_X1 U10867 ( .B1(n9649), .B2(n10023), .A(n9648), .ZN(n9650) );
  NAND2_X1 U10868 ( .A1(n9654), .A2(n9653), .ZN(n9733) );
  MUX2_X1 U10869 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9733), .S(n10042), .Z(
        P1_U3551) );
  NAND2_X1 U10870 ( .A1(n9655), .A2(n9719), .ZN(n9659) );
  MUX2_X1 U10871 ( .A(n9657), .B(n9656), .S(n10042), .Z(n9658) );
  OAI211_X1 U10872 ( .C1(n9660), .C2(n9721), .A(n9659), .B(n9658), .ZN(
        P1_U3550) );
  NAND2_X1 U10873 ( .A1(n9662), .A2(n9661), .ZN(n9734) );
  MUX2_X1 U10874 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9734), .S(n10042), .Z(
        n9663) );
  AOI21_X1 U10875 ( .B1(n9719), .B2(n9736), .A(n9663), .ZN(n9664) );
  OAI21_X1 U10876 ( .B1(n9738), .B2(n9721), .A(n9664), .ZN(P1_U3549) );
  NAND2_X1 U10877 ( .A1(n9666), .A2(n9665), .ZN(n9739) );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9739), .S(n10042), .Z(
        n9667) );
  AOI21_X1 U10879 ( .B1(n9719), .B2(n9741), .A(n9667), .ZN(n9668) );
  OAI21_X1 U10880 ( .B1(n9743), .B2(n9721), .A(n9668), .ZN(P1_U3548) );
  INV_X1 U10881 ( .A(n10026), .ZN(n9996) );
  AOI211_X1 U10882 ( .C1(n9724), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9672)
         );
  OAI21_X1 U10883 ( .B1(n9673), .B2(n9996), .A(n9672), .ZN(n9744) );
  MUX2_X1 U10884 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9744), .S(n10042), .Z(
        P1_U3547) );
  AOI211_X1 U10885 ( .C1(n9724), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9745)
         );
  MUX2_X1 U10886 ( .A(n9677), .B(n9745), .S(n10042), .Z(n9678) );
  OAI21_X1 U10887 ( .B1(n9748), .B2(n9721), .A(n9678), .ZN(P1_U3546) );
  AOI21_X1 U10888 ( .B1(n9724), .B2(n9680), .A(n9679), .ZN(n9681) );
  OAI211_X1 U10889 ( .C1(n9683), .C2(n9996), .A(n9682), .B(n9681), .ZN(n9749)
         );
  MUX2_X1 U10890 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9749), .S(n10042), .Z(
        P1_U3545) );
  NAND2_X1 U10891 ( .A1(n9685), .A2(n9684), .ZN(n9750) );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9750), .S(n10042), .Z(
        n9686) );
  AOI21_X1 U10893 ( .B1(n9719), .B2(n9752), .A(n9686), .ZN(n9687) );
  OAI21_X1 U10894 ( .B1(n9754), .B2(n9721), .A(n9687), .ZN(P1_U3544) );
  NAND2_X1 U10895 ( .A1(n9689), .A2(n9688), .ZN(n9755) );
  MUX2_X1 U10896 ( .A(n9755), .B(P1_REG1_REG_21__SCAN_IN), .S(n10039), .Z(
        n9690) );
  AOI21_X1 U10897 ( .B1(n9719), .B2(n9757), .A(n9690), .ZN(n9691) );
  OAI21_X1 U10898 ( .B1(n9759), .B2(n9721), .A(n9691), .ZN(P1_U3543) );
  INV_X1 U10899 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9695) );
  AOI211_X1 U10900 ( .C1(n9694), .C2(n10026), .A(n9693), .B(n9692), .ZN(n9760)
         );
  MUX2_X1 U10901 ( .A(n9695), .B(n9760), .S(n10042), .Z(n9696) );
  OAI21_X1 U10902 ( .B1(n9763), .B2(n9715), .A(n9696), .ZN(P1_U3542) );
  NAND2_X1 U10903 ( .A1(n9698), .A2(n9697), .ZN(n9764) );
  MUX2_X1 U10904 ( .A(n9764), .B(P1_REG1_REG_19__SCAN_IN), .S(n10039), .Z(
        n9699) );
  AOI21_X1 U10905 ( .B1(n9719), .B2(n9766), .A(n9699), .ZN(n9700) );
  OAI21_X1 U10906 ( .B1(n9768), .B2(n9721), .A(n9700), .ZN(P1_U3541) );
  AOI211_X1 U10907 ( .C1(n9724), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9769)
         );
  MUX2_X1 U10908 ( .A(n9704), .B(n9769), .S(n10042), .Z(n9705) );
  OAI21_X1 U10909 ( .B1(n9772), .B2(n9721), .A(n9705), .ZN(P1_U3540) );
  NAND2_X1 U10910 ( .A1(n9707), .A2(n9706), .ZN(n9773) );
  MUX2_X1 U10911 ( .A(n9773), .B(P1_REG1_REG_17__SCAN_IN), .S(n10039), .Z(
        n9708) );
  AOI21_X1 U10912 ( .B1(n9719), .B2(n9775), .A(n9708), .ZN(n9709) );
  OAI21_X1 U10913 ( .B1(n9777), .B2(n9721), .A(n9709), .ZN(P1_U3539) );
  AOI211_X1 U10914 ( .C1(n9712), .C2(n10026), .A(n9711), .B(n9710), .ZN(n9778)
         );
  MUX2_X1 U10915 ( .A(n9713), .B(n9778), .S(n10042), .Z(n9714) );
  OAI21_X1 U10916 ( .B1(n4479), .B2(n9715), .A(n9714), .ZN(P1_U3538) );
  NAND2_X1 U10917 ( .A1(n9717), .A2(n9716), .ZN(n9782) );
  MUX2_X1 U10918 ( .A(n9782), .B(P1_REG1_REG_15__SCAN_IN), .S(n10039), .Z(
        n9718) );
  AOI21_X1 U10919 ( .B1(n9719), .B2(n9784), .A(n9718), .ZN(n9720) );
  OAI21_X1 U10920 ( .B1(n9788), .B2(n9721), .A(n9720), .ZN(P1_U3537) );
  AOI21_X1 U10921 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9725) );
  OAI211_X1 U10922 ( .C1(n9728), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9789)
         );
  MUX2_X1 U10923 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9789), .S(n10042), .Z(
        P1_U3536) );
  INV_X1 U10924 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U10925 ( .A(n9730), .B(n9729), .S(n10030), .Z(n9731) );
  OAI21_X1 U10926 ( .B1(n9732), .B2(n9781), .A(n9731), .ZN(P1_U3520) );
  MUX2_X1 U10927 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9733), .S(n10030), .Z(
        P1_U3519) );
  MUX2_X1 U10928 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9734), .S(n10030), .Z(
        n9735) );
  AOI21_X1 U10929 ( .B1(n9785), .B2(n9736), .A(n9735), .ZN(n9737) );
  OAI21_X1 U10930 ( .B1(n9738), .B2(n9787), .A(n9737), .ZN(P1_U3517) );
  MUX2_X1 U10931 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9739), .S(n10030), .Z(
        n9740) );
  AOI21_X1 U10932 ( .B1(n9785), .B2(n9741), .A(n9740), .ZN(n9742) );
  OAI21_X1 U10933 ( .B1(n9743), .B2(n9787), .A(n9742), .ZN(P1_U3516) );
  MUX2_X1 U10934 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9744), .S(n10030), .Z(
        P1_U3515) );
  INV_X1 U10935 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9746) );
  MUX2_X1 U10936 ( .A(n9746), .B(n9745), .S(n10030), .Z(n9747) );
  OAI21_X1 U10937 ( .B1(n9748), .B2(n9787), .A(n9747), .ZN(P1_U3514) );
  MUX2_X1 U10938 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9749), .S(n10030), .Z(
        P1_U3513) );
  MUX2_X1 U10939 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9750), .S(n10030), .Z(
        n9751) );
  AOI21_X1 U10940 ( .B1(n9785), .B2(n9752), .A(n9751), .ZN(n9753) );
  OAI21_X1 U10941 ( .B1(n9754), .B2(n9787), .A(n9753), .ZN(P1_U3512) );
  MUX2_X1 U10942 ( .A(n9755), .B(P1_REG0_REG_21__SCAN_IN), .S(n10028), .Z(
        n9756) );
  AOI21_X1 U10943 ( .B1(n9785), .B2(n9757), .A(n9756), .ZN(n9758) );
  OAI21_X1 U10944 ( .B1(n9759), .B2(n9787), .A(n9758), .ZN(P1_U3511) );
  INV_X1 U10945 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9761) );
  MUX2_X1 U10946 ( .A(n9761), .B(n9760), .S(n10030), .Z(n9762) );
  OAI21_X1 U10947 ( .B1(n9763), .B2(n9781), .A(n9762), .ZN(P1_U3510) );
  MUX2_X1 U10948 ( .A(n9764), .B(P1_REG0_REG_19__SCAN_IN), .S(n10028), .Z(
        n9765) );
  AOI21_X1 U10949 ( .B1(n9785), .B2(n9766), .A(n9765), .ZN(n9767) );
  OAI21_X1 U10950 ( .B1(n9768), .B2(n9787), .A(n9767), .ZN(P1_U3509) );
  INV_X1 U10951 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U10952 ( .A(n9770), .B(n9769), .S(n10030), .Z(n9771) );
  OAI21_X1 U10953 ( .B1(n9772), .B2(n9787), .A(n9771), .ZN(P1_U3507) );
  MUX2_X1 U10954 ( .A(n9773), .B(P1_REG0_REG_17__SCAN_IN), .S(n10028), .Z(
        n9774) );
  AOI21_X1 U10955 ( .B1(n9785), .B2(n9775), .A(n9774), .ZN(n9776) );
  OAI21_X1 U10956 ( .B1(n9777), .B2(n9787), .A(n9776), .ZN(P1_U3504) );
  INV_X1 U10957 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9779) );
  MUX2_X1 U10958 ( .A(n9779), .B(n9778), .S(n10030), .Z(n9780) );
  OAI21_X1 U10959 ( .B1(n4479), .B2(n9781), .A(n9780), .ZN(P1_U3501) );
  MUX2_X1 U10960 ( .A(n9782), .B(P1_REG0_REG_15__SCAN_IN), .S(n10028), .Z(
        n9783) );
  AOI21_X1 U10961 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9786) );
  OAI21_X1 U10962 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(P1_U3498) );
  MUX2_X1 U10963 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9789), .S(n10030), .Z(
        P1_U3495) );
  MUX2_X1 U10964 ( .A(P1_D_REG_0__SCAN_IN), .B(n9790), .S(n9992), .Z(P1_U3439)
         );
  NOR4_X1 U10965 ( .A1(n4648), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9791), .ZN(n9793) );
  AOI21_X1 U10966 ( .B1(n9794), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9793), .ZN(
        n9795) );
  OAI21_X1 U10967 ( .B1(n9796), .B2(n9800), .A(n9795), .ZN(P1_U3324) );
  OAI222_X1 U10968 ( .A1(n9800), .A2(n9799), .B1(n5577), .B2(P1_U3086), .C1(
        n9798), .C2(n9797), .ZN(P1_U3326) );
  MUX2_X1 U10969 ( .A(n9801), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI22_X1 U10970 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(P1_U3086), .ZN(n9812) );
  OAI211_X1 U10971 ( .C1(n9804), .C2(n9803), .A(n9945), .B(n9802), .ZN(n9811)
         );
  OAI211_X1 U10972 ( .C1(n9807), .C2(n9806), .A(n9941), .B(n9805), .ZN(n9810)
         );
  NAND2_X1 U10973 ( .A1(n9943), .A2(n9808), .ZN(n9809) );
  NAND4_X1 U10974 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(
        P1_U3250) );
  AOI22_X1 U10975 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_8__SCAN_IN), .B2(P1_U3086), .ZN(n9823) );
  OAI211_X1 U10976 ( .C1(n9815), .C2(n9814), .A(n9941), .B(n9813), .ZN(n9822)
         );
  OAI211_X1 U10977 ( .C1(n9818), .C2(n9817), .A(n9945), .B(n9816), .ZN(n9821)
         );
  NAND2_X1 U10978 ( .A1(n9943), .A2(n9819), .ZN(n9820) );
  NAND4_X1 U10979 ( .A1(n9823), .A2(n9822), .A3(n9821), .A4(n9820), .ZN(
        P1_U3251) );
  AOI21_X1 U10980 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9828) );
  OR2_X1 U10981 ( .A1(n9828), .A2(n9827), .ZN(n9835) );
  AOI21_X1 U10982 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n9833) );
  OR2_X1 U10983 ( .A1(n9833), .A2(n9832), .ZN(n9834) );
  OAI211_X1 U10984 ( .C1(n9837), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9838)
         );
  INV_X1 U10985 ( .A(n9838), .ZN(n9840) );
  OAI211_X1 U10986 ( .C1(n9950), .C2(n9841), .A(n9840), .B(n9839), .ZN(
        P1_U3252) );
  OAI21_X1 U10987 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9853) );
  AOI21_X1 U10988 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9848) );
  OAI21_X1 U10989 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  AOI21_X1 U10990 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9854) );
  OAI21_X1 U10991 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(P1_U3217) );
  XNOR2_X1 U10992 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10993 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U10994 ( .A1(n4296), .A2(n10031), .ZN(n9859) );
  NOR2_X1 U10995 ( .A1(n9857), .A2(n9859), .ZN(n9858) );
  MUX2_X1 U10996 ( .A(n9859), .B(n9858), .S(P1_IR_REG_0__SCAN_IN), .Z(n9862)
         );
  INV_X1 U10997 ( .A(n9860), .ZN(n9861) );
  OR2_X1 U10998 ( .A1(n9862), .A2(n9861), .ZN(n9864) );
  AOI22_X1 U10999 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9863) );
  OAI21_X1 U11000 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(P1_U3243) );
  AOI22_X1 U11001 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_5__SCAN_IN), .B2(P1_U3086), .ZN(n9877) );
  INV_X1 U11002 ( .A(n9866), .ZN(n9867) );
  NAND2_X1 U11003 ( .A1(n9943), .A2(n9867), .ZN(n9876) );
  OAI211_X1 U11004 ( .C1(n9870), .C2(n9869), .A(n9941), .B(n9868), .ZN(n9875)
         );
  OAI211_X1 U11005 ( .C1(n9873), .C2(n9872), .A(n9945), .B(n9871), .ZN(n9874)
         );
  NAND4_X1 U11006 ( .A1(n9877), .A2(n9876), .A3(n9875), .A4(n9874), .ZN(
        P1_U3248) );
  OAI21_X1 U11007 ( .B1(n9950), .B2(n9879), .A(n9878), .ZN(n9880) );
  AOI21_X1 U11008 ( .B1(n9881), .B2(n9943), .A(n9880), .ZN(n9890) );
  OAI211_X1 U11009 ( .C1(n9884), .C2(n9883), .A(n9945), .B(n9882), .ZN(n9889)
         );
  OAI211_X1 U11010 ( .C1(n9887), .C2(n9886), .A(n9941), .B(n9885), .ZN(n9888)
         );
  NAND3_X1 U11011 ( .A1(n9890), .A2(n9889), .A3(n9888), .ZN(P1_U3249) );
  AOI22_X1 U11012 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(P1_U3086), .ZN(n9901) );
  NAND2_X1 U11013 ( .A1(n9943), .A2(n9891), .ZN(n9900) );
  OAI211_X1 U11014 ( .C1(n9894), .C2(n9893), .A(n9941), .B(n9892), .ZN(n9899)
         );
  OAI211_X1 U11015 ( .C1(n9897), .C2(n9896), .A(n9945), .B(n9895), .ZN(n9898)
         );
  NAND4_X1 U11016 ( .A1(n9901), .A2(n9900), .A3(n9899), .A4(n9898), .ZN(
        P1_U3254) );
  AOI22_X1 U11017 ( .A1(n9924), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(
        P1_REG3_REG_13__SCAN_IN), .B2(P1_U3086), .ZN(n9912) );
  NAND2_X1 U11018 ( .A1(n9943), .A2(n9902), .ZN(n9911) );
  OAI211_X1 U11019 ( .C1(n9905), .C2(n9904), .A(n9941), .B(n9903), .ZN(n9910)
         );
  OAI211_X1 U11020 ( .C1(n9908), .C2(n9907), .A(n9945), .B(n9906), .ZN(n9909)
         );
  NAND4_X1 U11021 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(
        P1_U3256) );
  AOI22_X1 U11022 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(P1_U3086), .ZN(n9923) );
  NAND2_X1 U11023 ( .A1(n9943), .A2(n9913), .ZN(n9922) );
  OAI211_X1 U11024 ( .C1(n9916), .C2(n9915), .A(n9945), .B(n9914), .ZN(n9921)
         );
  OAI211_X1 U11025 ( .C1(n9919), .C2(n9918), .A(n9941), .B(n9917), .ZN(n9920)
         );
  NAND4_X1 U11026 ( .A1(n9923), .A2(n9922), .A3(n9921), .A4(n9920), .ZN(
        P1_U3257) );
  AOI22_X1 U11027 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9924), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(P1_U3086), .ZN(n9933) );
  NAND2_X1 U11028 ( .A1(n9943), .A2(n9925), .ZN(n9932) );
  OAI211_X1 U11029 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9927), .A(n9941), .B(
        n9926), .ZN(n9931) );
  OAI211_X1 U11030 ( .C1(P1_REG2_REG_15__SCAN_IN), .C2(n9929), .A(n9945), .B(
        n9928), .ZN(n9930) );
  NAND4_X1 U11031 ( .A1(n9933), .A2(n9932), .A3(n9931), .A4(n9930), .ZN(
        P1_U3258) );
  OAI21_X1 U11032 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9946) );
  NAND2_X1 U11033 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  NAND2_X1 U11034 ( .A1(n9940), .A2(n9939), .ZN(n9942) );
  AOI222_X1 U11035 ( .A1(n9946), .A2(n9945), .B1(n9944), .B2(n9943), .C1(n9942), .C2(n9941), .ZN(n9948) );
  OAI211_X1 U11036 ( .C1(n9950), .C2(n9949), .A(n9948), .B(n9947), .ZN(
        P1_U3260) );
  XNOR2_X1 U11037 ( .A(n4370), .B(n9954), .ZN(n10027) );
  OAI21_X1 U11038 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9955) );
  XNOR2_X1 U11039 ( .A(n9955), .B(n9954), .ZN(n9958) );
  OAI22_X1 U11040 ( .A1(n9958), .A2(n9995), .B1(n9957), .B2(n9956), .ZN(n10025) );
  OAI22_X1 U11041 ( .A1(n4456), .A2(n9961), .B1(n9978), .B2(n9960), .ZN(n9962)
         );
  OR2_X1 U11042 ( .A1(n10025), .A2(n9962), .ZN(n9963) );
  AOI22_X1 U11043 ( .A1(n10027), .A2(n9964), .B1(n9984), .B2(n9963), .ZN(n9973) );
  OAI211_X1 U11044 ( .C1(n4456), .C2(n5951), .A(n9967), .B(n9966), .ZN(n10022)
         );
  NAND2_X1 U11045 ( .A1(n9969), .A2(n9968), .ZN(n10021) );
  AOI21_X1 U11046 ( .B1(n10022), .B2(n10021), .A(n9970), .ZN(n9971) );
  INV_X1 U11047 ( .A(n9971), .ZN(n9972) );
  OAI211_X1 U11048 ( .C1(n9984), .C2(n9974), .A(n9973), .B(n9972), .ZN(
        P1_U3284) );
  INV_X1 U11049 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9986) );
  NOR2_X1 U11050 ( .A1(n9976), .A2(n9975), .ZN(n9997) );
  INV_X1 U11051 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9979) );
  INV_X1 U11052 ( .A(n9998), .ZN(n9977) );
  OAI21_X1 U11053 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(n9982) );
  NOR2_X1 U11054 ( .A1(n9994), .A2(n9980), .ZN(n9981) );
  AOI211_X1 U11055 ( .C1(n9997), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9985)
         );
  AOI22_X1 U11056 ( .A1(n9987), .A2(n9986), .B1(n9985), .B2(n9984), .ZN(
        P1_U3293) );
  NOR2_X1 U11057 ( .A1(n9992), .A2(n9988), .ZN(P1_U3294) );
  AND2_X1 U11058 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9993), .ZN(P1_U3295) );
  NOR2_X1 U11059 ( .A1(n9992), .A2(n9989), .ZN(P1_U3296) );
  AND2_X1 U11060 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9993), .ZN(P1_U3297) );
  AND2_X1 U11061 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9993), .ZN(P1_U3298) );
  NOR2_X1 U11062 ( .A1(n9992), .A2(n9990), .ZN(P1_U3299) );
  AND2_X1 U11063 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9993), .ZN(P1_U3300) );
  AND2_X1 U11064 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9993), .ZN(P1_U3301) );
  AND2_X1 U11065 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9993), .ZN(P1_U3302) );
  AND2_X1 U11066 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9993), .ZN(P1_U3303) );
  AND2_X1 U11067 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9993), .ZN(P1_U3304) );
  NOR2_X1 U11068 ( .A1(n9992), .A2(n9991), .ZN(P1_U3305) );
  AND2_X1 U11069 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9993), .ZN(P1_U3306) );
  AND2_X1 U11070 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9993), .ZN(P1_U3307) );
  AND2_X1 U11071 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9993), .ZN(P1_U3308) );
  AND2_X1 U11072 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9993), .ZN(P1_U3309) );
  AND2_X1 U11073 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9993), .ZN(P1_U3310) );
  AND2_X1 U11074 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9993), .ZN(P1_U3311) );
  AND2_X1 U11075 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9993), .ZN(P1_U3312) );
  AND2_X1 U11076 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9993), .ZN(P1_U3313) );
  AND2_X1 U11077 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9993), .ZN(P1_U3314) );
  AND2_X1 U11078 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9993), .ZN(P1_U3315) );
  AND2_X1 U11079 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9993), .ZN(P1_U3316) );
  AND2_X1 U11080 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9993), .ZN(P1_U3317) );
  AND2_X1 U11081 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9993), .ZN(P1_U3318) );
  AND2_X1 U11082 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9993), .ZN(P1_U3319) );
  AND2_X1 U11083 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9993), .ZN(P1_U3320) );
  AND2_X1 U11084 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9993), .ZN(P1_U3321) );
  AND2_X1 U11085 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9993), .ZN(P1_U3322) );
  AND2_X1 U11086 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9993), .ZN(P1_U3323) );
  AOI21_X1 U11087 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9999) );
  NOR3_X1 U11088 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10032) );
  INV_X1 U11089 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11090 ( .A1(n10030), .A2(n10032), .B1(n10000), .B2(n10028), .ZN(
        P1_U3453) );
  OAI21_X1 U11091 ( .B1(n5991), .B2(n10023), .A(n10001), .ZN(n10002) );
  AOI21_X1 U11092 ( .B1(n10003), .B2(n10016), .A(n10002), .ZN(n10004) );
  AND2_X1 U11093 ( .A1(n10005), .A2(n10004), .ZN(n10034) );
  INV_X1 U11094 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U11095 ( .A1(n10030), .A2(n10034), .B1(n10006), .B2(n10028), .ZN(
        P1_U3456) );
  OAI21_X1 U11096 ( .B1(n10008), .B2(n10023), .A(n10007), .ZN(n10010) );
  AOI211_X1 U11097 ( .C1(n10026), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10036) );
  INV_X1 U11098 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11099 ( .A1(n10030), .A2(n10036), .B1(n10012), .B2(n10028), .ZN(
        P1_U3468) );
  OAI21_X1 U11100 ( .B1(n10014), .B2(n10023), .A(n10013), .ZN(n10015) );
  AOI21_X1 U11101 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(n10018) );
  AND2_X1 U11102 ( .A1(n10019), .A2(n10018), .ZN(n10038) );
  INV_X1 U11103 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11104 ( .A1(n10030), .A2(n10038), .B1(n10020), .B2(n10028), .ZN(
        P1_U3474) );
  OAI211_X1 U11105 ( .C1(n4456), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10024) );
  AOI211_X1 U11106 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10041) );
  INV_X1 U11107 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U11108 ( .A1(n10030), .A2(n10041), .B1(n10029), .B2(n10028), .ZN(
        P1_U3480) );
  AOI22_X1 U11109 ( .A1(n10042), .A2(n10032), .B1(n10031), .B2(n10039), .ZN(
        P1_U3522) );
  AOI22_X1 U11110 ( .A1(n10042), .A2(n10034), .B1(n10033), .B2(n10039), .ZN(
        P1_U3523) );
  AOI22_X1 U11111 ( .A1(n10042), .A2(n10036), .B1(n10035), .B2(n10039), .ZN(
        P1_U3527) );
  AOI22_X1 U11112 ( .A1(n10042), .A2(n10038), .B1(n10037), .B2(n10039), .ZN(
        P1_U3529) );
  AOI22_X1 U11113 ( .A1(n10042), .A2(n10041), .B1(n10040), .B2(n10039), .ZN(
        P1_U3531) );
  NAND3_X1 U11114 ( .A1(n10044), .A2(n4378), .A3(n10043), .ZN(n10045) );
  NAND2_X1 U11115 ( .A1(n10046), .A2(n10045), .ZN(n10051) );
  AOI222_X1 U11116 ( .A1(n10051), .A2(n10050), .B1(P2_ADDR_REG_8__SCAN_IN), 
        .B2(n10049), .C1(n10048), .C2(n10047), .ZN(n10065) );
  AOI21_X1 U11117 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n10056) );
  OR2_X1 U11118 ( .A1(n10056), .A2(n10055), .ZN(n10063) );
  OAI21_X1 U11119 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10061) );
  NAND2_X1 U11120 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  NAND4_X1 U11121 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        P2_U3190) );
  AOI22_X1 U11122 ( .A1(n10121), .A2(n5026), .B1(n10066), .B2(n10119), .ZN(
        P2_U3390) );
  NOR2_X1 U11123 ( .A1(n10067), .A2(n10108), .ZN(n10069) );
  AOI211_X1 U11124 ( .C1(n10080), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10122) );
  AOI22_X1 U11125 ( .A1(n10121), .A2(n5012), .B1(n10122), .B2(n10119), .ZN(
        P2_U3393) );
  OAI22_X1 U11126 ( .A1(n10072), .A2(n10113), .B1(n10071), .B2(n10108), .ZN(
        n10074) );
  NOR2_X1 U11127 ( .A1(n10074), .A2(n10073), .ZN(n10123) );
  AOI22_X1 U11128 ( .A1(n10121), .A2(n10075), .B1(n10123), .B2(n10119), .ZN(
        P2_U3399) );
  NOR2_X1 U11129 ( .A1(n10076), .A2(n10108), .ZN(n10078) );
  AOI211_X1 U11130 ( .C1(n10080), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10125) );
  AOI22_X1 U11131 ( .A1(n10121), .A2(n5078), .B1(n10125), .B2(n10119), .ZN(
        P2_U3402) );
  INV_X1 U11132 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U11133 ( .A1(n10083), .A2(n10082), .B1(n10118), .B2(n10081), .ZN(
        n10084) );
  AND2_X1 U11134 ( .A1(n10085), .A2(n10084), .ZN(n10126) );
  AOI22_X1 U11135 ( .A1(n10121), .A2(n10086), .B1(n10126), .B2(n10119), .ZN(
        P2_U3405) );
  INV_X1 U11136 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10092) );
  INV_X1 U11137 ( .A(n10087), .ZN(n10091) );
  OAI22_X1 U11138 ( .A1(n10089), .A2(n10113), .B1(n10088), .B2(n10108), .ZN(
        n10090) );
  NOR2_X1 U11139 ( .A1(n10091), .A2(n10090), .ZN(n10127) );
  AOI22_X1 U11140 ( .A1(n10121), .A2(n10092), .B1(n10127), .B2(n10119), .ZN(
        P2_U3408) );
  INV_X1 U11141 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10097) );
  OAI22_X1 U11142 ( .A1(n10094), .A2(n10102), .B1(n10093), .B2(n10108), .ZN(
        n10095) );
  NOR2_X1 U11143 ( .A1(n10096), .A2(n10095), .ZN(n10128) );
  AOI22_X1 U11144 ( .A1(n10121), .A2(n10097), .B1(n10128), .B2(n10119), .ZN(
        P2_U3411) );
  OAI22_X1 U11145 ( .A1(n10099), .A2(n10113), .B1(n10098), .B2(n10108), .ZN(
        n10100) );
  NOR2_X1 U11146 ( .A1(n10101), .A2(n10100), .ZN(n10130) );
  AOI22_X1 U11147 ( .A1(n10121), .A2(n5138), .B1(n10130), .B2(n10119), .ZN(
        P2_U3414) );
  INV_X1 U11148 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10107) );
  NOR2_X1 U11149 ( .A1(n10103), .A2(n10102), .ZN(n10105) );
  AOI211_X1 U11150 ( .C1(n10118), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        n10131) );
  AOI22_X1 U11151 ( .A1(n10121), .A2(n10107), .B1(n10131), .B2(n10119), .ZN(
        P2_U3417) );
  OAI22_X1 U11152 ( .A1(n10110), .A2(n10113), .B1(n10109), .B2(n10108), .ZN(
        n10111) );
  NOR2_X1 U11153 ( .A1(n10112), .A2(n10111), .ZN(n10132) );
  AOI22_X1 U11154 ( .A1(n10121), .A2(n5168), .B1(n10132), .B2(n10119), .ZN(
        P2_U3420) );
  INV_X1 U11155 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U11156 ( .A1(n10114), .A2(n10113), .ZN(n10116) );
  AOI211_X1 U11157 ( .C1(n10118), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10134) );
  AOI22_X1 U11158 ( .A1(n10121), .A2(n10120), .B1(n10134), .B2(n10119), .ZN(
        P2_U3423) );
  AOI22_X1 U11159 ( .A1(n10135), .A2(n10122), .B1(n6553), .B2(n10133), .ZN(
        P2_U3460) );
  AOI22_X1 U11160 ( .A1(n10135), .A2(n10123), .B1(n5054), .B2(n10133), .ZN(
        P2_U3462) );
  AOI22_X1 U11161 ( .A1(n10135), .A2(n10125), .B1(n10124), .B2(n10133), .ZN(
        P2_U3463) );
  AOI22_X1 U11162 ( .A1(n10135), .A2(n10126), .B1(n4569), .B2(n10133), .ZN(
        P2_U3464) );
  AOI22_X1 U11163 ( .A1(n10135), .A2(n10127), .B1(n6588), .B2(n10133), .ZN(
        P2_U3465) );
  AOI22_X1 U11164 ( .A1(n10135), .A2(n10128), .B1(n4576), .B2(n10133), .ZN(
        P2_U3466) );
  AOI22_X1 U11165 ( .A1(n10135), .A2(n10130), .B1(n10129), .B2(n10133), .ZN(
        P2_U3467) );
  AOI22_X1 U11166 ( .A1(n10135), .A2(n10131), .B1(n6931), .B2(n10133), .ZN(
        P2_U3468) );
  AOI22_X1 U11167 ( .A1(n10135), .A2(n10132), .B1(n7495), .B2(n10133), .ZN(
        P2_U3469) );
  AOI22_X1 U11168 ( .A1(n10135), .A2(n10134), .B1(n7505), .B2(n10133), .ZN(
        P2_U3470) );
  NOR2_X1 U11169 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  XOR2_X1 U11170 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10138), .Z(ADD_1068_U5) );
  XOR2_X1 U11171 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11172 ( .A1(n10140), .A2(n10139), .ZN(n10141) );
  XOR2_X1 U11173 ( .A(n10141), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11174 ( .A(n10143), .B(n10142), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11175 ( .A(n10145), .B(n10144), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11176 ( .A(n10147), .B(n10146), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11177 ( .A(n10149), .B(n10148), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11178 ( .A(n10151), .B(n10150), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11179 ( .A(n10153), .B(n10152), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11180 ( .A(n10155), .B(n10154), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11181 ( .A(n10157), .B(n10156), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11182 ( .A(n10159), .B(n10158), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11183 ( .A(n10161), .B(n10160), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11184 ( .A(n10163), .B(n10162), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11185 ( .A(n10165), .B(n10164), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11186 ( .A(n10167), .B(n10166), .ZN(ADD_1068_U48) );
  XOR2_X1 U11187 ( .A(n10169), .B(n10168), .Z(ADD_1068_U54) );
  XOR2_X1 U11188 ( .A(n10171), .B(n10170), .Z(ADD_1068_U53) );
  XNOR2_X1 U11189 ( .A(n10173), .B(n10172), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4818 ( .A(n6101), .Z(n6305) );
endmodule

