

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579;

  NOR2_X1 U3657 ( .A1(n6409), .A2(n3695), .ZN(n6403) );
  OR2_X1 U3658 ( .A1(n4703), .A2(n4702), .ZN(n6170) );
  OR2_X1 U3659 ( .A1(n6317), .A2(n6316), .ZN(n6319) );
  INV_X4 U3660 ( .A(n3633), .ZN(n6426) );
  OAI21_X1 U3661 ( .B1(n5084), .B2(n4330), .A(n4157), .ZN(n4935) );
  INV_X1 U3662 ( .A(n4086), .ZN(n4056) );
  CLKBUF_X2 U3663 ( .A(n3906), .Z(n4005) );
  CLKBUF_X2 U3664 ( .A(n3895), .Z(n4719) );
  CLKBUF_X2 U3665 ( .A(n3868), .Z(n4720) );
  CLKBUF_X2 U3666 ( .A(n3941), .Z(n4482) );
  BUF_X1 U3667 ( .A(n3964), .Z(n4665) );
  NAND4_X2 U3668 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3970)
         );
  AND4_X1 U3669 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3849)
         );
  AND2_X1 U3670 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5050) );
  INV_X1 U3672 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U3673 ( .A1(n3970), .A2(n3974), .ZN(n4754) );
  BUF_X1 U3674 ( .A(n4769), .Z(n3631) );
  OAI21_X1 U3675 ( .B1(n5066), .B2(STATE2_REG_0__SCAN_IN), .A(n4116), .ZN(
        n4117) );
  INV_X1 U3676 ( .A(n4741), .ZN(n4870) );
  XNOR2_X1 U3677 ( .A(n4616), .B(n4235), .ZN(n4607) );
  INV_X1 U3678 ( .A(n4856), .ZN(n4947) );
  NAND2_X1 U3679 ( .A1(n4616), .A2(n4619), .ZN(n4628) );
  OR2_X1 U3680 ( .A1(n4070), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4062) );
  AND4_X1 U3681 ( .A1(n3830), .A2(n3828), .A3(n3831), .A4(n3829), .ZN(n3965)
         );
  NAND2_X1 U3682 ( .A1(n3628), .A2(n3649), .ZN(n6304) );
  NAND2_X1 U3683 ( .A1(n6219), .A2(n6220), .ZN(n6209) );
  NAND2_X1 U3684 ( .A1(n3956), .A2(n3636), .ZN(n4979) );
  INV_X1 U3685 ( .A(n4763), .ZN(n5302) );
  INV_X1 U3686 ( .A(n3628), .ZN(n6059) );
  INV_X1 U3687 ( .A(n5109), .ZN(n3929) );
  XNOR2_X1 U3688 ( .A(n6353), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6486)
         );
  OAI22_X1 U3689 ( .A1(n6403), .A2(n6386), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6396), .ZN(n6387) );
  OR2_X1 U3690 ( .A1(n3999), .A2(n5038), .ZN(n3623) );
  NAND2_X1 U3691 ( .A1(n4118), .A2(n4117), .ZN(n4145) );
  INV_X1 U3692 ( .A(n3626), .ZN(n6424) );
  OAI21_X2 U3694 ( .B1(n6439), .B2(n6442), .A(n6440), .ZN(n6431) );
  NAND2_X2 U3695 ( .A1(n4636), .A2(n6091), .ZN(n6439) );
  XNOR2_X2 U3696 ( .A(n4614), .B(n6890), .ZN(n5617) );
  NAND2_X2 U3698 ( .A1(n5031), .A2(n4104), .ZN(n5066) );
  AND2_X1 U3700 ( .A1(n6310), .A2(n6300), .ZN(n6756) );
  NAND2_X1 U3701 ( .A1(n5631), .A2(n5630), .ZN(n6048) );
  NAND2_X1 U3702 ( .A1(n4013), .A2(n4012), .ZN(n4083) );
  BUF_X2 U3703 ( .A(n4769), .Z(n3630) );
  INV_X2 U3704 ( .A(n3970), .ZN(n4750) );
  AND2_X2 U3705 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6146)
         );
  AND2_X2 U3706 ( .A1(n3651), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5053)
         );
  INV_X2 U3707 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3887) );
  INV_X1 U3708 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U3709 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  OAI21_X1 U3710 ( .B1(n6816), .B2(n6383), .A(n6382), .ZN(n6411) );
  NAND2_X1 U3711 ( .A1(n4551), .A2(n4886), .ZN(n6119) );
  NAND2_X1 U3712 ( .A1(n6381), .A2(n6817), .ZN(n6816) );
  OAI21_X1 U3713 ( .B1(n3626), .B2(n3643), .A(n3676), .ZN(n6374) );
  AND2_X2 U3714 ( .A1(n6280), .A2(n3678), .ZN(n6219) );
  AND2_X1 U3715 ( .A1(n4882), .A2(n3647), .ZN(n4883) );
  OAI21_X1 U3716 ( .B1(n6023), .B2(n6024), .A(n4630), .ZN(n4633) );
  NAND2_X1 U3717 ( .A1(n6015), .A2(n6014), .ZN(n6023) );
  NAND2_X1 U3718 ( .A1(n4627), .A2(n4626), .ZN(n6015) );
  NAND2_X1 U3719 ( .A1(n6175), .A2(n4947), .ZN(n6173) );
  AND2_X2 U3720 ( .A1(n6058), .A2(n6060), .ZN(n3628) );
  NAND2_X1 U3721 ( .A1(n4337), .A2(n4336), .ZN(n6058) );
  NAND2_X1 U3722 ( .A1(n6123), .A2(n4880), .ZN(n6175) );
  CLKBUF_X1 U3723 ( .A(n6250), .Z(n6276) );
  AND2_X1 U3724 ( .A1(n5558), .A2(n3666), .ZN(n3671) );
  BUF_X4 U3725 ( .A(n4628), .Z(n3633) );
  NAND2_X1 U3726 ( .A1(n6756), .A2(n6755), .ZN(n6758) );
  AND2_X1 U3727 ( .A1(n4913), .A2(n4935), .ZN(n5369) );
  NAND2_X1 U3728 ( .A1(n4125), .A2(n4124), .ZN(n4913) );
  NAND2_X1 U3729 ( .A1(n4565), .A2(n4977), .ZN(n6774) );
  NAND2_X1 U3730 ( .A1(n4994), .A2(n4121), .ZN(n4915) );
  AOI21_X1 U3731 ( .B1(n5087), .B2(n4694), .A(n4573), .ZN(n6775) );
  NAND2_X1 U3732 ( .A1(n4564), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4977)
         );
  NAND2_X1 U3733 ( .A1(n4144), .A2(n3692), .ZN(n4196) );
  INV_X1 U3734 ( .A(n4145), .ZN(n4144) );
  NAND2_X1 U3735 ( .A1(n4807), .A2(n4806), .ZN(n6062) );
  CLKBUF_X2 U3736 ( .A(n5083), .Z(n3632) );
  AND2_X1 U3737 ( .A1(n4146), .A2(n3693), .ZN(n3692) );
  INV_X1 U3738 ( .A(n6048), .ZN(n4807) );
  CLKBUF_X1 U3739 ( .A(n5037), .Z(n7359) );
  OAI21_X1 U3740 ( .B1(n4087), .B2(n4086), .A(n4085), .ZN(n4118) );
  AOI21_X1 U3741 ( .B1(n4055), .B2(n4064), .A(n4617), .ZN(n4086) );
  NAND2_X1 U3742 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  AND2_X1 U3743 ( .A1(n4092), .A2(n4091), .ZN(n4100) );
  INV_X1 U3744 ( .A(n4089), .ZN(n3624) );
  NAND2_X1 U3745 ( .A1(n4781), .A2(n4780), .ZN(n5252) );
  NAND3_X1 U3746 ( .A1(n4768), .A2(n4762), .A3(n3658), .ZN(n4938) );
  NAND2_X1 U3747 ( .A1(n4982), .A2(n5302), .ZN(n3658) );
  NOR2_X1 U3748 ( .A1(n6046), .A2(n6047), .ZN(n4806) );
  CLKBUF_X1 U3749 ( .A(n4921), .Z(n5040) );
  NAND2_X1 U3750 ( .A1(n4757), .A2(n4756), .ZN(n4760) );
  INV_X1 U3751 ( .A(n4170), .ZN(n3693) );
  NOR2_X1 U3752 ( .A1(n4051), .A2(n7224), .ZN(n4617) );
  OR2_X1 U3753 ( .A1(n4011), .A2(n4010), .ZN(n4553) );
  OR2_X1 U3754 ( .A1(n4047), .A2(n4046), .ZN(n4561) );
  OR2_X1 U3755 ( .A1(n4028), .A2(n4027), .ZN(n4620) );
  OR2_X1 U3756 ( .A1(n4015), .A2(n7224), .ZN(n4664) );
  AND2_X2 U3757 ( .A1(n3970), .A2(n4665), .ZN(n4694) );
  INV_X2 U3758 ( .A(n4754), .ZN(n4765) );
  OR2_X1 U3759 ( .A1(n3969), .A2(n4015), .ZN(n4943) );
  NAND2_X1 U3760 ( .A1(n5109), .A2(n4750), .ZN(n6003) );
  AND2_X1 U3761 ( .A1(n4015), .A2(n4014), .ZN(n4686) );
  NAND4_X2 U3762 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3964)
         );
  NAND2_X1 U3763 ( .A1(n3639), .A2(n3635), .ZN(n3974) );
  AND4_X2 U3764 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n4068)
         );
  INV_X2 U3765 ( .A(n3965), .ZN(n3625) );
  NAND4_X2 U3766 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3962)
         );
  AND4_X1 U3767 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  NAND2_X2 U3768 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6829), .ZN(n6713) );
  AND4_X1 U3769 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3928)
         );
  AND4_X1 U3770 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3831)
         );
  AND4_X1 U3771 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(n3953)
         );
  AND4_X1 U3772 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3886)
         );
  AND4_X1 U3773 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3851)
         );
  AND4_X1 U3774 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3861)
         );
  INV_X2 U3775 ( .A(n6791), .ZN(n6818) );
  AND4_X1 U3776 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3830)
         );
  AND4_X1 U3777 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3926)
         );
  AND4_X1 U3778 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3811)
         );
  AND4_X1 U3779 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3885)
         );
  AND4_X1 U3780 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3927)
         );
  AND4_X1 U3781 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  AND4_X1 U3782 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3809)
         );
  AND4_X1 U3783 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AND4_X1 U3784 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  AND4_X1 U3785 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3884)
         );
  AND4_X1 U3786 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3952)
         );
  NAND2_X2 U3787 ( .A1(n6829), .A2(n6830), .ZN(n6719) );
  AND4_X1 U3788 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3848)
         );
  AND4_X1 U3789 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  AND4_X1 U3790 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  AND4_X1 U3791 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3883)
         );
  AND4_X1 U3792 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3954)
         );
  AND4_X1 U3793 ( .A1(n3799), .A2(n3798), .A3(n3797), .A4(n3796), .ZN(n3810)
         );
  BUF_X2 U3794 ( .A(n3894), .Z(n4718) );
  BUF_X2 U3795 ( .A(n3867), .Z(n4728) );
  BUF_X2 U3796 ( .A(n4016), .Z(n4017) );
  BUF_X2 U3797 ( .A(n3878), .Z(n4443) );
  BUF_X2 U3798 ( .A(n3905), .Z(n4726) );
  BUF_X2 U3799 ( .A(n3873), .Z(n4465) );
  AND2_X2 U3800 ( .A1(n5054), .A2(n6146), .ZN(n3919) );
  AND2_X2 U3801 ( .A1(n5053), .A2(n6146), .ZN(n3936) );
  INV_X2 U3802 ( .A(n7246), .ZN(n6829) );
  AND2_X2 U3803 ( .A1(n5054), .A2(n5078), .ZN(n3868) );
  BUF_X2 U3804 ( .A(n3931), .Z(n4727) );
  AND2_X2 U3805 ( .A1(n5053), .A2(n6147), .ZN(n3905) );
  AND2_X2 U3806 ( .A1(n5054), .A2(n5049), .ZN(n3941) );
  AND2_X2 U3807 ( .A1(n6146), .A2(n5048), .ZN(n3867) );
  AND2_X2 U3808 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5049) );
  NOR2_X2 U3809 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5078) );
  INV_X4 U3810 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3707) );
  NOR2_X2 U3811 ( .A1(n6431), .A2(n3627), .ZN(n3626) );
  AND2_X1 U3812 ( .A1(n3633), .A2(n6606), .ZN(n3627) );
  NAND2_X1 U3813 ( .A1(n3632), .A2(n4694), .ZN(n3675) );
  XNOR2_X1 U3814 ( .A(n4196), .B(n4207), .ZN(n4589) );
  NAND2_X1 U3815 ( .A1(n3663), .A2(n3661), .ZN(n5237) );
  OR2_X1 U3816 ( .A1(n6774), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4575)
         );
  NAND2_X1 U3817 ( .A1(n4068), .A2(n3964), .ZN(n4944) );
  NAND2_X2 U3818 ( .A1(n3860), .A2(n3861), .ZN(n5364) );
  AOI21_X1 U3819 ( .B1(n4552), .B2(n4551), .A(n4746), .ZN(n6198) );
  XNOR2_X1 U3820 ( .A(n4088), .B(n4089), .ZN(n5089) );
  NAND2_X1 U3821 ( .A1(n3981), .A2(n4091), .ZN(n4088) );
  OAI21_X1 U3822 ( .B1(n4585), .B2(n4330), .A(n4183), .ZN(n5370) );
  NOR2_X2 U3823 ( .A1(n6411), .A2(n6410), .ZN(n6409) );
  INV_X4 U3824 ( .A(n3962), .ZN(n3963) );
  AND2_X4 U3825 ( .A1(n4057), .A2(n5364), .ZN(n3966) );
  INV_X2 U3826 ( .A(n4068), .ZN(n4057) );
  NOR2_X2 U3827 ( .A1(n6746), .A2(n5543), .ZN(n5631) );
  AND2_X2 U3828 ( .A1(n6366), .A2(n4644), .ZN(n6357) );
  AND2_X4 U3829 ( .A1(n3712), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5054)
         );
  AND2_X1 U3830 ( .A1(n5054), .A2(n5049), .ZN(n3629) );
  NOR2_X4 U3831 ( .A1(n5247), .A2(n5251), .ZN(n5249) );
  OAI22_X2 U3832 ( .A1(n4648), .A2(n4861), .B1(n6426), .B2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4649) );
  OAI21_X2 U3835 ( .B1(n6374), .B2(n6375), .A(n4643), .ZN(n6366) );
  XNOR2_X2 U3836 ( .A(n5623), .B(n4334), .ZN(n6044) );
  AND2_X2 U3837 ( .A1(n6221), .A2(n6222), .ZN(n6223) );
  NOR3_X4 U3838 ( .A1(n6250), .A2(n6252), .A3(n6235), .ZN(n6222) );
  INV_X4 U3839 ( .A(n4765), .ZN(n4856) );
  NOR2_X2 U3840 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  NAND2_X1 U3841 ( .A1(n3929), .A2(n4969), .ZN(n4769) );
  NOR2_X4 U3842 ( .A1(n6304), .A2(n6306), .ZN(n6297) );
  NOR2_X4 U3843 ( .A1(n6291), .A2(n6408), .ZN(n6280) );
  OR2_X1 U3844 ( .A1(n4234), .A2(n5455), .ZN(n4195) );
  NOR2_X1 U3845 ( .A1(n5109), .A2(n7224), .ZN(n4014) );
  CLKBUF_X1 U3846 ( .A(n4057), .Z(n4749) );
  NAND2_X1 U3847 ( .A1(n4885), .A2(n3691), .ZN(n3690) );
  INV_X1 U3848 ( .A(n6211), .ZN(n3691) );
  NOR2_X1 U3849 ( .A1(n4749), .A2(n3887), .ZN(n4366) );
  INV_X1 U3850 ( .A(n4223), .ZN(n4221) );
  AND2_X1 U3851 ( .A1(n4990), .A2(n4985), .ZN(n6093) );
  INV_X1 U3852 ( .A(n4694), .ZN(n4747) );
  CLKBUF_X1 U3853 ( .A(n4901), .Z(n6164) );
  AND2_X1 U3854 ( .A1(n3887), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4869) );
  NAND2_X1 U3855 ( .A1(n3689), .A2(n3964), .ZN(n3688) );
  NAND2_X1 U3856 ( .A1(n3625), .A2(n3963), .ZN(n3689) );
  NAND2_X1 U3857 ( .A1(n3625), .A2(n3687), .ZN(n3686) );
  AOI21_X1 U3858 ( .B1(n4944), .B2(n3974), .A(n3970), .ZN(n3988) );
  AND2_X1 U3859 ( .A1(n4169), .A2(n4168), .ZN(n4170) );
  AND2_X1 U3860 ( .A1(n4220), .A2(n4219), .ZN(n4223) );
  OR2_X1 U3861 ( .A1(n4234), .A2(n5431), .ZN(n4220) );
  NAND2_X1 U3862 ( .A1(n5109), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4105) );
  NAND2_X1 U3863 ( .A1(n4105), .A2(n4664), .ZN(n4700) );
  AND2_X1 U3864 ( .A1(n6244), .A2(n3681), .ZN(n3680) );
  NOR2_X1 U3865 ( .A1(n6275), .A2(n3682), .ZN(n3681) );
  INV_X1 U3866 ( .A(n6281), .ZN(n3682) );
  INV_X1 U3867 ( .A(n4366), .ZN(n4330) );
  INV_X1 U3868 ( .A(n4841), .ZN(n4848) );
  NAND2_X1 U3869 ( .A1(n5302), .A2(n4856), .ZN(n4841) );
  AOI21_X1 U3870 ( .B1(n7216), .B2(n7211), .A(n6108), .ZN(n5097) );
  OR2_X1 U3871 ( .A1(n7169), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4707) );
  OR2_X1 U3872 ( .A1(n7139), .A2(n7075), .ZN(n7074) );
  OR2_X1 U3873 ( .A1(n4874), .A2(n6346), .ZN(n4875) );
  OR2_X1 U3874 ( .A1(n4534), .A2(n4533), .ZN(n4543) );
  OAI21_X1 U3875 ( .B1(n6377), .B2(n5289), .A(n4524), .ZN(n6234) );
  AOI21_X1 U3876 ( .B1(n4598), .B2(n4366), .A(n4232), .ZN(n5251) );
  CLKBUF_X1 U3877 ( .A(n5249), .Z(n5250) );
  NAND2_X1 U3878 ( .A1(n4205), .A2(n4204), .ZN(n5000) );
  AOI21_X1 U3879 ( .B1(n6118), .B2(n4069), .A(n3887), .ZN(n4911) );
  NAND2_X1 U3880 ( .A1(n4911), .A2(n4910), .ZN(n4909) );
  INV_X1 U3881 ( .A(n4949), .ZN(n6176) );
  NAND2_X1 U3882 ( .A1(n3657), .A2(n3656), .ZN(n6568) );
  INV_X1 U3883 ( .A(n6289), .ZN(n3656) );
  INV_X1 U3884 ( .A(n6758), .ZN(n3657) );
  NOR2_X2 U3885 ( .A1(n6319), .A2(n6308), .ZN(n6310) );
  NOR2_X2 U3886 ( .A1(n5252), .A2(n5253), .ZN(n5324) );
  NAND2_X1 U3887 ( .A1(n6786), .A2(n4588), .ZN(n3663) );
  INV_X1 U3888 ( .A(n6786), .ZN(n3665) );
  INV_X1 U3889 ( .A(n4917), .ZN(n4768) );
  CLKBUF_X1 U3890 ( .A(n4903), .Z(n4904) );
  NAND2_X1 U3891 ( .A1(n3957), .A2(n3966), .ZN(n4972) );
  INV_X1 U3892 ( .A(n4979), .ZN(n3957) );
  AND2_X1 U3893 ( .A1(n4968), .A2(n7221), .ZN(n4990) );
  AND2_X1 U3894 ( .A1(n3631), .A2(n4856), .ZN(n4949) );
  OR2_X1 U3895 ( .A1(n4234), .A2(n5155), .ZN(n4054) );
  NAND2_X1 U3896 ( .A1(n3959), .A2(n4750), .ZN(n5039) );
  NOR2_X2 U3897 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5097), .ZN(n5413) );
  INV_X1 U3898 ( .A(n6118), .ZN(n7371) );
  AND2_X1 U3899 ( .A1(n6170), .A2(n4971), .ZN(n7194) );
  OR2_X1 U3900 ( .A1(n6838), .A2(n5291), .ZN(n6941) );
  OR2_X1 U3901 ( .A1(n6908), .A2(n5290), .ZN(n5291) );
  NAND2_X1 U3902 ( .A1(n6773), .A2(n6141), .ZN(n6320) );
  AND2_X1 U3903 ( .A1(n4753), .A2(n7221), .ZN(n6773) );
  INV_X1 U3904 ( .A(n5364), .ZN(n6141) );
  INV_X1 U3905 ( .A(n6198), .ZN(n4716) );
  OR2_X1 U3906 ( .A1(n4884), .A2(n4885), .ZN(n4886) );
  INV_X1 U3907 ( .A(n6822), .ZN(n6801) );
  XNOR2_X1 U3908 ( .A(n4867), .B(n6104), .ZN(n6485) );
  NAND2_X1 U3909 ( .A1(n5327), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U3910 ( .A1(n3968), .A2(n5109), .ZN(n3996) );
  OAI21_X1 U3911 ( .B1(n4068), .B2(n3964), .A(n5364), .ZN(n3969) );
  NAND2_X1 U3912 ( .A1(n4654), .A2(n4653), .ZN(n4684) );
  INV_X1 U3913 ( .A(n4682), .ZN(n4653) );
  INV_X1 U3914 ( .A(n4683), .ZN(n4654) );
  XNOR2_X1 U3915 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4659) );
  AOI21_X1 U3916 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n7361), .A(n4656), 
        .ZN(n4657) );
  AND2_X1 U3917 ( .A1(n4660), .A2(n4659), .ZN(n4656) );
  OR2_X1 U3918 ( .A1(n4218), .A2(n4217), .ZN(n4609) );
  OR2_X1 U3919 ( .A1(n4193), .A2(n4192), .ZN(n4600) );
  OR2_X1 U3920 ( .A1(n4167), .A2(n4166), .ZN(n4590) );
  AOI21_X1 U3921 ( .B1(n3986), .B2(n3974), .A(n4750), .ZN(n3987) );
  AOI22_X1 U3922 ( .A1(n3895), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3896) );
  AND2_X1 U3923 ( .A1(n4686), .A2(n4694), .ZN(n4701) );
  NAND2_X1 U3924 ( .A1(n7161), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4540) );
  AND2_X1 U3925 ( .A1(n4177), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4197)
         );
  AND3_X1 U3926 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .A3(PHYADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4149) );
  OR2_X1 U3927 ( .A1(n4141), .A2(n4140), .ZN(n4578) );
  NAND2_X1 U3928 ( .A1(n3974), .A2(n5109), .ZN(n4955) );
  INV_X1 U3929 ( .A(n4686), .ZN(n4234) );
  AND2_X2 U3930 ( .A1(n5050), .A2(n5049), .ZN(n3946) );
  AND2_X1 U3931 ( .A1(n4095), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4126)
         );
  INV_X1 U3932 ( .A(n4554), .ZN(n4569) );
  NAND2_X1 U3933 ( .A1(n4357), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4374)
         );
  INV_X1 U3934 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U3935 ( .A1(n4131), .A2(n4130), .ZN(n5029) );
  AND2_X1 U3936 ( .A1(n4834), .A2(n4833), .ZN(n6283) );
  AND2_X1 U3937 ( .A1(n4785), .A2(n4784), .ZN(n5253) );
  NAND2_X1 U3938 ( .A1(n5016), .A2(n5015), .ZN(n5361) );
  OR2_X1 U3939 ( .A1(n5039), .A2(n5014), .ZN(n5015) );
  AND2_X1 U3940 ( .A1(n4924), .A2(n6006), .ZN(n6652) );
  AOI21_X1 U3941 ( .B1(n6348), .B2(n4550), .A(n4745), .ZN(n4868) );
  OR2_X1 U3942 ( .A1(n3705), .A2(n3704), .ZN(n4874) );
  AOI22_X1 U3943 ( .A1(n6124), .A2(n4550), .B1(n4549), .B2(n4548), .ZN(n4885)
         );
  AOI22_X1 U3944 ( .A1(n6226), .A2(n4550), .B1(n4532), .B2(n4531), .ZN(n6220)
         );
  NOR2_X1 U3945 ( .A1(n4510), .A2(n6247), .ZN(n4515) );
  AND2_X1 U3946 ( .A1(n3680), .A2(n3679), .ZN(n3678) );
  INV_X1 U3947 ( .A(n6234), .ZN(n3679) );
  NAND2_X1 U3948 ( .A1(n4481), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4500)
         );
  NOR2_X1 U3949 ( .A1(n4419), .A2(n3701), .ZN(n4423) );
  AND2_X1 U3950 ( .A1(n4423), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4442)
         );
  AND2_X1 U3951 ( .A1(n4441), .A2(n6299), .ZN(n3683) );
  NOR2_X1 U3952 ( .A1(n4374), .A2(n3700), .ZN(n4389) );
  INV_X1 U3953 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U3954 ( .A1(n4389), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4419)
         );
  CLKBUF_X1 U3955 ( .A(n6304), .Z(n6305) );
  NAND2_X1 U3956 ( .A1(n4331), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4342)
         );
  NOR2_X1 U3957 ( .A1(n4272), .A2(n5551), .ZN(n4298) );
  NAND2_X1 U3958 ( .A1(n4256), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4272)
         );
  NOR2_X1 U3959 ( .A1(n4251), .A2(n3699), .ZN(n4256) );
  NAND2_X1 U3960 ( .A1(n4236), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4251)
         );
  AND2_X1 U3961 ( .A1(n4197), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4236)
         );
  OAI21_X1 U3962 ( .B1(n5137), .B2(n4330), .A(n4120), .ZN(n4916) );
  NAND2_X1 U3963 ( .A1(n4061), .A2(n4060), .ZN(n4996) );
  NAND2_X1 U3964 ( .A1(n6357), .A2(n4645), .ZN(n4888) );
  INV_X1 U3965 ( .A(n3677), .ZN(n3676) );
  OAI21_X1 U3966 ( .B1(n3634), .B2(n3643), .A(n4642), .ZN(n3677) );
  NOR2_X2 U3967 ( .A1(n6566), .A2(n6283), .ZN(n6282) );
  AND2_X1 U3968 ( .A1(n4828), .A2(n4827), .ZN(n6289) );
  AND2_X1 U3969 ( .A1(n4824), .A2(n4823), .ZN(n6755) );
  AND2_X1 U3970 ( .A1(n4816), .A2(n4815), .ZN(n6316) );
  AND2_X1 U3971 ( .A1(n4813), .A2(n4812), .ZN(n6259) );
  AND2_X1 U3972 ( .A1(n4810), .A2(n4809), .ZN(n6061) );
  NAND2_X1 U3973 ( .A1(n6082), .A2(n6083), .ZN(n3673) );
  AND2_X1 U3974 ( .A1(n4805), .A2(n4804), .ZN(n6047) );
  NOR2_X1 U3975 ( .A1(n4618), .A2(n4747), .ZN(n4619) );
  NAND2_X1 U3976 ( .A1(n3671), .A2(n3672), .ZN(n3668) );
  NOR2_X1 U3977 ( .A1(n6921), .A2(n6093), .ZN(n6589) );
  NAND2_X1 U3978 ( .A1(n3653), .A2(n3652), .ZN(n6746) );
  INV_X1 U3979 ( .A(n6749), .ZN(n3652) );
  INV_X1 U3980 ( .A(n6748), .ZN(n3653) );
  NAND2_X1 U3981 ( .A1(n5318), .A2(n5319), .ZN(n6748) );
  INV_X1 U3982 ( .A(n5003), .ZN(n4780) );
  NAND2_X1 U3983 ( .A1(n4576), .A2(n4575), .ZN(n6780) );
  NOR2_X2 U3984 ( .A1(n4938), .A2(n4937), .ZN(n6768) );
  AND2_X1 U3985 ( .A1(n4940), .A2(n4958), .ZN(n6166) );
  OR2_X1 U3986 ( .A1(n6589), .A2(n5241), .ZN(n6473) );
  AND2_X1 U3987 ( .A1(n4988), .A2(n4987), .ZN(n6587) );
  AND2_X1 U3988 ( .A1(n4559), .A2(n4560), .ZN(n3674) );
  CLKBUF_X1 U3989 ( .A(n5089), .Z(n5090) );
  NAND2_X1 U3990 ( .A1(n4099), .A2(n4098), .ZN(n4101) );
  NAND2_X2 U3991 ( .A1(n4119), .A2(n4145), .ZN(n5137) );
  OR2_X1 U3992 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  AND2_X2 U3993 ( .A1(n3650), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6147)
         );
  AND2_X1 U3994 ( .A1(n3991), .A2(n4665), .ZN(n7161) );
  INV_X1 U3995 ( .A(n6170), .ZN(n6004) );
  AND2_X1 U3996 ( .A1(n5137), .A2(n3632), .ZN(n5332) );
  AND2_X1 U3997 ( .A1(n5158), .A2(n5258), .ZN(n7401) );
  OR2_X1 U3998 ( .A1(n7368), .A2(n7371), .ZN(n7373) );
  NOR2_X1 U3999 ( .A1(n7359), .A2(n7426), .ZN(n5336) );
  CLKBUF_X2 U4000 ( .A(n3965), .Z(n5403) );
  OR2_X1 U4001 ( .A1(n7213), .A2(n5097), .ZN(n5410) );
  INV_X1 U4002 ( .A(n4126), .ZN(n5093) );
  NAND2_X1 U4003 ( .A1(n7214), .A2(n3887), .ZN(n7426) );
  NAND2_X1 U4004 ( .A1(n3887), .A2(n7413), .ZN(n5289) );
  INV_X1 U4005 ( .A(n7249), .ZN(n5286) );
  CLKBUF_X1 U4006 ( .A(n4569), .Z(n4570) );
  NOR2_X1 U4007 ( .A1(n5304), .A2(n5299), .ZN(n7139) );
  AND2_X1 U4008 ( .A1(n6941), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7144) );
  AND2_X1 U4009 ( .A1(n5295), .A2(n5294), .ZN(n7133) );
  NAND2_X1 U4010 ( .A1(n3658), .A2(n4762), .ZN(n4918) );
  INV_X1 U4011 ( .A(n6320), .ZN(n6769) );
  INV_X1 U4012 ( .A(n6142), .ZN(n7437) );
  AND2_X1 U4013 ( .A1(n6142), .A2(n5366), .ZN(n7438) );
  NOR2_X2 U4015 ( .A1(n7434), .A2(n7438), .ZN(n6343) );
  NAND2_X1 U4016 ( .A1(n7249), .A2(n5362), .ZN(n7329) );
  CLKBUF_X2 U4017 ( .A(n7327), .Z(n7330) );
  XNOR2_X1 U4018 ( .A(n4746), .B(n4868), .ZN(n6356) );
  INV_X1 U4020 ( .A(n6174), .ZN(n3654) );
  NAND2_X1 U4021 ( .A1(n6173), .A2(n3697), .ZN(n3655) );
  NAND2_X1 U4022 ( .A1(n6357), .A2(n3633), .ZN(n6358) );
  OR3_X1 U4023 ( .A1(n6357), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n3633), 
        .ZN(n6359) );
  OR2_X1 U4024 ( .A1(n6571), .A2(n6476), .ZN(n6551) );
  CLKBUF_X1 U4025 ( .A(n6431), .Z(n6433) );
  INV_X1 U4026 ( .A(n6870), .ZN(n6471) );
  NAND2_X1 U4027 ( .A1(n5616), .A2(n5617), .ZN(n3670) );
  NAND2_X1 U4028 ( .A1(n6787), .A2(n4588), .ZN(n5239) );
  NAND2_X1 U4029 ( .A1(n4990), .A2(n4981), .ZN(n6884) );
  INV_X1 U4030 ( .A(n6473), .ZN(n6866) );
  INV_X1 U4031 ( .A(n6467), .ZN(n6603) );
  AND2_X1 U4032 ( .A1(n4990), .A2(n4975), .ZN(n6915) );
  INV_X1 U4033 ( .A(n6884), .ZN(n6917) );
  NAND2_X2 U4034 ( .A1(n4067), .A2(n4066), .ZN(n6118) );
  INV_X1 U4035 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7412) );
  INV_X1 U4036 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U4037 ( .A1(n5082), .A2(n5081), .ZN(n6647) );
  INV_X1 U4038 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3651) );
  INV_X1 U4039 ( .A(n5428), .ZN(n5411) );
  INV_X1 U4040 ( .A(n5185), .ZN(n7558) );
  INV_X1 U4041 ( .A(n7373), .ZN(n7551) );
  INV_X1 U4042 ( .A(n7433), .ZN(n5600) );
  AND2_X1 U4043 ( .A1(n6818), .A2(DATAI_24_), .ZN(n7422) );
  INV_X1 U4044 ( .A(n7456), .ZN(n5592) );
  INV_X1 U4045 ( .A(n7472), .ZN(n5584) );
  AND2_X1 U4046 ( .A1(n6818), .A2(DATAI_26_), .ZN(n7468) );
  INV_X1 U4047 ( .A(n7488), .ZN(n5604) );
  AND2_X1 U4048 ( .A1(n6818), .A2(DATAI_27_), .ZN(n7484) );
  INV_X1 U4049 ( .A(n5511), .ZN(n7501) );
  INV_X1 U4050 ( .A(n7504), .ZN(n5580) );
  INV_X1 U4051 ( .A(n7520), .ZN(n5611) );
  AND2_X1 U4052 ( .A1(n6818), .A2(DATAI_29_), .ZN(n7517) );
  INV_X1 U4053 ( .A(n7536), .ZN(n5588) );
  AND2_X1 U4054 ( .A1(n6818), .A2(DATAI_30_), .ZN(n7532) );
  AND2_X1 U4055 ( .A1(n5099), .A2(n7371), .ZN(n5496) );
  INV_X1 U4056 ( .A(n7578), .ZN(n5596) );
  AND2_X1 U4057 ( .A1(n6818), .A2(DATAI_31_), .ZN(n7574) );
  AND2_X1 U4058 ( .A1(n4705), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7221) );
  INV_X1 U4059 ( .A(n7221), .ZN(n7206) );
  INV_X1 U4060 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U4061 ( .A1(STATE_REG_1__SCAN_IN), .A2(n7240), .ZN(n7246) );
  OR2_X1 U4062 ( .A1(n6500), .A2(n6320), .ZN(n4882) );
  OAI21_X1 U4063 ( .B1(n6485), .B2(n6804), .A(n3637), .ZN(U2955) );
  OAI21_X1 U4064 ( .B1(n6514), .B2(n6804), .A(n4892), .ZN(n4893) );
  AOI21_X1 U4065 ( .B1(n6801), .B2(n6124), .A(n4891), .ZN(n4892) );
  INV_X1 U4066 ( .A(n3862), .ZN(n4022) );
  NAND2_X1 U4067 ( .A1(n3665), .A2(n4586), .ZN(n6787) );
  NAND2_X1 U4068 ( .A1(n3633), .A2(n6457), .ZN(n3634) );
  NAND2_X1 U4069 ( .A1(n6280), .A2(n6281), .ZN(n6274) );
  NAND2_X1 U4070 ( .A1(n6280), .A2(n3680), .ZN(n6233) );
  NAND2_X1 U4071 ( .A1(n6297), .A2(n6299), .ZN(n6298) );
  AND4_X1 U4072 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3635)
         );
  AND3_X1 U4073 ( .A1(n4969), .A2(n5403), .A3(n3687), .ZN(n3636) );
  AND2_X1 U4074 ( .A1(n4879), .A2(n4878), .ZN(n3637) );
  INV_X1 U4075 ( .A(n3684), .ZN(n5315) );
  INV_X1 U4076 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3650) );
  AND2_X1 U4077 ( .A1(n6280), .A2(n3681), .ZN(n6243) );
  NAND2_X1 U4078 ( .A1(n3628), .A2(n4373), .ZN(n6256) );
  AND2_X1 U4079 ( .A1(n4969), .A2(n5109), .ZN(n3638) );
  AND4_X1 U4080 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3639)
         );
  AND2_X1 U4081 ( .A1(n6394), .A2(n4638), .ZN(n6381) );
  AND4_X1 U4082 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n5071), .ZN(n3640)
         );
  INV_X1 U4083 ( .A(n4588), .ZN(n3664) );
  AND2_X1 U4084 ( .A1(n4616), .A2(n4225), .ZN(n4598) );
  OR2_X1 U4085 ( .A1(n6209), .A2(n3690), .ZN(n4551) );
  INV_X1 U4086 ( .A(n3659), .ZN(n6251) );
  NOR2_X1 U4087 ( .A1(n6250), .A2(n6252), .ZN(n3659) );
  OR2_X1 U4088 ( .A1(n5109), .A2(n3970), .ZN(n4554) );
  AND2_X1 U4089 ( .A1(n6223), .A2(n6208), .ZN(n6120) );
  AND2_X1 U4090 ( .A1(n3696), .A2(n4635), .ZN(n3641) );
  INV_X1 U4091 ( .A(n4615), .ZN(n3672) );
  NOR2_X2 U4092 ( .A1(n7414), .A2(n6118), .ZN(n3642) );
  AND2_X1 U4093 ( .A1(n5541), .A2(n5627), .ZN(n5622) );
  NAND2_X1 U4094 ( .A1(n4641), .A2(n4638), .ZN(n3643) );
  NAND2_X1 U4095 ( .A1(n3673), .A2(n4635), .ZN(n6090) );
  NAND2_X1 U4096 ( .A1(n3670), .A2(n4615), .ZN(n5557) );
  OR2_X1 U4097 ( .A1(n4552), .A2(n3690), .ZN(n3644) );
  NAND2_X1 U4098 ( .A1(n5249), .A2(n5322), .ZN(n3684) );
  AND2_X1 U4099 ( .A1(n5627), .A2(n5625), .ZN(n3645) );
  AND2_X1 U4100 ( .A1(n4271), .A2(n5317), .ZN(n3646) );
  INV_X1 U4101 ( .A(n6804), .ZN(n6819) );
  AND2_X1 U4102 ( .A1(n5324), .A2(n5325), .ZN(n5318) );
  INV_X1 U4103 ( .A(n3974), .ZN(n4969) );
  OR2_X1 U4104 ( .A1(n4881), .A2(n6773), .ZN(n3647) );
  OR2_X1 U4105 ( .A1(n6773), .A2(n6188), .ZN(n3648) );
  NAND2_X1 U4106 ( .A1(n4996), .A2(n4995), .ZN(n4994) );
  NAND2_X1 U4107 ( .A1(n3675), .A2(n3674), .ZN(n4976) );
  NAND2_X1 U4108 ( .A1(n7194), .A2(n7221), .ZN(n6804) );
  INV_X1 U4109 ( .A(n4146), .ZN(n5094) );
  NAND2_X1 U4110 ( .A1(n4143), .A2(n4142), .ZN(n4146) );
  AND2_X1 U4111 ( .A1(n4388), .A2(n4373), .ZN(n3649) );
  OR2_X1 U4112 ( .A1(n7426), .A2(n6833), .ZN(n6791) );
  NOR2_X4 U4113 ( .A1(n6829), .A2(n6651), .ZN(n7229) );
  XNOR2_X2 U4114 ( .A(n3655), .B(n3654), .ZN(n6494) );
  NAND2_X1 U4115 ( .A1(n3660), .A2(n6781), .ZN(n4582) );
  NAND3_X1 U4116 ( .A1(n4576), .A2(n4575), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n3660) );
  NAND2_X1 U4117 ( .A1(n6780), .A2(n4770), .ZN(n4581) );
  INV_X1 U4118 ( .A(n3662), .ZN(n3661) );
  OAI21_X1 U4119 ( .B1(n3664), .B2(n4586), .A(n5238), .ZN(n3662) );
  NAND2_X1 U4120 ( .A1(n5616), .A2(n3671), .ZN(n3669) );
  NAND2_X1 U4121 ( .A1(n4615), .A2(n3667), .ZN(n3666) );
  INV_X1 U4122 ( .A(n5617), .ZN(n3667) );
  NAND3_X1 U4123 ( .A1(n3669), .A2(n3668), .A3(n4625), .ZN(n6009) );
  NAND2_X1 U4124 ( .A1(n3673), .A2(n3641), .ZN(n4636) );
  NAND2_X1 U4125 ( .A1(n3675), .A2(n4559), .ZN(n4564) );
  NAND2_X1 U4126 ( .A1(n3626), .A2(n3634), .ZN(n6394) );
  AND2_X2 U4127 ( .A1(n5048), .A2(n5049), .ZN(n3931) );
  AND2_X2 U4128 ( .A1(n5048), .A2(n5078), .ZN(n3895) );
  AND2_X2 U4129 ( .A1(n6147), .A2(n5048), .ZN(n3873) );
  NOR2_X4 U4130 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U4131 ( .A1(n6297), .A2(n3683), .ZN(n6293) );
  INV_X1 U4132 ( .A(n6293), .ZN(n4462) );
  NAND2_X1 U4133 ( .A1(n5541), .A2(n3645), .ZN(n5623) );
  NAND2_X1 U4134 ( .A1(n6044), .A2(n6045), .ZN(n4337) );
  NAND3_X1 U4135 ( .A1(n5249), .A2(n5322), .A3(n5317), .ZN(n5316) );
  NAND3_X1 U4136 ( .A1(n5249), .A2(n5322), .A3(n3646), .ZN(n5540) );
  NAND2_X1 U4137 ( .A1(n3685), .A2(n4748), .ZN(n3967) );
  NAND4_X1 U4138 ( .A1(n4068), .A2(n5364), .A3(n3965), .A4(n3962), .ZN(n4748)
         );
  NAND3_X1 U4139 ( .A1(n3688), .A2(n3966), .A3(n3686), .ZN(n3685) );
  NOR2_X1 U4140 ( .A1(n6209), .A2(n6211), .ZN(n4884) );
  NAND2_X1 U4141 ( .A1(n4144), .A2(n4146), .ZN(n4171) );
  INV_X1 U4142 ( .A(n4196), .ZN(n4208) );
  NAND2_X1 U4143 ( .A1(n4706), .A2(n6819), .ZN(n4715) );
  INV_X1 U4144 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6412) );
  INV_X1 U4145 ( .A(n6003), .ZN(n3956) );
  INV_X1 U4146 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3701) );
  AND2_X1 U4147 ( .A1(n3625), .A2(n4665), .ZN(n3694) );
  INV_X1 U4148 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4560) );
  AND2_X1 U4149 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3695)
         );
  NAND2_X1 U4150 ( .A1(n3633), .A2(n6455), .ZN(n3696) );
  INV_X1 U4151 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4152 ( .A1(n6123), .A2(n4857), .ZN(n3697) );
  INV_X1 U4153 ( .A(n3920), .ZN(n3751) );
  OR2_X1 U4154 ( .A1(n3977), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3698)
         );
  NOR2_X1 U4155 ( .A1(n4754), .A2(n4664), .ZN(n3975) );
  OR2_X1 U4156 ( .A1(n4234), .A2(n5449), .ZN(n4169) );
  NAND2_X1 U4157 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7417), .ZN(n4670) );
  AND2_X1 U4158 ( .A1(n4673), .A2(n4651), .ZN(n4683) );
  INV_X1 U4159 ( .A(n6258), .ZN(n4373) );
  OR2_X1 U4160 ( .A1(n4115), .A2(n4114), .ZN(n4566) );
  OR2_X1 U4161 ( .A1(n4671), .A2(n4670), .ZN(n4673) );
  NAND2_X1 U4162 ( .A1(n4684), .A2(n4655), .ZN(n4660) );
  INV_X1 U4163 ( .A(n6753), .ZN(n4441) );
  INV_X1 U4164 ( .A(n6313), .ZN(n4388) );
  INV_X1 U4165 ( .A(n6294), .ZN(n4461) );
  OR2_X1 U4166 ( .A1(n5623), .A2(n4335), .ZN(n4336) );
  OR2_X1 U4167 ( .A1(n4525), .A2(n4526), .ZN(n4534) );
  NAND2_X1 U4168 ( .A1(n6141), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U4169 ( .A1(n5237), .A2(n4597), .ZN(n5383) );
  AND2_X1 U4170 ( .A1(n7161), .A2(n4970), .ZN(n5045) );
  INV_X1 U4171 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4338) );
  INV_X1 U4172 ( .A(n5004), .ZN(n4781) );
  INV_X1 U4173 ( .A(n5397), .ZN(n4271) );
  NAND2_X1 U4174 ( .A1(n5083), .A2(n4366), .ZN(n4061) );
  NAND2_X1 U4175 ( .A1(n4515), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4525)
         );
  NOR2_X1 U4176 ( .A1(n4302), .A2(n7040), .ZN(n4331) );
  NAND2_X1 U4177 ( .A1(n4863), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4864) );
  INV_X1 U4178 ( .A(n3632), .ZN(n5258) );
  OR2_X1 U4179 ( .A1(n6239), .A2(n6130), .ZN(n6214) );
  NAND2_X1 U4180 ( .A1(n4442), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4463)
         );
  NOR2_X1 U4181 ( .A1(n4342), .A2(n4338), .ZN(n4357) );
  INV_X1 U4182 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U4183 ( .A1(n6941), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5304) );
  AND2_X1 U4184 ( .A1(n4797), .A2(n4796), .ZN(n5543) );
  NAND2_X1 U4185 ( .A1(n4298), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4302)
         );
  AND2_X1 U4186 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4177)
         );
  AND2_X1 U4187 ( .A1(n6804), .A2(n4708), .ZN(n4711) );
  INV_X1 U4188 ( .A(n3946), .ZN(n5058) );
  NAND2_X1 U4189 ( .A1(n4171), .A2(n4147), .ZN(n5084) );
  NOR2_X1 U4190 ( .A1(n5084), .A2(n5177), .ZN(n7387) );
  INV_X1 U4191 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7417) );
  AND2_X1 U4192 ( .A1(n5259), .A2(n5258), .ZN(n7348) );
  AND2_X1 U4193 ( .A1(n7164), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4705) );
  AND2_X1 U4194 ( .A1(n6170), .A2(n4905), .ZN(n7249) );
  INV_X1 U4195 ( .A(READY_N), .ZN(n7250) );
  OAI21_X1 U4196 ( .B1(n6494), .B2(n7152), .A(n6195), .ZN(n6196) );
  OR2_X1 U4197 ( .A1(n4500), .A2(n3702), .ZN(n4510) );
  NOR2_X1 U4198 ( .A1(n4463), .A2(n6412), .ZN(n4481) );
  XNOR2_X1 U4199 ( .A(n4875), .B(n6184), .ZN(n5295) );
  INV_X1 U4200 ( .A(n7130), .ZN(n7155) );
  INV_X1 U4201 ( .A(n7094), .ZN(n7086) );
  NOR2_X2 U4202 ( .A1(n5304), .A2(n5303), .ZN(n7125) );
  INV_X1 U4203 ( .A(n6773), .ZN(n6311) );
  AND2_X1 U4204 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  OAI21_X1 U4205 ( .B1(n5361), .B2(n5360), .A(n7221), .ZN(n5363) );
  INV_X1 U4206 ( .A(n6813), .ZN(n7336) );
  INV_X1 U4207 ( .A(n4711), .ZN(n6448) );
  AND2_X1 U4208 ( .A1(n4990), .A2(n6166), .ZN(n6870) );
  AND2_X1 U4209 ( .A1(n4990), .A2(n7159), .ZN(n6921) );
  INV_X1 U4210 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7164) );
  NOR2_X1 U4211 ( .A1(n6004), .A2(n7214), .ZN(n6108) );
  INV_X1 U4212 ( .A(n5144), .ZN(n7573) );
  AND3_X1 U4213 ( .A1(n5332), .A2(n6118), .A3(n5084), .ZN(n5608) );
  AND2_X1 U4214 ( .A1(n7401), .A2(n6118), .ZN(n7564) );
  AND2_X1 U4215 ( .A1(n7401), .A2(n7371), .ZN(n7565) );
  INV_X1 U4216 ( .A(n5522), .ZN(n5503) );
  AND2_X1 U4217 ( .A1(n7387), .A2(n7371), .ZN(n7556) );
  INV_X1 U4218 ( .A(n5346), .ZN(n7545) );
  AND2_X1 U4219 ( .A1(n7348), .A2(n6118), .ZN(n7538) );
  AND2_X1 U4220 ( .A1(n7348), .A2(n7371), .ZN(n7539) );
  AND2_X1 U4221 ( .A1(n6818), .A2(DATAI_25_), .ZN(n7453) );
  AND2_X1 U4222 ( .A1(n6818), .A2(DATAI_28_), .ZN(n7500) );
  AND2_X1 U4223 ( .A1(n5099), .A2(n6118), .ZN(n5533) );
  INV_X1 U4224 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7240) );
  OR2_X1 U4225 ( .A1(n7426), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U4226 ( .A1(n5286), .A2(n5285), .ZN(n6838) );
  INV_X1 U4227 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7413) );
  INV_X1 U4228 ( .A(n7125), .ZN(n7152) );
  INV_X1 U4229 ( .A(n7144), .ZN(n7122) );
  INV_X1 U4230 ( .A(n7145), .ZN(n7120) );
  OR2_X1 U4231 ( .A1(n5295), .A2(n5293), .ZN(n7130) );
  INV_X1 U4232 ( .A(n7133), .ZN(n7157) );
  NAND2_X1 U4233 ( .A1(n5363), .A2(n7329), .ZN(n6142) );
  NAND2_X1 U4234 ( .A1(n6652), .A2(n3929), .ZN(n5284) );
  INV_X1 U4235 ( .A(n6652), .ZN(n6670) );
  NAND2_X2 U4236 ( .A1(n6170), .A2(n4922), .ZN(n7333) );
  NAND2_X1 U4237 ( .A1(n6448), .A2(n5008), .ZN(n6822) );
  INV_X1 U4238 ( .A(n6915), .ZN(n6619) );
  OR2_X1 U4239 ( .A1(n6160), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6924) );
  INV_X1 U4240 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7361) );
  INV_X1 U4241 ( .A(n7420), .ZN(n7579) );
  OR2_X1 U4242 ( .A1(n5178), .A2(n6118), .ZN(n5522) );
  AOI22_X1 U4243 ( .A1(n7377), .A2(n7384), .B1(n7376), .B2(n7375), .ZN(n7555)
         );
  AND2_X1 U4244 ( .A1(n7408), .A2(n5096), .ZN(n5494) );
  OAI21_X1 U4245 ( .B1(n4716), .B2(n6315), .A(n4883), .ZN(U2830) );
  INV_X1 U4246 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3702) );
  INV_X1 U4247 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6247) );
  INV_X1 U4248 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4526) );
  INV_X1 U4249 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4533) );
  INV_X1 U4250 ( .A(n4543), .ZN(n3703) );
  NAND2_X1 U4251 ( .A1(n3703), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3705)
         );
  INV_X1 U4252 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4253 ( .A1(n3705), .A2(n3704), .ZN(n3706) );
  NAND2_X1 U4254 ( .A1(n4874), .A2(n3706), .ZN(n6199) );
  INV_X1 U4255 ( .A(n3936), .ZN(n4490) );
  INV_X2 U4256 ( .A(n4490), .ZN(n4721) );
  AOI22_X1 U4257 ( .A1(n4721), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4726), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3711) );
  AND2_X4 U4258 ( .A1(n5053), .A2(n5049), .ZN(n3894) );
  AOI22_X1 U4259 ( .A1(n4728), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3710) );
  AND2_X2 U4260 ( .A1(n6146), .A2(n5050), .ZN(n3862) );
  AOI22_X1 U4261 ( .A1(n4448), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3709) );
  AND2_X2 U4262 ( .A1(n5078), .A2(n5050), .ZN(n3906) );
  INV_X2 U4263 ( .A(n5058), .ZN(n4470) );
  AOI22_X1 U4264 ( .A1(n4005), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4265 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3718)
         );
  AND2_X4 U4266 ( .A1(n5054), .A2(n6147), .ZN(n4016) );
  AND2_X4 U4267 ( .A1(n6147), .A2(n5050), .ZN(n3920) );
  INV_X2 U4268 ( .A(n3751), .ZN(n4487) );
  AOI22_X1 U4269 ( .A1(n4016), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4270 ( .A1(n3868), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3715) );
  AND2_X2 U4271 ( .A1(n5053), .A2(n5078), .ZN(n3878) );
  AOI22_X1 U4272 ( .A1(n4465), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3714) );
  INV_X1 U4273 ( .A(n3919), .ZN(n4000) );
  INV_X2 U4274 ( .A(n4000), .ZN(n4717) );
  AOI22_X1 U4275 ( .A1(n4717), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4276 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  NOR2_X1 U4277 ( .A1(n3718), .A2(n3717), .ZN(n4736) );
  AOI22_X1 U4278 ( .A1(n4017), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4279 ( .A1(n4720), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4280 ( .A1(n4719), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4281 ( .A1(n4005), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4282 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3728)
         );
  INV_X2 U4283 ( .A(n4022), .ZN(n4448) );
  AOI22_X1 U4284 ( .A1(n4717), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4285 ( .A1(n4482), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4286 ( .A1(n4726), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4287 ( .A1(n4721), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4288 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  NOR2_X1 U4289 ( .A1(n3728), .A2(n3727), .ZN(n4546) );
  AOI22_X1 U4290 ( .A1(n4721), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4291 ( .A1(n4717), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4292 ( .A1(n4726), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4293 ( .A1(n4728), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4294 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3738)
         );
  AOI22_X1 U4295 ( .A1(n4017), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4296 ( .A1(n4720), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4297 ( .A1(n4465), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4298 ( .A1(n4487), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4299 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3737)
         );
  NOR2_X1 U4300 ( .A1(n3738), .A2(n3737), .ZN(n4529) );
  AOI22_X1 U4301 ( .A1(n4448), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4302 ( .A1(n4720), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4303 ( .A1(n4726), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4304 ( .A1(n4719), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4305 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3748)
         );
  AOI22_X1 U4306 ( .A1(n4017), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4717), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4307 ( .A1(n4482), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4308 ( .A1(n4721), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4309 ( .A1(n4005), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3743) );
  NAND4_X1 U4310 ( .A1(n3746), .A2(n3745), .A3(n3744), .A4(n3743), .ZN(n3747)
         );
  NOR2_X1 U4311 ( .A1(n3748), .A2(n3747), .ZN(n4508) );
  INV_X1 U4312 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3749) );
  NOR2_X1 U4313 ( .A1(n4022), .A2(n3749), .ZN(n3753) );
  INV_X1 U4314 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5188) );
  INV_X1 U4315 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3750) );
  OAI22_X1 U4316 ( .A1(n4000), .A2(n5188), .B1(n3751), .B2(n3750), .ZN(n3752)
         );
  AOI211_X1 U4317 ( .C1(INSTQUEUE_REG_9__7__SCAN_IN), .C2(n4017), .A(n3753), 
        .B(n3752), .ZN(n3761) );
  AOI22_X1 U4318 ( .A1(n4719), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4319 ( .A1(n4720), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4320 ( .A1(n4482), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4321 ( .A1(n4721), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4322 ( .A1(n4718), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4323 ( .A1(n4726), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3754) );
  AND4_X1 U4324 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NAND4_X1 U4325 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n4503)
         );
  AOI22_X1 U4326 ( .A1(n4017), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4327 ( .A1(n4717), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4328 ( .A1(n4720), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4329 ( .A1(n4719), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3762) );
  NAND4_X1 U4330 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3771)
         );
  AOI22_X1 U4331 ( .A1(n4482), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4332 ( .A1(n4721), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4333 ( .A1(n4718), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4334 ( .A1(n4726), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3766) );
  NAND4_X1 U4335 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3770)
         );
  OR2_X1 U4336 ( .A1(n3771), .A2(n3770), .ZN(n4502) );
  NAND2_X1 U4337 ( .A1(n4503), .A2(n4502), .ZN(n4509) );
  NOR2_X1 U4338 ( .A1(n4508), .A2(n4509), .ZN(n4519) );
  AOI22_X1 U4339 ( .A1(n4017), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4340 ( .A1(n4717), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4341 ( .A1(n4720), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4342 ( .A1(n4719), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4343 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3781)
         );
  AOI22_X1 U4344 ( .A1(n4482), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4345 ( .A1(n4721), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4346 ( .A1(n4718), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4347 ( .A1(n4726), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4348 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  OR2_X1 U4349 ( .A1(n3781), .A2(n3780), .ZN(n4520) );
  NAND2_X1 U4350 ( .A1(n4519), .A2(n4520), .ZN(n4528) );
  NOR2_X1 U4351 ( .A1(n4529), .A2(n4528), .ZN(n4537) );
  AOI22_X1 U4352 ( .A1(n4016), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4353 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4717), .B1(n4487), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4354 ( .A1(n4720), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4355 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4719), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4356 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AOI22_X1 U4357 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4465), .B1(n4482), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4358 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4721), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4359 ( .A1(n4718), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4360 ( .A1(n4726), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4361 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  OR2_X1 U4362 ( .A1(n3791), .A2(n3790), .ZN(n4536) );
  NAND2_X1 U4363 ( .A1(n4537), .A2(n4536), .ZN(n4545) );
  OR2_X1 U4364 ( .A1(n4546), .A2(n4545), .ZN(n4735) );
  XNOR2_X1 U4365 ( .A(n4736), .B(n4735), .ZN(n3890) );
  NAND2_X1 U4366 ( .A1(n3905), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U4367 ( .A1(n3936), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U4368 ( .A1(n3878), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3793) );
  NAND2_X1 U4369 ( .A1(n3906), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3792)
         );
  NAND2_X1 U4370 ( .A1(n3867), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4371 ( .A1(n3868), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3798) );
  NAND2_X1 U4372 ( .A1(n3895), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4373 ( .A1(n3931), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4374 ( .A1(n4016), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4375 ( .A1(n3862), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3802)
         );
  NAND2_X1 U4376 ( .A1(n3919), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4377 ( .A1(n3920), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4378 ( .A1(n3873), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4379 ( .A1(n3629), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3806) );
  NAND2_X1 U4380 ( .A1(n3894), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3805)
         );
  NAND2_X1 U4381 ( .A1(n3946), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3804)
         );
  NAND2_X1 U4382 ( .A1(n3936), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4383 ( .A1(n3905), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3814)
         );
  NAND2_X1 U4384 ( .A1(n3878), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3813) );
  NAND2_X1 U4385 ( .A1(n3906), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3812)
         );
  NAND2_X1 U4386 ( .A1(n3862), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3819)
         );
  NAND2_X1 U4387 ( .A1(n4016), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4388 ( .A1(n3919), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4389 ( .A1(n3920), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3816)
         );
  NAND2_X1 U4390 ( .A1(n3867), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3823) );
  NAND2_X1 U4391 ( .A1(n3868), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4392 ( .A1(n3895), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4393 ( .A1(n3931), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3820) );
  NAND2_X1 U4394 ( .A1(n3873), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4395 ( .A1(n3941), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4396 ( .A1(n3894), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3825)
         );
  NAND2_X1 U4397 ( .A1(n3946), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3824)
         );
  NAND2_X1 U4398 ( .A1(n3862), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3835)
         );
  NAND2_X1 U4399 ( .A1(n4016), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4400 ( .A1(n3868), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3833) );
  NAND2_X1 U4401 ( .A1(n3895), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4402 ( .A1(n3919), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4403 ( .A1(n3920), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3838)
         );
  NAND2_X1 U4404 ( .A1(n3867), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4405 ( .A1(n3931), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4407 ( .A1(n3941), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3843) );
  NAND2_X1 U4408 ( .A1(n3936), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4409 ( .A1(n3894), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3841)
         );
  NAND2_X1 U4410 ( .A1(n3878), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3840) );
  NAND2_X1 U4411 ( .A1(n3905), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3847)
         );
  NAND2_X1 U4412 ( .A1(n3946), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3846)
         );
  NAND2_X1 U4413 ( .A1(n3873), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4414 ( .A1(n3906), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3844)
         );
  AOI22_X1 U4415 ( .A1(n3919), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4416 ( .A1(n3941), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4417 ( .A1(n3905), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4418 ( .A1(n3868), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4419 ( .A1(n3873), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4420 ( .A1(n3936), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4421 ( .A1(n4016), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4422 ( .A1(n3906), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3946), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3856) );
  INV_X1 U4423 ( .A(n4748), .ZN(n3991) );
  NAND2_X1 U4424 ( .A1(n3862), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U4425 ( .A1(n4016), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U4426 ( .A1(n3919), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4427 ( .A1(n3920), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3863)
         );
  NAND2_X1 U4428 ( .A1(n3867), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U4429 ( .A1(n3868), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4430 ( .A1(n3895), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3870) );
  NAND2_X1 U4431 ( .A1(n3931), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4432 ( .A1(n3873), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3877) );
  NAND2_X1 U4433 ( .A1(n3941), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U4434 ( .A1(n3894), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3875)
         );
  NAND2_X1 U4435 ( .A1(n3946), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3874)
         );
  NAND2_X1 U4436 ( .A1(n3905), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3882)
         );
  NAND2_X1 U4437 ( .A1(n3936), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U4438 ( .A1(n3878), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U4439 ( .A1(n3906), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3879)
         );
  INV_X2 U4440 ( .A(n5289), .ZN(n4550) );
  AOI21_X1 U4441 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n3887), .A(n4550), 
        .ZN(n3889) );
  NAND2_X1 U4442 ( .A1(n4870), .A2(EAX_REG_29__SCAN_IN), .ZN(n3888) );
  OAI211_X1 U4443 ( .C1(n3890), .C2(n4540), .A(n3889), .B(n3888), .ZN(n3891)
         );
  OAI21_X1 U4444 ( .B1(n6199), .B2(n5289), .A(n3891), .ZN(n4552) );
  INV_X1 U4445 ( .A(n3969), .ZN(n3892) );
  OAI21_X1 U4446 ( .B1(n3962), .B2(n4944), .A(n3892), .ZN(n4948) );
  AND2_X1 U4447 ( .A1(n4944), .A2(n4015), .ZN(n3893) );
  NOR2_X2 U4448 ( .A1(n4948), .A2(n3893), .ZN(n3986) );
  AOI22_X1 U4449 ( .A1(n3919), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4450 ( .A1(n3868), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4451 ( .A1(n3936), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4452 ( .A1(n4016), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4453 ( .A1(n3941), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4454 ( .A1(n3905), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3878), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4455 ( .A1(n3906), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3946), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U4456 ( .A1(n5403), .A2(n3974), .ZN(n4555) );
  NOR2_X1 U4457 ( .A1(n4555), .A2(n4665), .ZN(n3904) );
  NAND2_X1 U4458 ( .A1(n3986), .A2(n3904), .ZN(n4921) );
  INV_X1 U4459 ( .A(n4921), .ZN(n3930) );
  NAND2_X1 U4460 ( .A1(n3905), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3910)
         );
  NAND2_X1 U4461 ( .A1(n3936), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U4462 ( .A1(n3878), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4463 ( .A1(n3906), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3907)
         );
  NAND2_X1 U4464 ( .A1(n3868), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3914) );
  NAND2_X1 U4465 ( .A1(n3867), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3913) );
  NAND2_X1 U4466 ( .A1(n3895), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3912) );
  NAND2_X1 U4467 ( .A1(n3931), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4468 ( .A1(n3873), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U4469 ( .A1(n3941), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3917) );
  NAND2_X1 U4470 ( .A1(n3894), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3916)
         );
  NAND2_X1 U4471 ( .A1(n3946), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3915)
         );
  NAND2_X1 U4472 ( .A1(n3862), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3924)
         );
  NAND2_X1 U4473 ( .A1(n4016), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U4474 ( .A1(n3919), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4475 ( .A1(n3920), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3921)
         );
  AND4_X4 U4476 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n5109)
         );
  NAND2_X1 U4477 ( .A1(n3930), .A2(n3929), .ZN(n4903) );
  NAND2_X1 U4478 ( .A1(n4016), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4479 ( .A1(n3919), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4480 ( .A1(n3920), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3933)
         );
  NAND2_X1 U4481 ( .A1(n3931), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3932) );
  NAND2_X1 U4482 ( .A1(n3905), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3940)
         );
  NAND2_X1 U4483 ( .A1(n3868), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4484 ( .A1(n3936), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U4485 ( .A1(n3878), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3937) );
  NAND2_X1 U4486 ( .A1(n3862), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3945)
         );
  NAND2_X1 U4487 ( .A1(n3941), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U4488 ( .A1(n3867), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3943) );
  NAND2_X1 U4489 ( .A1(n3895), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3942) );
  NAND2_X1 U4490 ( .A1(n3873), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3950) );
  NAND2_X1 U4491 ( .A1(n3894), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3949)
         );
  NAND2_X1 U4492 ( .A1(n3906), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3948)
         );
  NAND2_X1 U4493 ( .A1(n3946), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3947)
         );
  XNOR2_X1 U4494 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n7237) );
  INV_X1 U4495 ( .A(n7237), .ZN(n3955) );
  NOR2_X1 U4496 ( .A1(n3970), .A2(n3955), .ZN(n3971) );
  NAND2_X1 U4497 ( .A1(n3966), .A2(n3963), .ZN(n4980) );
  INV_X1 U4498 ( .A(n4980), .ZN(n3958) );
  NAND3_X1 U4499 ( .A1(n3638), .A2(n3694), .A3(n3958), .ZN(n4901) );
  INV_X1 U4500 ( .A(n4901), .ZN(n3959) );
  OAI211_X1 U4501 ( .C1(n4903), .C2(n3971), .A(n4972), .B(n5039), .ZN(n3960)
         );
  NAND2_X1 U4502 ( .A1(n3960), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3978) );
  INV_X1 U4503 ( .A(n3978), .ZN(n3961) );
  NAND2_X1 U4504 ( .A1(n7164), .A2(n7214), .ZN(n7169) );
  NAND2_X1 U4505 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5121) );
  OAI21_X1 U4506 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n5121), .ZN(n5342) );
  OAI22_X1 U4507 ( .A1(n4707), .A2(n5342), .B1(n4705), .B2(n7412), .ZN(n3977)
         );
  NAND2_X1 U4508 ( .A1(n3961), .A2(n3698), .ZN(n3981) );
  NAND2_X1 U4509 ( .A1(n3967), .A2(n3988), .ZN(n3968) );
  NAND2_X1 U4510 ( .A1(n4943), .A2(n4569), .ZN(n3993) );
  INV_X1 U4511 ( .A(n3971), .ZN(n3972) );
  AOI21_X1 U4512 ( .B1(n3687), .B2(n3972), .A(n4555), .ZN(n3973) );
  NAND4_X1 U4513 ( .A1(n3996), .A2(n3993), .A3(n3986), .A4(n3973), .ZN(n3976)
         );
  AOI21_X2 U4514 ( .B1(n3976), .B2(STATE2_REG_0__SCAN_IN), .A(n3975), .ZN(
        n3982) );
  OR2_X1 U4515 ( .A1(n3982), .A2(n3707), .ZN(n3980) );
  INV_X1 U4516 ( .A(n3977), .ZN(n3979) );
  NAND3_X1 U4517 ( .A1(n3980), .A2(n3979), .A3(n3978), .ZN(n4091) );
  INV_X1 U4518 ( .A(n3982), .ZN(n4093) );
  NAND2_X1 U4519 ( .A1(n4093), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3985) );
  INV_X1 U4520 ( .A(n4705), .ZN(n4128) );
  INV_X1 U4521 ( .A(n4707), .ZN(n4129) );
  MUX2_X1 U4522 ( .A(n4128), .B(n4129), .S(n7417), .Z(n3983) );
  INV_X1 U4523 ( .A(n3983), .ZN(n3984) );
  NAND2_X1 U4524 ( .A1(n3985), .A2(n3984), .ZN(n4033) );
  INV_X1 U4525 ( .A(n3987), .ZN(n3995) );
  INV_X1 U4526 ( .A(n3988), .ZN(n3989) );
  NAND2_X1 U4527 ( .A1(n3989), .A2(n5403), .ZN(n3990) );
  NAND2_X1 U4528 ( .A1(n3990), .A2(n3929), .ZN(n3994) );
  OR2_X1 U4529 ( .A1(n7169), .A2(n7224), .ZN(n7207) );
  INV_X1 U4530 ( .A(n7207), .ZN(n3992) );
  NAND2_X1 U4531 ( .A1(n3991), .A2(n3638), .ZN(n5071) );
  NAND2_X1 U4532 ( .A1(n3995), .A2(n3640), .ZN(n3999) );
  INV_X1 U4533 ( .A(n3996), .ZN(n3997) );
  NAND2_X1 U4534 ( .A1(n4694), .A2(n3963), .ZN(n4956) );
  NAND2_X1 U4535 ( .A1(n3997), .A2(n4956), .ZN(n4983) );
  NAND3_X1 U4536 ( .A1(n4765), .A2(n3963), .A3(n4665), .ZN(n3998) );
  NAND2_X1 U4537 ( .A1(n4983), .A2(n3998), .ZN(n5038) );
  AND2_X2 U4538 ( .A1(n4033), .A2(n3623), .ZN(n4089) );
  NAND2_X1 U4539 ( .A1(n5089), .A2(n7224), .ZN(n4013) );
  INV_X1 U4540 ( .A(n4664), .ZN(n4030) );
  AOI22_X1 U4541 ( .A1(n4017), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4542 ( .A1(n4717), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4543 ( .A1(n4482), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4544 ( .A1(n3867), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4545 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4011)
         );
  AOI22_X1 U4546 ( .A1(n4721), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4726), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4547 ( .A1(n4465), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4548 ( .A1(n4720), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4549 ( .A1(n4005), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4550 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  NAND2_X1 U4551 ( .A1(n4030), .A2(n4553), .ZN(n4012) );
  INV_X1 U4552 ( .A(n4553), .ZN(n4032) );
  INV_X1 U4553 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5152) );
  OR2_X1 U4554 ( .A1(n4234), .A2(n5152), .ZN(n4031) );
  AOI22_X1 U4555 ( .A1(n4017), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4556 ( .A1(n4482), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4557 ( .A1(n4720), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4558 ( .A1(n3894), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4559 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4028)
         );
  AOI22_X1 U4560 ( .A1(n4717), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4561 ( .A1(n4721), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4562 ( .A1(n3873), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4563 ( .A1(n4726), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4564 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  INV_X1 U4565 ( .A(n4620), .ZN(n4029) );
  NAND2_X1 U4566 ( .A1(n4030), .A2(n4029), .ZN(n4037) );
  OAI211_X1 U4567 ( .C1(n4032), .C2(n4105), .A(n4031), .B(n4037), .ZN(n4084)
         );
  INV_X1 U4569 ( .A(n4033), .ZN(n4035) );
  INV_X1 U4570 ( .A(n3623), .ZN(n4034) );
  NAND2_X1 U4571 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  NAND2_X1 U4572 ( .A1(n3624), .A2(n4036), .ZN(n4070) );
  INV_X1 U4573 ( .A(n4037), .ZN(n4049) );
  NAND2_X1 U4574 ( .A1(n3963), .A2(n4620), .ZN(n4051) );
  AOI22_X1 U4575 ( .A1(n4717), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4576 ( .A1(n4482), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4577 ( .A1(n4720), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4578 ( .A1(n4443), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U4579 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U4580 ( .A1(n4017), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4581 ( .A1(n4721), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4726), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4582 ( .A1(n3867), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4583 ( .A1(n3894), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U4584 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  INV_X1 U4585 ( .A(n4561), .ZN(n4048) );
  MUX2_X1 U4586 ( .A(n4049), .B(n4617), .S(n4048), .Z(n4065) );
  INV_X1 U4587 ( .A(n4065), .ZN(n4050) );
  NAND2_X1 U4588 ( .A1(n4062), .A2(n4050), .ZN(n4055) );
  INV_X1 U4589 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5155) );
  AOI21_X1 U4590 ( .B1(n5109), .B2(n4561), .A(n7224), .ZN(n4052) );
  AND2_X1 U4591 ( .A1(n4052), .A2(n4051), .ZN(n4053) );
  NAND2_X1 U4592 ( .A1(n4054), .A2(n4053), .ZN(n4064) );
  AOI22_X1 U4594 ( .A1(n4870), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n3887), .ZN(n4059) );
  AND2_X1 U4595 ( .A1(n3966), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4148) );
  NAND2_X1 U4596 ( .A1(n4148), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4058) );
  AND2_X1 U4597 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  NAND2_X1 U4598 ( .A1(n4062), .A2(n4064), .ZN(n4063) );
  NAND2_X1 U4599 ( .A1(n4063), .A2(n4050), .ZN(n4067) );
  NAND2_X1 U4600 ( .A1(n4065), .A2(n4064), .ZN(n4066) );
  AND2_X1 U4601 ( .A1(n4068), .A2(n5364), .ZN(n4069) );
  OR2_X1 U4603 ( .A1(n5092), .A2(n4330), .ZN(n4074) );
  AOI22_X1 U4604 ( .A1(n4870), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n3887), .ZN(n4072) );
  NAND2_X1 U4605 ( .A1(n4148), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4071) );
  AND2_X1 U4606 ( .A1(n4072), .A2(n4071), .ZN(n4073) );
  NAND2_X1 U4607 ( .A1(n4074), .A2(n4073), .ZN(n4910) );
  INV_X1 U4608 ( .A(n4910), .ZN(n4075) );
  NAND2_X1 U4609 ( .A1(n4075), .A2(n4550), .ZN(n4076) );
  NAND2_X1 U4610 ( .A1(n4909), .A2(n4076), .ZN(n4995) );
  NAND2_X1 U4611 ( .A1(n4148), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4082) );
  INV_X1 U4612 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5313) );
  INV_X1 U4613 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6930) );
  NOR2_X1 U4614 ( .A1(n5313), .A2(n6930), .ZN(n4150) );
  AOI21_X1 U4615 ( .B1(n5313), .B2(n6930), .A(n4150), .ZN(n4077) );
  INV_X1 U4616 ( .A(n4077), .ZN(n6938) );
  NAND2_X1 U4617 ( .A1(n6938), .A2(n4550), .ZN(n4079) );
  NAND2_X1 U4618 ( .A1(n4869), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4078)
         );
  NAND2_X1 U4619 ( .A1(n4079), .A2(n4078), .ZN(n4080) );
  AOI21_X1 U4620 ( .B1(n4870), .B2(EAX_REG_2__SCAN_IN), .A(n4080), .ZN(n4081)
         );
  AND2_X1 U4621 ( .A1(n4082), .A2(n4081), .ZN(n4121) );
  NAND2_X1 U4622 ( .A1(n4083), .A2(n4084), .ZN(n4085) );
  INV_X1 U4623 ( .A(n4088), .ZN(n4090) );
  NAND2_X1 U4624 ( .A1(n4090), .A2(n3624), .ZN(n4092) );
  NAND2_X1 U4626 ( .A1(n4094), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4099) );
  INV_X1 U4627 ( .A(n5121), .ZN(n4095) );
  NAND2_X1 U4628 ( .A1(n5121), .A2(n5327), .ZN(n4096) );
  NAND2_X1 U4629 ( .A1(n5093), .A2(n4096), .ZN(n5142) );
  OAI22_X1 U4630 ( .A1(n5142), .A2(n4707), .B1(n4705), .B2(n5327), .ZN(n4097)
         );
  INV_X1 U4631 ( .A(n4097), .ZN(n4098) );
  INV_X1 U4632 ( .A(n4100), .ZN(n4103) );
  INV_X1 U4633 ( .A(n4101), .ZN(n4102) );
  AOI22_X1 U4634 ( .A1(n4017), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4635 ( .A1(n4717), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4636 ( .A1(n4720), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4637 ( .A1(n4719), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U4638 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4115)
         );
  AOI22_X1 U4639 ( .A1(n4482), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4640 ( .A1(n4721), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4641 ( .A1(n4718), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U4642 ( .A1(n4726), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U4643 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4114)
         );
  AOI22_X1 U4644 ( .A1(n4686), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4700), 
        .B2(n4566), .ZN(n4116) );
  INV_X1 U4645 ( .A(n4869), .ZN(n4120) );
  NAND2_X1 U4646 ( .A1(n4915), .A2(n4916), .ZN(n4125) );
  INV_X1 U4647 ( .A(n4994), .ZN(n4123) );
  INV_X1 U4648 ( .A(n4121), .ZN(n4122) );
  NAND2_X1 U4649 ( .A1(n4123), .A2(n4122), .ZN(n4124) );
  NAND2_X1 U4650 ( .A1(n4094), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4131) );
  NAND2_X1 U4651 ( .A1(n4126), .A2(n7361), .ZN(n5199) );
  NAND2_X1 U4652 ( .A1(n5093), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4127) );
  NAND2_X1 U4653 ( .A1(n5199), .A2(n4127), .ZN(n5341) );
  AOI22_X1 U4654 ( .A1(n5341), .A2(n4129), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4128), .ZN(n4130) );
  XNOR2_X1 U4655 ( .A(n5031), .B(n5029), .ZN(n5037) );
  NAND2_X1 U4656 ( .A1(n5037), .A2(n7224), .ZN(n4143) );
  AOI22_X1 U4657 ( .A1(n4017), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4658 ( .A1(n4717), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4659 ( .A1(n4720), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4660 ( .A1(n4719), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4132) );
  NAND4_X1 U4661 ( .A1(n4135), .A2(n4134), .A3(n4133), .A4(n4132), .ZN(n4141)
         );
  AOI22_X1 U4662 ( .A1(n4482), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U4663 ( .A1(n4721), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4664 ( .A1(n4718), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U4665 ( .A1(n4726), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4136) );
  NAND4_X1 U4666 ( .A1(n4139), .A2(n4138), .A3(n4137), .A4(n4136), .ZN(n4140)
         );
  AOI22_X1 U4667 ( .A1(n4686), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4700), 
        .B2(n4578), .ZN(n4142) );
  NAND2_X1 U4668 ( .A1(n4145), .A2(n5094), .ZN(n4147) );
  INV_X1 U4669 ( .A(n4148), .ZN(n4176) );
  INV_X1 U4670 ( .A(n4149), .ZN(n4179) );
  INV_X1 U4671 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4152) );
  INV_X1 U4672 ( .A(n4150), .ZN(n4151) );
  NAND2_X1 U4673 ( .A1(n4152), .A2(n4151), .ZN(n4153) );
  NAND2_X1 U4674 ( .A1(n4179), .A2(n4153), .ZN(n6951) );
  AOI22_X1 U4675 ( .A1(n6951), .A2(n4550), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U4676 ( .A1(n4870), .A2(EAX_REG_3__SCAN_IN), .ZN(n4154) );
  OAI211_X1 U4677 ( .C1(n4176), .C2(n3712), .A(n4155), .B(n4154), .ZN(n4156)
         );
  INV_X1 U4678 ( .A(n4156), .ZN(n4157) );
  INV_X1 U4679 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5449) );
  AOI22_X1 U4680 ( .A1(n4448), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U4681 ( .A1(n4482), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U4682 ( .A1(n4487), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4683 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4717), .B1(n4719), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U4684 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4167)
         );
  AOI22_X1 U4685 ( .A1(n4721), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4686 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4465), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4687 ( .A1(n4726), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4688 ( .A1(n4017), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U4689 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4166)
         );
  NAND2_X1 U4690 ( .A1(n4700), .A2(n4590), .ZN(n4168) );
  NAND2_X1 U4691 ( .A1(n4171), .A2(n4170), .ZN(n4172) );
  NAND2_X1 U4692 ( .A1(n4196), .A2(n4172), .ZN(n4585) );
  INV_X1 U4693 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U4694 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4174)
         );
  NAND2_X1 U4695 ( .A1(n4870), .A2(EAX_REG_4__SCAN_IN), .ZN(n4173) );
  OAI211_X1 U4696 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4173), .ZN(n4182)
         );
  INV_X1 U4697 ( .A(n4177), .ZN(n4199) );
  INV_X1 U4698 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U4699 ( .A1(n4179), .A2(n4178), .ZN(n4180) );
  NAND2_X1 U4700 ( .A1(n4199), .A2(n4180), .ZN(n6966) );
  AND2_X1 U4701 ( .A1(n6966), .A2(n4550), .ZN(n4181) );
  AOI21_X1 U4702 ( .B1(n4182), .B2(n5289), .A(n4181), .ZN(n4183) );
  NAND2_X1 U4703 ( .A1(n5369), .A2(n5370), .ZN(n5001) );
  INV_X1 U4704 ( .A(n5001), .ZN(n4206) );
  INV_X1 U4705 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5455) );
  AOI22_X1 U4706 ( .A1(n4017), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4707 ( .A1(n4717), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4708 ( .A1(n4720), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4709 ( .A1(n4719), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U4710 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4193)
         );
  AOI22_X1 U4711 ( .A1(n4482), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U4712 ( .A1(n4721), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U4713 ( .A1(n4718), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4714 ( .A1(n4726), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4188) );
  NAND4_X1 U4715 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4192)
         );
  NAND2_X1 U4716 ( .A1(n4700), .A2(n4600), .ZN(n4194) );
  NAND2_X1 U4717 ( .A1(n4195), .A2(n4194), .ZN(n4207) );
  NAND2_X1 U4718 ( .A1(n4589), .A2(n4366), .ZN(n4205) );
  INV_X1 U4719 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4202) );
  INV_X1 U4720 ( .A(n4197), .ZN(n4226) );
  INV_X1 U4721 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4198) );
  NAND2_X1 U4722 ( .A1(n4199), .A2(n4198), .ZN(n4200) );
  NAND2_X1 U4723 ( .A1(n4226), .A2(n4200), .ZN(n6972) );
  AOI22_X1 U4724 ( .A1(n6972), .A2(n4550), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4201) );
  OAI21_X1 U4725 ( .B1(n4741), .B2(n4202), .A(n4201), .ZN(n4203) );
  INV_X1 U4726 ( .A(n4203), .ZN(n4204) );
  NAND2_X1 U4727 ( .A1(n4206), .A2(n5000), .ZN(n5247) );
  NAND2_X1 U4728 ( .A1(n4208), .A2(n4207), .ZN(n4224) );
  INV_X1 U4729 ( .A(n4224), .ZN(n4222) );
  INV_X1 U4730 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5431) );
  AOI22_X1 U4731 ( .A1(n4017), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U4732 ( .A1(n4717), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U4733 ( .A1(n4720), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U4734 ( .A1(n4719), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4209) );
  NAND4_X1 U4735 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4218)
         );
  AOI22_X1 U4736 ( .A1(n4482), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U4737 ( .A1(n4721), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U4738 ( .A1(n4718), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U4739 ( .A1(n4726), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U4740 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  NAND2_X1 U4741 ( .A1(n4700), .A2(n4609), .ZN(n4219) );
  NAND2_X1 U4742 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  INV_X1 U4743 ( .A(n4236), .ZN(n4228) );
  INV_X1 U4744 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4229) );
  NAND2_X1 U4745 ( .A1(n4226), .A2(n4229), .ZN(n4227) );
  NAND2_X1 U4746 ( .A1(n4228), .A2(n4227), .ZN(n6985) );
  INV_X1 U4747 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4230) );
  OAI22_X1 U4748 ( .A1(n4741), .A2(n4230), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4229), .ZN(n4231) );
  MUX2_X1 U4749 ( .A(n6985), .B(n4231), .S(n5289), .Z(n4232) );
  NAND2_X1 U4750 ( .A1(n4700), .A2(n4620), .ZN(n4233) );
  OAI21_X1 U4751 ( .B1(n4234), .B2(n3749), .A(n4233), .ZN(n4235) );
  NAND2_X1 U4752 ( .A1(n4607), .A2(n4366), .ZN(n4240) );
  NAND2_X1 U4753 ( .A1(n4870), .A2(EAX_REG_7__SCAN_IN), .ZN(n4238) );
  OAI21_X1 U4754 ( .B1(n4236), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4251), 
        .ZN(n6994) );
  AOI22_X1 U4755 ( .A1(n6994), .A2(n4550), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4237) );
  AND2_X1 U4756 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  NAND2_X1 U4757 ( .A1(n4240), .A2(n4239), .ZN(n5322) );
  AOI22_X1 U4758 ( .A1(n4717), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U4759 ( .A1(n4482), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U4760 ( .A1(n4721), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4726), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U4761 ( .A1(n4718), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4241) );
  NAND4_X1 U4762 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(n4250)
         );
  AOI22_X1 U4763 ( .A1(n4017), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U4764 ( .A1(n4487), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U4765 ( .A1(n4720), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U4766 ( .A1(n4443), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4245) );
  NAND4_X1 U4767 ( .A1(n4248), .A2(n4247), .A3(n4246), .A4(n4245), .ZN(n4249)
         );
  NOR2_X1 U4768 ( .A1(n4250), .A2(n4249), .ZN(n4255) );
  NAND2_X1 U4769 ( .A1(n4870), .A2(EAX_REG_8__SCAN_IN), .ZN(n4254) );
  XNOR2_X1 U4770 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4251), .ZN(n7009) );
  INV_X1 U4771 ( .A(n7009), .ZN(n4252) );
  AOI22_X1 U4772 ( .A1(n4869), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4550), 
        .B2(n4252), .ZN(n4253) );
  OAI211_X1 U4773 ( .C1(n4255), .C2(n4330), .A(n4254), .B(n4253), .ZN(n5317)
         );
  XNOR2_X1 U4774 ( .A(n4256), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U4775 ( .A1(n4728), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4260) );
  AOI22_X1 U4776 ( .A1(n4721), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4259) );
  AOI22_X1 U4777 ( .A1(n4448), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U4778 ( .A1(n4726), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4257) );
  NAND4_X1 U4779 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), .ZN(n4266)
         );
  AOI22_X1 U4780 ( .A1(n4017), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U4781 ( .A1(n4720), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4782 ( .A1(n4717), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U4783 ( .A1(n4465), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4261) );
  NAND4_X1 U4784 ( .A1(n4264), .A2(n4263), .A3(n4262), .A4(n4261), .ZN(n4265)
         );
  OAI21_X1 U4785 ( .B1(n4266), .B2(n4265), .A(n4366), .ZN(n4269) );
  NAND2_X1 U4786 ( .A1(n4870), .A2(EAX_REG_9__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U4787 ( .A1(n4869), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4267)
         );
  NAND3_X1 U4788 ( .A1(n4269), .A2(n4268), .A3(n4267), .ZN(n4270) );
  AOI21_X1 U4789 ( .B1(n7019), .B2(n4550), .A(n4270), .ZN(n5397) );
  XNOR2_X1 U4790 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4272), .ZN(n6020)
         );
  INV_X1 U4791 ( .A(n6020), .ZN(n4287) );
  AOI22_X1 U4792 ( .A1(n4717), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4793 ( .A1(n4720), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4794 ( .A1(n4721), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U4795 ( .A1(n4719), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4273) );
  NAND4_X1 U4796 ( .A1(n4276), .A2(n4275), .A3(n4274), .A4(n4273), .ZN(n4282)
         );
  AOI22_X1 U4797 ( .A1(n4017), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U4798 ( .A1(n4482), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U4799 ( .A1(n4465), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U4800 ( .A1(n4726), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4277) );
  NAND4_X1 U4801 ( .A1(n4280), .A2(n4279), .A3(n4278), .A4(n4277), .ZN(n4281)
         );
  OAI21_X1 U4802 ( .B1(n4282), .B2(n4281), .A(n4366), .ZN(n4285) );
  NAND2_X1 U4803 ( .A1(n4870), .A2(EAX_REG_10__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U4804 ( .A1(n4869), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4283)
         );
  NAND3_X1 U4805 ( .A1(n4285), .A2(n4284), .A3(n4283), .ZN(n4286) );
  AOI21_X1 U4806 ( .B1(n4287), .B2(n4550), .A(n4286), .ZN(n5539) );
  AOI22_X1 U4807 ( .A1(n4448), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U4808 ( .A1(n4482), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4290) );
  AOI22_X1 U4809 ( .A1(n4720), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4289) );
  AOI22_X1 U4810 ( .A1(n4726), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4288) );
  NAND4_X1 U4811 ( .A1(n4291), .A2(n4290), .A3(n4289), .A4(n4288), .ZN(n4297)
         );
  AOI22_X1 U4812 ( .A1(n4017), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4717), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4813 ( .A1(n4721), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4294) );
  AOI22_X1 U4814 ( .A1(n4728), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U4815 ( .A1(n4718), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4292) );
  NAND4_X1 U4816 ( .A1(n4295), .A2(n4294), .A3(n4293), .A4(n4292), .ZN(n4296)
         );
  NOR2_X1 U4817 ( .A1(n4297), .A2(n4296), .ZN(n4301) );
  XNOR2_X1 U4818 ( .A(n4298), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n7032)
         );
  NAND2_X1 U4819 ( .A1(n7032), .A2(n4550), .ZN(n4300) );
  AOI22_X1 U4820 ( .A1(n4870), .A2(EAX_REG_11__SCAN_IN), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4299) );
  OAI211_X1 U4821 ( .C1(n4301), .C2(n4330), .A(n4300), .B(n4299), .ZN(n5627)
         );
  XNOR2_X1 U4822 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4302), .ZN(n7042)
         );
  NAND2_X1 U4823 ( .A1(n7042), .A2(n4550), .ZN(n4306) );
  INV_X1 U4824 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4304) );
  OAI21_X1 U4825 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n7413), .A(n3887), 
        .ZN(n4303) );
  OAI21_X1 U4826 ( .B1(n4741), .B2(n4304), .A(n4303), .ZN(n4305) );
  NAND2_X1 U4827 ( .A1(n4306), .A2(n4305), .ZN(n4318) );
  AOI22_X1 U4828 ( .A1(n4726), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U4829 ( .A1(n4482), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U4830 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4487), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U4831 ( .A1(n4465), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4307) );
  NAND4_X1 U4832 ( .A1(n4310), .A2(n4309), .A3(n4308), .A4(n4307), .ZN(n4316)
         );
  AOI22_X1 U4833 ( .A1(n4016), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U4834 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4717), .B1(n4720), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U4835 ( .A1(n4728), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4836 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4721), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4311) );
  NAND4_X1 U4837 ( .A1(n4314), .A2(n4313), .A3(n4312), .A4(n4311), .ZN(n4315)
         );
  OAI21_X1 U4838 ( .B1(n4316), .B2(n4315), .A(n4366), .ZN(n4317) );
  NAND2_X1 U4839 ( .A1(n4318), .A2(n4317), .ZN(n5625) );
  AOI22_X1 U4840 ( .A1(n4016), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4841 ( .A1(n4717), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4842 ( .A1(n4720), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U4843 ( .A1(n4719), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4319) );
  NAND4_X1 U4844 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4328)
         );
  AOI22_X1 U4845 ( .A1(n4482), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4846 ( .A1(n4721), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4847 ( .A1(n4718), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U4848 ( .A1(n4726), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U4849 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4327)
         );
  NOR2_X1 U4850 ( .A1(n4328), .A2(n4327), .ZN(n4329) );
  NOR2_X1 U4851 ( .A1(n4330), .A2(n4329), .ZN(n4334) );
  XNOR2_X1 U4852 ( .A(n4331), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6085)
         );
  NAND2_X1 U4853 ( .A1(n6085), .A2(n4550), .ZN(n4333) );
  AOI22_X1 U4854 ( .A1(n4870), .A2(EAX_REG_13__SCAN_IN), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U4855 ( .A1(n4333), .A2(n4332), .ZN(n6045) );
  INV_X1 U4856 ( .A(n4334), .ZN(n4335) );
  INV_X1 U4857 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4341) );
  AOI21_X1 U4858 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n4338), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4339) );
  INV_X1 U4859 ( .A(n4339), .ZN(n4340) );
  OAI21_X1 U4860 ( .B1(n4741), .B2(n4341), .A(n4340), .ZN(n4344) );
  XNOR2_X1 U4861 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4342), .ZN(n7055)
         );
  NAND2_X1 U4862 ( .A1(n7055), .A2(n4550), .ZN(n4343) );
  NAND2_X1 U4863 ( .A1(n4344), .A2(n4343), .ZN(n4356) );
  AOI22_X1 U4864 ( .A1(n4448), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4865 ( .A1(n4465), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U4866 ( .A1(n4721), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4867 ( .A1(n4005), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4345) );
  NAND4_X1 U4868 ( .A1(n4348), .A2(n4347), .A3(n4346), .A4(n4345), .ZN(n4354)
         );
  AOI22_X1 U4869 ( .A1(n4017), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U4870 ( .A1(n4728), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4726), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4351) );
  AOI22_X1 U4871 ( .A1(n4717), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4872 ( .A1(n4720), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4349) );
  NAND4_X1 U4873 ( .A1(n4352), .A2(n4351), .A3(n4350), .A4(n4349), .ZN(n4353)
         );
  OAI21_X1 U4874 ( .B1(n4354), .B2(n4353), .A(n4366), .ZN(n4355) );
  NAND2_X1 U4875 ( .A1(n4356), .A2(n4355), .ZN(n6060) );
  XOR2_X1 U4876 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4357), .Z(n6266) );
  INV_X1 U4877 ( .A(n6266), .ZN(n6445) );
  AOI22_X1 U4878 ( .A1(n4448), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U4879 ( .A1(n4717), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U4880 ( .A1(n4721), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4881 ( .A1(n4465), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4358) );
  NAND4_X1 U4882 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4368)
         );
  AOI22_X1 U4883 ( .A1(n4482), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4884 ( .A1(n4016), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4885 ( .A1(n4720), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U4886 ( .A1(n4726), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4362) );
  NAND4_X1 U4887 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4367)
         );
  OAI21_X1 U4888 ( .B1(n4368), .B2(n4367), .A(n4366), .ZN(n4371) );
  NAND2_X1 U4889 ( .A1(n4870), .A2(EAX_REG_15__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U4890 ( .A1(n4869), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4369)
         );
  NAND3_X1 U4891 ( .A1(n4371), .A2(n4370), .A3(n4369), .ZN(n4372) );
  AOI21_X1 U4892 ( .B1(n6445), .B2(n4550), .A(n4372), .ZN(n6258) );
  XNOR2_X1 U4893 ( .A(n4374), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7068)
         );
  INV_X1 U4894 ( .A(n7068), .ZN(n6435) );
  AOI22_X1 U4895 ( .A1(n4016), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4896 ( .A1(n4465), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4897 ( .A1(n4721), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U4898 ( .A1(n4482), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4375) );
  NAND4_X1 U4899 ( .A1(n4378), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4384)
         );
  AOI22_X1 U4900 ( .A1(n4717), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4901 ( .A1(n4720), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U4902 ( .A1(n4726), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4380) );
  AOI22_X1 U4903 ( .A1(n4728), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4379) );
  NAND4_X1 U4904 ( .A1(n4382), .A2(n4381), .A3(n4380), .A4(n4379), .ZN(n4383)
         );
  NOR2_X1 U4905 ( .A1(n4384), .A2(n4383), .ZN(n4386) );
  AOI22_X1 U4906 ( .A1(n4870), .A2(EAX_REG_16__SCAN_IN), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U4907 ( .B1(n4540), .B2(n4386), .A(n4385), .ZN(n4387) );
  AOI21_X1 U4908 ( .B1(n6435), .B2(n4550), .A(n4387), .ZN(n6313) );
  OR2_X1 U4909 ( .A1(n4389), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4390)
         );
  NAND2_X1 U4910 ( .A1(n4390), .A2(n4419), .ZN(n7082) );
  AOI22_X1 U4911 ( .A1(n4017), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U4912 ( .A1(n4717), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U4913 ( .A1(n4465), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4914 ( .A1(n4718), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4391) );
  NAND4_X1 U4915 ( .A1(n4394), .A2(n4393), .A3(n4392), .A4(n4391), .ZN(n4400)
         );
  AOI22_X1 U4916 ( .A1(n4482), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U4917 ( .A1(n4721), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4918 ( .A1(n4720), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4919 ( .A1(n4726), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4395) );
  NAND4_X1 U4920 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(n4399)
         );
  NOR2_X1 U4921 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  NOR2_X1 U4922 ( .A1(n4540), .A2(n4401), .ZN(n4405) );
  INV_X1 U4923 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U4924 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4402)
         );
  OAI211_X1 U4925 ( .C1(n4741), .C2(n4403), .A(n5289), .B(n4402), .ZN(n4404)
         );
  OAI22_X1 U4926 ( .A1(n7082), .A2(n5289), .B1(n4405), .B2(n4404), .ZN(n6306)
         );
  NAND2_X1 U4927 ( .A1(n4540), .A2(n5289), .ZN(n4495) );
  AOI22_X1 U4928 ( .A1(n4017), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U4929 ( .A1(n4726), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4407)
         );
  NAND2_X1 U4930 ( .A1(n4487), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4406) );
  AND3_X1 U4931 ( .A1(n4407), .A2(n4406), .A3(n5289), .ZN(n4410) );
  AOI22_X1 U4932 ( .A1(n4728), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U4933 ( .A1(n4465), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U4934 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4417)
         );
  AOI22_X1 U4935 ( .A1(n4448), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4936 ( .A1(n4717), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4937 ( .A1(n4721), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4938 ( .A1(n4443), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U4939 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4416)
         );
  OR2_X1 U4940 ( .A1(n4417), .A2(n4416), .ZN(n4418) );
  NAND2_X1 U4941 ( .A1(n4495), .A2(n4418), .ZN(n4422) );
  AOI22_X1 U4942 ( .A1(n4870), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3887), .ZN(n4421) );
  XNOR2_X1 U4943 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4419), .ZN(n7090)
         );
  AND2_X1 U4944 ( .A1(n7090), .A2(n4550), .ZN(n4420) );
  AOI21_X1 U4945 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n6299) );
  INV_X1 U4946 ( .A(n4442), .ZN(n4425) );
  OR2_X1 U4947 ( .A1(n4423), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4424)
         );
  NAND2_X1 U4948 ( .A1(n4425), .A2(n4424), .ZN(n7104) );
  AOI22_X1 U4949 ( .A1(n4720), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4429) );
  AOI22_X1 U4950 ( .A1(n4482), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4951 ( .A1(n4721), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U4952 ( .A1(n4448), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4426) );
  NAND4_X1 U4953 ( .A1(n4429), .A2(n4428), .A3(n4427), .A4(n4426), .ZN(n4435)
         );
  AOI22_X1 U4954 ( .A1(n4016), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U4955 ( .A1(n4717), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4956 ( .A1(n4726), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U4957 ( .A1(n4718), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4430) );
  NAND4_X1 U4958 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4434)
         );
  NOR2_X1 U4959 ( .A1(n4435), .A2(n4434), .ZN(n4436) );
  NOR2_X1 U4960 ( .A1(n4540), .A2(n4436), .ZN(n4440) );
  INV_X1 U4961 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U4962 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4437)
         );
  OAI211_X1 U4963 ( .C1(n4741), .C2(n4438), .A(n5289), .B(n4437), .ZN(n4439)
         );
  OAI22_X1 U4964 ( .A1(n7104), .A2(n5289), .B1(n4440), .B2(n4439), .ZN(n6753)
         );
  INV_X1 U4965 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n7117) );
  XNOR2_X1 U4966 ( .A(n4442), .B(n7117), .ZN(n7114) );
  NAND2_X1 U4967 ( .A1(n7114), .A2(n4550), .ZN(n4460) );
  AOI22_X1 U4968 ( .A1(n4016), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U4969 ( .A1(n4721), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4487), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U4970 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4465), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U4971 ( .A1(n4727), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4444) );
  NAND4_X1 U4972 ( .A1(n4447), .A2(n4446), .A3(n4445), .A4(n4444), .ZN(n4456)
         );
  AOI22_X1 U4973 ( .A1(n4448), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U4974 ( .A1(n4717), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U4975 ( .A1(n4726), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4449)
         );
  AND3_X1 U4976 ( .A1(n4450), .A2(n4449), .A3(n5289), .ZN(n4453) );
  AOI22_X1 U4977 ( .A1(n4718), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U4978 ( .A1(n4482), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4451) );
  NAND4_X1 U4979 ( .A1(n4454), .A2(n4453), .A3(n4452), .A4(n4451), .ZN(n4455)
         );
  OAI21_X1 U4980 ( .B1(n4456), .B2(n4455), .A(n4495), .ZN(n4458) );
  AOI22_X1 U4981 ( .A1(n4870), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3887), .ZN(n4457) );
  NAND2_X1 U4982 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U4983 ( .A1(n4460), .A2(n4459), .ZN(n6294) );
  NAND2_X1 U4984 ( .A1(n4462), .A2(n4461), .ZN(n6291) );
  AND2_X1 U4985 ( .A1(n4463), .A2(n6412), .ZN(n4464) );
  OR2_X1 U4986 ( .A1(n4464), .A2(n4481), .ZN(n7128) );
  AOI22_X1 U4987 ( .A1(n4017), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U4988 ( .A1(n4465), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4468) );
  AOI22_X1 U4989 ( .A1(n3941), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U4990 ( .A1(n4487), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4466) );
  NAND4_X1 U4991 ( .A1(n4469), .A2(n4468), .A3(n4467), .A4(n4466), .ZN(n4476)
         );
  AOI22_X1 U4992 ( .A1(n4717), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U4993 ( .A1(n4721), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U4994 ( .A1(n4728), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U4995 ( .A1(n4726), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U4996 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4475)
         );
  NOR2_X1 U4997 ( .A1(n4476), .A2(n4475), .ZN(n4479) );
  OAI21_X1 U4998 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6412), .A(n5289), .ZN(
        n4477) );
  AOI21_X1 U4999 ( .B1(n4870), .B2(EAX_REG_21__SCAN_IN), .A(n4477), .ZN(n4478)
         );
  OAI21_X1 U5000 ( .B1(n4540), .B2(n4479), .A(n4478), .ZN(n4480) );
  OAI21_X1 U5001 ( .B1(n7128), .B2(n5289), .A(n4480), .ZN(n6408) );
  INV_X1 U5002 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6404) );
  XNOR2_X1 U5003 ( .A(n4481), .B(n6404), .ZN(n7134) );
  AOI22_X1 U5004 ( .A1(n4870), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n3887), .ZN(n4499) );
  AOI22_X1 U5005 ( .A1(n4717), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4482), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5006 ( .A1(n4728), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5007 ( .A1(n4448), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5008 ( .A1(n4727), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4483) );
  NAND4_X1 U5009 ( .A1(n4486), .A2(n4485), .A3(n4484), .A4(n4483), .ZN(n4497)
         );
  INV_X1 U5010 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5434) );
  AOI22_X1 U5011 ( .A1(n4726), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4489) );
  AOI21_X1 U5012 ( .B1(n4487), .B2(INSTQUEUE_REG_1__6__SCAN_IN), .A(n4550), 
        .ZN(n4488) );
  OAI211_X1 U5013 ( .C1(n4490), .C2(n5434), .A(n4489), .B(n4488), .ZN(n4491)
         );
  INV_X1 U5014 ( .A(n4491), .ZN(n4494) );
  AOI22_X1 U5015 ( .A1(n4017), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4465), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U5016 ( .A1(n4720), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4492) );
  NAND3_X1 U5017 ( .A1(n4494), .A2(n4493), .A3(n4492), .ZN(n4496) );
  OAI21_X1 U5018 ( .B1(n4497), .B2(n4496), .A(n4495), .ZN(n4498) );
  AOI22_X1 U5019 ( .A1(n7134), .A2(n4550), .B1(n4499), .B2(n4498), .ZN(n6281)
         );
  INV_X1 U5020 ( .A(n4500), .ZN(n4501) );
  OAI21_X1 U5021 ( .B1(n4501), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4510), 
        .ZN(n7158) );
  INV_X1 U5022 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4506) );
  INV_X1 U5023 ( .A(n4540), .ZN(n4743) );
  OAI211_X1 U5024 ( .C1(n4503), .C2(n4502), .A(n4743), .B(n4509), .ZN(n4505)
         );
  AOI21_X1 U5025 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n3887), .A(n4550), 
        .ZN(n4504) );
  OAI211_X1 U5026 ( .C1(n4741), .C2(n4506), .A(n4505), .B(n4504), .ZN(n4507)
         );
  OAI21_X1 U5027 ( .B1(n7158), .B2(n5289), .A(n4507), .ZN(n6275) );
  XNOR2_X1 U5028 ( .A(n4509), .B(n4508), .ZN(n4514) );
  INV_X1 U5029 ( .A(n4510), .ZN(n4511) );
  XNOR2_X1 U5030 ( .A(n4511), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6390)
         );
  NAND2_X1 U5031 ( .A1(n6390), .A2(n4550), .ZN(n4513) );
  AOI22_X1 U5032 ( .A1(n4870), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4869), .ZN(n4512) );
  OAI211_X1 U5033 ( .C1(n4514), .C2(n4540), .A(n4513), .B(n4512), .ZN(n6244)
         );
  INV_X1 U5034 ( .A(n4515), .ZN(n4517) );
  INV_X1 U5035 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5036 ( .A1(n4517), .A2(n4516), .ZN(n4518) );
  NAND2_X1 U5037 ( .A1(n4525), .A2(n4518), .ZN(n6377) );
  XNOR2_X1 U5038 ( .A(n4520), .B(n4519), .ZN(n4523) );
  OAI21_X1 U5039 ( .B1(n7413), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n3887), 
        .ZN(n4522) );
  NAND2_X1 U5040 ( .A1(n4870), .A2(EAX_REG_25__SCAN_IN), .ZN(n4521) );
  OAI211_X1 U5041 ( .C1(n4540), .C2(n4523), .A(n4522), .B(n4521), .ZN(n4524)
         );
  XNOR2_X1 U5042 ( .A(n4525), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6226)
         );
  AOI21_X1 U5043 ( .B1(n4526), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4527) );
  AOI21_X1 U5044 ( .B1(n4870), .B2(EAX_REG_26__SCAN_IN), .A(n4527), .ZN(n4532)
         );
  XOR2_X1 U5045 ( .A(n4529), .B(n4528), .Z(n4530) );
  NAND2_X1 U5046 ( .A1(n4530), .A2(n4743), .ZN(n4531) );
  NAND2_X1 U5047 ( .A1(n4534), .A2(n4533), .ZN(n4535) );
  NAND2_X1 U5048 ( .A1(n4543), .A2(n4535), .ZN(n6362) );
  XNOR2_X1 U5049 ( .A(n4537), .B(n4536), .ZN(n4541) );
  AOI21_X1 U5050 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n3887), .A(n4550), 
        .ZN(n4539) );
  NAND2_X1 U5051 ( .A1(n4870), .A2(EAX_REG_27__SCAN_IN), .ZN(n4538) );
  OAI211_X1 U5052 ( .C1(n4541), .C2(n4540), .A(n4539), .B(n4538), .ZN(n4542)
         );
  OAI21_X1 U5053 ( .B1(n6362), .B2(n5289), .A(n4542), .ZN(n6211) );
  XNOR2_X1 U5054 ( .A(n4543), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6124)
         );
  INV_X1 U5055 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6127) );
  NOR2_X1 U5056 ( .A1(n6127), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4544) );
  AOI211_X1 U5057 ( .C1(n4870), .C2(EAX_REG_28__SCAN_IN), .A(n4550), .B(n4544), 
        .ZN(n4549) );
  XOR2_X1 U5058 ( .A(n4546), .B(n4545), .Z(n4547) );
  NAND2_X1 U5059 ( .A1(n4547), .A2(n4743), .ZN(n4548) );
  NOR2_X1 U5060 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7164), .ZN(n5287) );
  NAND2_X1 U5061 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5287), .ZN(n6833) );
  NAND2_X1 U5062 ( .A1(n4561), .A2(n4553), .ZN(n4567) );
  OAI21_X1 U5063 ( .B1(n4561), .B2(n4553), .A(n4567), .ZN(n4557) );
  INV_X1 U5064 ( .A(n4555), .ZN(n4556) );
  OAI211_X1 U5065 ( .C1(n4557), .C2(n4554), .A(n4556), .B(n4665), .ZN(n4558)
         );
  INV_X1 U5066 ( .A(n4558), .ZN(n4559) );
  OAI21_X1 U5067 ( .B1(n4554), .B2(n4561), .A(n4955), .ZN(n4562) );
  INV_X1 U5068 ( .A(n4562), .ZN(n4563) );
  OAI21_X1 U5069 ( .B1(n6118), .B2(n4747), .A(n4563), .ZN(n5009) );
  AND2_X1 U5070 ( .A1(n5009), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5010)
         );
  NAND2_X1 U5071 ( .A1(n4976), .A2(n5010), .ZN(n4565) );
  NAND2_X1 U5072 ( .A1(n6774), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4574)
         );
  INV_X1 U5073 ( .A(n5137), .ZN(n5087) );
  INV_X1 U5074 ( .A(n4566), .ZN(n4568) );
  NAND2_X1 U5075 ( .A1(n4567), .A2(n4568), .ZN(n4577) );
  OAI21_X1 U5076 ( .B1(n4568), .B2(n4567), .A(n4577), .ZN(n4571) );
  NAND2_X1 U5077 ( .A1(n4571), .A2(n4570), .ZN(n4572) );
  NAND2_X1 U5078 ( .A1(n4572), .A2(n4955), .ZN(n4573) );
  NAND2_X1 U5079 ( .A1(n4574), .A2(n6775), .ZN(n4576) );
  INV_X1 U5080 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4770) );
  INV_X1 U5081 ( .A(n5084), .ZN(n5333) );
  NAND2_X1 U5082 ( .A1(n4577), .A2(n4578), .ZN(n4592) );
  OAI211_X1 U5083 ( .C1(n4578), .C2(n4577), .A(n4592), .B(n4570), .ZN(n4579)
         );
  INV_X1 U5084 ( .A(n4579), .ZN(n4580) );
  AOI21_X1 U5085 ( .B1(n5333), .B2(n4694), .A(n4580), .ZN(n6781) );
  NAND2_X1 U5086 ( .A1(n4582), .A2(n4581), .ZN(n6786) );
  XNOR2_X1 U5087 ( .A(n4592), .B(n4590), .ZN(n4583) );
  NAND2_X1 U5088 ( .A1(n4583), .A2(n4570), .ZN(n4584) );
  OAI21_X2 U5089 ( .B1(n4585), .B2(n4747), .A(n4584), .ZN(n4587) );
  XNOR2_X1 U5090 ( .A(n4587), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6785)
         );
  INV_X1 U5091 ( .A(n6785), .ZN(n4586) );
  NAND2_X1 U5092 ( .A1(n4587), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4588)
         );
  NAND2_X1 U5093 ( .A1(n4589), .A2(n4694), .ZN(n4595) );
  INV_X1 U5094 ( .A(n4590), .ZN(n4591) );
  OR2_X1 U5095 ( .A1(n4592), .A2(n4591), .ZN(n4599) );
  XNOR2_X1 U5096 ( .A(n4599), .B(n4600), .ZN(n4593) );
  NAND2_X1 U5097 ( .A1(n4593), .A2(n4570), .ZN(n4594) );
  NAND2_X1 U5098 ( .A1(n4595), .A2(n4594), .ZN(n4596) );
  INV_X1 U5099 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5240) );
  XNOR2_X1 U5100 ( .A(n4596), .B(n5240), .ZN(n5238) );
  NAND2_X1 U5101 ( .A1(n4596), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4597)
         );
  INV_X1 U5102 ( .A(n4598), .ZN(n4604) );
  INV_X1 U5103 ( .A(n4599), .ZN(n4601) );
  NAND2_X1 U5104 ( .A1(n4601), .A2(n4600), .ZN(n4608) );
  XNOR2_X1 U5105 ( .A(n4608), .B(n4609), .ZN(n4602) );
  NAND2_X1 U5106 ( .A1(n4602), .A2(n4570), .ZN(n4603) );
  OAI21_X1 U5107 ( .B1(n4604), .B2(n4747), .A(n4603), .ZN(n4605) );
  OR2_X1 U5108 ( .A1(n4605), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5384)
         );
  NAND2_X1 U5109 ( .A1(n5383), .A2(n5384), .ZN(n4606) );
  NAND2_X1 U5110 ( .A1(n4605), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5385)
         );
  NAND2_X1 U5111 ( .A1(n4606), .A2(n5385), .ZN(n5616) );
  NAND2_X1 U5112 ( .A1(n4607), .A2(n4694), .ZN(n4613) );
  INV_X1 U5113 ( .A(n4608), .ZN(n4610) );
  NAND2_X1 U5114 ( .A1(n4610), .A2(n4609), .ZN(n4622) );
  XNOR2_X1 U5115 ( .A(n4622), .B(n4620), .ZN(n4611) );
  NAND2_X1 U5116 ( .A1(n4611), .A2(n4570), .ZN(n4612) );
  INV_X1 U5117 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U5118 ( .A1(n4614), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4615)
         );
  INV_X1 U5119 ( .A(n4617), .ZN(n4618) );
  NAND2_X1 U5120 ( .A1(n4570), .A2(n4620), .ZN(n4621) );
  OR2_X1 U5121 ( .A1(n4622), .A2(n4621), .ZN(n4623) );
  NAND2_X1 U5122 ( .A1(n4628), .A2(n4623), .ZN(n4624) );
  INV_X1 U5123 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5561) );
  XNOR2_X1 U5124 ( .A(n4624), .B(n5561), .ZN(n5558) );
  NAND2_X1 U5125 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4625)
         );
  XNOR2_X1 U5126 ( .A(n3633), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6010)
         );
  NAND2_X1 U5127 ( .A1(n6009), .A2(n6010), .ZN(n4627) );
  NAND2_X1 U5128 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4626)
         );
  INV_X1 U5129 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U5130 ( .A1(n3633), .A2(n4794), .ZN(n6014) );
  INV_X1 U5131 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6904) );
  AND2_X1 U5132 ( .A1(n3633), .A2(n6904), .ZN(n6024) );
  INV_X1 U5133 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4631) );
  OR2_X1 U5134 ( .A1(n3633), .A2(n6904), .ZN(n6067) );
  OR2_X1 U5135 ( .A1(n3633), .A2(n4794), .ZN(n6022) );
  OAI211_X1 U5136 ( .C1(n3633), .C2(n4631), .A(n6067), .B(n6022), .ZN(n4629)
         );
  INV_X1 U5137 ( .A(n4629), .ZN(n4630) );
  NAND2_X1 U5138 ( .A1(n3633), .A2(n4631), .ZN(n4632) );
  NAND2_X1 U5139 ( .A1(n4633), .A2(n4632), .ZN(n6082) );
  XNOR2_X1 U5140 ( .A(n3633), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6083)
         );
  INV_X1 U5141 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5142 ( .A1(n3633), .A2(n4634), .ZN(n4635) );
  NAND2_X1 U5143 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6091) );
  INV_X1 U5144 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6612) );
  NOR2_X1 U5145 ( .A1(n3633), .A2(n6612), .ZN(n6442) );
  NAND2_X1 U5146 ( .A1(n3633), .A2(n6612), .ZN(n6440) );
  INV_X1 U5147 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5148 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6457) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6912) );
  INV_X1 U5150 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6596) );
  NAND3_X1 U5151 ( .A1(n6606), .A2(n6912), .A3(n6596), .ZN(n4637) );
  NAND2_X1 U5152 ( .A1(n6426), .A2(n4637), .ZN(n4638) );
  NOR2_X1 U5153 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6579) );
  NOR2_X1 U5154 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6384) );
  INV_X1 U5155 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4639) );
  INV_X1 U5156 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4837) );
  NAND4_X1 U5157 ( .A1(n6579), .A2(n6384), .A3(n4639), .A4(n4837), .ZN(n4640)
         );
  NAND2_X1 U5158 ( .A1(n6426), .A2(n4640), .ZN(n4641) );
  AND2_X1 U5159 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6578) );
  AND2_X1 U5160 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U5161 ( .A1(n6578), .A2(n6475), .ZN(n6393) );
  NAND2_X1 U5162 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U5163 ( .B1(n6393), .B2(n6477), .A(n3633), .ZN(n4642) );
  INV_X1 U5164 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6537) );
  XNOR2_X1 U5165 ( .A(n3633), .B(n6537), .ZN(n6375) );
  NAND2_X1 U5166 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4643) );
  INV_X1 U5167 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U5168 ( .A1(n3633), .A2(n6526), .ZN(n4644) );
  INV_X1 U5169 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U5170 ( .A1(n3633), .A2(n6508), .ZN(n4645) );
  INV_X1 U5171 ( .A(n4888), .ZN(n4648) );
  NAND2_X1 U5172 ( .A1(n6426), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4647) );
  NOR2_X1 U5173 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4646) );
  OR2_X1 U5174 ( .A1(n3633), .A2(n4646), .ZN(n4887) );
  NAND2_X1 U5175 ( .A1(n4647), .A2(n4887), .ZN(n4861) );
  INV_X1 U5176 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4854) );
  XNOR2_X1 U5177 ( .A(n3633), .B(n4854), .ZN(n4860) );
  XNOR2_X1 U5178 ( .A(n4649), .B(n4860), .ZN(n6504) );
  INV_X1 U5179 ( .A(n6504), .ZN(n4706) );
  NAND2_X1 U5180 ( .A1(n7412), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5181 ( .A1(n3707), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U5182 ( .A1(n4651), .A2(n4650), .ZN(n4671) );
  NAND2_X1 U5183 ( .A1(n3651), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U5184 ( .A1(n4655), .A2(n4652), .ZN(n4682) );
  AOI222_X1 U5185 ( .A1(n4657), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n4657), .B2(n4175), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n4175), 
        .ZN(n4900) );
  AND2_X1 U5186 ( .A1(n4657), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4658)
         );
  NAND2_X1 U5187 ( .A1(n4658), .A2(n4175), .ZN(n4898) );
  XNOR2_X1 U5188 ( .A(n4660), .B(n4659), .ZN(n4897) );
  INV_X1 U5189 ( .A(n4897), .ZN(n4661) );
  AOI21_X1 U5190 ( .B1(n4898), .B2(n4661), .A(n4686), .ZN(n4698) );
  OAI21_X1 U5191 ( .B1(n7417), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n4670), 
        .ZN(n4662) );
  INV_X1 U5192 ( .A(n4662), .ZN(n4663) );
  AOI21_X1 U5193 ( .B1(n4663), .B2(n4700), .A(n4701), .ZN(n4669) );
  OAI21_X1 U5194 ( .B1(n4664), .B2(n3687), .A(n4663), .ZN(n4667) );
  NAND2_X1 U5195 ( .A1(n4750), .A2(n4665), .ZN(n4666) );
  NAND2_X1 U5196 ( .A1(n6003), .A2(n4666), .ZN(n4688) );
  AOI21_X1 U5197 ( .B1(n3929), .B2(n4667), .A(n4688), .ZN(n4668) );
  NOR2_X1 U5198 ( .A1(n4669), .A2(n4668), .ZN(n4681) );
  INV_X1 U5199 ( .A(n4701), .ZN(n4675) );
  NAND2_X1 U5200 ( .A1(n4671), .A2(n4670), .ZN(n4672) );
  NAND2_X1 U5201 ( .A1(n4673), .A2(n4672), .ZN(n4895) );
  NOR2_X1 U5202 ( .A1(n4895), .A2(n7224), .ZN(n4676) );
  INV_X1 U5203 ( .A(n4676), .ZN(n4674) );
  NAND2_X1 U5204 ( .A1(n4675), .A2(n4674), .ZN(n4680) );
  INV_X1 U5205 ( .A(n4700), .ZN(n4689) );
  NAND2_X1 U5206 ( .A1(n4681), .A2(n4676), .ZN(n4678) );
  AOI21_X1 U5207 ( .B1(n4686), .B2(n4895), .A(n3687), .ZN(n4677) );
  OAI211_X1 U5208 ( .C1(n4689), .C2(n4750), .A(n4678), .B(n4677), .ZN(n4679)
         );
  OAI21_X1 U5209 ( .B1(n4681), .B2(n4680), .A(n4679), .ZN(n4691) );
  NAND2_X1 U5210 ( .A1(n4683), .A2(n4682), .ZN(n4685) );
  NAND2_X1 U5211 ( .A1(n4685), .A2(n4684), .ZN(n4896) );
  AOI21_X1 U5212 ( .B1(n4686), .B2(n4896), .A(n4688), .ZN(n4687) );
  NOR2_X1 U5213 ( .A1(n4691), .A2(n4687), .ZN(n4693) );
  INV_X1 U5214 ( .A(n4688), .ZN(n4690) );
  AOI211_X1 U5215 ( .C1(n4691), .C2(n4690), .A(n4689), .B(n4896), .ZN(n4692)
         );
  AOI211_X1 U5216 ( .C1(n4694), .C2(n4897), .A(n4693), .B(n4692), .ZN(n4697)
         );
  INV_X1 U5217 ( .A(n4898), .ZN(n4695) );
  AOI22_X1 U5218 ( .A1(n4695), .A2(n4701), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7224), .ZN(n4696) );
  OAI21_X1 U5219 ( .B1(n4698), .B2(n4697), .A(n4696), .ZN(n4699) );
  AOI21_X1 U5220 ( .B1(n4700), .B2(n4900), .A(n4699), .ZN(n4703) );
  AND2_X1 U5221 ( .A1(n4900), .A2(n4701), .ZN(n4702) );
  NOR2_X1 U5222 ( .A1(n4980), .A2(n3687), .ZN(n4704) );
  NOR2_X1 U5223 ( .A1(n4555), .A2(n5109), .ZN(n4958) );
  AND2_X1 U5224 ( .A1(n4704), .A2(n4958), .ZN(n4971) );
  NAND2_X1 U5225 ( .A1(n4707), .A2(n7426), .ZN(n6839) );
  NAND2_X1 U5226 ( .A1(n6839), .A2(n7224), .ZN(n4708) );
  NAND2_X1 U5227 ( .A1(n7224), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5228 ( .A1(n7413), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5229 ( .A1(n4710), .A2(n4709), .ZN(n5008) );
  INV_X2 U5230 ( .A(n6924), .ZN(n6908) );
  AND2_X1 U5231 ( .A1(n6908), .A2(REIP_REG_29__SCAN_IN), .ZN(n6498) );
  AOI21_X1 U5232 ( .B1(n4711), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6498), 
        .ZN(n4712) );
  OAI21_X1 U5233 ( .B1(n6199), .B2(n6822), .A(n4712), .ZN(n4713) );
  INV_X1 U5234 ( .A(n4713), .ZN(n4714) );
  OAI211_X1 U5235 ( .C1(n4716), .C2(n6791), .A(n4715), .B(n4714), .ZN(U2957)
         );
  XNOR2_X1 U5236 ( .A(n4874), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6348)
         );
  AOI22_X1 U5237 ( .A1(n4717), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5238 ( .A1(n4465), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5239 ( .A1(n4720), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U5240 ( .A1(n4721), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4005), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4722) );
  NAND4_X1 U5241 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4734)
         );
  AOI22_X1 U5242 ( .A1(n4017), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4448), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5243 ( .A1(n4726), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4443), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5244 ( .A1(n4728), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5245 ( .A1(n3941), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4470), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4729) );
  NAND4_X1 U5246 ( .A1(n4732), .A2(n4731), .A3(n4730), .A4(n4729), .ZN(n4733)
         );
  NOR2_X1 U5247 ( .A1(n4734), .A2(n4733), .ZN(n4738) );
  NOR2_X1 U5248 ( .A1(n4736), .A2(n4735), .ZN(n4737) );
  XNOR2_X1 U5249 ( .A(n4738), .B(n4737), .ZN(n4744) );
  INV_X1 U5250 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U5251 ( .A1(n3887), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4739)
         );
  OAI211_X1 U5252 ( .C1(n4741), .C2(n4740), .A(n4739), .B(n5289), .ZN(n4742)
         );
  AOI21_X1 U5253 ( .B1(n4744), .B2(n4743), .A(n4742), .ZN(n4745) );
  NOR2_X1 U5254 ( .A1(n4748), .A2(n4747), .ZN(n4940) );
  NAND2_X1 U5255 ( .A1(n6004), .A2(n6166), .ZN(n5025) );
  NAND3_X1 U5256 ( .A1(n6141), .A2(n3963), .A3(n4749), .ZN(n5359) );
  INV_X1 U5257 ( .A(n5359), .ZN(n4751) );
  OR2_X2 U5258 ( .A1(n4750), .A2(n5109), .ZN(n4763) );
  NAND3_X1 U5259 ( .A1(n3636), .A2(n4751), .A3(n5302), .ZN(n4752) );
  NAND2_X1 U5260 ( .A1(n5025), .A2(n4752), .ZN(n4753) );
  NAND2_X2 U5261 ( .A1(n6773), .A2(n5364), .ZN(n6315) );
  NAND2_X1 U5262 ( .A1(n3630), .A2(n4560), .ZN(n4755) );
  OAI211_X1 U5263 ( .C1(n4763), .C2(EBX_REG_1__SCAN_IN), .A(n4755), .B(n4856), 
        .ZN(n4757) );
  INV_X1 U5264 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U5265 ( .A1(n4765), .A2(n5311), .ZN(n4756) );
  NAND2_X1 U5266 ( .A1(n3631), .A2(EBX_REG_0__SCAN_IN), .ZN(n4759) );
  INV_X1 U5267 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U5268 ( .A1(n4856), .A2(n5377), .ZN(n4758) );
  NAND2_X1 U5269 ( .A1(n4759), .A2(n4758), .ZN(n4907) );
  XNOR2_X1 U5270 ( .A(n4760), .B(n4907), .ZN(n4982) );
  INV_X1 U5271 ( .A(n4760), .ZN(n4761) );
  NAND2_X1 U5272 ( .A1(n4761), .A2(n4907), .ZN(n4762) );
  INV_X1 U5273 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U5274 ( .A1(n3630), .A2(n6878), .ZN(n4764) );
  OAI211_X1 U5275 ( .C1(n4763), .C2(EBX_REG_2__SCAN_IN), .A(n4764), .B(n4856), 
        .ZN(n4767) );
  INV_X1 U5276 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U5277 ( .A1(n4765), .A2(n6926), .ZN(n4766) );
  AND2_X1 U5278 ( .A1(n4767), .A2(n4766), .ZN(n4917) );
  MUX2_X1 U5279 ( .A(n4841), .B(n4856), .S(EBX_REG_3__SCAN_IN), .Z(n4772) );
  NAND2_X1 U5280 ( .A1(n4949), .A2(n4770), .ZN(n4771) );
  NAND2_X1 U5281 ( .A1(n4772), .A2(n4771), .ZN(n4937) );
  INV_X1 U5282 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4773) );
  NAND2_X1 U5283 ( .A1(n3630), .A2(n4773), .ZN(n4774) );
  OAI211_X1 U5284 ( .C1(n4763), .C2(EBX_REG_4__SCAN_IN), .A(n4774), .B(n4856), 
        .ZN(n4776) );
  INV_X1 U5285 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U5286 ( .A1(n4947), .A2(n6772), .ZN(n4775) );
  NAND2_X1 U5287 ( .A1(n4776), .A2(n4775), .ZN(n6766) );
  NAND2_X1 U5288 ( .A1(n6768), .A2(n6766), .ZN(n5004) );
  INV_X1 U5289 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U5290 ( .A1(n4848), .A2(n6969), .ZN(n4779) );
  NAND2_X1 U5291 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4777)
         );
  OAI211_X1 U5292 ( .C1(n4763), .C2(EBX_REG_5__SCAN_IN), .A(n3631), .B(n4777), 
        .ZN(n4778) );
  NAND2_X1 U5293 ( .A1(n4779), .A2(n4778), .ZN(n5003) );
  INV_X1 U5294 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U5295 ( .A1(n3630), .A2(n4782), .ZN(n4783) );
  OAI211_X1 U5296 ( .C1(n4763), .C2(EBX_REG_6__SCAN_IN), .A(n4783), .B(n4856), 
        .ZN(n4785) );
  INV_X1 U5297 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U5298 ( .A1(n4947), .A2(n6980), .ZN(n4784) );
  MUX2_X1 U5299 ( .A(n4848), .B(n4765), .S(EBX_REG_7__SCAN_IN), .Z(n4787) );
  NOR2_X1 U5300 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4786)
         );
  NOR2_X1 U5301 ( .A1(n4787), .A2(n4786), .ZN(n5325) );
  NAND2_X1 U5302 ( .A1(n3631), .A2(n5561), .ZN(n4788) );
  OAI211_X1 U5303 ( .C1(n4763), .C2(EBX_REG_8__SCAN_IN), .A(n4788), .B(n4856), 
        .ZN(n4790) );
  INV_X1 U5304 ( .A(EBX_REG_8__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U5305 ( .A1(n4947), .A2(n7006), .ZN(n4789) );
  NAND2_X1 U5306 ( .A1(n4790), .A2(n4789), .ZN(n5319) );
  INV_X1 U5307 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U5308 ( .A1(n4848), .A2(n6751), .ZN(n4793) );
  NAND2_X1 U5309 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4791)
         );
  OAI211_X1 U5310 ( .C1(n4763), .C2(EBX_REG_9__SCAN_IN), .A(n3630), .B(n4791), 
        .ZN(n4792) );
  NAND2_X1 U5311 ( .A1(n4793), .A2(n4792), .ZN(n6749) );
  NAND2_X1 U5312 ( .A1(n3631), .A2(n4794), .ZN(n4795) );
  OAI211_X1 U5313 ( .C1(n4763), .C2(EBX_REG_10__SCAN_IN), .A(n4795), .B(n4856), 
        .ZN(n4797) );
  INV_X1 U5314 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U5315 ( .A1(n4947), .A2(n5548), .ZN(n4796) );
  MUX2_X1 U5316 ( .A(n4848), .B(n4947), .S(EBX_REG_11__SCAN_IN), .Z(n4799) );
  NOR2_X1 U5317 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4798)
         );
  NOR2_X1 U5318 ( .A1(n4799), .A2(n4798), .ZN(n5630) );
  MUX2_X1 U5319 ( .A(n4841), .B(n4856), .S(EBX_REG_13__SCAN_IN), .Z(n4801) );
  NAND2_X1 U5320 ( .A1(n4949), .A2(n4634), .ZN(n4800) );
  NAND2_X1 U5321 ( .A1(n4801), .A2(n4800), .ZN(n6046) );
  NAND2_X1 U5322 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U5323 ( .A1(n3630), .A2(n4802), .ZN(n4803) );
  OAI21_X1 U5324 ( .B1(n4763), .B2(EBX_REG_12__SCAN_IN), .A(n4803), .ZN(n4805)
         );
  OR2_X1 U5325 ( .A1(n4856), .A2(EBX_REG_12__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U5326 ( .A1(n3631), .A2(n6455), .ZN(n4808) );
  OAI211_X1 U5327 ( .C1(n4763), .C2(EBX_REG_14__SCAN_IN), .A(n4808), .B(n4856), 
        .ZN(n4810) );
  INV_X1 U5328 ( .A(EBX_REG_14__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U5329 ( .A1(n4947), .A2(n7058), .ZN(n4809) );
  NOR2_X2 U5330 ( .A1(n6062), .A2(n6061), .ZN(n6260) );
  INV_X1 U5331 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U5332 ( .A1(n4848), .A2(n6765), .ZN(n4813) );
  NAND2_X1 U5333 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4811) );
  OAI211_X1 U5334 ( .C1(n4763), .C2(EBX_REG_15__SCAN_IN), .A(n3630), .B(n4811), 
        .ZN(n4812) );
  NAND2_X1 U5335 ( .A1(n6260), .A2(n6259), .ZN(n6317) );
  NAND2_X1 U5336 ( .A1(n3631), .A2(n6606), .ZN(n4814) );
  OAI211_X1 U5337 ( .C1(n4763), .C2(EBX_REG_16__SCAN_IN), .A(n4814), .B(n4856), 
        .ZN(n4816) );
  INV_X1 U5338 ( .A(EBX_REG_16__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U5339 ( .A1(n4947), .A2(n7071), .ZN(n4815) );
  MUX2_X1 U5340 ( .A(n4841), .B(n4856), .S(EBX_REG_17__SCAN_IN), .Z(n4818) );
  NAND2_X1 U5341 ( .A1(n4949), .A2(n6912), .ZN(n4817) );
  NAND2_X1 U5342 ( .A1(n4818), .A2(n4817), .ZN(n6308) );
  NAND2_X1 U5343 ( .A1(n3630), .A2(n6596), .ZN(n4819) );
  OAI211_X1 U5344 ( .C1(n4763), .C2(EBX_REG_18__SCAN_IN), .A(n4819), .B(n4856), 
        .ZN(n4821) );
  INV_X1 U5345 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U5346 ( .A1(n4947), .A2(n7093), .ZN(n4820) );
  NAND2_X1 U5347 ( .A1(n4821), .A2(n4820), .ZN(n6300) );
  INV_X1 U5348 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U5349 ( .A1(n4848), .A2(n6760), .ZN(n4824) );
  NAND2_X1 U5350 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4822) );
  OAI211_X1 U5351 ( .C1(n4763), .C2(EBX_REG_19__SCAN_IN), .A(n3631), .B(n4822), 
        .ZN(n4823) );
  NAND2_X1 U5352 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U5353 ( .A1(n3630), .A2(n4825), .ZN(n4826) );
  OAI21_X1 U5354 ( .B1(n4763), .B2(EBX_REG_20__SCAN_IN), .A(n4826), .ZN(n4828)
         );
  OR2_X1 U5355 ( .A1(n4856), .A2(EBX_REG_20__SCAN_IN), .ZN(n4827) );
  INV_X1 U5356 ( .A(EBX_REG_21__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U5357 ( .A1(n4848), .A2(n7121), .ZN(n4831) );
  NAND2_X1 U5358 ( .A1(n4856), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4829) );
  OAI211_X1 U5359 ( .C1(n4763), .C2(EBX_REG_21__SCAN_IN), .A(n3631), .B(n4829), 
        .ZN(n4830) );
  NAND2_X1 U5360 ( .A1(n4831), .A2(n4830), .ZN(n6569) );
  OR2_X2 U5361 ( .A1(n6568), .A2(n6569), .ZN(n6566) );
  INV_X1 U5362 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U5363 ( .A1(n3630), .A2(n6401), .ZN(n4832) );
  OAI211_X1 U5364 ( .C1(n4763), .C2(EBX_REG_22__SCAN_IN), .A(n4832), .B(n4856), 
        .ZN(n4834) );
  INV_X1 U5365 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5366 ( .A1(n4947), .A2(n6286), .ZN(n4833) );
  MUX2_X1 U5367 ( .A(n4848), .B(n4947), .S(EBX_REG_23__SCAN_IN), .Z(n4836) );
  NOR2_X1 U5368 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4835)
         );
  NOR2_X1 U5369 ( .A1(n4836), .A2(n4835), .ZN(n6277) );
  NAND2_X1 U5370 ( .A1(n6282), .A2(n6277), .ZN(n6250) );
  NAND2_X1 U5371 ( .A1(n3631), .A2(n4837), .ZN(n4838) );
  OAI211_X1 U5372 ( .C1(n4763), .C2(EBX_REG_24__SCAN_IN), .A(n4838), .B(n4856), 
        .ZN(n4840) );
  INV_X1 U5373 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U5374 ( .A1(n4765), .A2(n6246), .ZN(n4839) );
  AND2_X1 U5375 ( .A1(n4840), .A2(n4839), .ZN(n6252) );
  MUX2_X1 U5376 ( .A(n4841), .B(n4856), .S(EBX_REG_25__SCAN_IN), .Z(n4843) );
  NAND2_X1 U5377 ( .A1(n4949), .A2(n6537), .ZN(n4842) );
  NAND2_X1 U5378 ( .A1(n4843), .A2(n4842), .ZN(n6235) );
  NAND2_X1 U5379 ( .A1(n3630), .A2(n6526), .ZN(n4844) );
  OAI211_X1 U5380 ( .C1(n4763), .C2(EBX_REG_26__SCAN_IN), .A(n4844), .B(n4856), 
        .ZN(n4847) );
  INV_X1 U5381 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U5382 ( .A1(n4947), .A2(n4845), .ZN(n4846) );
  NAND2_X1 U5383 ( .A1(n4847), .A2(n4846), .ZN(n6221) );
  MUX2_X1 U5384 ( .A(n4848), .B(n4947), .S(EBX_REG_27__SCAN_IN), .Z(n4850) );
  NOR2_X1 U5385 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4849)
         );
  NOR2_X1 U5386 ( .A1(n4850), .A2(n4849), .ZN(n6208) );
  INV_X1 U5387 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U5388 ( .A1(n3631), .A2(n6507), .ZN(n4851) );
  OAI211_X1 U5389 ( .C1(n4763), .C2(EBX_REG_28__SCAN_IN), .A(n4851), .B(n4856), 
        .ZN(n4853) );
  OR2_X1 U5390 ( .A1(n4856), .A2(EBX_REG_28__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5391 ( .A1(n4853), .A2(n4852), .ZN(n6121) );
  AND2_X2 U5392 ( .A1(n6120), .A2(n6121), .ZN(n6123) );
  INV_X1 U5393 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U5394 ( .A1(n4949), .A2(n4854), .B1(n5302), .B2(n4881), .ZN(n4857)
         );
  NAND2_X1 U5395 ( .A1(n4857), .A2(n4856), .ZN(n4855) );
  OAI21_X1 U5396 ( .B1(EBX_REG_29__SCAN_IN), .B2(n4856), .A(n4855), .ZN(n4880)
         );
  OAI22_X1 U5397 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n4763), .ZN(n6174) );
  INV_X1 U5398 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6188) );
  OAI21_X1 U5399 ( .B1(n6494), .B2(n6320), .A(n3648), .ZN(n4858) );
  INV_X1 U5400 ( .A(n4858), .ZN(n4859) );
  OAI21_X1 U5401 ( .B1(n6356), .B2(n6315), .A(n4859), .ZN(U2829) );
  AOI21_X1 U5402 ( .B1(n4888), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4860), 
        .ZN(n4866) );
  AND2_X1 U5403 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U5404 ( .A1(n6506), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U5405 ( .A1(n3633), .A2(n6488), .ZN(n4862) );
  AOI21_X2 U5406 ( .B1(n6357), .B2(n4862), .A(n4861), .ZN(n6350) );
  NAND2_X1 U5407 ( .A1(n6350), .A2(n4854), .ZN(n6349) );
  AND2_X1 U5408 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5409 ( .A1(n6349), .A2(n4864), .ZN(n4865) );
  NAND2_X1 U5410 ( .A1(n4866), .A2(n4865), .ZN(n4867) );
  INV_X1 U5411 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U5412 ( .A1(n4746), .A2(n4868), .ZN(n4873) );
  AOI22_X1 U5413 ( .A1(n4870), .A2(EAX_REG_31__SCAN_IN), .B1(n4869), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4871) );
  INV_X1 U5414 ( .A(n4871), .ZN(n4872) );
  XNOR2_X2 U5415 ( .A(n4873), .B(n4872), .ZN(n6172) );
  NAND2_X1 U5416 ( .A1(n6172), .A2(n6818), .ZN(n4879) );
  INV_X1 U5417 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6346) );
  INV_X1 U5418 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6184) );
  INV_X1 U5419 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U5420 ( .A1(n6924), .A2(n6718), .ZN(n6480) );
  AOI21_X1 U5421 ( .B1(n4711), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6480), 
        .ZN(n4876) );
  OAI21_X1 U5422 ( .B1(n5295), .B2(n6822), .A(n4876), .ZN(n4877) );
  INV_X1 U5423 ( .A(n4877), .ZN(n4878) );
  OAI21_X1 U5424 ( .B1(n6123), .B2(n4880), .A(n6175), .ZN(n6500) );
  NOR2_X1 U5425 ( .A1(n6119), .A2(n6791), .ZN(n4894) );
  NAND2_X1 U5426 ( .A1(n4888), .A2(n4887), .ZN(n4890) );
  XNOR2_X1 U5427 ( .A(n3633), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4889)
         );
  XNOR2_X1 U5428 ( .A(n4890), .B(n4889), .ZN(n6514) );
  NAND2_X1 U5429 ( .A1(n6908), .A2(REIP_REG_28__SCAN_IN), .ZN(n6505) );
  OAI21_X1 U5430 ( .B1(n6448), .B2(n6127), .A(n6505), .ZN(n4891) );
  OR2_X1 U5431 ( .A1(n4894), .A2(n4893), .ZN(U2958) );
  NOR3_X1 U5432 ( .A1(n4897), .A2(n4896), .A3(n4895), .ZN(n4899) );
  OAI21_X1 U5433 ( .B1(n4900), .B2(n4899), .A(n4898), .ZN(n6165) );
  NOR2_X1 U5434 ( .A1(n6164), .A2(n7206), .ZN(n4902) );
  NAND2_X1 U5435 ( .A1(n6165), .A2(n4902), .ZN(n5285) );
  INV_X1 U5436 ( .A(n5285), .ZN(n4906) );
  INV_X1 U5437 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7248) );
  NOR2_X1 U5438 ( .A1(n4904), .A2(n7206), .ZN(n4905) );
  OAI211_X1 U5439 ( .C1(n4906), .C2(n7248), .A(n5286), .B(n6160), .ZN(U2788)
         );
  INV_X1 U5440 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U5441 ( .A1(n4949), .A2(n6151), .ZN(n4908) );
  AND2_X1 U5442 ( .A1(n4908), .A2(n4907), .ZN(n6916) );
  INV_X1 U5443 ( .A(n6916), .ZN(n4912) );
  OAI21_X1 U5444 ( .B1(n4911), .B2(n4910), .A(n4909), .ZN(n5381) );
  OAI222_X1 U5445 ( .A1(n4912), .A2(n6320), .B1(n5377), .B2(n6773), .C1(n5381), 
        .C2(n6315), .ZN(U2859) );
  INV_X1 U5446 ( .A(n4913), .ZN(n4914) );
  OAI21_X1 U5447 ( .B1(n4916), .B2(n4915), .A(n4914), .ZN(n6931) );
  NAND2_X1 U5448 ( .A1(n4918), .A2(n4917), .ZN(n4919) );
  AND2_X1 U5449 ( .A1(n4938), .A2(n4919), .ZN(n6935) );
  AOI22_X1 U5450 ( .A1(n6769), .A2(n6935), .B1(EBX_REG_2__SCAN_IN), .B2(n6311), 
        .ZN(n4920) );
  OAI21_X1 U5451 ( .B1(n6931), .B2(n6315), .A(n4920), .ZN(U2857) );
  OR2_X1 U5452 ( .A1(n5040), .A2(n4554), .ZN(n7202) );
  NOR2_X1 U5453 ( .A1(n7202), .A2(n7206), .ZN(n4922) );
  NOR2_X1 U5454 ( .A1(n6164), .A2(n4750), .ZN(n7159) );
  NAND3_X1 U5455 ( .A1(n6170), .A2(n7221), .A3(n7159), .ZN(n4923) );
  NAND2_X1 U5456 ( .A1(n7333), .A2(n4923), .ZN(n4924) );
  OR2_X1 U5457 ( .A1(n7237), .A2(STATE_REG_0__SCAN_IN), .ZN(n6831) );
  INV_X1 U5458 ( .A(n6831), .ZN(n6006) );
  NAND2_X1 U5459 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5287), .ZN(n7200) );
  INV_X2 U5460 ( .A(n7200), .ZN(n6668) );
  NOR2_X4 U5461 ( .A1(n6668), .A2(n6652), .ZN(n6649) );
  AOI22_X1 U5462 ( .A1(n6668), .A2(UWORD_REG_7__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4925) );
  OAI21_X1 U5463 ( .B1(n4506), .B2(n5284), .A(n4925), .ZN(U2900) );
  INV_X1 U5464 ( .A(EAX_REG_29__SCAN_IN), .ZN(n7321) );
  AOI22_X1 U5465 ( .A1(n6668), .A2(UWORD_REG_13__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4926) );
  OAI21_X1 U5466 ( .B1(n7321), .B2(n5284), .A(n4926), .ZN(U2894) );
  INV_X1 U5467 ( .A(EAX_REG_24__SCAN_IN), .ZN(n7292) );
  AOI22_X1 U5468 ( .A1(n6668), .A2(UWORD_REG_8__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4927) );
  OAI21_X1 U5469 ( .B1(n7292), .B2(n5284), .A(n4927), .ZN(U2899) );
  INV_X1 U5470 ( .A(EAX_REG_27__SCAN_IN), .ZN(n7310) );
  AOI22_X1 U5471 ( .A1(n6668), .A2(UWORD_REG_11__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4928) );
  OAI21_X1 U5472 ( .B1(n7310), .B2(n5284), .A(n4928), .ZN(U2896) );
  INV_X1 U5473 ( .A(EAX_REG_28__SCAN_IN), .ZN(n7316) );
  AOI22_X1 U5474 ( .A1(n6668), .A2(UWORD_REG_12__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4929) );
  OAI21_X1 U5475 ( .B1(n7316), .B2(n5284), .A(n4929), .ZN(U2895) );
  INV_X1 U5476 ( .A(EAX_REG_25__SCAN_IN), .ZN(n7298) );
  AOI22_X1 U5477 ( .A1(n6668), .A2(UWORD_REG_9__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4930) );
  OAI21_X1 U5478 ( .B1(n7298), .B2(n5284), .A(n4930), .ZN(U2898) );
  INV_X1 U5479 ( .A(EAX_REG_26__SCAN_IN), .ZN(n7304) );
  AOI22_X1 U5480 ( .A1(n6668), .A2(UWORD_REG_10__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4931) );
  OAI21_X1 U5481 ( .B1(n7304), .B2(n5284), .A(n4931), .ZN(U2897) );
  INV_X1 U5482 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7279) );
  AOI22_X1 U5483 ( .A1(n6668), .A2(UWORD_REG_5__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4932) );
  OAI21_X1 U5484 ( .B1(n7279), .B2(n5284), .A(n4932), .ZN(U2902) );
  INV_X1 U5485 ( .A(EAX_REG_20__SCAN_IN), .ZN(n7274) );
  AOI22_X1 U5486 ( .A1(n6668), .A2(UWORD_REG_4__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4933) );
  OAI21_X1 U5487 ( .B1(n7274), .B2(n5284), .A(n4933), .ZN(U2903) );
  INV_X1 U5488 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7284) );
  AOI22_X1 U5489 ( .A1(n6668), .A2(UWORD_REG_6__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4934) );
  OAI21_X1 U5490 ( .B1(n7284), .B2(n5284), .A(n4934), .ZN(U2901) );
  INV_X1 U5491 ( .A(n4935), .ZN(n4936) );
  XNOR2_X1 U5492 ( .A(n4913), .B(n4936), .ZN(n6944) );
  INV_X1 U5493 ( .A(n6944), .ZN(n5368) );
  AOI21_X1 U5494 ( .B1(n4938), .B2(n4937), .A(n6768), .ZN(n6939) );
  AOI22_X1 U5495 ( .A1(n6769), .A2(n6939), .B1(EBX_REG_3__SCAN_IN), .B2(n6311), 
        .ZN(n4939) );
  OAI21_X1 U5496 ( .B1(n5368), .B2(n6315), .A(n4939), .ZN(U2856) );
  INV_X1 U5497 ( .A(n4940), .ZN(n4967) );
  NAND2_X1 U5498 ( .A1(n4750), .A2(n6831), .ZN(n5298) );
  NAND2_X1 U5499 ( .A1(n5298), .A2(n7250), .ZN(n5017) );
  OAI21_X1 U5500 ( .B1(n3966), .B2(n5109), .A(n5403), .ZN(n4941) );
  OAI21_X1 U5501 ( .B1(n5040), .B2(n5017), .A(n4941), .ZN(n4942) );
  NAND2_X1 U5502 ( .A1(n6170), .A2(n4942), .ZN(n4966) );
  NAND2_X1 U5503 ( .A1(n4943), .A2(n3929), .ZN(n4945) );
  MUX2_X1 U5504 ( .A(n4554), .B(n4945), .S(n4944), .Z(n4954) );
  AOI21_X1 U5505 ( .B1(n3966), .B2(n5109), .A(n5403), .ZN(n4946) );
  AOI21_X1 U5506 ( .B1(n4948), .B2(n4947), .A(n4946), .ZN(n4952) );
  NAND2_X1 U5507 ( .A1(n5109), .A2(n3970), .ZN(n6005) );
  OR2_X1 U5508 ( .A1(n6005), .A2(n3625), .ZN(n5021) );
  NAND2_X1 U5509 ( .A1(n4949), .A2(n5021), .ZN(n4950) );
  NAND2_X1 U5510 ( .A1(n4950), .A2(n4555), .ZN(n4951) );
  AND2_X1 U5511 ( .A1(n4952), .A2(n4951), .ZN(n4953) );
  NAND2_X1 U5512 ( .A1(n4954), .A2(n4953), .ZN(n5041) );
  OAI21_X1 U5513 ( .B1(n4956), .B2(n4955), .A(n5071), .ZN(n4957) );
  NOR2_X1 U5514 ( .A1(n5041), .A2(n4957), .ZN(n4984) );
  INV_X1 U5515 ( .A(n7161), .ZN(n4960) );
  INV_X1 U5516 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U5517 ( .A1(n4960), .A2(n4959), .ZN(n4961) );
  NAND2_X1 U5518 ( .A1(n4984), .A2(n4961), .ZN(n4962) );
  NAND2_X1 U5519 ( .A1(n4962), .A2(n6164), .ZN(n5022) );
  NAND2_X1 U5520 ( .A1(n7250), .A2(n6165), .ZN(n5014) );
  INV_X1 U5521 ( .A(n5014), .ZN(n4963) );
  OAI211_X1 U5522 ( .C1(n4750), .C2(n6006), .A(n3625), .B(n4963), .ZN(n4964)
         );
  AND2_X1 U5523 ( .A1(n5022), .A2(n4964), .ZN(n4965) );
  OAI211_X1 U5524 ( .C1(n6170), .C2(n4967), .A(n4966), .B(n4965), .ZN(n4968)
         );
  NOR2_X1 U5525 ( .A1(n6003), .A2(n4969), .ZN(n4970) );
  NOR2_X1 U5526 ( .A1(n5045), .A2(n4971), .ZN(n6163) );
  OAI21_X1 U5527 ( .B1(n4972), .B2(n3963), .A(n5039), .ZN(n4973) );
  INV_X1 U5528 ( .A(n4973), .ZN(n4974) );
  OAI211_X1 U5529 ( .C1(n4904), .C2(n4750), .A(n6163), .B(n4974), .ZN(n4975)
         );
  NAND2_X1 U5530 ( .A1(n4976), .A2(n4977), .ZN(n4978) );
  XOR2_X1 U5531 ( .A(n5010), .B(n4978), .Z(n5118) );
  OAI21_X1 U5532 ( .B1(n4979), .B2(n4980), .A(n7202), .ZN(n4981) );
  XNOR2_X1 U5533 ( .A(n4982), .B(n5302), .ZN(n4998) );
  NAND2_X1 U5534 ( .A1(n4984), .A2(n4983), .ZN(n4985) );
  NAND2_X1 U5535 ( .A1(n6093), .A2(n6151), .ZN(n4988) );
  INV_X1 U5536 ( .A(n4990), .ZN(n4986) );
  NAND2_X1 U5537 ( .A1(n4986), .A2(n6924), .ZN(n4987) );
  INV_X1 U5538 ( .A(n6587), .ZN(n4989) );
  AOI21_X1 U5539 ( .B1(n6870), .B2(n6151), .A(n4989), .ZN(n6918) );
  NAND2_X1 U5540 ( .A1(n6908), .A2(REIP_REG_1__SCAN_IN), .ZN(n5113) );
  OAI21_X1 U5541 ( .B1(n6918), .B2(n4560), .A(n5113), .ZN(n4992) );
  NAND2_X1 U5542 ( .A1(n6589), .A2(n6471), .ZN(n6467) );
  NOR2_X1 U5543 ( .A1(n6921), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5241)
         );
  NOR3_X1 U5544 ( .A1(n6603), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5241), 
        .ZN(n4991) );
  AOI211_X1 U5545 ( .C1(n6917), .C2(n4998), .A(n4992), .B(n4991), .ZN(n4993)
         );
  OAI21_X1 U5546 ( .B1(n6619), .B2(n5118), .A(n4993), .ZN(U3017) );
  OR2_X1 U5547 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  NAND2_X1 U5548 ( .A1(n4994), .A2(n4997), .ZN(n5373) );
  AOI22_X1 U5549 ( .A1(n6769), .A2(n4998), .B1(EBX_REG_1__SCAN_IN), .B2(n6311), 
        .ZN(n4999) );
  OAI21_X1 U5550 ( .B1(n6315), .B2(n5373), .A(n4999), .ZN(U2858) );
  INV_X1 U5551 ( .A(n5000), .ZN(n5002) );
  XNOR2_X1 U5552 ( .A(n5002), .B(n5001), .ZN(n6971) );
  NAND2_X1 U5553 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NAND2_X1 U5554 ( .A1(n5252), .A2(n5005), .ZN(n6968) );
  INV_X1 U5555 ( .A(n6968), .ZN(n5006) );
  AOI22_X1 U5556 ( .A1(n6769), .A2(n5006), .B1(EBX_REG_5__SCAN_IN), .B2(n6311), 
        .ZN(n5007) );
  OAI21_X1 U5557 ( .B1(n6971), .B2(n6315), .A(n5007), .ZN(U2854) );
  OAI21_X1 U5558 ( .B1(n4711), .B2(n5008), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5013) );
  INV_X1 U5559 ( .A(n5009), .ZN(n5011) );
  AOI21_X1 U5560 ( .B1(n5011), .B2(n6151), .A(n5010), .ZN(n6914) );
  AOI22_X1 U5561 ( .A1(n6819), .A2(n6914), .B1(n6908), .B2(REIP_REG_0__SCAN_IN), .ZN(n5012) );
  OAI211_X1 U5562 ( .C1(n5381), .C2(n6791), .A(n5013), .B(n5012), .ZN(U2986)
         );
  NAND2_X1 U5563 ( .A1(n6170), .A2(n5045), .ZN(n5016) );
  INV_X1 U5564 ( .A(n5361), .ZN(n5027) );
  NAND2_X1 U5565 ( .A1(n4904), .A2(n6831), .ZN(n5020) );
  INV_X1 U5566 ( .A(n7159), .ZN(n5018) );
  AOI21_X1 U5567 ( .B1(n5018), .B2(n5040), .A(n5017), .ZN(n5019) );
  AND2_X1 U5568 ( .A1(n5020), .A2(n5019), .ZN(n5024) );
  NAND2_X1 U5569 ( .A1(n5022), .A2(n5021), .ZN(n5023) );
  AOI21_X1 U5570 ( .B1(n6170), .B2(n5024), .A(n5023), .ZN(n5026) );
  NAND3_X1 U5571 ( .A1(n5027), .A2(n5026), .A3(n5025), .ZN(n7175) );
  MUX2_X1 U5572 ( .A(n7175), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5028) );
  INV_X1 U5573 ( .A(n5028), .ZN(n5034) );
  INV_X1 U5574 ( .A(n5029), .ZN(n5030) );
  NOR2_X1 U5575 ( .A1(n5031), .A2(n5030), .ZN(n5032) );
  XNOR2_X1 U5576 ( .A(n5032), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6960)
         );
  OR2_X1 U5577 ( .A1(n5039), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5033) );
  NOR2_X1 U5578 ( .A1(n6960), .A2(n5033), .ZN(n7170) );
  AOI21_X1 U5579 ( .B1(n5034), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n7170), 
        .ZN(n7198) );
  INV_X1 U5580 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7192) );
  NAND2_X1 U5581 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7192), .ZN(n5035) );
  OAI21_X1 U5582 ( .B1(n7175), .B2(STATE2_REG_1__SCAN_IN), .A(n5035), .ZN(
        n5036) );
  NAND2_X1 U5583 ( .A1(n5036), .A2(n5050), .ZN(n5077) );
  INV_X1 U5584 ( .A(n5038), .ZN(n5044) );
  NAND3_X1 U5585 ( .A1(n5040), .A2(n5039), .A3(n4979), .ZN(n5042) );
  NOR2_X1 U5586 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  NAND2_X1 U5587 ( .A1(n5044), .A2(n5043), .ZN(n5067) );
  NAND2_X1 U5588 ( .A1(n7359), .A2(n5067), .ZN(n5065) );
  NAND2_X1 U5589 ( .A1(n7159), .A2(n3707), .ZN(n6149) );
  INV_X1 U5590 ( .A(n5045), .ZN(n5047) );
  INV_X1 U5591 ( .A(n6166), .ZN(n5046) );
  NAND2_X1 U5592 ( .A1(n5047), .A2(n5046), .ZN(n5068) );
  MUX2_X1 U5593 ( .A(n5048), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5049), 
        .Z(n5051) );
  NOR2_X1 U5594 ( .A1(n5051), .A2(n5050), .ZN(n5052) );
  NAND2_X1 U5595 ( .A1(n5068), .A2(n5052), .ZN(n5062) );
  INV_X1 U5596 ( .A(n5053), .ZN(n5056) );
  NAND2_X1 U5597 ( .A1(n5054), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U5598 ( .A1(n5056), .A2(n5055), .ZN(n5060) );
  INV_X1 U5599 ( .A(n5048), .ZN(n5057) );
  OAI211_X1 U5600 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n5049), .A(n5058), .B(n5057), .ZN(n6621) );
  NOR2_X1 U5601 ( .A1(n5071), .A2(n6621), .ZN(n5059) );
  AOI21_X1 U5602 ( .B1(n7159), .B2(n5060), .A(n5059), .ZN(n5061) );
  OAI211_X1 U5603 ( .C1(n6149), .C2(n3712), .A(n5062), .B(n5061), .ZN(n5063)
         );
  INV_X1 U5604 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U5605 ( .A1(n5065), .A2(n5064), .ZN(n7174) );
  INV_X1 U5606 ( .A(n5067), .ZN(n7160) );
  INV_X1 U5607 ( .A(n5068), .ZN(n5070) );
  XNOR2_X1 U5608 ( .A(n5049), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5069)
         );
  MUX2_X1 U5609 ( .A(n5071), .B(n5070), .S(n5069), .Z(n5074) );
  NAND2_X1 U5610 ( .A1(n7159), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5072) );
  MUX2_X1 U5611 ( .A(n5072), .B(n6149), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n5073) );
  AND2_X1 U5612 ( .A1(n5074), .A2(n5073), .ZN(n5075) );
  OAI21_X1 U5613 ( .B1(n5066), .B2(n7160), .A(n5075), .ZN(n7176) );
  NAND4_X1 U5614 ( .A1(n7175), .A2(n7164), .A3(n7174), .A4(n7176), .ZN(n5076)
         );
  NAND2_X1 U5615 ( .A1(n5077), .A2(n5076), .ZN(n7196) );
  INV_X1 U5616 ( .A(n5078), .ZN(n5079) );
  NAND2_X1 U5617 ( .A1(n7196), .A2(n5079), .ZN(n6111) );
  NAND3_X1 U5618 ( .A1(n7198), .A2(n7192), .A3(n6111), .ZN(n5080) );
  NAND2_X1 U5619 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n7211) );
  INV_X1 U5620 ( .A(n7211), .ZN(n6112) );
  NAND2_X1 U5621 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6112), .ZN(n7212) );
  INV_X1 U5622 ( .A(n7212), .ZN(n6835) );
  NAND2_X1 U5623 ( .A1(n5080), .A2(n6835), .ZN(n5082) );
  NAND2_X1 U5624 ( .A1(n7164), .A2(n3887), .ZN(n7216) );
  INV_X1 U5625 ( .A(n5413), .ZN(n5081) );
  INV_X1 U5626 ( .A(n7359), .ZN(n6942) );
  OAI21_X1 U5627 ( .B1(n7164), .B2(STATE2_REG_3__SCAN_IN), .A(n6647), .ZN(
        n6113) );
  INV_X1 U5628 ( .A(n7426), .ZN(n7415) );
  NAND2_X1 U5629 ( .A1(n6647), .A2(n7415), .ZN(n6117) );
  NOR2_X1 U5630 ( .A1(n5137), .A2(n4146), .ZN(n5158) );
  NAND2_X1 U5631 ( .A1(n5158), .A2(n3632), .ZN(n5178) );
  NOR2_X1 U5632 ( .A1(n5178), .A2(n7413), .ZN(n5198) );
  AND2_X1 U5633 ( .A1(n3632), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5119) );
  AOI21_X1 U5634 ( .B1(n5087), .B2(n5119), .A(n5084), .ZN(n5085) );
  NOR2_X1 U5635 ( .A1(n5198), .A2(n5085), .ZN(n5086) );
  OAI222_X1 U5636 ( .A1(n6647), .A2(n7361), .B1(n6942), .B2(n6113), .C1(n6117), 
        .C2(n5086), .ZN(U3462) );
  XNOR2_X1 U5637 ( .A(n5087), .B(n5119), .ZN(n5088) );
  OAI222_X1 U5638 ( .A1(n5088), .A2(n6117), .B1(n5066), .B2(n6113), .C1(n5327), 
        .C2(n6647), .ZN(U3463) );
  XNOR2_X1 U5639 ( .A(n3632), .B(STATEBS16_REG_SCAN_IN), .ZN(n5091) );
  INV_X1 U5640 ( .A(n5090), .ZN(n6150) );
  OAI222_X1 U5641 ( .A1(n6647), .A2(n7412), .B1(n6117), .B2(n5091), .C1(n6150), 
        .C2(n6113), .ZN(U3464) );
  OAI21_X1 U5642 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n7214), .A(n5413), 
        .ZN(n7424) );
  INV_X1 U5643 ( .A(n7424), .ZN(n7408) );
  INV_X1 U5644 ( .A(n5092), .ZN(n7363) );
  AND2_X1 U5645 ( .A1(n7359), .A2(n7363), .ZN(n7388) );
  NOR2_X1 U5646 ( .A1(n5066), .A2(n6150), .ZN(n5200) );
  NOR2_X1 U5647 ( .A1(n5093), .A2(n7361), .ZN(n5489) );
  AOI21_X1 U5648 ( .B1(n7388), .B2(n5200), .A(n5489), .ZN(n5098) );
  NOR2_X1 U5649 ( .A1(n5137), .A2(n5094), .ZN(n5259) );
  AND2_X1 U5650 ( .A1(n5259), .A2(n3632), .ZN(n5099) );
  NOR2_X1 U5651 ( .A1(n7426), .A2(STATEBS16_REG_SCAN_IN), .ZN(n7372) );
  INV_X1 U5652 ( .A(n7372), .ZN(n7400) );
  OAI21_X1 U5653 ( .B1(n5099), .B2(n6791), .A(n7400), .ZN(n5095) );
  NAND3_X1 U5654 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n5256) );
  AOI22_X1 U5655 ( .A1(n5098), .A2(n5095), .B1(n7426), .B2(n5256), .ZN(n5096)
         );
  INV_X1 U5656 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U5657 ( .A1(n6818), .A2(DATAI_19_), .ZN(n5211) );
  INV_X1 U5658 ( .A(n5211), .ZN(n7485) );
  NAND2_X1 U5659 ( .A1(n7224), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7213) );
  NOR2_X2 U5660 ( .A1(n5410), .A2(n4969), .ZN(n7483) );
  AOI22_X1 U5661 ( .A1(n7485), .A2(n5496), .B1(n7483), .B2(n5489), .ZN(n5101)
         );
  NAND2_X1 U5662 ( .A1(DATAI_3_), .A2(n5413), .ZN(n7488) );
  OAI22_X1 U5663 ( .A1(n5098), .A2(n7426), .B1(n5256), .B2(n3887), .ZN(n5490)
         );
  AOI22_X1 U5664 ( .A1(n5604), .A2(n5490), .B1(n7484), .B2(n5533), .ZN(n5100)
         );
  OAI211_X1 U5665 ( .C1(n5494), .C2(n5102), .A(n5101), .B(n5100), .ZN(U3143)
         );
  INV_X1 U5666 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U5667 ( .A1(n6818), .A2(DATAI_23_), .ZN(n5208) );
  INV_X1 U5668 ( .A(n5208), .ZN(n7572) );
  NOR2_X2 U5669 ( .A1(n5410), .A2(n6141), .ZN(n7571) );
  AOI22_X1 U5670 ( .A1(n7572), .A2(n5496), .B1(n7571), .B2(n5489), .ZN(n5104)
         );
  NAND2_X1 U5671 ( .A1(DATAI_7_), .A2(n5413), .ZN(n7578) );
  AOI22_X1 U5672 ( .A1(n5596), .A2(n5490), .B1(n7574), .B2(n5533), .ZN(n5103)
         );
  OAI211_X1 U5673 ( .C1(n5494), .C2(n5105), .A(n5104), .B(n5103), .ZN(U3147)
         );
  INV_X1 U5674 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U5675 ( .A1(n6818), .A2(DATAI_17_), .ZN(n5214) );
  INV_X1 U5676 ( .A(n5214), .ZN(n7452) );
  NOR2_X2 U5677 ( .A1(n5410), .A2(n4750), .ZN(n7451) );
  AOI22_X1 U5678 ( .A1(n7452), .A2(n5496), .B1(n7451), .B2(n5489), .ZN(n5107)
         );
  NAND2_X1 U5679 ( .A1(DATAI_1_), .A2(n5413), .ZN(n7456) );
  AOI22_X1 U5680 ( .A1(n5592), .A2(n5490), .B1(n7453), .B2(n5533), .ZN(n5106)
         );
  OAI211_X1 U5681 ( .C1(n5494), .C2(n5108), .A(n5107), .B(n5106), .ZN(U3141)
         );
  INV_X1 U5682 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5683 ( .A1(n6818), .A2(DATAI_16_), .ZN(n5217) );
  INV_X1 U5684 ( .A(n5217), .ZN(n7430) );
  NOR2_X2 U5685 ( .A1(n5410), .A2(n5109), .ZN(n7421) );
  AOI22_X1 U5686 ( .A1(n7430), .A2(n5496), .B1(n7421), .B2(n5489), .ZN(n5111)
         );
  NAND2_X1 U5687 ( .A1(DATAI_0_), .A2(n5413), .ZN(n7433) );
  AOI22_X1 U5688 ( .A1(n5600), .A2(n5490), .B1(n7422), .B2(n5533), .ZN(n5110)
         );
  OAI211_X1 U5689 ( .C1(n5494), .C2(n5112), .A(n5111), .B(n5110), .ZN(U3140)
         );
  NAND2_X1 U5690 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5114)
         );
  NAND2_X1 U5691 ( .A1(n5114), .A2(n5113), .ZN(n5116) );
  NOR2_X1 U5692 ( .A1(n5373), .A2(n6791), .ZN(n5115) );
  AOI211_X1 U5693 ( .C1(n6801), .C2(n5313), .A(n5116), .B(n5115), .ZN(n5117)
         );
  OAI21_X1 U5694 ( .B1(n6804), .B2(n5118), .A(n5117), .ZN(U2985) );
  NAND3_X1 U5695 ( .A1(n5332), .A2(n7371), .A3(n5084), .ZN(n5428) );
  NAND3_X1 U5696 ( .A1(n5084), .A2(n5119), .A3(n5137), .ZN(n5120) );
  NAND2_X1 U5697 ( .A1(n5120), .A2(n7415), .ZN(n5124) );
  NOR2_X1 U5698 ( .A1(n5092), .A2(n7359), .ZN(n7419) );
  AND2_X1 U5699 ( .A1(n5090), .A2(n5066), .ZN(n7360) );
  NOR2_X1 U5700 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7411) );
  INV_X1 U5701 ( .A(n7411), .ZN(n5134) );
  NOR2_X1 U5702 ( .A1(n5134), .A2(n5121), .ZN(n5425) );
  AOI21_X1 U5703 ( .B1(n7419), .B2(n7360), .A(n5425), .ZN(n5125) );
  INV_X1 U5704 ( .A(n5125), .ZN(n5123) );
  NAND2_X1 U5705 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7411), .ZN(n5572) );
  AOI21_X1 U5706 ( .B1(n7426), .B2(n5572), .A(n7424), .ZN(n5122) );
  OAI21_X1 U5707 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n5424) );
  OAI22_X1 U5708 ( .A1(n5125), .A2(n5124), .B1(n3887), .B2(n5572), .ZN(n5423)
         );
  AOI22_X1 U5709 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5424), .B1(n5600), 
        .B2(n5423), .ZN(n5127) );
  AOI22_X1 U5710 ( .A1(n7421), .A2(n5425), .B1(n7422), .B2(n5608), .ZN(n5126)
         );
  OAI211_X1 U5711 ( .C1(n5217), .C2(n5428), .A(n5127), .B(n5126), .ZN(U3044)
         );
  AOI22_X1 U5712 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5424), .B1(n5592), 
        .B2(n5423), .ZN(n5129) );
  AOI22_X1 U5713 ( .A1(n7451), .A2(n5425), .B1(n7453), .B2(n5608), .ZN(n5128)
         );
  OAI211_X1 U5714 ( .C1(n5214), .C2(n5428), .A(n5129), .B(n5128), .ZN(U3045)
         );
  AOI22_X1 U5715 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5424), .B1(n5604), 
        .B2(n5423), .ZN(n5131) );
  AOI22_X1 U5716 ( .A1(n7483), .A2(n5425), .B1(n7484), .B2(n5608), .ZN(n5130)
         );
  OAI211_X1 U5717 ( .C1(n5211), .C2(n5428), .A(n5131), .B(n5130), .ZN(U3047)
         );
  AOI22_X1 U5718 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5424), .B1(n5596), 
        .B2(n5423), .ZN(n5133) );
  AOI22_X1 U5719 ( .A1(n7571), .A2(n5425), .B1(n7574), .B2(n5608), .ZN(n5132)
         );
  OAI211_X1 U5720 ( .C1(n5208), .C2(n5428), .A(n5133), .B(n5132), .ZN(U3051)
         );
  NOR3_X2 U5721 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n5134), .ZN(n5495) );
  INV_X1 U5722 ( .A(n5495), .ZN(n5136) );
  INV_X1 U5723 ( .A(n5342), .ZN(n5135) );
  NOR2_X1 U5724 ( .A1(n5341), .A2(n5135), .ZN(n5143) );
  NOR2_X1 U5725 ( .A1(n5143), .A2(n3887), .ZN(n5218) );
  OR2_X1 U5726 ( .A1(n5142), .A2(n3887), .ZN(n5340) );
  NAND2_X1 U5727 ( .A1(n5413), .A2(n5340), .ZN(n7379) );
  AOI211_X1 U5728 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5136), .A(n5218), .B(
        n7379), .ZN(n5141) );
  AND2_X1 U5729 ( .A1(n5066), .A2(n6150), .ZN(n7418) );
  INV_X1 U5730 ( .A(n7418), .ZN(n5184) );
  NAND2_X1 U5731 ( .A1(n5184), .A2(n7372), .ZN(n5180) );
  NAND2_X1 U5732 ( .A1(n7359), .A2(n7415), .ZN(n5345) );
  INV_X1 U5733 ( .A(n5345), .ZN(n5161) );
  NOR2_X1 U5734 ( .A1(n7418), .A2(n7426), .ZN(n5179) );
  INV_X1 U5735 ( .A(n5496), .ZN(n5139) );
  NAND2_X1 U5736 ( .A1(n5137), .A2(n5258), .ZN(n5177) );
  INV_X1 U5737 ( .A(n5177), .ZN(n5138) );
  NAND2_X1 U5738 ( .A1(n5138), .A2(n5084), .ZN(n7414) );
  OR2_X1 U5739 ( .A1(n7414), .A2(n7371), .ZN(n5144) );
  OAI211_X1 U5740 ( .C1(n5161), .C2(n5179), .A(n5139), .B(n5144), .ZN(n5140)
         );
  AND3_X1 U5741 ( .A1(n5141), .A2(n5180), .A3(n5140), .ZN(n5501) );
  AOI22_X1 U5742 ( .A1(n7574), .A2(n5496), .B1(n7571), .B2(n5495), .ZN(n5146)
         );
  INV_X1 U5743 ( .A(n5336), .ZN(n5579) );
  NAND2_X1 U5744 ( .A1(n5142), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5576) );
  INV_X1 U5745 ( .A(n5143), .ZN(n5224) );
  OAI22_X1 U5746 ( .A1(n5579), .A2(n5184), .B1(n5576), .B2(n5224), .ZN(n5497)
         );
  AOI22_X1 U5747 ( .A1(n5596), .A2(n5497), .B1(n7572), .B2(n7573), .ZN(n5145)
         );
  OAI211_X1 U5748 ( .C1(n5501), .C2(n3749), .A(n5146), .B(n5145), .ZN(U3027)
         );
  INV_X1 U5749 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5149) );
  AOI22_X1 U5750 ( .A1(n7484), .A2(n5496), .B1(n7483), .B2(n5495), .ZN(n5148)
         );
  AOI22_X1 U5751 ( .A1(n5604), .A2(n5497), .B1(n7485), .B2(n7573), .ZN(n5147)
         );
  OAI211_X1 U5752 ( .C1(n5501), .C2(n5149), .A(n5148), .B(n5147), .ZN(U3023)
         );
  AOI22_X1 U5753 ( .A1(n7453), .A2(n5496), .B1(n7451), .B2(n5495), .ZN(n5151)
         );
  AOI22_X1 U5754 ( .A1(n5592), .A2(n5497), .B1(n7452), .B2(n7573), .ZN(n5150)
         );
  OAI211_X1 U5755 ( .C1(n5501), .C2(n5152), .A(n5151), .B(n5150), .ZN(U3021)
         );
  AOI22_X1 U5756 ( .A1(n7422), .A2(n5496), .B1(n7421), .B2(n5495), .ZN(n5154)
         );
  AOI22_X1 U5757 ( .A1(n5600), .A2(n5497), .B1(n7430), .B2(n7573), .ZN(n5153)
         );
  OAI211_X1 U5758 ( .C1(n5501), .C2(n5155), .A(n5154), .B(n5153), .ZN(U3020)
         );
  NAND3_X1 U5759 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(n7361), .ZN(n5203) );
  NOR2_X1 U5760 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5203), .ZN(n5477)
         );
  INV_X1 U5761 ( .A(n5477), .ZN(n5157) );
  OR2_X1 U5762 ( .A1(n5342), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5577)
         );
  INV_X1 U5763 ( .A(n5577), .ZN(n5156) );
  NOR2_X1 U5764 ( .A1(n5156), .A2(n3887), .ZN(n5574) );
  NAND2_X1 U5765 ( .A1(n5413), .A2(n5576), .ZN(n5328) );
  AOI211_X1 U5766 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5157), .A(n5574), .B(
        n5328), .ZN(n5163) );
  NOR2_X1 U5767 ( .A1(n5200), .A2(n7426), .ZN(n5262) );
  NOR2_X2 U5768 ( .A1(n5178), .A2(n7371), .ZN(n5518) );
  INV_X1 U5769 ( .A(n5518), .ZN(n5160) );
  INV_X1 U5770 ( .A(n7565), .ZN(n5159) );
  OAI211_X1 U5771 ( .C1(n5161), .C2(n5262), .A(n5160), .B(n5159), .ZN(n5162)
         );
  OR2_X1 U5772 ( .A1(n5200), .A2(n7400), .ZN(n5264) );
  AND3_X1 U5773 ( .A1(n5163), .A2(n5162), .A3(n5264), .ZN(n5482) );
  INV_X1 U5774 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5166) );
  AOI22_X1 U5775 ( .A1(n7422), .A2(n7565), .B1(n7421), .B2(n5477), .ZN(n5165)
         );
  INV_X1 U5776 ( .A(n5200), .ZN(n5267) );
  OAI22_X1 U5777 ( .A1(n5579), .A2(n5267), .B1(n5577), .B2(n5340), .ZN(n5478)
         );
  AOI22_X1 U5778 ( .A1(n5600), .A2(n5478), .B1(n7430), .B2(n5518), .ZN(n5164)
         );
  OAI211_X1 U5779 ( .C1(n5482), .C2(n5166), .A(n5165), .B(n5164), .ZN(U3068)
         );
  INV_X1 U5780 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5169) );
  AOI22_X1 U5781 ( .A1(n7574), .A2(n7565), .B1(n7571), .B2(n5477), .ZN(n5168)
         );
  AOI22_X1 U5782 ( .A1(n5596), .A2(n5478), .B1(n5518), .B2(n7572), .ZN(n5167)
         );
  OAI211_X1 U5783 ( .C1(n5482), .C2(n5169), .A(n5168), .B(n5167), .ZN(U3075)
         );
  INV_X1 U5784 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5172) );
  AOI22_X1 U5785 ( .A1(n7484), .A2(n7565), .B1(n7483), .B2(n5477), .ZN(n5171)
         );
  AOI22_X1 U5786 ( .A1(n5604), .A2(n5478), .B1(n5518), .B2(n7485), .ZN(n5170)
         );
  OAI211_X1 U5787 ( .C1(n5482), .C2(n5172), .A(n5171), .B(n5170), .ZN(U3071)
         );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5175) );
  AOI22_X1 U5789 ( .A1(n7453), .A2(n7565), .B1(n7451), .B2(n5477), .ZN(n5174)
         );
  AOI22_X1 U5790 ( .A1(n5592), .A2(n5478), .B1(n5518), .B2(n7452), .ZN(n5173)
         );
  OAI211_X1 U5791 ( .C1(n5482), .C2(n5175), .A(n5174), .B(n5173), .ZN(U3069)
         );
  NOR3_X1 U5792 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7361), .ZN(n7391) );
  INV_X1 U5793 ( .A(n7391), .ZN(n7393) );
  NOR2_X1 U5794 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7393), .ZN(n5502)
         );
  INV_X1 U5795 ( .A(n5502), .ZN(n5176) );
  AOI21_X1 U5796 ( .B1(n5342), .B2(n5341), .A(n3887), .ZN(n5329) );
  AOI211_X1 U5797 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5176), .A(n5329), .B(
        n7379), .ZN(n5182) );
  NAND2_X1 U5798 ( .A1(n7387), .A2(n6118), .ZN(n5185) );
  OAI211_X1 U5799 ( .C1(n5336), .C2(n5179), .A(n5185), .B(n5522), .ZN(n5181)
         );
  AND3_X1 U5800 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n5508) );
  AOI22_X1 U5801 ( .A1(n5503), .A2(n7574), .B1(n7571), .B2(n5502), .ZN(n5187)
         );
  INV_X1 U5802 ( .A(n5576), .ZN(n7376) );
  NAND3_X1 U5803 ( .A1(n7376), .A2(n5342), .A3(n5341), .ZN(n5183) );
  OAI21_X1 U5804 ( .B1(n5184), .B2(n5345), .A(n5183), .ZN(n5504) );
  AOI22_X1 U5805 ( .A1(n5596), .A2(n5504), .B1(n7572), .B2(n7558), .ZN(n5186)
         );
  OAI211_X1 U5806 ( .C1(n5508), .C2(n5188), .A(n5187), .B(n5186), .ZN(U3091)
         );
  INV_X1 U5807 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U5808 ( .A1(n5503), .A2(n7422), .B1(n7421), .B2(n5502), .ZN(n5190)
         );
  AOI22_X1 U5809 ( .A1(n5600), .A2(n5504), .B1(n7430), .B2(n7558), .ZN(n5189)
         );
  OAI211_X1 U5810 ( .C1(n5508), .C2(n5191), .A(n5190), .B(n5189), .ZN(U3084)
         );
  INV_X1 U5811 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5194) );
  AOI22_X1 U5812 ( .A1(n5503), .A2(n7453), .B1(n7451), .B2(n5502), .ZN(n5193)
         );
  AOI22_X1 U5813 ( .A1(n5592), .A2(n5504), .B1(n7452), .B2(n7558), .ZN(n5192)
         );
  OAI211_X1 U5814 ( .C1(n5508), .C2(n5194), .A(n5193), .B(n5192), .ZN(U3085)
         );
  INV_X1 U5815 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5197) );
  AOI22_X1 U5816 ( .A1(n5503), .A2(n7484), .B1(n7483), .B2(n5502), .ZN(n5196)
         );
  AOI22_X1 U5817 ( .A1(n5604), .A2(n5504), .B1(n7485), .B2(n7558), .ZN(n5195)
         );
  OAI211_X1 U5818 ( .C1(n5508), .C2(n5197), .A(n5196), .B(n5195), .ZN(U3087)
         );
  NOR2_X1 U5819 ( .A1(n5198), .A2(n7426), .ZN(n5202) );
  INV_X1 U5820 ( .A(n5199), .ZN(n5517) );
  AOI21_X1 U5821 ( .B1(n7419), .B2(n5200), .A(n5517), .ZN(n5205) );
  AOI22_X1 U5822 ( .A1(n5202), .A2(n5205), .B1(n7426), .B2(n5203), .ZN(n5201)
         );
  NAND2_X1 U5823 ( .A1(n7408), .A2(n5201), .ZN(n5516) );
  INV_X1 U5824 ( .A(n5202), .ZN(n5204) );
  OAI22_X1 U5825 ( .A1(n5205), .A2(n5204), .B1(n3887), .B2(n5203), .ZN(n5515)
         );
  AOI22_X1 U5826 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5516), .B1(n5596), 
        .B2(n5515), .ZN(n5207) );
  AOI22_X1 U5827 ( .A1(n5518), .A2(n7574), .B1(n7571), .B2(n5517), .ZN(n5206)
         );
  OAI211_X1 U5828 ( .C1(n5522), .C2(n5208), .A(n5207), .B(n5206), .ZN(U3083)
         );
  AOI22_X1 U5829 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5516), .B1(n5604), 
        .B2(n5515), .ZN(n5210) );
  AOI22_X1 U5830 ( .A1(n5518), .A2(n7484), .B1(n7483), .B2(n5517), .ZN(n5209)
         );
  OAI211_X1 U5831 ( .C1(n5522), .C2(n5211), .A(n5210), .B(n5209), .ZN(U3079)
         );
  AOI22_X1 U5832 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5516), .B1(n5592), 
        .B2(n5515), .ZN(n5213) );
  AOI22_X1 U5833 ( .A1(n5518), .A2(n7453), .B1(n7451), .B2(n5517), .ZN(n5212)
         );
  OAI211_X1 U5834 ( .C1(n5522), .C2(n5214), .A(n5213), .B(n5212), .ZN(U3077)
         );
  AOI22_X1 U5835 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5516), .B1(n5600), 
        .B2(n5515), .ZN(n5216) );
  AOI22_X1 U5836 ( .A1(n5518), .A2(n7422), .B1(n7421), .B2(n5517), .ZN(n5215)
         );
  OAI211_X1 U5837 ( .C1(n5522), .C2(n5217), .A(n5216), .B(n5215), .ZN(U3076)
         );
  NOR3_X1 U5838 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5327), .ZN(n7403) );
  INV_X1 U5839 ( .A(n7403), .ZN(n7404) );
  NOR2_X1 U5840 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7404), .ZN(n5412)
         );
  INV_X1 U5841 ( .A(n5412), .ZN(n5219) );
  AOI211_X1 U5842 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5219), .A(n5218), .B(
        n5328), .ZN(n5223) );
  OR2_X1 U5843 ( .A1(n5066), .A2(n5090), .ZN(n7349) );
  NAND2_X1 U5844 ( .A1(n7349), .A2(n7415), .ZN(n5331) );
  NAND2_X1 U5845 ( .A1(n5345), .A2(n5331), .ZN(n5220) );
  NAND2_X1 U5846 ( .A1(n5428), .A2(n5220), .ZN(n5221) );
  OR2_X1 U5847 ( .A1(n7564), .A2(n5221), .ZN(n5222) );
  NAND2_X1 U5848 ( .A1(n7349), .A2(n7372), .ZN(n5338) );
  AND3_X1 U5849 ( .A1(n5223), .A2(n5222), .A3(n5338), .ZN(n5418) );
  INV_X1 U5850 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U5851 ( .A1(n7451), .A2(n5412), .B1(n5411), .B2(n7453), .ZN(n5226)
         );
  OAI22_X1 U5852 ( .A1(n5579), .A2(n7349), .B1(n5224), .B2(n5340), .ZN(n5414)
         );
  AOI22_X1 U5853 ( .A1(n5592), .A2(n5414), .B1(n7452), .B2(n7564), .ZN(n5225)
         );
  OAI211_X1 U5854 ( .C1(n5418), .C2(n5227), .A(n5226), .B(n5225), .ZN(U3053)
         );
  INV_X1 U5855 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5230) );
  AOI22_X1 U5856 ( .A1(n7483), .A2(n5412), .B1(n5411), .B2(n7484), .ZN(n5229)
         );
  AOI22_X1 U5857 ( .A1(n5604), .A2(n5414), .B1(n7485), .B2(n7564), .ZN(n5228)
         );
  OAI211_X1 U5858 ( .C1(n5418), .C2(n5230), .A(n5229), .B(n5228), .ZN(U3055)
         );
  INV_X1 U5859 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5233) );
  AOI22_X1 U5860 ( .A1(n7571), .A2(n5412), .B1(n5411), .B2(n7574), .ZN(n5232)
         );
  AOI22_X1 U5861 ( .A1(n5596), .A2(n5414), .B1(n7572), .B2(n7564), .ZN(n5231)
         );
  OAI211_X1 U5862 ( .C1(n5418), .C2(n5233), .A(n5232), .B(n5231), .ZN(U3059)
         );
  INV_X1 U5863 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5236) );
  AOI22_X1 U5864 ( .A1(n7421), .A2(n5412), .B1(n5411), .B2(n7422), .ZN(n5235)
         );
  AOI22_X1 U5865 ( .A1(n5600), .A2(n5414), .B1(n7430), .B2(n7564), .ZN(n5234)
         );
  OAI211_X1 U5866 ( .C1(n5418), .C2(n5236), .A(n5235), .B(n5234), .ZN(U3052)
         );
  OAI21_X1 U5867 ( .B1(n5239), .B2(n5238), .A(n5237), .ZN(n6792) );
  NAND2_X1 U5868 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6857) );
  OAI21_X1 U5869 ( .B1(n4560), .B2(n6151), .A(n6878), .ZN(n6867) );
  NAND2_X1 U5870 ( .A1(n6870), .A2(n6867), .ZN(n5389) );
  OR2_X1 U5871 ( .A1(n5240), .A2(n6857), .ZN(n5559) );
  NOR2_X1 U5872 ( .A1(n6878), .A2(n4560), .ZN(n6035) );
  OAI21_X1 U5873 ( .B1(n6589), .B2(n6035), .A(n6587), .ZN(n5560) );
  INV_X1 U5874 ( .A(n5560), .ZN(n6877) );
  OAI21_X1 U5875 ( .B1(n6867), .B2(n6471), .A(n6877), .ZN(n6862) );
  AOI21_X1 U5876 ( .B1(n6467), .B2(n5559), .A(n6862), .ZN(n5391) );
  AOI221_X1 U5877 ( .B1(n6857), .B2(n5240), .C1(n5389), .C2(n5240), .A(n5391), 
        .ZN(n5245) );
  NAND2_X1 U5878 ( .A1(n6866), .A2(n6035), .ZN(n5390) );
  NOR3_X1 U5879 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6857), .A3(n5390), 
        .ZN(n5244) );
  INV_X1 U5880 ( .A(REIP_REG_5__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U5881 ( .A1(n6884), .A2(n6968), .B1(n6924), .B2(n5242), .ZN(n5243)
         );
  NOR3_X1 U5882 ( .A1(n5245), .A2(n5244), .A3(n5243), .ZN(n5246) );
  OAI21_X1 U5883 ( .B1(n6619), .B2(n6792), .A(n5246), .ZN(U3013) );
  AOI21_X1 U5884 ( .B1(n5251), .B2(n5247), .A(n5250), .ZN(n6796) );
  INV_X1 U5885 ( .A(n6796), .ZN(n6986) );
  AOI21_X1 U5886 ( .B1(n5253), .B2(n5252), .A(n5324), .ZN(n5387) );
  AOI22_X1 U5887 ( .A1(n6769), .A2(n5387), .B1(EBX_REG_6__SCAN_IN), .B2(n6311), 
        .ZN(n5254) );
  OAI21_X1 U5888 ( .B1(n6986), .B2(n6315), .A(n5254), .ZN(U2853) );
  INV_X1 U5889 ( .A(EAX_REG_18__SCAN_IN), .ZN(n7263) );
  AOI22_X1 U5890 ( .A1(n6668), .A2(UWORD_REG_2__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5255) );
  OAI21_X1 U5891 ( .B1(n7263), .B2(n5284), .A(n5255), .ZN(U2905) );
  NOR2_X1 U5892 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5256), .ZN(n5532)
         );
  INV_X1 U5893 ( .A(n5532), .ZN(n5257) );
  OR2_X1 U5894 ( .A1(n5342), .A2(n7361), .ZN(n5266) );
  INV_X1 U5895 ( .A(n5266), .ZN(n7375) );
  NOR2_X1 U5896 ( .A1(n7375), .A2(n3887), .ZN(n7380) );
  AOI211_X1 U5897 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5257), .A(n7380), .B(
        n5328), .ZN(n5265) );
  INV_X1 U5898 ( .A(n7539), .ZN(n5261) );
  INV_X1 U5899 ( .A(n5533), .ZN(n5260) );
  OAI211_X1 U5900 ( .C1(n5336), .C2(n5262), .A(n5261), .B(n5260), .ZN(n5263)
         );
  AND3_X1 U5901 ( .A1(n5265), .A2(n5264), .A3(n5263), .ZN(n5538) );
  INV_X1 U5902 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U5903 ( .A1(n7453), .A2(n7539), .B1(n7451), .B2(n5532), .ZN(n5269)
         );
  OAI22_X1 U5904 ( .A1(n5267), .A2(n5345), .B1(n5340), .B2(n5266), .ZN(n5534)
         );
  AOI22_X1 U5905 ( .A1(n5592), .A2(n5534), .B1(n7452), .B2(n5533), .ZN(n5268)
         );
  OAI211_X1 U5906 ( .C1(n5538), .C2(n5270), .A(n5269), .B(n5268), .ZN(U3133)
         );
  INV_X1 U5907 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5273) );
  AOI22_X1 U5908 ( .A1(n7484), .A2(n7539), .B1(n7483), .B2(n5532), .ZN(n5272)
         );
  AOI22_X1 U5909 ( .A1(n5604), .A2(n5534), .B1(n7485), .B2(n5533), .ZN(n5271)
         );
  OAI211_X1 U5910 ( .C1(n5538), .C2(n5273), .A(n5272), .B(n5271), .ZN(U3135)
         );
  INV_X1 U5911 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5276) );
  AOI22_X1 U5912 ( .A1(n7574), .A2(n7539), .B1(n7571), .B2(n5532), .ZN(n5275)
         );
  AOI22_X1 U5913 ( .A1(n5596), .A2(n5534), .B1(n7572), .B2(n5533), .ZN(n5274)
         );
  OAI211_X1 U5914 ( .C1(n5538), .C2(n5276), .A(n5275), .B(n5274), .ZN(U3139)
         );
  INV_X1 U5915 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U5916 ( .A1(n7422), .A2(n7539), .B1(n7421), .B2(n5532), .ZN(n5278)
         );
  AOI22_X1 U5917 ( .A1(n5600), .A2(n5534), .B1(n7430), .B2(n5533), .ZN(n5277)
         );
  OAI211_X1 U5918 ( .C1(n5538), .C2(n5279), .A(n5278), .B(n5277), .ZN(U3132)
         );
  AOI22_X1 U5919 ( .A1(n6668), .A2(UWORD_REG_1__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U5920 ( .B1(n4403), .B2(n5284), .A(n5280), .ZN(U2906) );
  INV_X1 U5921 ( .A(EAX_REG_16__SCAN_IN), .ZN(n7253) );
  AOI22_X1 U5922 ( .A1(n6668), .A2(UWORD_REG_0__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5281) );
  OAI21_X1 U5923 ( .B1(n7253), .B2(n5284), .A(n5281), .ZN(U2907) );
  AOI22_X1 U5924 ( .A1(n6668), .A2(UWORD_REG_14__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5282) );
  OAI21_X1 U5925 ( .B1(n4740), .B2(n5284), .A(n5282), .ZN(U2893) );
  AOI22_X1 U5926 ( .A1(n6668), .A2(UWORD_REG_3__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5283) );
  OAI21_X1 U5927 ( .B1(n4438), .B2(n5284), .A(n5283), .ZN(U2904) );
  INV_X1 U5928 ( .A(n5287), .ZN(n5288) );
  NOR2_X1 U5929 ( .A1(n5289), .A2(n5288), .ZN(n7205) );
  NOR3_X1 U5930 ( .A1(n7224), .A2(n7214), .A3(n7216), .ZN(n7219) );
  OR2_X1 U5931 ( .A1(n7205), .A2(n7219), .ZN(n5290) );
  NAND2_X1 U5932 ( .A1(n6941), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5293) );
  INV_X1 U5933 ( .A(n5304), .ZN(n6181) );
  NAND2_X1 U5934 ( .A1(n6181), .A2(n3956), .ZN(n5292) );
  NAND2_X1 U5935 ( .A1(n7130), .A2(n5292), .ZN(n6974) );
  INV_X1 U5936 ( .A(n6974), .ZN(n6932) );
  INV_X1 U5937 ( .A(n5293), .ZN(n5294) );
  NOR2_X1 U5938 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n5300) );
  NAND2_X1 U5939 ( .A1(n6006), .A2(n5300), .ZN(n7203) );
  NOR2_X1 U5940 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5300), .ZN(n5296) );
  AOI22_X1 U5941 ( .A1(n4570), .A2(n7203), .B1(n5296), .B2(n3929), .ZN(n5297)
         );
  NOR2_X2 U5942 ( .A1(n5304), .A2(n5297), .ZN(n7145) );
  NAND3_X1 U5943 ( .A1(n5298), .A2(n3929), .A3(n5300), .ZN(n5299) );
  INV_X1 U5944 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5305) );
  INV_X1 U5945 ( .A(n5300), .ZN(n5301) );
  NAND3_X1 U5946 ( .A1(n5302), .A2(EBX_REG_31__SCAN_IN), .A3(n5301), .ZN(n5303) );
  AOI22_X1 U5947 ( .A1(n7139), .A2(n5305), .B1(n7125), .B2(n4982), .ZN(n5310)
         );
  INV_X1 U5948 ( .A(n6005), .ZN(n5306) );
  NAND2_X1 U5949 ( .A1(n6181), .A2(n5306), .ZN(n6961) );
  INV_X1 U5950 ( .A(n6941), .ZN(n7075) );
  AOI22_X1 U5951 ( .A1(n7144), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7075), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5307) );
  OAI21_X1 U5952 ( .B1(n6961), .B2(n6150), .A(n5307), .ZN(n5308) );
  INV_X1 U5953 ( .A(n5308), .ZN(n5309) );
  OAI211_X1 U5954 ( .C1(n5311), .C2(n7120), .A(n5310), .B(n5309), .ZN(n5312)
         );
  AOI21_X1 U5955 ( .B1(n7133), .B2(n5313), .A(n5312), .ZN(n5314) );
  OAI21_X1 U5956 ( .B1(n6932), .B2(n5373), .A(n5314), .ZN(U2826) );
  OAI21_X1 U5957 ( .B1(n5315), .B2(n5317), .A(n5316), .ZN(n7008) );
  OAI21_X1 U5958 ( .B1(n5318), .B2(n5319), .A(n6748), .ZN(n7005) );
  INV_X1 U5959 ( .A(n7005), .ZN(n5320) );
  AOI22_X1 U5960 ( .A1(n6769), .A2(n5320), .B1(EBX_REG_8__SCAN_IN), .B2(n6311), 
        .ZN(n5321) );
  OAI21_X1 U5961 ( .B1(n7008), .B2(n6315), .A(n5321), .ZN(U2851) );
  OAI21_X1 U5962 ( .B1(n5250), .B2(n5322), .A(n3684), .ZN(n6995) );
  INV_X1 U5963 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5326) );
  INV_X1 U5964 ( .A(n5318), .ZN(n5323) );
  OAI21_X1 U5965 ( .B1(n5325), .B2(n5324), .A(n5323), .ZN(n6991) );
  OAI222_X1 U5966 ( .A1(n6995), .A2(n6315), .B1(n5326), .B2(n6773), .C1(n6991), 
        .C2(n6320), .ZN(U2852) );
  NOR3_X1 U5967 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5327), .A3(n7361), 
        .ZN(n7355) );
  INV_X1 U5968 ( .A(n7355), .ZN(n7350) );
  NOR2_X1 U5969 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7350), .ZN(n5483)
         );
  INV_X1 U5970 ( .A(n5483), .ZN(n5330) );
  AOI211_X1 U5971 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5330), .A(n5329), .B(
        n5328), .ZN(n5339) );
  INV_X1 U5972 ( .A(n5331), .ZN(n5335) );
  INV_X1 U5973 ( .A(n7538), .ZN(n5334) );
  NAND2_X1 U5974 ( .A1(n5333), .A2(n5332), .ZN(n7368) );
  OR2_X1 U5975 ( .A1(n7368), .A2(n6118), .ZN(n5346) );
  OAI211_X1 U5976 ( .C1(n5336), .C2(n5335), .A(n5334), .B(n5346), .ZN(n5337)
         );
  AND3_X1 U5977 ( .A1(n5339), .A2(n5338), .A3(n5337), .ZN(n5488) );
  INV_X1 U5978 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5349) );
  AOI22_X1 U5979 ( .A1(n7430), .A2(n7538), .B1(n7421), .B2(n5483), .ZN(n5348)
         );
  INV_X1 U5980 ( .A(n5340), .ZN(n5343) );
  NAND3_X1 U5981 ( .A1(n5343), .A2(n5342), .A3(n5341), .ZN(n5344) );
  OAI21_X1 U5982 ( .B1(n5345), .B2(n7349), .A(n5344), .ZN(n5484) );
  AOI22_X1 U5983 ( .A1(n5600), .A2(n5484), .B1(n7422), .B2(n7545), .ZN(n5347)
         );
  OAI211_X1 U5984 ( .C1(n5488), .C2(n5349), .A(n5348), .B(n5347), .ZN(U3116)
         );
  INV_X1 U5985 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5352) );
  AOI22_X1 U5986 ( .A1(n7485), .A2(n7538), .B1(n7483), .B2(n5483), .ZN(n5351)
         );
  AOI22_X1 U5987 ( .A1(n5604), .A2(n5484), .B1(n7484), .B2(n7545), .ZN(n5350)
         );
  OAI211_X1 U5988 ( .C1(n5488), .C2(n5352), .A(n5351), .B(n5350), .ZN(U3119)
         );
  INV_X1 U5989 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5355) );
  AOI22_X1 U5990 ( .A1(n7572), .A2(n7538), .B1(n7571), .B2(n5483), .ZN(n5354)
         );
  AOI22_X1 U5991 ( .A1(n5596), .A2(n5484), .B1(n7574), .B2(n7545), .ZN(n5353)
         );
  OAI211_X1 U5992 ( .C1(n5488), .C2(n5355), .A(n5354), .B(n5353), .ZN(U3123)
         );
  INV_X1 U5993 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U5994 ( .A1(n7452), .A2(n7538), .B1(n7451), .B2(n5483), .ZN(n5357)
         );
  AOI22_X1 U5995 ( .A1(n5592), .A2(n5484), .B1(n7453), .B2(n7545), .ZN(n5356)
         );
  OAI211_X1 U5996 ( .C1(n5488), .C2(n5358), .A(n5357), .B(n5356), .ZN(U3117)
         );
  NOR2_X1 U5997 ( .A1(n4979), .A2(n5359), .ZN(n5360) );
  AND2_X1 U5998 ( .A1(n3970), .A2(n7250), .ZN(n5362) );
  AND2_X1 U5999 ( .A1(n3687), .A2(n5364), .ZN(n5366) );
  NOR2_X1 U6000 ( .A1(n5366), .A2(n3966), .ZN(n5365) );
  NAND2_X2 U6001 ( .A1(n6142), .A2(n5365), .ZN(n7335) );
  AND2_X1 U6002 ( .A1(n6142), .A2(n3966), .ZN(n7434) );
  INV_X1 U6003 ( .A(DATAI_2_), .ZN(n5367) );
  INV_X1 U6004 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7266) );
  OAI222_X1 U6005 ( .A1(n6931), .A2(n7335), .B1(n6343), .B2(n5367), .C1(n6142), 
        .C2(n7266), .ZN(U2889) );
  OAI222_X1 U6006 ( .A1(n6986), .A2(n7335), .B1(n6343), .B2(n7282), .C1(n6142), 
        .C2(n4230), .ZN(U2885) );
  INV_X1 U6007 ( .A(DATAI_7_), .ZN(n5849) );
  INV_X1 U6008 ( .A(EAX_REG_7__SCAN_IN), .ZN(n7290) );
  OAI222_X1 U6009 ( .A1(n6995), .A2(n7335), .B1(n6343), .B2(n5849), .C1(n6142), 
        .C2(n7290), .ZN(U2884) );
  INV_X1 U6010 ( .A(DATAI_8_), .ZN(n5851) );
  INV_X1 U6011 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7295) );
  OAI222_X1 U6012 ( .A1(n7008), .A2(n7335), .B1(n6343), .B2(n5851), .C1(n6142), 
        .C2(n7295), .ZN(U2883) );
  INV_X1 U6013 ( .A(DATAI_0_), .ZN(n7251) );
  INV_X1 U6014 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7256) );
  OAI222_X1 U6015 ( .A1(n5381), .A2(n7335), .B1(n7251), .B2(n6343), .C1(n6142), 
        .C2(n7256), .ZN(U2891) );
  INV_X1 U6016 ( .A(DATAI_3_), .ZN(n7267) );
  INV_X1 U6017 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7271) );
  OAI222_X1 U6018 ( .A1(n5368), .A2(n7335), .B1(n7267), .B2(n6343), .C1(n6142), 
        .C2(n7271), .ZN(U2888) );
  OR2_X1 U6019 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  AND2_X1 U6020 ( .A1(n5001), .A2(n5371), .ZN(n6964) );
  INV_X1 U6021 ( .A(n6964), .ZN(n5372) );
  INV_X1 U6022 ( .A(DATAI_4_), .ZN(n7272) );
  INV_X1 U6023 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7277) );
  OAI222_X1 U6024 ( .A1(n5372), .A2(n7335), .B1(n7272), .B2(n6343), .C1(n6142), 
        .C2(n7277), .ZN(U2887) );
  INV_X1 U6025 ( .A(DATAI_1_), .ZN(n7257) );
  INV_X1 U6026 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7261) );
  OAI222_X1 U6027 ( .A1(n5373), .A2(n7335), .B1(n7257), .B2(n6343), .C1(n6142), 
        .C2(n7261), .ZN(U2890) );
  NAND2_X1 U6028 ( .A1(n7157), .A2(n7122), .ZN(n5379) );
  INV_X1 U6029 ( .A(n6961), .ZN(n5374) );
  AOI22_X1 U6030 ( .A1(n5374), .A2(n7363), .B1(n7125), .B2(n6916), .ZN(n5376)
         );
  NAND2_X1 U6031 ( .A1(n7074), .A2(REIP_REG_0__SCAN_IN), .ZN(n5375) );
  OAI211_X1 U6032 ( .C1(n5377), .C2(n7120), .A(n5376), .B(n5375), .ZN(n5378)
         );
  AOI21_X1 U6033 ( .B1(n5379), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5378), 
        .ZN(n5380) );
  OAI21_X1 U6034 ( .B1(n6932), .B2(n5381), .A(n5380), .ZN(U2827) );
  INV_X1 U6035 ( .A(DATAI_5_), .ZN(n5382) );
  OAI222_X1 U6036 ( .A1(n7335), .A2(n6971), .B1(n6142), .B2(n4202), .C1(n5382), 
        .C2(n6343), .ZN(U2886) );
  NAND2_X1 U6037 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  XNOR2_X1 U6038 ( .A(n5383), .B(n5386), .ZN(n6797) );
  INV_X1 U6039 ( .A(n5387), .ZN(n6979) );
  INV_X1 U6040 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5388) );
  OAI22_X1 U6041 ( .A1(n6884), .A2(n6979), .B1(n6924), .B2(n5388), .ZN(n5395)
         );
  NAND2_X1 U6042 ( .A1(n5390), .A2(n5389), .ZN(n6880) );
  INV_X1 U6043 ( .A(n6880), .ZN(n6865) );
  NOR2_X1 U6044 ( .A1(n6865), .A2(n5559), .ZN(n5393) );
  INV_X1 U6045 ( .A(n5391), .ZN(n5392) );
  MUX2_X1 U6046 ( .A(n5393), .B(n5392), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n5394) );
  AOI211_X1 U6047 ( .C1(n6915), .C2(n6797), .A(n5395), .B(n5394), .ZN(n5396)
         );
  INV_X1 U6048 ( .A(n5396), .ZN(U3012) );
  XNOR2_X1 U6049 ( .A(n5316), .B(n5397), .ZN(n6745) );
  INV_X1 U6050 ( .A(DATAI_9_), .ZN(n7296) );
  INV_X1 U6051 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7301) );
  OAI222_X1 U6052 ( .A1(n7335), .A2(n6745), .B1(n7296), .B2(n6343), .C1(n6142), 
        .C2(n7301), .ZN(U2882) );
  INV_X1 U6053 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5400) );
  NOR2_X2 U6054 ( .A1(n5410), .A2(n4068), .ZN(n7531) );
  AOI22_X1 U6055 ( .A1(n7531), .A2(n5412), .B1(n5411), .B2(n7532), .ZN(n5399)
         );
  NAND2_X1 U6056 ( .A1(DATAI_6_), .A2(n5413), .ZN(n7536) );
  NAND2_X1 U6057 ( .A1(n6818), .A2(DATAI_22_), .ZN(n5446) );
  INV_X1 U6058 ( .A(n5446), .ZN(n7533) );
  AOI22_X1 U6059 ( .A1(n5588), .A2(n5414), .B1(n7533), .B2(n7564), .ZN(n5398)
         );
  OAI211_X1 U6060 ( .C1(n5418), .C2(n5400), .A(n5399), .B(n5398), .ZN(U3058)
         );
  AOI22_X1 U6061 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5424), .B1(n5588), 
        .B2(n5423), .ZN(n5402) );
  AOI22_X1 U6062 ( .A1(n7531), .A2(n5425), .B1(n7532), .B2(n5608), .ZN(n5401)
         );
  OAI211_X1 U6063 ( .C1(n5446), .C2(n5428), .A(n5402), .B(n5401), .ZN(U3050)
         );
  INV_X1 U6064 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5406) );
  NOR2_X2 U6065 ( .A1(n5410), .A2(n5403), .ZN(n7467) );
  AOI22_X1 U6066 ( .A1(n7467), .A2(n5412), .B1(n5411), .B2(n7468), .ZN(n5405)
         );
  NAND2_X1 U6067 ( .A1(DATAI_2_), .A2(n5413), .ZN(n7472) );
  NAND2_X1 U6068 ( .A1(n6818), .A2(DATAI_18_), .ZN(n5521) );
  INV_X1 U6069 ( .A(n5521), .ZN(n7469) );
  AOI22_X1 U6070 ( .A1(n5584), .A2(n5414), .B1(n7469), .B2(n7564), .ZN(n5404)
         );
  OAI211_X1 U6071 ( .C1(n5418), .C2(n5406), .A(n5405), .B(n5404), .ZN(U3054)
         );
  INV_X1 U6072 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5409) );
  NOR2_X2 U6073 ( .A1(n5410), .A2(n3687), .ZN(n7515) );
  AOI22_X1 U6074 ( .A1(n7515), .A2(n5412), .B1(n5411), .B2(n7517), .ZN(n5408)
         );
  NAND2_X1 U6075 ( .A1(DATAI_5_), .A2(n5413), .ZN(n7520) );
  NAND2_X1 U6076 ( .A1(n6818), .A2(DATAI_21_), .ZN(n5514) );
  INV_X1 U6077 ( .A(n5514), .ZN(n7516) );
  AOI22_X1 U6078 ( .A1(n5611), .A2(n5414), .B1(n7516), .B2(n7564), .ZN(n5407)
         );
  OAI211_X1 U6079 ( .C1(n5418), .C2(n5409), .A(n5408), .B(n5407), .ZN(U3057)
         );
  INV_X1 U6080 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5417) );
  NOR2_X2 U6081 ( .A1(n5410), .A2(n3963), .ZN(n7499) );
  AOI22_X1 U6082 ( .A1(n7499), .A2(n5412), .B1(n5411), .B2(n7500), .ZN(n5416)
         );
  NAND2_X1 U6083 ( .A1(DATAI_4_), .A2(n5413), .ZN(n7504) );
  NAND2_X1 U6084 ( .A1(n6818), .A2(DATAI_20_), .ZN(n5511) );
  AOI22_X1 U6085 ( .A1(n5580), .A2(n5414), .B1(n7501), .B2(n7564), .ZN(n5415)
         );
  OAI211_X1 U6086 ( .C1(n5418), .C2(n5417), .A(n5416), .B(n5415), .ZN(U3056)
         );
  AOI22_X1 U6087 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5424), .B1(n5584), 
        .B2(n5423), .ZN(n5420) );
  AOI22_X1 U6088 ( .A1(n7467), .A2(n5425), .B1(n7468), .B2(n5608), .ZN(n5419)
         );
  OAI211_X1 U6089 ( .C1(n5521), .C2(n5428), .A(n5420), .B(n5419), .ZN(U3046)
         );
  AOI22_X1 U6090 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5424), .B1(n5611), 
        .B2(n5423), .ZN(n5422) );
  AOI22_X1 U6091 ( .A1(n7515), .A2(n5425), .B1(n7517), .B2(n5608), .ZN(n5421)
         );
  OAI211_X1 U6092 ( .C1(n5514), .C2(n5428), .A(n5422), .B(n5421), .ZN(U3049)
         );
  AOI22_X1 U6093 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5424), .B1(n5580), 
        .B2(n5423), .ZN(n5427) );
  AOI22_X1 U6094 ( .A1(n7499), .A2(n5425), .B1(n7500), .B2(n5608), .ZN(n5426)
         );
  OAI211_X1 U6095 ( .C1(n5511), .C2(n5428), .A(n5427), .B(n5426), .ZN(U3048)
         );
  AOI22_X1 U6096 ( .A1(n7532), .A2(n5496), .B1(n7531), .B2(n5495), .ZN(n5430)
         );
  AOI22_X1 U6097 ( .A1(n5588), .A2(n5497), .B1(n7533), .B2(n7573), .ZN(n5429)
         );
  OAI211_X1 U6098 ( .C1(n5501), .C2(n5431), .A(n5430), .B(n5429), .ZN(U3026)
         );
  AOI22_X1 U6099 ( .A1(n7533), .A2(n7538), .B1(n7531), .B2(n5483), .ZN(n5433)
         );
  AOI22_X1 U6100 ( .A1(n5588), .A2(n5484), .B1(n7532), .B2(n7545), .ZN(n5432)
         );
  OAI211_X1 U6101 ( .C1(n5488), .C2(n5434), .A(n5433), .B(n5432), .ZN(U3122)
         );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5437) );
  AOI22_X1 U6103 ( .A1(n7532), .A2(n7565), .B1(n7531), .B2(n5477), .ZN(n5436)
         );
  AOI22_X1 U6104 ( .A1(n5588), .A2(n5478), .B1(n5518), .B2(n7533), .ZN(n5435)
         );
  OAI211_X1 U6105 ( .C1(n5482), .C2(n5437), .A(n5436), .B(n5435), .ZN(U3074)
         );
  INV_X1 U6106 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5440) );
  AOI22_X1 U6107 ( .A1(n7533), .A2(n5496), .B1(n7531), .B2(n5489), .ZN(n5439)
         );
  AOI22_X1 U6108 ( .A1(n5588), .A2(n5490), .B1(n7532), .B2(n5533), .ZN(n5438)
         );
  OAI211_X1 U6109 ( .C1(n5494), .C2(n5440), .A(n5439), .B(n5438), .ZN(U3146)
         );
  INV_X1 U6110 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5443) );
  AOI22_X1 U6111 ( .A1(n5503), .A2(n7532), .B1(n7531), .B2(n5502), .ZN(n5442)
         );
  AOI22_X1 U6112 ( .A1(n5588), .A2(n5504), .B1(n7533), .B2(n7558), .ZN(n5441)
         );
  OAI211_X1 U6113 ( .C1(n5508), .C2(n5443), .A(n5442), .B(n5441), .ZN(U3090)
         );
  AOI22_X1 U6114 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5516), .B1(n5588), 
        .B2(n5515), .ZN(n5445) );
  AOI22_X1 U6115 ( .A1(n5518), .A2(n7532), .B1(n7531), .B2(n5517), .ZN(n5444)
         );
  OAI211_X1 U6116 ( .C1(n5522), .C2(n5446), .A(n5445), .B(n5444), .ZN(U3082)
         );
  AOI22_X1 U6117 ( .A1(n7500), .A2(n5496), .B1(n7499), .B2(n5495), .ZN(n5448)
         );
  AOI22_X1 U6118 ( .A1(n5580), .A2(n5497), .B1(n7501), .B2(n7573), .ZN(n5447)
         );
  OAI211_X1 U6119 ( .C1(n5501), .C2(n5449), .A(n5448), .B(n5447), .ZN(U3024)
         );
  INV_X1 U6120 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5452) );
  AOI22_X1 U6121 ( .A1(n7501), .A2(n7538), .B1(n7499), .B2(n5483), .ZN(n5451)
         );
  AOI22_X1 U6122 ( .A1(n5580), .A2(n5484), .B1(n7500), .B2(n7545), .ZN(n5450)
         );
  OAI211_X1 U6123 ( .C1(n5488), .C2(n5452), .A(n5451), .B(n5450), .ZN(U3120)
         );
  AOI22_X1 U6124 ( .A1(n7517), .A2(n5496), .B1(n7515), .B2(n5495), .ZN(n5454)
         );
  AOI22_X1 U6125 ( .A1(n5611), .A2(n5497), .B1(n7516), .B2(n7573), .ZN(n5453)
         );
  OAI211_X1 U6126 ( .C1(n5501), .C2(n5455), .A(n5454), .B(n5453), .ZN(U3025)
         );
  INV_X1 U6127 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5458) );
  AOI22_X1 U6128 ( .A1(n7517), .A2(n7565), .B1(n7515), .B2(n5477), .ZN(n5457)
         );
  AOI22_X1 U6129 ( .A1(n5611), .A2(n5478), .B1(n5518), .B2(n7516), .ZN(n5456)
         );
  OAI211_X1 U6130 ( .C1(n5482), .C2(n5458), .A(n5457), .B(n5456), .ZN(U3073)
         );
  INV_X1 U6131 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5461) );
  AOI22_X1 U6132 ( .A1(n7516), .A2(n5496), .B1(n7515), .B2(n5489), .ZN(n5460)
         );
  AOI22_X1 U6133 ( .A1(n5611), .A2(n5490), .B1(n7517), .B2(n5533), .ZN(n5459)
         );
  OAI211_X1 U6134 ( .C1(n5494), .C2(n5461), .A(n5460), .B(n5459), .ZN(U3145)
         );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5464) );
  AOI22_X1 U6136 ( .A1(n7516), .A2(n7538), .B1(n7515), .B2(n5483), .ZN(n5463)
         );
  AOI22_X1 U6137 ( .A1(n5611), .A2(n5484), .B1(n7517), .B2(n7545), .ZN(n5462)
         );
  OAI211_X1 U6138 ( .C1(n5488), .C2(n5464), .A(n5463), .B(n5462), .ZN(U3121)
         );
  INV_X1 U6139 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5467) );
  AOI22_X1 U6140 ( .A1(n7501), .A2(n5496), .B1(n7499), .B2(n5489), .ZN(n5466)
         );
  AOI22_X1 U6141 ( .A1(n5580), .A2(n5490), .B1(n7500), .B2(n5533), .ZN(n5465)
         );
  OAI211_X1 U6142 ( .C1(n5494), .C2(n5467), .A(n5466), .B(n5465), .ZN(U3144)
         );
  INV_X1 U6143 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5470) );
  AOI22_X1 U6144 ( .A1(n5503), .A2(n7517), .B1(n7515), .B2(n5502), .ZN(n5469)
         );
  AOI22_X1 U6145 ( .A1(n5611), .A2(n5504), .B1(n7516), .B2(n7558), .ZN(n5468)
         );
  OAI211_X1 U6146 ( .C1(n5508), .C2(n5470), .A(n5469), .B(n5468), .ZN(U3089)
         );
  INV_X1 U6147 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5473) );
  AOI22_X1 U6148 ( .A1(n7500), .A2(n7565), .B1(n7499), .B2(n5477), .ZN(n5472)
         );
  AOI22_X1 U6149 ( .A1(n5580), .A2(n5478), .B1(n5518), .B2(n7501), .ZN(n5471)
         );
  OAI211_X1 U6150 ( .C1(n5482), .C2(n5473), .A(n5472), .B(n5471), .ZN(U3072)
         );
  INV_X1 U6151 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5476) );
  AOI22_X1 U6152 ( .A1(n5503), .A2(n7500), .B1(n7499), .B2(n5502), .ZN(n5475)
         );
  AOI22_X1 U6153 ( .A1(n5580), .A2(n5504), .B1(n7501), .B2(n7558), .ZN(n5474)
         );
  OAI211_X1 U6154 ( .C1(n5508), .C2(n5476), .A(n5475), .B(n5474), .ZN(U3088)
         );
  INV_X1 U6155 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5481) );
  AOI22_X1 U6156 ( .A1(n7468), .A2(n7565), .B1(n7467), .B2(n5477), .ZN(n5480)
         );
  AOI22_X1 U6157 ( .A1(n5584), .A2(n5478), .B1(n5518), .B2(n7469), .ZN(n5479)
         );
  OAI211_X1 U6158 ( .C1(n5482), .C2(n5481), .A(n5480), .B(n5479), .ZN(U3070)
         );
  INV_X1 U6159 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5487) );
  AOI22_X1 U6160 ( .A1(n7469), .A2(n7538), .B1(n7467), .B2(n5483), .ZN(n5486)
         );
  AOI22_X1 U6161 ( .A1(n5584), .A2(n5484), .B1(n7468), .B2(n7545), .ZN(n5485)
         );
  OAI211_X1 U6162 ( .C1(n5488), .C2(n5487), .A(n5486), .B(n5485), .ZN(U3118)
         );
  INV_X1 U6163 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5493) );
  AOI22_X1 U6164 ( .A1(n7469), .A2(n5496), .B1(n7467), .B2(n5489), .ZN(n5492)
         );
  AOI22_X1 U6165 ( .A1(n5584), .A2(n5490), .B1(n7468), .B2(n5533), .ZN(n5491)
         );
  OAI211_X1 U6166 ( .C1(n5494), .C2(n5493), .A(n5492), .B(n5491), .ZN(U3142)
         );
  INV_X1 U6167 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5500) );
  AOI22_X1 U6168 ( .A1(n7468), .A2(n5496), .B1(n7467), .B2(n5495), .ZN(n5499)
         );
  AOI22_X1 U6169 ( .A1(n5584), .A2(n5497), .B1(n7469), .B2(n7573), .ZN(n5498)
         );
  OAI211_X1 U6170 ( .C1(n5501), .C2(n5500), .A(n5499), .B(n5498), .ZN(U3022)
         );
  INV_X1 U6171 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5507) );
  AOI22_X1 U6172 ( .A1(n5503), .A2(n7468), .B1(n7467), .B2(n5502), .ZN(n5506)
         );
  AOI22_X1 U6173 ( .A1(n5584), .A2(n5504), .B1(n7469), .B2(n7558), .ZN(n5505)
         );
  OAI211_X1 U6174 ( .C1(n5508), .C2(n5507), .A(n5506), .B(n5505), .ZN(U3086)
         );
  AOI22_X1 U6175 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5516), .B1(n5580), 
        .B2(n5515), .ZN(n5510) );
  AOI22_X1 U6176 ( .A1(n5518), .A2(n7500), .B1(n7499), .B2(n5517), .ZN(n5509)
         );
  OAI211_X1 U6177 ( .C1(n5522), .C2(n5511), .A(n5510), .B(n5509), .ZN(U3080)
         );
  AOI22_X1 U6178 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5516), .B1(n5611), 
        .B2(n5515), .ZN(n5513) );
  AOI22_X1 U6179 ( .A1(n5518), .A2(n7517), .B1(n7515), .B2(n5517), .ZN(n5512)
         );
  OAI211_X1 U6180 ( .C1(n5522), .C2(n5514), .A(n5513), .B(n5512), .ZN(U3081)
         );
  AOI22_X1 U6181 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5516), .B1(n5584), 
        .B2(n5515), .ZN(n5520) );
  AOI22_X1 U6182 ( .A1(n5518), .A2(n7468), .B1(n7467), .B2(n5517), .ZN(n5519)
         );
  OAI211_X1 U6183 ( .C1(n5522), .C2(n5521), .A(n5520), .B(n5519), .ZN(U3078)
         );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5525) );
  AOI22_X1 U6185 ( .A1(n7532), .A2(n7539), .B1(n7531), .B2(n5532), .ZN(n5524)
         );
  AOI22_X1 U6186 ( .A1(n5588), .A2(n5534), .B1(n7533), .B2(n5533), .ZN(n5523)
         );
  OAI211_X1 U6187 ( .C1(n5538), .C2(n5525), .A(n5524), .B(n5523), .ZN(U3138)
         );
  INV_X1 U6188 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5528) );
  AOI22_X1 U6189 ( .A1(n7517), .A2(n7539), .B1(n7515), .B2(n5532), .ZN(n5527)
         );
  AOI22_X1 U6190 ( .A1(n5611), .A2(n5534), .B1(n7516), .B2(n5533), .ZN(n5526)
         );
  OAI211_X1 U6191 ( .C1(n5538), .C2(n5528), .A(n5527), .B(n5526), .ZN(U3137)
         );
  INV_X1 U6192 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5531) );
  AOI22_X1 U6193 ( .A1(n7500), .A2(n7539), .B1(n7499), .B2(n5532), .ZN(n5530)
         );
  AOI22_X1 U6194 ( .A1(n5580), .A2(n5534), .B1(n7501), .B2(n5533), .ZN(n5529)
         );
  OAI211_X1 U6195 ( .C1(n5538), .C2(n5531), .A(n5530), .B(n5529), .ZN(U3136)
         );
  INV_X1 U6196 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5537) );
  AOI22_X1 U6197 ( .A1(n7468), .A2(n7539), .B1(n7467), .B2(n5532), .ZN(n5536)
         );
  AOI22_X1 U6198 ( .A1(n5584), .A2(n5534), .B1(n7469), .B2(n5533), .ZN(n5535)
         );
  OAI211_X1 U6199 ( .C1(n5538), .C2(n5537), .A(n5536), .B(n5535), .ZN(U3134)
         );
  AND2_X1 U6200 ( .A1(n5540), .A2(n5539), .ZN(n5542) );
  OR2_X1 U6201 ( .A1(n5542), .A2(n5541), .ZN(n6017) );
  AND2_X1 U6202 ( .A1(n6746), .A2(n5543), .ZN(n5544) );
  OR2_X1 U6203 ( .A1(n5544), .A2(n5631), .ZN(n6039) );
  INV_X1 U6204 ( .A(n6039), .ZN(n5545) );
  AOI22_X1 U6205 ( .A1(n6769), .A2(n5545), .B1(EBX_REG_10__SCAN_IN), .B2(n6311), .ZN(n5546) );
  OAI21_X1 U6206 ( .B1(n6017), .B2(n6315), .A(n5546), .ZN(U2849) );
  INV_X1 U6207 ( .A(n7139), .ZN(n7147) );
  NAND3_X1 U6208 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U6209 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n6983) );
  NAND2_X1 U6210 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n6998) );
  NOR3_X1 U6211 ( .A1(n6953), .A2(n6983), .A3(n6998), .ZN(n7004) );
  NAND2_X1 U6212 ( .A1(n7004), .A2(REIP_REG_8__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U6213 ( .A1(n7139), .A2(n7014), .ZN(n5547) );
  AND2_X1 U6214 ( .A1(n5547), .A2(n6941), .ZN(n7017) );
  OAI21_X1 U6215 ( .B1(REIP_REG_9__SCAN_IN), .B2(n7147), .A(n7017), .ZN(n5554)
         );
  OAI22_X1 U6216 ( .A1(n7120), .A2(n5548), .B1(n7152), .B2(n6039), .ZN(n5553)
         );
  INV_X1 U6217 ( .A(n6160), .ZN(n5549) );
  NAND2_X1 U6218 ( .A1(n6941), .A2(n5549), .ZN(n7094) );
  INV_X1 U6219 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6681) );
  NOR2_X1 U6220 ( .A1(n7014), .A2(n6681), .ZN(n6051) );
  INV_X1 U6221 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6683) );
  NAND3_X1 U6222 ( .A1(n7139), .A2(n6051), .A3(n6683), .ZN(n5550) );
  OAI211_X1 U6223 ( .C1(n7122), .C2(n5551), .A(n7094), .B(n5550), .ZN(n5552)
         );
  AOI211_X1 U6224 ( .C1(REIP_REG_10__SCAN_IN), .C2(n5554), .A(n5553), .B(n5552), .ZN(n5556) );
  NAND2_X1 U6225 ( .A1(n7133), .A2(n6020), .ZN(n5555) );
  OAI211_X1 U6226 ( .C1(n6017), .C2(n7130), .A(n5556), .B(n5555), .ZN(U2817)
         );
  XNOR2_X1 U6227 ( .A(n5557), .B(n5558), .ZN(n5570) );
  NAND2_X1 U6228 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6032) );
  NOR2_X1 U6229 ( .A1(n4782), .A2(n5559), .ZN(n6881) );
  INV_X1 U6230 ( .A(n6881), .ZN(n6031) );
  AOI211_X1 U6231 ( .C1(n5561), .C2(n6890), .A(n6865), .B(n6031), .ZN(n5564)
         );
  NAND2_X1 U6232 ( .A1(n6908), .A2(REIP_REG_8__SCAN_IN), .ZN(n5566) );
  OAI21_X1 U6233 ( .B1(n6884), .B2(n7005), .A(n5566), .ZN(n5563) );
  OAI22_X1 U6234 ( .A1(n6862), .A2(n6031), .B1(n5560), .B2(n6467), .ZN(n6889)
         );
  NOR2_X1 U6235 ( .A1(n6889), .A2(n5561), .ZN(n5562) );
  AOI211_X1 U6236 ( .C1(n6032), .C2(n5564), .A(n5563), .B(n5562), .ZN(n5565)
         );
  OAI21_X1 U6237 ( .B1(n6619), .B2(n5570), .A(n5565), .ZN(U3010) );
  INV_X1 U6238 ( .A(DATAI_10_), .ZN(n7302) );
  INV_X1 U6239 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7307) );
  OAI222_X1 U6240 ( .A1(n6017), .A2(n7335), .B1(n7302), .B2(n6343), .C1(n6142), 
        .C2(n7307), .ZN(U2881) );
  OAI21_X1 U6241 ( .B1(n6448), .B2(n3699), .A(n5566), .ZN(n5568) );
  NOR2_X1 U6242 ( .A1(n7008), .A2(n6791), .ZN(n5567) );
  AOI211_X1 U6243 ( .C1(n6801), .C2(n7009), .A(n5568), .B(n5567), .ZN(n5569)
         );
  OAI21_X1 U6244 ( .B1(n6804), .B2(n5570), .A(n5569), .ZN(U2978) );
  INV_X1 U6245 ( .A(n7360), .ZN(n5578) );
  OAI21_X1 U6246 ( .B1(n3642), .B2(n5608), .A(n7400), .ZN(n5571) );
  OAI21_X1 U6247 ( .B1(n7359), .B2(n5578), .A(n5571), .ZN(n5573) );
  NOR2_X1 U6248 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5572), .ZN(n5609)
         );
  AOI21_X1 U6249 ( .B1(n5573), .B2(n7214), .A(n5609), .ZN(n5575) );
  NOR3_X2 U6250 ( .A1(n5575), .A2(n7379), .A3(n5574), .ZN(n5615) );
  INV_X1 U6251 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5583) );
  AOI22_X1 U6252 ( .A1(n7499), .A2(n5609), .B1(n7501), .B2(n5608), .ZN(n5582)
         );
  OAI22_X1 U6253 ( .A1(n5579), .A2(n5578), .B1(n5577), .B2(n5576), .ZN(n5610)
         );
  AOI22_X1 U6254 ( .A1(n5580), .A2(n5610), .B1(n7500), .B2(n3642), .ZN(n5581)
         );
  OAI211_X1 U6255 ( .C1(n5615), .C2(n5583), .A(n5582), .B(n5581), .ZN(U3040)
         );
  INV_X1 U6256 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5587) );
  AOI22_X1 U6257 ( .A1(n7467), .A2(n5609), .B1(n7469), .B2(n5608), .ZN(n5586)
         );
  AOI22_X1 U6258 ( .A1(n5584), .A2(n5610), .B1(n7468), .B2(n3642), .ZN(n5585)
         );
  OAI211_X1 U6259 ( .C1(n5615), .C2(n5587), .A(n5586), .B(n5585), .ZN(U3038)
         );
  INV_X1 U6260 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5591) );
  AOI22_X1 U6261 ( .A1(n7531), .A2(n5609), .B1(n7533), .B2(n5608), .ZN(n5590)
         );
  AOI22_X1 U6262 ( .A1(n5588), .A2(n5610), .B1(n7532), .B2(n3642), .ZN(n5589)
         );
  OAI211_X1 U6263 ( .C1(n5615), .C2(n5591), .A(n5590), .B(n5589), .ZN(U3042)
         );
  INV_X1 U6264 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5595) );
  AOI22_X1 U6265 ( .A1(n7451), .A2(n5609), .B1(n7452), .B2(n5608), .ZN(n5594)
         );
  AOI22_X1 U6266 ( .A1(n5592), .A2(n5610), .B1(n7453), .B2(n3642), .ZN(n5593)
         );
  OAI211_X1 U6267 ( .C1(n5615), .C2(n5595), .A(n5594), .B(n5593), .ZN(U3037)
         );
  INV_X1 U6268 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5599) );
  AOI22_X1 U6269 ( .A1(n7571), .A2(n5609), .B1(n7572), .B2(n5608), .ZN(n5598)
         );
  AOI22_X1 U6270 ( .A1(n5596), .A2(n5610), .B1(n7574), .B2(n3642), .ZN(n5597)
         );
  OAI211_X1 U6271 ( .C1(n5615), .C2(n5599), .A(n5598), .B(n5597), .ZN(U3043)
         );
  INV_X1 U6272 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5603) );
  AOI22_X1 U6273 ( .A1(n7421), .A2(n5609), .B1(n7430), .B2(n5608), .ZN(n5602)
         );
  AOI22_X1 U6274 ( .A1(n5600), .A2(n5610), .B1(n7422), .B2(n3642), .ZN(n5601)
         );
  OAI211_X1 U6275 ( .C1(n5615), .C2(n5603), .A(n5602), .B(n5601), .ZN(U3036)
         );
  INV_X1 U6276 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5607) );
  AOI22_X1 U6277 ( .A1(n7483), .A2(n5609), .B1(n7485), .B2(n5608), .ZN(n5606)
         );
  AOI22_X1 U6278 ( .A1(n5604), .A2(n5610), .B1(n7484), .B2(n3642), .ZN(n5605)
         );
  OAI211_X1 U6279 ( .C1(n5615), .C2(n5607), .A(n5606), .B(n5605), .ZN(U3039)
         );
  INV_X1 U6280 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5614) );
  AOI22_X1 U6281 ( .A1(n7515), .A2(n5609), .B1(n7516), .B2(n5608), .ZN(n5613)
         );
  AOI22_X1 U6282 ( .A1(n5611), .A2(n5610), .B1(n7517), .B2(n3642), .ZN(n5612)
         );
  OAI211_X1 U6283 ( .C1(n5615), .C2(n5614), .A(n5613), .B(n5612), .ZN(U3041)
         );
  XOR2_X1 U6284 ( .A(n5616), .B(n5617), .Z(n6887) );
  NAND2_X1 U6285 ( .A1(n6887), .A2(n6819), .ZN(n5621) );
  NAND2_X1 U6286 ( .A1(n6908), .A2(REIP_REG_7__SCAN_IN), .ZN(n6883) );
  INV_X1 U6287 ( .A(n6883), .ZN(n5619) );
  NOR2_X1 U6288 ( .A1(n6822), .A2(n6994), .ZN(n5618) );
  AOI211_X1 U6289 ( .C1(n4711), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5619), 
        .B(n5618), .ZN(n5620) );
  OAI211_X1 U6290 ( .C1(n6791), .C2(n6995), .A(n5621), .B(n5620), .ZN(U2979)
         );
  OAI21_X1 U6291 ( .B1(n5622), .B2(n5625), .A(n5623), .ZN(n6800) );
  XOR2_X1 U6292 ( .A(n6047), .B(n6048), .Z(n7038) );
  AOI22_X1 U6293 ( .A1(n7038), .A2(n6769), .B1(EBX_REG_12__SCAN_IN), .B2(n6311), .ZN(n5626) );
  OAI21_X1 U6294 ( .B1(n6800), .B2(n6315), .A(n5626), .ZN(U2847) );
  INV_X1 U6295 ( .A(n5627), .ZN(n5629) );
  INV_X1 U6296 ( .A(n5541), .ZN(n5628) );
  AOI21_X1 U6297 ( .B1(n5629), .B2(n5628), .A(n5622), .ZN(n7034) );
  INV_X1 U6298 ( .A(n7034), .ZN(n5633) );
  INV_X1 U6299 ( .A(DATAI_11_), .ZN(n7308) );
  INV_X1 U6300 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7313) );
  OAI222_X1 U6301 ( .A1(n5633), .A2(n7335), .B1(n7308), .B2(n6343), .C1(n6142), 
        .C2(n7313), .ZN(U2880) );
  INV_X1 U6302 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5632) );
  OAI21_X1 U6303 ( .B1(n5631), .B2(n5630), .A(n6048), .ZN(n6897) );
  OAI222_X1 U6304 ( .A1(n5633), .A2(n6315), .B1(n5632), .B2(n6773), .C1(n6320), 
        .C2(n6897), .ZN(U2848) );
  INV_X1 U6305 ( .A(DATAI_12_), .ZN(n7314) );
  OAI222_X1 U6306 ( .A1(n6800), .A2(n7335), .B1(n7314), .B2(n6343), .C1(n6142), 
        .C2(n4304), .ZN(U2879) );
  INV_X1 U6307 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6645) );
  XNOR2_X1 U6308 ( .A(n6645), .B(keyinput_127), .ZN(n6001) );
  XOR2_X1 U6309 ( .A(DATAI_26_), .B(keyinput_5), .Z(n5637) );
  XNOR2_X1 U6310 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n5636) );
  XNOR2_X1 U6311 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n5635) );
  XNOR2_X1 U6312 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n5634) );
  NOR4_X1 U6313 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n5650)
         );
  XOR2_X1 U6314 ( .A(DATAI_31_), .B(keyinput_0), .Z(n5640) );
  XOR2_X1 U6315 ( .A(DATAI_30_), .B(keyinput_1), .Z(n5639) );
  XNOR2_X1 U6316 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n5638) );
  AOI21_X1 U6317 ( .B1(n5640), .B2(n5639), .A(n5638), .ZN(n5643) );
  XOR2_X1 U6318 ( .A(DATAI_27_), .B(keyinput_4), .Z(n5642) );
  XNOR2_X1 U6319 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n5641) );
  NAND3_X1 U6320 ( .A1(n5643), .A2(n5642), .A3(n5641), .ZN(n5649) );
  XOR2_X1 U6321 ( .A(DATAI_21_), .B(keyinput_10), .Z(n5647) );
  XOR2_X1 U6322 ( .A(DATAI_22_), .B(keyinput_9), .Z(n5646) );
  XOR2_X1 U6323 ( .A(DATAI_20_), .B(keyinput_11), .Z(n5645) );
  XOR2_X1 U6324 ( .A(DATAI_19_), .B(keyinput_12), .Z(n5644) );
  NAND4_X1 U6325 ( .A1(n5647), .A2(n5646), .A3(n5645), .A4(n5644), .ZN(n5648)
         );
  AOI21_X1 U6326 ( .B1(n5650), .B2(n5649), .A(n5648), .ZN(n5653) );
  XOR2_X1 U6327 ( .A(DATAI_18_), .B(keyinput_13), .Z(n5652) );
  XNOR2_X1 U6328 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n5651) );
  OAI21_X1 U6329 ( .B1(n5653), .B2(n5652), .A(n5651), .ZN(n5656) );
  XNOR2_X1 U6330 ( .A(DATAI_16_), .B(keyinput_15), .ZN(n5655) );
  XNOR2_X1 U6331 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n5654) );
  NAND3_X1 U6332 ( .A1(n5656), .A2(n5655), .A3(n5654), .ZN(n5659) );
  XOR2_X1 U6333 ( .A(DATAI_14_), .B(keyinput_17), .Z(n5658) );
  XOR2_X1 U6334 ( .A(DATAI_13_), .B(keyinput_18), .Z(n5657) );
  AOI21_X1 U6335 ( .B1(n5659), .B2(n5658), .A(n5657), .ZN(n5665) );
  XOR2_X1 U6336 ( .A(DATAI_12_), .B(keyinput_19), .Z(n5664) );
  XOR2_X1 U6337 ( .A(DATAI_10_), .B(keyinput_21), .Z(n5662) );
  XOR2_X1 U6338 ( .A(DATAI_11_), .B(keyinput_20), .Z(n5661) );
  XNOR2_X1 U6339 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n5660) );
  NOR3_X1 U6340 ( .A1(n5662), .A2(n5661), .A3(n5660), .ZN(n5663) );
  OAI21_X1 U6341 ( .B1(n5665), .B2(n5664), .A(n5663), .ZN(n5672) );
  XOR2_X1 U6342 ( .A(keyinput_24), .B(DATAI_7_), .Z(n5671) );
  XOR2_X1 U6343 ( .A(DATAI_6_), .B(keyinput_25), .Z(n5670) );
  XOR2_X1 U6344 ( .A(DATAI_4_), .B(keyinput_27), .Z(n5668) );
  XNOR2_X1 U6345 ( .A(keyinput_23), .B(DATAI_8_), .ZN(n5667) );
  XNOR2_X1 U6346 ( .A(keyinput_26), .B(DATAI_5_), .ZN(n5666) );
  NOR3_X1 U6347 ( .A1(n5668), .A2(n5667), .A3(n5666), .ZN(n5669) );
  NAND4_X1 U6348 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n5675)
         );
  XOR2_X1 U6349 ( .A(DATAI_2_), .B(keyinput_29), .Z(n5674) );
  XNOR2_X1 U6350 ( .A(keyinput_28), .B(DATAI_3_), .ZN(n5673) );
  NAND3_X1 U6351 ( .A1(n5675), .A2(n5674), .A3(n5673), .ZN(n5678) );
  XNOR2_X1 U6352 ( .A(keyinput_30), .B(DATAI_1_), .ZN(n5677) );
  XOR2_X1 U6353 ( .A(DATAI_0_), .B(keyinput_31), .Z(n5676) );
  AOI21_X1 U6354 ( .B1(n5678), .B2(n5677), .A(n5676), .ZN(n5684) );
  XOR2_X1 U6355 ( .A(keyinput_32), .B(MEMORYFETCH_REG_SCAN_IN), .Z(n5683) );
  XOR2_X1 U6356 ( .A(keyinput_33), .B(NA_N), .Z(n5681) );
  XNOR2_X1 U6357 ( .A(n7250), .B(keyinput_35), .ZN(n5680) );
  INV_X1 U6358 ( .A(BS16_N), .ZN(n6624) );
  XNOR2_X1 U6359 ( .A(n6624), .B(keyinput_34), .ZN(n5679) );
  NOR3_X1 U6360 ( .A1(n5681), .A2(n5680), .A3(n5679), .ZN(n5682) );
  OAI21_X1 U6361 ( .B1(n5684), .B2(n5683), .A(n5682), .ZN(n5687) );
  XOR2_X1 U6362 ( .A(keyinput_37), .B(READREQUEST_REG_SCAN_IN), .Z(n5686) );
  XNOR2_X1 U6363 ( .A(keyinput_36), .B(HOLD), .ZN(n5685) );
  NAND3_X1 U6364 ( .A1(n5687), .A2(n5686), .A3(n5685), .ZN(n5690) );
  INV_X1 U6365 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6650) );
  XNOR2_X1 U6366 ( .A(n6650), .B(keyinput_38), .ZN(n5689) );
  INV_X1 U6367 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6824) );
  XNOR2_X1 U6368 ( .A(n6824), .B(keyinput_39), .ZN(n5688) );
  NAND3_X1 U6369 ( .A1(n5690), .A2(n5689), .A3(n5688), .ZN(n5693) );
  XNOR2_X1 U6370 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .ZN(n5692) );
  XNOR2_X1 U6371 ( .A(keyinput_41), .B(D_C_N_REG_SCAN_IN), .ZN(n5691) );
  NAND3_X1 U6372 ( .A1(n5693), .A2(n5692), .A3(n5691), .ZN(n5696) );
  XNOR2_X1 U6373 ( .A(n7413), .B(keyinput_43), .ZN(n5695) );
  XOR2_X1 U6374 ( .A(keyinput_42), .B(REQUESTPENDING_REG_SCAN_IN), .Z(n5694)
         );
  NAND3_X1 U6375 ( .A1(n5696), .A2(n5695), .A3(n5694), .ZN(n5704) );
  XOR2_X1 U6376 ( .A(keyinput_48), .B(BYTEENABLE_REG_1__SCAN_IN), .Z(n5703) );
  XOR2_X1 U6377 ( .A(keyinput_47), .B(BYTEENABLE_REG_0__SCAN_IN), .Z(n5702) );
  XOR2_X1 U6378 ( .A(keyinput_44), .B(MORE_REG_SCAN_IN), .Z(n5700) );
  XNOR2_X1 U6379 ( .A(keyinput_45), .B(FLUSH_REG_SCAN_IN), .ZN(n5699) );
  XNOR2_X1 U6380 ( .A(keyinput_49), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n5698)
         );
  XNOR2_X1 U6381 ( .A(keyinput_46), .B(W_R_N_REG_SCAN_IN), .ZN(n5697) );
  NOR4_X1 U6382 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n5701)
         );
  NAND4_X1 U6383 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), .ZN(n5707)
         );
  INV_X1 U6384 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6721) );
  XNOR2_X1 U6385 ( .A(n6721), .B(keyinput_50), .ZN(n5706) );
  XOR2_X1 U6386 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n5705) );
  NAND3_X1 U6387 ( .A1(n5707), .A2(n5706), .A3(n5705), .ZN(n5710) );
  XNOR2_X1 U6388 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .ZN(n5709) );
  XNOR2_X1 U6389 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n5708) );
  NAND3_X1 U6390 ( .A1(n5710), .A2(n5709), .A3(n5708), .ZN(n5714) );
  XOR2_X1 U6391 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .Z(n5713) );
  XOR2_X1 U6392 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .Z(n5712) );
  XNOR2_X1 U6393 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .ZN(n5711) );
  NAND4_X1 U6394 ( .A1(n5714), .A2(n5713), .A3(n5712), .A4(n5711), .ZN(n5718)
         );
  XOR2_X1 U6395 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .Z(n5717) );
  XOR2_X1 U6396 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .Z(n5716) );
  XOR2_X1 U6397 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .Z(n5715) );
  NAND4_X1 U6398 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .ZN(n5722)
         );
  XOR2_X1 U6399 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .Z(n5721) );
  XNOR2_X1 U6400 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n5720) );
  XNOR2_X1 U6401 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n5719) );
  NAND4_X1 U6402 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n5725)
         );
  XNOR2_X1 U6403 ( .A(keyinput_63), .B(REIP_REG_19__SCAN_IN), .ZN(n5724) );
  XOR2_X1 U6404 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .Z(n5723) );
  AOI21_X1 U6405 ( .B1(n5725), .B2(n5724), .A(n5723), .ZN(n5728) );
  XOR2_X1 U6406 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n5727) );
  XNOR2_X1 U6407 ( .A(keyinput_65), .B(REIP_REG_17__SCAN_IN), .ZN(n5726) );
  NOR3_X1 U6408 ( .A1(n5728), .A2(n5727), .A3(n5726), .ZN(n5731) );
  INV_X1 U6409 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6720) );
  XNOR2_X1 U6410 ( .A(n6720), .B(keyinput_67), .ZN(n5730) );
  XNOR2_X1 U6411 ( .A(keyinput_68), .B(BE_N_REG_2__SCAN_IN), .ZN(n5729) );
  OAI21_X1 U6412 ( .B1(n5731), .B2(n5730), .A(n5729), .ZN(n5734) );
  XNOR2_X1 U6413 ( .A(keyinput_70), .B(BE_N_REG_0__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U6414 ( .A(keyinput_69), .B(BE_N_REG_1__SCAN_IN), .ZN(n5732) );
  NAND3_X1 U6415 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n5737) );
  XNOR2_X1 U6416 ( .A(keyinput_71), .B(ADDRESS_REG_29__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U6417 ( .A(keyinput_72), .B(ADDRESS_REG_28__SCAN_IN), .ZN(n5735) );
  AOI21_X1 U6418 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n5744) );
  XOR2_X1 U6419 ( .A(keyinput_76), .B(ADDRESS_REG_24__SCAN_IN), .Z(n5741) );
  INV_X1 U6420 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6707) );
  XNOR2_X1 U6421 ( .A(n6707), .B(keyinput_75), .ZN(n5740) );
  XNOR2_X1 U6422 ( .A(keyinput_74), .B(ADDRESS_REG_26__SCAN_IN), .ZN(n5739) );
  XNOR2_X1 U6423 ( .A(keyinput_73), .B(ADDRESS_REG_27__SCAN_IN), .ZN(n5738) );
  NAND4_X1 U6424 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), .ZN(n5743)
         );
  XNOR2_X1 U6425 ( .A(keyinput_77), .B(ADDRESS_REG_23__SCAN_IN), .ZN(n5742) );
  OAI21_X1 U6426 ( .B1(n5744), .B2(n5743), .A(n5742), .ZN(n5747) );
  INV_X1 U6427 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6701) );
  XNOR2_X1 U6428 ( .A(n6701), .B(keyinput_78), .ZN(n5746) );
  INV_X1 U6429 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6700) );
  XNOR2_X1 U6430 ( .A(n6700), .B(keyinput_79), .ZN(n5745) );
  AOI21_X1 U6431 ( .B1(n5747), .B2(n5746), .A(n5745), .ZN(n5750) );
  INV_X1 U6432 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6698) );
  XNOR2_X1 U6433 ( .A(n6698), .B(keyinput_80), .ZN(n5749) );
  INV_X1 U6434 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6697) );
  XNOR2_X1 U6435 ( .A(n6697), .B(keyinput_81), .ZN(n5748) );
  NOR3_X1 U6436 ( .A1(n5750), .A2(n5749), .A3(n5748), .ZN(n5754) );
  XOR2_X1 U6437 ( .A(keyinput_82), .B(ADDRESS_REG_18__SCAN_IN), .Z(n5753) );
  XNOR2_X1 U6438 ( .A(keyinput_84), .B(ADDRESS_REG_16__SCAN_IN), .ZN(n5752) );
  XNOR2_X1 U6439 ( .A(keyinput_83), .B(ADDRESS_REG_17__SCAN_IN), .ZN(n5751) );
  NOR4_X1 U6440 ( .A1(n5754), .A2(n5753), .A3(n5752), .A4(n5751), .ZN(n5757)
         );
  XNOR2_X1 U6441 ( .A(keyinput_86), .B(ADDRESS_REG_14__SCAN_IN), .ZN(n5756) );
  XNOR2_X1 U6442 ( .A(keyinput_85), .B(ADDRESS_REG_15__SCAN_IN), .ZN(n5755) );
  NOR3_X1 U6443 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(n5761) );
  XOR2_X1 U6444 ( .A(keyinput_88), .B(ADDRESS_REG_12__SCAN_IN), .Z(n5760) );
  XNOR2_X1 U6445 ( .A(keyinput_89), .B(ADDRESS_REG_11__SCAN_IN), .ZN(n5759) );
  XNOR2_X1 U6446 ( .A(keyinput_87), .B(ADDRESS_REG_13__SCAN_IN), .ZN(n5758) );
  NOR4_X1 U6447 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n5765)
         );
  INV_X1 U6448 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6682) );
  XNOR2_X1 U6449 ( .A(n6682), .B(keyinput_92), .ZN(n5764) );
  INV_X1 U6450 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6685) );
  XNOR2_X1 U6451 ( .A(n6685), .B(keyinput_90), .ZN(n5763) );
  XNOR2_X1 U6452 ( .A(keyinput_91), .B(ADDRESS_REG_9__SCAN_IN), .ZN(n5762) );
  NOR4_X1 U6453 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n5768)
         );
  INV_X1 U6454 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6680) );
  XNOR2_X1 U6455 ( .A(n6680), .B(keyinput_93), .ZN(n5767) );
  XNOR2_X1 U6456 ( .A(keyinput_94), .B(ADDRESS_REG_6__SCAN_IN), .ZN(n5766) );
  NOR3_X1 U6457 ( .A1(n5768), .A2(n5767), .A3(n5766), .ZN(n5771) );
  INV_X1 U6458 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6676) );
  XNOR2_X1 U6459 ( .A(n6676), .B(keyinput_96), .ZN(n5770) );
  XNOR2_X1 U6460 ( .A(keyinput_95), .B(ADDRESS_REG_5__SCAN_IN), .ZN(n5769) );
  NOR3_X1 U6461 ( .A1(n5771), .A2(n5770), .A3(n5769), .ZN(n5774) );
  INV_X1 U6462 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6675) );
  XNOR2_X1 U6463 ( .A(n6675), .B(keyinput_97), .ZN(n5773) );
  XNOR2_X1 U6464 ( .A(keyinput_98), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n5772) );
  NOR3_X1 U6465 ( .A1(n5774), .A2(n5773), .A3(n5772), .ZN(n5777) );
  XNOR2_X1 U6466 ( .A(keyinput_100), .B(ADDRESS_REG_0__SCAN_IN), .ZN(n5776) );
  XNOR2_X1 U6467 ( .A(keyinput_99), .B(ADDRESS_REG_1__SCAN_IN), .ZN(n5775) );
  NOR3_X1 U6468 ( .A1(n5777), .A2(n5776), .A3(n5775), .ZN(n5781) );
  XNOR2_X1 U6469 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .ZN(n5780) );
  XNOR2_X1 U6470 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .ZN(n5779) );
  XNOR2_X1 U6471 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .ZN(n5778) );
  OAI211_X1 U6472 ( .C1(n5781), .C2(n5780), .A(n5779), .B(n5778), .ZN(n5789)
         );
  XOR2_X1 U6473 ( .A(keyinput_104), .B(DATAWIDTH_REG_0__SCAN_IN), .Z(n5785) );
  INV_X1 U6474 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6626) );
  XNOR2_X1 U6475 ( .A(n6626), .B(keyinput_106), .ZN(n5784) );
  INV_X1 U6476 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7228) );
  XNOR2_X1 U6477 ( .A(n7228), .B(keyinput_105), .ZN(n5783) );
  INV_X1 U6478 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6627) );
  XNOR2_X1 U6479 ( .A(n6627), .B(keyinput_107), .ZN(n5782) );
  NOR4_X1 U6480 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5788)
         );
  XNOR2_X1 U6481 ( .A(keyinput_109), .B(DATAWIDTH_REG_5__SCAN_IN), .ZN(n5787)
         );
  XNOR2_X1 U6482 ( .A(keyinput_108), .B(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5786)
         );
  NAND4_X1 U6483 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n5795)
         );
  XNOR2_X1 U6484 ( .A(keyinput_110), .B(DATAWIDTH_REG_6__SCAN_IN), .ZN(n5794)
         );
  XOR2_X1 U6485 ( .A(keyinput_112), .B(DATAWIDTH_REG_8__SCAN_IN), .Z(n5792) );
  INV_X1 U6486 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6632) );
  XNOR2_X1 U6487 ( .A(n6632), .B(keyinput_113), .ZN(n5791) );
  XNOR2_X1 U6488 ( .A(keyinput_111), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n5790)
         );
  NAND3_X1 U6489 ( .A1(n5792), .A2(n5791), .A3(n5790), .ZN(n5793) );
  AOI21_X1 U6490 ( .B1(n5795), .B2(n5794), .A(n5793), .ZN(n5799) );
  INV_X1 U6491 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U6492 ( .A(n6633), .B(keyinput_115), .ZN(n5798) );
  XNOR2_X1 U6493 ( .A(keyinput_114), .B(DATAWIDTH_REG_10__SCAN_IN), .ZN(n5797)
         );
  XNOR2_X1 U6494 ( .A(keyinput_116), .B(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5796)
         );
  NOR4_X1 U6495 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(n5802)
         );
  XNOR2_X1 U6496 ( .A(keyinput_117), .B(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5801)
         );
  XNOR2_X1 U6497 ( .A(keyinput_118), .B(DATAWIDTH_REG_14__SCAN_IN), .ZN(n5800)
         );
  NOR3_X1 U6498 ( .A1(n5802), .A2(n5801), .A3(n5800), .ZN(n5805) );
  INV_X1 U6499 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6638) );
  XNOR2_X1 U6500 ( .A(n6638), .B(keyinput_120), .ZN(n5804) );
  XNOR2_X1 U6501 ( .A(keyinput_119), .B(DATAWIDTH_REG_15__SCAN_IN), .ZN(n5803)
         );
  NOR3_X1 U6502 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n5808) );
  INV_X1 U6503 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6640) );
  XNOR2_X1 U6504 ( .A(n6640), .B(keyinput_122), .ZN(n5807) );
  INV_X1 U6505 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6639) );
  XNOR2_X1 U6506 ( .A(n6639), .B(keyinput_121), .ZN(n5806) );
  NOR3_X1 U6507 ( .A1(n5808), .A2(n5807), .A3(n5806), .ZN(n5814) );
  XNOR2_X1 U6508 ( .A(keyinput_123), .B(DATAWIDTH_REG_19__SCAN_IN), .ZN(n5813)
         );
  INV_X1 U6509 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6643) );
  XNOR2_X1 U6510 ( .A(n6643), .B(keyinput_125), .ZN(n5811) );
  XNOR2_X1 U6511 ( .A(keyinput_124), .B(DATAWIDTH_REG_20__SCAN_IN), .ZN(n5810)
         );
  XNOR2_X1 U6512 ( .A(keyinput_126), .B(DATAWIDTH_REG_22__SCAN_IN), .ZN(n5809)
         );
  NOR3_X1 U6513 ( .A1(n5811), .A2(n5810), .A3(n5809), .ZN(n5812) );
  OAI21_X1 U6514 ( .B1(n5814), .B2(n5813), .A(n5812), .ZN(n6000) );
  XNOR2_X1 U6515 ( .A(DATAWIDTH_REG_23__SCAN_IN), .B(keyinput_255), .ZN(n5999)
         );
  XNOR2_X1 U6516 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n5818) );
  XNOR2_X1 U6517 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n5817) );
  XNOR2_X1 U6518 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n5816) );
  XNOR2_X1 U6519 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n5815) );
  NOR4_X1 U6520 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n5832)
         );
  XOR2_X1 U6521 ( .A(DATAI_31_), .B(keyinput_128), .Z(n5821) );
  XOR2_X1 U6522 ( .A(DATAI_30_), .B(keyinput_129), .Z(n5820) );
  XNOR2_X1 U6523 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n5819) );
  AOI21_X1 U6524 ( .B1(n5821), .B2(n5820), .A(n5819), .ZN(n5824) );
  XOR2_X1 U6525 ( .A(DATAI_27_), .B(keyinput_132), .Z(n5823) );
  XNOR2_X1 U6526 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n5822) );
  NAND3_X1 U6527 ( .A1(n5824), .A2(n5823), .A3(n5822), .ZN(n5831) );
  INV_X1 U6528 ( .A(keyinput_138), .ZN(n5825) );
  XNOR2_X1 U6529 ( .A(n5825), .B(DATAI_21_), .ZN(n5829) );
  XNOR2_X1 U6530 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n5828) );
  XNOR2_X1 U6531 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n5827) );
  XNOR2_X1 U6532 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n5826) );
  NAND4_X1 U6533 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(n5830)
         );
  AOI21_X1 U6534 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5835) );
  XOR2_X1 U6535 ( .A(DATAI_18_), .B(keyinput_141), .Z(n5834) );
  XOR2_X1 U6536 ( .A(DATAI_17_), .B(keyinput_142), .Z(n5833) );
  OAI21_X1 U6537 ( .B1(n5835), .B2(n5834), .A(n5833), .ZN(n5838) );
  XOR2_X1 U6538 ( .A(DATAI_16_), .B(keyinput_143), .Z(n5837) );
  XNOR2_X1 U6539 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n5836) );
  NAND3_X1 U6540 ( .A1(n5838), .A2(n5837), .A3(n5836), .ZN(n5841) );
  XOR2_X1 U6541 ( .A(DATAI_14_), .B(keyinput_145), .Z(n5840) );
  XNOR2_X1 U6542 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n5839) );
  AOI21_X1 U6543 ( .B1(n5841), .B2(n5840), .A(n5839), .ZN(n5847) );
  XOR2_X1 U6544 ( .A(DATAI_12_), .B(keyinput_147), .Z(n5846) );
  XOR2_X1 U6545 ( .A(DATAI_9_), .B(keyinput_150), .Z(n5844) );
  XOR2_X1 U6546 ( .A(DATAI_11_), .B(keyinput_148), .Z(n5843) );
  XNOR2_X1 U6547 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n5842) );
  NOR3_X1 U6548 ( .A1(n5844), .A2(n5843), .A3(n5842), .ZN(n5845) );
  OAI21_X1 U6549 ( .B1(n5847), .B2(n5846), .A(n5845), .ZN(n5855) );
  OAI22_X1 U6550 ( .A1(n5849), .A2(keyinput_152), .B1(keyinput_154), .B2(
        DATAI_5_), .ZN(n5848) );
  AOI221_X1 U6551 ( .B1(n5849), .B2(keyinput_152), .C1(DATAI_5_), .C2(
        keyinput_154), .A(n5848), .ZN(n5854) );
  XOR2_X1 U6552 ( .A(DATAI_6_), .B(keyinput_153), .Z(n5853) );
  OAI22_X1 U6553 ( .A1(n5851), .A2(keyinput_151), .B1(DATAI_4_), .B2(
        keyinput_155), .ZN(n5850) );
  AOI221_X1 U6554 ( .B1(n5851), .B2(keyinput_151), .C1(keyinput_155), .C2(
        DATAI_4_), .A(n5850), .ZN(n5852) );
  NAND4_X1 U6555 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n5858)
         );
  XOR2_X1 U6556 ( .A(DATAI_3_), .B(keyinput_156), .Z(n5857) );
  XOR2_X1 U6557 ( .A(DATAI_2_), .B(keyinput_157), .Z(n5856) );
  NAND3_X1 U6558 ( .A1(n5858), .A2(n5857), .A3(n5856), .ZN(n5861) );
  XNOR2_X1 U6559 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n5860) );
  XNOR2_X1 U6560 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n5859) );
  AOI21_X1 U6561 ( .B1(n5861), .B2(n5860), .A(n5859), .ZN(n5863) );
  XOR2_X1 U6562 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_160), .Z(n5862) );
  NOR2_X1 U6563 ( .A1(n5863), .A2(n5862), .ZN(n5867) );
  XNOR2_X1 U6564 ( .A(n7250), .B(keyinput_163), .ZN(n5866) );
  XNOR2_X1 U6565 ( .A(n6624), .B(keyinput_162), .ZN(n5865) );
  XNOR2_X1 U6566 ( .A(NA_N), .B(keyinput_161), .ZN(n5864) );
  NOR4_X1 U6567 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n5870)
         );
  XOR2_X1 U6568 ( .A(HOLD), .B(keyinput_164), .Z(n5869) );
  XNOR2_X1 U6569 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_165), .ZN(n5868)
         );
  NOR3_X1 U6570 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n5873) );
  XNOR2_X1 U6571 ( .A(n6650), .B(keyinput_166), .ZN(n5872) );
  XNOR2_X1 U6572 ( .A(n6824), .B(keyinput_167), .ZN(n5871) );
  NOR3_X1 U6573 ( .A1(n5873), .A2(n5872), .A3(n5871), .ZN(n5876) );
  INV_X1 U6574 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7247) );
  XNOR2_X1 U6575 ( .A(n7247), .B(keyinput_168), .ZN(n5875) );
  INV_X1 U6576 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U6577 ( .A(n6826), .B(keyinput_169), .ZN(n5874) );
  NOR3_X1 U6578 ( .A1(n5876), .A2(n5875), .A3(n5874), .ZN(n5879) );
  XOR2_X1 U6579 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_170), .Z(n5878)
         );
  XNOR2_X1 U6580 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_171), .ZN(n5877) );
  NOR3_X1 U6581 ( .A1(n5879), .A2(n5878), .A3(n5877), .ZN(n5887) );
  XNOR2_X1 U6582 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_173), .ZN(n5886) );
  XNOR2_X1 U6583 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_177), .ZN(n5885)
         );
  XOR2_X1 U6584 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_176), .Z(n5883)
         );
  XOR2_X1 U6585 ( .A(MORE_REG_SCAN_IN), .B(keyinput_172), .Z(n5882) );
  XOR2_X1 U6586 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_174), .Z(n5881) );
  XOR2_X1 U6587 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_175), .Z(n5880)
         );
  NAND4_X1 U6588 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n5884)
         );
  NOR4_X1 U6589 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n5890)
         );
  XNOR2_X1 U6590 ( .A(n6721), .B(keyinput_178), .ZN(n5889) );
  XOR2_X1 U6591 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .Z(n5888) );
  NOR3_X1 U6592 ( .A1(n5890), .A2(n5889), .A3(n5888), .ZN(n5893) );
  INV_X1 U6593 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6716) );
  XNOR2_X1 U6594 ( .A(n6716), .B(keyinput_180), .ZN(n5892) );
  XOR2_X1 U6595 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .Z(n5891) );
  NOR3_X1 U6596 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n5897) );
  XOR2_X1 U6597 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .Z(n5896) );
  XOR2_X1 U6598 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .Z(n5895) );
  XNOR2_X1 U6599 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n5894) );
  NOR4_X1 U6600 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(n5901)
         );
  XOR2_X1 U6601 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .Z(n5900) );
  XNOR2_X1 U6602 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .ZN(n5899) );
  XNOR2_X1 U6603 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n5898) );
  NOR4_X1 U6604 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5905)
         );
  XOR2_X1 U6605 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .Z(n5904) );
  XNOR2_X1 U6606 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .ZN(n5903) );
  XNOR2_X1 U6607 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .ZN(n5902) );
  NOR4_X1 U6608 ( .A1(n5905), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(n5908)
         );
  XOR2_X1 U6609 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n5907) );
  XNOR2_X1 U6610 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .ZN(n5906) );
  OAI21_X1 U6611 ( .B1(n5908), .B2(n5907), .A(n5906), .ZN(n5911) );
  XOR2_X1 U6612 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .Z(n5910) );
  XOR2_X1 U6613 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .Z(n5909) );
  NAND3_X1 U6614 ( .A1(n5911), .A2(n5910), .A3(n5909), .ZN(n5914) );
  XNOR2_X1 U6615 ( .A(n6720), .B(keyinput_195), .ZN(n5913) );
  INV_X1 U6616 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6733) );
  XNOR2_X1 U6617 ( .A(n6733), .B(keyinput_196), .ZN(n5912) );
  AOI21_X1 U6618 ( .B1(n5914), .B2(n5913), .A(n5912), .ZN(n5917) );
  XNOR2_X1 U6619 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_197), .ZN(n5916) );
  XNOR2_X1 U6620 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_198), .ZN(n5915) );
  NOR3_X1 U6621 ( .A1(n5917), .A2(n5916), .A3(n5915), .ZN(n5920) );
  XNOR2_X1 U6622 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_199), .ZN(n5919)
         );
  XNOR2_X1 U6623 ( .A(ADDRESS_REG_28__SCAN_IN), .B(keyinput_200), .ZN(n5918)
         );
  OAI21_X1 U6624 ( .B1(n5920), .B2(n5919), .A(n5918), .ZN(n5927) );
  XNOR2_X1 U6625 ( .A(n6707), .B(keyinput_203), .ZN(n5924) );
  XNOR2_X1 U6626 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_204), .ZN(n5923)
         );
  XNOR2_X1 U6627 ( .A(ADDRESS_REG_27__SCAN_IN), .B(keyinput_201), .ZN(n5922)
         );
  XNOR2_X1 U6628 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_202), .ZN(n5921)
         );
  NOR4_X1 U6629 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n5926)
         );
  INV_X1 U6630 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6704) );
  XNOR2_X1 U6631 ( .A(n6704), .B(keyinput_205), .ZN(n5925) );
  AOI21_X1 U6632 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5930) );
  XNOR2_X1 U6633 ( .A(ADDRESS_REG_22__SCAN_IN), .B(keyinput_206), .ZN(n5929)
         );
  XNOR2_X1 U6634 ( .A(n6700), .B(keyinput_207), .ZN(n5928) );
  OAI21_X1 U6635 ( .B1(n5930), .B2(n5929), .A(n5928), .ZN(n5933) );
  XNOR2_X1 U6636 ( .A(n6697), .B(keyinput_209), .ZN(n5932) );
  XNOR2_X1 U6637 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_208), .ZN(n5931)
         );
  NAND3_X1 U6638 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(n5937) );
  XOR2_X1 U6639 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_212), .Z(n5936) );
  XNOR2_X1 U6640 ( .A(ADDRESS_REG_17__SCAN_IN), .B(keyinput_211), .ZN(n5935)
         );
  XNOR2_X1 U6641 ( .A(ADDRESS_REG_18__SCAN_IN), .B(keyinput_210), .ZN(n5934)
         );
  NAND4_X1 U6642 ( .A1(n5937), .A2(n5936), .A3(n5935), .A4(n5934), .ZN(n5940)
         );
  XNOR2_X1 U6643 ( .A(ADDRESS_REG_15__SCAN_IN), .B(keyinput_213), .ZN(n5939)
         );
  XNOR2_X1 U6644 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_214), .ZN(n5938)
         );
  NAND3_X1 U6645 ( .A1(n5940), .A2(n5939), .A3(n5938), .ZN(n5944) );
  XOR2_X1 U6646 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_216), .Z(n5943) );
  XOR2_X1 U6647 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_215), .Z(n5942) );
  XOR2_X1 U6648 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_217), .Z(n5941) );
  NAND4_X1 U6649 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5948)
         );
  XNOR2_X1 U6650 ( .A(n6685), .B(keyinput_218), .ZN(n5947) );
  XNOR2_X1 U6651 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_220), .ZN(n5946) );
  XNOR2_X1 U6652 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_219), .ZN(n5945) );
  NAND4_X1 U6653 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n5951)
         );
  XNOR2_X1 U6654 ( .A(n6680), .B(keyinput_221), .ZN(n5950) );
  XNOR2_X1 U6655 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_222), .ZN(n5949) );
  NAND3_X1 U6656 ( .A1(n5951), .A2(n5950), .A3(n5949), .ZN(n5954) );
  XNOR2_X1 U6657 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_224), .ZN(n5953) );
  XNOR2_X1 U6658 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_223), .ZN(n5952) );
  NAND3_X1 U6659 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n5957) );
  XOR2_X1 U6660 ( .A(ADDRESS_REG_2__SCAN_IN), .B(keyinput_226), .Z(n5956) );
  XNOR2_X1 U6661 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_225), .ZN(n5955) );
  NAND3_X1 U6662 ( .A1(n5957), .A2(n5956), .A3(n5955), .ZN(n5960) );
  XOR2_X1 U6663 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_227), .Z(n5959) );
  XOR2_X1 U6664 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_228), .Z(n5958) );
  NAND3_X1 U6665 ( .A1(n5960), .A2(n5959), .A3(n5958), .ZN(n5964) );
  XNOR2_X1 U6666 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_229), .ZN(n5963) );
  XNOR2_X1 U6667 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_230), .ZN(n5962) );
  XNOR2_X1 U6668 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_231), .ZN(n5961) );
  AOI211_X1 U6669 ( .C1(n5964), .C2(n5963), .A(n5962), .B(n5961), .ZN(n5972)
         );
  XNOR2_X1 U6670 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_237), .ZN(n5971)
         );
  XNOR2_X1 U6671 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .ZN(n5970)
         );
  XNOR2_X1 U6672 ( .A(n6627), .B(keyinput_235), .ZN(n5968) );
  XNOR2_X1 U6673 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_232), .ZN(n5967)
         );
  XNOR2_X1 U6674 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_236), .ZN(n5966)
         );
  XNOR2_X1 U6675 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_234), .ZN(n5965)
         );
  NAND4_X1 U6676 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n5969)
         );
  NOR4_X1 U6677 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n5978)
         );
  INV_X1 U6678 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6630) );
  XNOR2_X1 U6679 ( .A(n6630), .B(keyinput_238), .ZN(n5977) );
  XNOR2_X1 U6680 ( .A(n6632), .B(keyinput_241), .ZN(n5975) );
  XNOR2_X1 U6681 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_240), .ZN(n5974)
         );
  XNOR2_X1 U6682 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_239), .ZN(n5973)
         );
  NOR3_X1 U6683 ( .A1(n5975), .A2(n5974), .A3(n5973), .ZN(n5976) );
  OAI21_X1 U6684 ( .B1(n5978), .B2(n5977), .A(n5976), .ZN(n5982) );
  XOR2_X1 U6685 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_242), .Z(n5981)
         );
  XNOR2_X1 U6686 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_243), .ZN(n5980)
         );
  XNOR2_X1 U6687 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_244), .ZN(n5979)
         );
  NAND4_X1 U6688 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5985)
         );
  XNOR2_X1 U6689 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_245), .ZN(n5984)
         );
  XNOR2_X1 U6690 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_246), .ZN(n5983)
         );
  NAND3_X1 U6691 ( .A1(n5985), .A2(n5984), .A3(n5983), .ZN(n5988) );
  XNOR2_X1 U6692 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_247), .ZN(n5987)
         );
  XNOR2_X1 U6693 ( .A(DATAWIDTH_REG_16__SCAN_IN), .B(keyinput_248), .ZN(n5986)
         );
  NAND3_X1 U6694 ( .A1(n5988), .A2(n5987), .A3(n5986), .ZN(n5991) );
  XNOR2_X1 U6695 ( .A(DATAWIDTH_REG_18__SCAN_IN), .B(keyinput_250), .ZN(n5990)
         );
  XNOR2_X1 U6696 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_249), .ZN(n5989)
         );
  NAND3_X1 U6697 ( .A1(n5991), .A2(n5990), .A3(n5989), .ZN(n5997) );
  XNOR2_X1 U6698 ( .A(DATAWIDTH_REG_19__SCAN_IN), .B(keyinput_251), .ZN(n5996)
         );
  XNOR2_X1 U6699 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_253), .ZN(n5994)
         );
  XNOR2_X1 U6700 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_254), .ZN(n5993)
         );
  XNOR2_X1 U6701 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_252), .ZN(n5992)
         );
  NAND3_X1 U6702 ( .A1(n5994), .A2(n5993), .A3(n5992), .ZN(n5995) );
  AOI21_X1 U6703 ( .B1(n5997), .B2(n5996), .A(n5995), .ZN(n5998) );
  AOI211_X1 U6704 ( .C1(n6001), .C2(n6000), .A(n5999), .B(n5998), .ZN(n6008)
         );
  NAND2_X1 U6705 ( .A1(n6165), .A2(n3959), .ZN(n6002) );
  AOI22_X1 U6706 ( .A1(n6004), .A2(n6003), .B1(n4904), .B2(n6002), .ZN(n6823)
         );
  AND2_X1 U6707 ( .A1(n4554), .A2(n6005), .ZN(n6161) );
  OAI21_X1 U6708 ( .B1(n6161), .B2(n6006), .A(n7250), .ZN(n6836) );
  NAND2_X1 U6709 ( .A1(n6823), .A2(n6836), .ZN(n7190) );
  NAND2_X1 U6710 ( .A1(n7190), .A2(n7221), .ZN(n6171) );
  AOI21_X1 U6711 ( .B1(n6171), .B2(FLUSH_REG_SCAN_IN), .A(n6819), .ZN(n6007)
         );
  XNOR2_X1 U6712 ( .A(n6008), .B(n6007), .ZN(U2793) );
  XOR2_X1 U6713 ( .A(n6009), .B(n6010), .Z(n6893) );
  NAND2_X1 U6714 ( .A1(n6893), .A2(n6819), .ZN(n6013) );
  NOR2_X1 U6715 ( .A1(n6924), .A2(n6681), .ZN(n6891) );
  NOR2_X1 U6716 ( .A1(n6822), .A2(n7019), .ZN(n6011) );
  AOI211_X1 U6717 ( .C1(n4711), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6891), 
        .B(n6011), .ZN(n6012) );
  OAI211_X1 U6718 ( .C1(n6745), .C2(n6791), .A(n6013), .B(n6012), .ZN(U2977)
         );
  NAND2_X1 U6719 ( .A1(n6022), .A2(n6014), .ZN(n6016) );
  XOR2_X1 U6720 ( .A(n6016), .B(n6015), .Z(n6033) );
  NAND2_X1 U6721 ( .A1(n6908), .A2(REIP_REG_10__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U6722 ( .B1(n6448), .B2(n5551), .A(n6038), .ZN(n6019) );
  NOR2_X1 U6723 ( .A1(n6017), .A2(n6791), .ZN(n6018) );
  AOI211_X1 U6724 ( .C1(n6801), .C2(n6020), .A(n6019), .B(n6018), .ZN(n6021)
         );
  OAI21_X1 U6725 ( .B1(n6033), .B2(n6804), .A(n6021), .ZN(U2976) );
  NAND2_X1 U6726 ( .A1(n6023), .A2(n6022), .ZN(n6027) );
  INV_X1 U6727 ( .A(n6067), .ZN(n6025) );
  NOR2_X1 U6728 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U6729 ( .A1(n6027), .A2(n6026), .ZN(n6068) );
  OAI21_X1 U6730 ( .B1(n6027), .B2(n6026), .A(n6068), .ZN(n6900) );
  NAND2_X1 U6731 ( .A1(n6908), .A2(REIP_REG_11__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U6732 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6028)
         );
  OAI211_X1 U6733 ( .C1(n6822), .C2(n7032), .A(n6898), .B(n6028), .ZN(n6029)
         );
  AOI21_X1 U6734 ( .B1(n7034), .B2(n6818), .A(n6029), .ZN(n6030) );
  OAI21_X1 U6735 ( .B1(n6900), .B2(n6804), .A(n6030), .ZN(U2975) );
  NAND2_X1 U6736 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U6737 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6073), .ZN(n6043) );
  NOR2_X1 U6738 ( .A1(n6032), .A2(n6031), .ZN(n6034) );
  NAND2_X1 U6739 ( .A1(n6034), .A2(n6880), .ZN(n6896) );
  OR2_X1 U6740 ( .A1(n6033), .A2(n6619), .ZN(n6042) );
  NAND2_X1 U6741 ( .A1(n6034), .A2(n6867), .ZN(n6072) );
  INV_X1 U6742 ( .A(n6589), .ZN(n6036) );
  NAND2_X1 U6743 ( .A1(n6035), .A2(n6034), .ZN(n6071) );
  AOI22_X1 U6744 ( .A1(n6870), .A2(n6072), .B1(n6036), .B2(n6071), .ZN(n6037)
         );
  NAND2_X1 U6745 ( .A1(n6037), .A2(n6587), .ZN(n6892) );
  OAI21_X1 U6746 ( .B1(n6884), .B2(n6039), .A(n6038), .ZN(n6040) );
  AOI21_X1 U6747 ( .B1(n6892), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6040), 
        .ZN(n6041) );
  OAI211_X1 U6748 ( .C1(n6043), .C2(n6896), .A(n6042), .B(n6041), .ZN(U3008)
         );
  XNOR2_X1 U6749 ( .A(n6044), .B(n6045), .ZN(n6089) );
  INV_X1 U6750 ( .A(n6085), .ZN(n6056) );
  OAI21_X1 U6751 ( .B1(n6048), .B2(n6047), .A(n6046), .ZN(n6049) );
  NAND2_X1 U6752 ( .A1(n6049), .A2(n6062), .ZN(n6847) );
  AOI21_X1 U6753 ( .B1(n7144), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7086), 
        .ZN(n6050) );
  OAI21_X1 U6754 ( .B1(n7152), .B2(n6847), .A(n6050), .ZN(n6055) );
  NAND2_X1 U6755 ( .A1(n6051), .A2(REIP_REG_10__SCAN_IN), .ZN(n7027) );
  INV_X1 U6756 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U6757 ( .A1(n7027), .A2(n7029), .ZN(n6125) );
  OAI21_X1 U6758 ( .B1(n7147), .B2(n6125), .A(n6941), .ZN(n7039) );
  AOI22_X1 U6759 ( .A1(EBX_REG_13__SCAN_IN), .A2(n7145), .B1(
        REIP_REG_13__SCAN_IN), .B2(n7039), .ZN(n6053) );
  AND2_X1 U6760 ( .A1(n7139), .A2(n6125), .ZN(n7072) );
  NAND2_X1 U6761 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n7048) );
  OAI211_X1 U6762 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n7072), .B(n7048), .ZN(n6052) );
  NAND2_X1 U6763 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  AOI211_X1 U6764 ( .C1(n7133), .C2(n6056), .A(n6055), .B(n6054), .ZN(n6057)
         );
  OAI21_X1 U6765 ( .B1(n6089), .B2(n7130), .A(n6057), .ZN(U2814) );
  OAI21_X1 U6766 ( .B1(n6058), .B2(n6060), .A(n6059), .ZN(n7053) );
  INV_X1 U6767 ( .A(n6260), .ZN(n6064) );
  NAND2_X1 U6768 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U6769 ( .A1(n6064), .A2(n6063), .ZN(n7052) );
  INV_X1 U6770 ( .A(n7052), .ZN(n6065) );
  AOI22_X1 U6771 ( .A1(n6065), .A2(n6769), .B1(EBX_REG_14__SCAN_IN), .B2(n6311), .ZN(n6066) );
  OAI21_X1 U6772 ( .B1(n7053), .B2(n6315), .A(n6066), .ZN(U2845) );
  NAND2_X1 U6773 ( .A1(n6068), .A2(n6067), .ZN(n6070) );
  XNOR2_X1 U6774 ( .A(n3633), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6069)
         );
  XNOR2_X1 U6775 ( .A(n6070), .B(n6069), .ZN(n6805) );
  AOI22_X1 U6776 ( .A1(n7038), .A2(n6917), .B1(n6908), .B2(
        REIP_REG_12__SCAN_IN), .ZN(n6079) );
  AOI21_X1 U6777 ( .B1(n6467), .B2(n6073), .A(n6892), .ZN(n6905) );
  INV_X1 U6778 ( .A(n6905), .ZN(n6077) );
  NOR2_X1 U6779 ( .A1(n6071), .A2(n6073), .ZN(n6453) );
  NAND2_X1 U6780 ( .A1(n6866), .A2(n6453), .ZN(n6593) );
  NAND2_X1 U6781 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6094) );
  INV_X1 U6782 ( .A(n6094), .ZN(n6096) );
  AOI21_X1 U6783 ( .B1(n6593), .B2(n6471), .A(n6096), .ZN(n6076) );
  NOR2_X1 U6784 ( .A1(n6073), .A2(n6072), .ZN(n6460) );
  NAND2_X1 U6785 ( .A1(n6870), .A2(n6460), .ZN(n6098) );
  NAND2_X1 U6786 ( .A1(n6593), .A2(n6098), .ZN(n6906) );
  AOI21_X1 U6787 ( .B1(n6906), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6074) );
  INV_X1 U6788 ( .A(n6074), .ZN(n6075) );
  OAI21_X1 U6789 ( .B1(n6077), .B2(n6076), .A(n6075), .ZN(n6078) );
  OAI211_X1 U6790 ( .C1(n6805), .C2(n6619), .A(n6079), .B(n6078), .ZN(U3006)
         );
  INV_X1 U6791 ( .A(DATAI_14_), .ZN(n6080) );
  OAI222_X1 U6792 ( .A1(n7053), .A2(n7335), .B1(n6343), .B2(n6080), .C1(n6142), 
        .C2(n4341), .ZN(U2877) );
  INV_X1 U6793 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7324) );
  INV_X1 U6794 ( .A(DATAI_13_), .ZN(n7319) );
  OAI222_X1 U6795 ( .A1(n6142), .A2(n7324), .B1(n7319), .B2(n6343), .C1(n7335), 
        .C2(n6089), .ZN(U2878) );
  INV_X1 U6796 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6081) );
  OAI222_X1 U6797 ( .A1(n6847), .A2(n6320), .B1(n6315), .B2(n6089), .C1(n6081), 
        .C2(n6773), .ZN(U2846) );
  XNOR2_X1 U6798 ( .A(n6082), .B(n6083), .ZN(n6851) );
  NAND2_X1 U6799 ( .A1(n6851), .A2(n6819), .ZN(n6088) );
  INV_X1 U6800 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6084) );
  NOR2_X1 U6801 ( .A1(n6924), .A2(n6084), .ZN(n6848) );
  NOR2_X1 U6802 ( .A1(n6822), .A2(n6085), .ZN(n6086) );
  AOI211_X1 U6803 ( .C1(n4711), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6848), 
        .B(n6086), .ZN(n6087) );
  OAI211_X1 U6804 ( .C1(n6089), .C2(n6791), .A(n6088), .B(n6087), .ZN(U2973)
         );
  NAND2_X1 U6805 ( .A1(n3696), .A2(n6091), .ZN(n6092) );
  XNOR2_X1 U6806 ( .A(n6090), .B(n6092), .ZN(n6452) );
  NAND2_X1 U6807 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6096), .ZN(n6454) );
  INV_X1 U6808 ( .A(n6093), .ZN(n6097) );
  NAND2_X1 U6809 ( .A1(n6471), .A2(n6097), .ZN(n6919) );
  AOI22_X1 U6810 ( .A1(n6921), .A2(n6454), .B1(n6919), .B2(n6094), .ZN(n6095)
         );
  NAND2_X1 U6811 ( .A1(n6905), .A2(n6095), .ZN(n6850) );
  NAND2_X1 U6812 ( .A1(n6096), .A2(n4634), .ZN(n6854) );
  AOI21_X1 U6813 ( .B1(n6098), .B2(n6097), .A(n6854), .ZN(n6099) );
  OR2_X1 U6814 ( .A1(n6850), .A2(n6099), .ZN(n6102) );
  INV_X1 U6815 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6689) );
  OAI22_X1 U6816 ( .A1(n7052), .A2(n6884), .B1(n6689), .B2(n6924), .ZN(n6101)
         );
  INV_X1 U6817 ( .A(n6906), .ZN(n6855) );
  NOR3_X1 U6818 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6855), .A3(n6454), 
        .ZN(n6100) );
  AOI211_X1 U6819 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6102), .A(n6101), .B(n6100), .ZN(n6103) );
  OAI21_X1 U6820 ( .B1(n6452), .B2(n6619), .A(n6103), .ZN(U3004) );
  AOI22_X1 U6821 ( .A1(n7175), .A2(n7221), .B1(FLUSH_REG_SCAN_IN), .B2(n6835), 
        .ZN(n7173) );
  NAND2_X1 U6822 ( .A1(n7173), .A2(n7213), .ZN(n7171) );
  INV_X1 U6823 ( .A(n7171), .ZN(n6158) );
  INV_X1 U6824 ( .A(n7169), .ZN(n6155) );
  AOI22_X1 U6825 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6104), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4560), .ZN(n6153) );
  NOR3_X1 U6826 ( .A1(n7164), .A2(n6151), .A3(n6153), .ZN(n6107) );
  INV_X1 U6827 ( .A(n5049), .ZN(n6105) );
  INV_X1 U6828 ( .A(n6108), .ZN(n7217) );
  NOR3_X1 U6829 ( .A1(n6105), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n7217), 
        .ZN(n6106) );
  AOI211_X1 U6830 ( .C1(n7176), .C2(n6155), .A(n6107), .B(n6106), .ZN(n6110)
         );
  OAI21_X1 U6831 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7217), .A(n7171), 
        .ZN(n7166) );
  AOI21_X1 U6832 ( .B1(n3707), .B2(n6108), .A(n7166), .ZN(n6109) );
  OAI22_X1 U6833 ( .A1(n6158), .A2(n6110), .B1(n6109), .B2(n3651), .ZN(U3459)
         );
  NAND3_X1 U6834 ( .A1(n7198), .A2(n6112), .A3(n6111), .ZN(n7223) );
  INV_X1 U6835 ( .A(n7223), .ZN(n6115) );
  OAI22_X1 U6836 ( .A1(n6647), .A2(n7417), .B1(n6113), .B2(n5092), .ZN(n6114)
         );
  AOI21_X1 U6837 ( .B1(n6115), .B2(n6647), .A(n6114), .ZN(n6116) );
  OAI21_X1 U6838 ( .B1(n6118), .B2(n6117), .A(n6116), .ZN(U3465) );
  NOR2_X1 U6839 ( .A1(n6120), .A2(n6121), .ZN(n6122) );
  NOR2_X1 U6840 ( .A1(n6123), .A2(n6122), .ZN(n6511) );
  INV_X1 U6841 ( .A(n6124), .ZN(n6134) );
  INV_X1 U6842 ( .A(n7074), .ZN(n7106) );
  INV_X1 U6843 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6712) );
  INV_X1 U6844 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6710) );
  NOR2_X1 U6845 ( .A1(n6712), .A2(n6710), .ZN(n6126) );
  INV_X1 U6846 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6702) );
  INV_X1 U6847 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6699) );
  NAND3_X1 U6848 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .ZN(n6262) );
  INV_X1 U6849 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7061) );
  INV_X1 U6850 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7059) );
  NOR3_X1 U6851 ( .A1(n6262), .A2(n7061), .A3(n7059), .ZN(n7073) );
  NAND3_X1 U6852 ( .A1(n6125), .A2(n7073), .A3(REIP_REG_17__SCAN_IN), .ZN(
        n7083) );
  NAND3_X1 U6853 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n7119) );
  NOR3_X1 U6854 ( .A1(n6699), .A2(n7083), .A3(n7119), .ZN(n7138) );
  NAND2_X1 U6855 ( .A1(REIP_REG_22__SCAN_IN), .A2(n7138), .ZN(n7146) );
  NOR3_X1 U6856 ( .A1(n7075), .A2(n6702), .A3(n7146), .ZN(n6245) );
  NAND2_X1 U6857 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6245), .ZN(n6236) );
  NAND2_X1 U6858 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6130) );
  OAI21_X1 U6859 ( .B1(n6236), .B2(n6130), .A(n7074), .ZN(n6212) );
  OAI21_X1 U6860 ( .B1(n7106), .B2(n6126), .A(n6212), .ZN(n6204) );
  INV_X1 U6861 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6138) );
  OAI22_X1 U6862 ( .A1(n7120), .A2(n6138), .B1(n6127), .B2(n7122), .ZN(n6132)
         );
  INV_X1 U6863 ( .A(n7146), .ZN(n6128) );
  AND2_X1 U6864 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6128), .ZN(n6129) );
  AND2_X1 U6865 ( .A1(n7139), .A2(n6129), .ZN(n6249) );
  NAND2_X1 U6866 ( .A1(n6249), .A2(REIP_REG_24__SCAN_IN), .ZN(n6239) );
  NOR3_X1 U6867 ( .A1(n6214), .A2(REIP_REG_28__SCAN_IN), .A3(n6710), .ZN(n6131) );
  AOI211_X1 U6868 ( .C1(REIP_REG_28__SCAN_IN), .C2(n6204), .A(n6132), .B(n6131), .ZN(n6133) );
  OAI21_X1 U6869 ( .B1(n6134), .B2(n7157), .A(n6133), .ZN(n6135) );
  AOI21_X1 U6870 ( .B1(n6511), .B2(n7125), .A(n6135), .ZN(n6136) );
  OAI21_X1 U6871 ( .B1(n6119), .B2(n7130), .A(n6136), .ZN(U2799) );
  INV_X1 U6872 ( .A(n6511), .ZN(n6137) );
  OAI222_X1 U6873 ( .A1(n6315), .A2(n6119), .B1(n6138), .B2(n6773), .C1(n6137), 
        .C2(n6320), .ZN(U2831) );
  AOI22_X1 U6874 ( .A1(n7434), .A2(DATAI_28_), .B1(n7437), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U6875 ( .A1(n7438), .A2(DATAI_12_), .ZN(n6139) );
  OAI211_X1 U6876 ( .C1(n6119), .C2(n7335), .A(n6140), .B(n6139), .ZN(U2863)
         );
  NAND2_X1 U6877 ( .A1(n6172), .A2(n6143), .ZN(n6145) );
  AOI22_X1 U6878 ( .A1(n7434), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7437), .ZN(n6144) );
  NAND2_X1 U6879 ( .A1(n6145), .A2(n6144), .ZN(U2860) );
  OAI21_X1 U6880 ( .B1(n6146), .B2(n6147), .A(n7161), .ZN(n6148) );
  OAI211_X1 U6881 ( .C1(n6150), .C2(n7160), .A(n6149), .B(n6148), .ZN(n7180)
         );
  NOR2_X1 U6882 ( .A1(n7164), .A2(n6151), .ZN(n6154) );
  NOR2_X1 U6883 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n7217), .ZN(n6152)
         );
  AOI222_X1 U6884 ( .A1(n7180), .A2(n6155), .B1(n6154), .B2(n6153), .C1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6152), .ZN(n6157) );
  INV_X1 U6885 ( .A(n7166), .ZN(n6156) );
  OAI22_X1 U6886 ( .A1(n6158), .A2(n6157), .B1(n3707), .B2(n6156), .ZN(U3460)
         );
  INV_X1 U6887 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6159) );
  NAND2_X1 U6888 ( .A1(n6160), .A2(n6159), .ZN(n6162) );
  MUX2_X1 U6889 ( .A(n6162), .B(n6161), .S(n6838), .Z(U3474) );
  AND2_X1 U6890 ( .A1(n4904), .A2(n6163), .ZN(n6169) );
  OR2_X1 U6891 ( .A1(n6165), .A2(n6164), .ZN(n6168) );
  NAND2_X1 U6892 ( .A1(n6170), .A2(n6166), .ZN(n6167) );
  OAI211_X1 U6893 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(n7193)
         );
  MUX2_X1 U6894 ( .A(n7193), .B(MORE_REG_SCAN_IN), .S(n6171), .Z(U3471) );
  INV_X1 U6895 ( .A(n6172), .ZN(n6187) );
  OAI21_X1 U6896 ( .B1(n6175), .B2(n6174), .A(n6173), .ZN(n6178) );
  OAI22_X1 U6897 ( .A1(n6176), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4763), .ZN(n6177) );
  XNOR2_X1 U6898 ( .A(n6178), .B(n6177), .ZN(n6482) );
  NOR3_X1 U6899 ( .A1(n6214), .A2(n6710), .A3(n6712), .ZN(n6189) );
  NAND3_X1 U6900 ( .A1(n6189), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U6901 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n6179) );
  AOI21_X1 U6902 ( .B1(n7139), .B2(n6179), .A(n6204), .ZN(n6193) );
  MUX2_X1 U6903 ( .A(n6180), .B(n6193), .S(REIP_REG_31__SCAN_IN), .Z(n6183) );
  NAND4_X1 U6904 ( .A1(n6181), .A2(n4570), .A3(EBX_REG_31__SCAN_IN), .A4(n7203), .ZN(n6182) );
  OAI211_X1 U6905 ( .C1(n6184), .C2(n7122), .A(n6183), .B(n6182), .ZN(n6185)
         );
  AOI21_X1 U6906 ( .B1(n6482), .B2(n7125), .A(n6185), .ZN(n6186) );
  OAI21_X1 U6907 ( .B1(n6187), .B2(n7130), .A(n6186), .ZN(U2796) );
  OAI22_X1 U6908 ( .A1(n7120), .A2(n6188), .B1(n6346), .B2(n7122), .ZN(n6191)
         );
  INV_X1 U6909 ( .A(n6189), .ZN(n6201) );
  INV_X1 U6910 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6715) );
  NOR3_X1 U6911 ( .A1(n6201), .A2(REIP_REG_30__SCAN_IN), .A3(n6715), .ZN(n6190) );
  AOI211_X1 U6912 ( .C1(n7133), .C2(n6348), .A(n6191), .B(n6190), .ZN(n6192)
         );
  OAI21_X1 U6913 ( .B1(n6193), .B2(n6716), .A(n6192), .ZN(n6194) );
  INV_X1 U6914 ( .A(n6194), .ZN(n6195) );
  INV_X1 U6915 ( .A(n6196), .ZN(n6197) );
  OAI21_X1 U6916 ( .B1(n6356), .B2(n7130), .A(n6197), .ZN(U2797) );
  NAND2_X1 U6917 ( .A1(n6198), .A2(n7155), .ZN(n6206) );
  NOR2_X1 U6918 ( .A1(n7157), .A2(n6199), .ZN(n6203) );
  AOI22_X1 U6919 ( .A1(n7145), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7144), .ZN(n6200) );
  OAI21_X1 U6920 ( .B1(n6201), .B2(REIP_REG_29__SCAN_IN), .A(n6200), .ZN(n6202) );
  AOI211_X1 U6921 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6204), .A(n6203), .B(n6202), .ZN(n6205) );
  OAI211_X1 U6922 ( .C1(n7152), .C2(n6500), .A(n6206), .B(n6205), .ZN(U2798)
         );
  INV_X1 U6923 ( .A(n6120), .ZN(n6207) );
  OAI21_X1 U6924 ( .B1(n6208), .B2(n6223), .A(n6207), .ZN(n6519) );
  AOI21_X1 U6926 ( .B1(n6211), .B2(n6210), .A(n4884), .ZN(n6364) );
  NAND2_X1 U6927 ( .A1(n6364), .A2(n7155), .ZN(n6218) );
  INV_X1 U6928 ( .A(n6212), .ZN(n6227) );
  AOI22_X1 U6929 ( .A1(n7145), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n7144), .ZN(n6213) );
  OAI21_X1 U6930 ( .B1(n6214), .B2(REIP_REG_27__SCAN_IN), .A(n6213), .ZN(n6216) );
  NOR2_X1 U6931 ( .A1(n7157), .A2(n6362), .ZN(n6215) );
  AOI211_X1 U6932 ( .C1(n6227), .C2(REIP_REG_27__SCAN_IN), .A(n6216), .B(n6215), .ZN(n6217) );
  OAI211_X1 U6933 ( .C1(n7152), .C2(n6519), .A(n6218), .B(n6217), .ZN(U2800)
         );
  OAI21_X1 U6934 ( .B1(n6219), .B2(n6220), .A(n6210), .ZN(n6368) );
  INV_X1 U6935 ( .A(n6221), .ZN(n6225) );
  INV_X1 U6936 ( .A(n6222), .ZN(n6224) );
  AOI21_X1 U6937 ( .B1(n6225), .B2(n6224), .A(n6223), .ZN(n6530) );
  INV_X1 U6938 ( .A(n6226), .ZN(n6370) );
  AOI22_X1 U6939 ( .A1(n7145), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n7144), .ZN(n6230) );
  INV_X1 U6940 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U6941 ( .A1(n6239), .A2(n6706), .ZN(n6228) );
  OAI21_X1 U6942 ( .B1(n6228), .B2(REIP_REG_26__SCAN_IN), .A(n6227), .ZN(n6229) );
  OAI211_X1 U6943 ( .C1(n7157), .C2(n6370), .A(n6230), .B(n6229), .ZN(n6231)
         );
  AOI21_X1 U6944 ( .B1(n6530), .B2(n7125), .A(n6231), .ZN(n6232) );
  OAI21_X1 U6945 ( .B1(n6368), .B2(n7130), .A(n6232), .ZN(U2801) );
  AOI21_X1 U6946 ( .B1(n6234), .B2(n6233), .A(n6219), .ZN(n6379) );
  INV_X1 U6947 ( .A(n6379), .ZN(n6334) );
  AOI21_X1 U6948 ( .B1(n6235), .B2(n6251), .A(n6222), .ZN(n6539) );
  NOR2_X1 U6949 ( .A1(n7157), .A2(n6377), .ZN(n6241) );
  AOI22_X1 U6950 ( .A1(n7145), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n7144), .ZN(n6238) );
  NAND3_X1 U6951 ( .A1(n7074), .A2(REIP_REG_25__SCAN_IN), .A3(n6236), .ZN(
        n6237) );
  OAI211_X1 U6952 ( .C1(n6239), .C2(REIP_REG_25__SCAN_IN), .A(n6238), .B(n6237), .ZN(n6240) );
  AOI211_X1 U6953 ( .C1(n6539), .C2(n7125), .A(n6241), .B(n6240), .ZN(n6242)
         );
  OAI21_X1 U6954 ( .B1(n6334), .B2(n7130), .A(n6242), .ZN(U2802) );
  OAI21_X1 U6955 ( .B1(n6243), .B2(n6244), .A(n6233), .ZN(n6388) );
  NOR2_X1 U6956 ( .A1(n7106), .A2(n6245), .ZN(n7148) );
  INV_X1 U6957 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6703) );
  OAI22_X1 U6958 ( .A1(n6247), .A2(n7122), .B1(n6246), .B2(n7120), .ZN(n6248)
         );
  AOI221_X1 U6959 ( .B1(n7148), .B2(REIP_REG_24__SCAN_IN), .C1(n6249), .C2(
        n6703), .A(n6248), .ZN(n6255) );
  AOI21_X1 U6960 ( .B1(n6252), .B2(n6276), .A(n3659), .ZN(n6547) );
  INV_X1 U6961 ( .A(n6390), .ZN(n6253) );
  AOI22_X1 U6962 ( .A1(n6547), .A2(n7125), .B1(n6253), .B2(n7133), .ZN(n6254)
         );
  OAI211_X1 U6963 ( .C1(n6388), .C2(n7130), .A(n6255), .B(n6254), .ZN(U2803)
         );
  INV_X1 U6964 ( .A(n6256), .ZN(n6257) );
  AOI21_X1 U6965 ( .B1(n6258), .B2(n6059), .A(n6257), .ZN(n6763) );
  INV_X1 U6966 ( .A(n6763), .ZN(n6345) );
  OR2_X1 U6967 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  NAND2_X1 U6968 ( .A1(n6317), .A2(n6261), .ZN(n6761) );
  OAI22_X1 U6969 ( .A1(n7120), .A2(n6765), .B1(n7152), .B2(n6761), .ZN(n6265)
         );
  INV_X1 U6970 ( .A(n7072), .ZN(n7047) );
  OR2_X1 U6971 ( .A1(n6262), .A2(n7047), .ZN(n7063) );
  AOI21_X1 U6972 ( .B1(n6262), .B2(n7074), .A(n7039), .ZN(n7060) );
  AOI21_X1 U6973 ( .B1(n7144), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7086), 
        .ZN(n6263) );
  OAI221_X1 U6974 ( .B1(REIP_REG_15__SCAN_IN), .B2(n7063), .C1(n7059), .C2(
        n7060), .A(n6263), .ZN(n6264) );
  AOI211_X1 U6975 ( .C1(n6266), .C2(n7133), .A(n6265), .B(n6264), .ZN(n6267)
         );
  OAI21_X1 U6976 ( .B1(n6345), .B2(n7130), .A(n6267), .ZN(U2812) );
  INV_X1 U6977 ( .A(n6482), .ZN(n6269) );
  INV_X1 U6978 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6268) );
  OAI22_X1 U6979 ( .A1(n6269), .A2(n6320), .B1(n6773), .B2(n6268), .ZN(U2828)
         );
  INV_X1 U6980 ( .A(n6364), .ZN(n6329) );
  INV_X1 U6981 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6270) );
  OAI222_X1 U6982 ( .A1(n6315), .A2(n6329), .B1(n6270), .B2(n6773), .C1(n6519), 
        .C2(n6320), .ZN(U2832) );
  AOI22_X1 U6983 ( .A1(n6530), .A2(n6769), .B1(EBX_REG_26__SCAN_IN), .B2(n6311), .ZN(n6271) );
  OAI21_X1 U6984 ( .B1(n6368), .B2(n6315), .A(n6271), .ZN(U2833) );
  AOI22_X1 U6985 ( .A1(n6539), .A2(n6769), .B1(EBX_REG_25__SCAN_IN), .B2(n6311), .ZN(n6272) );
  OAI21_X1 U6986 ( .B1(n6334), .B2(n6315), .A(n6272), .ZN(U2834) );
  AOI22_X1 U6987 ( .A1(n6547), .A2(n6769), .B1(EBX_REG_24__SCAN_IN), .B2(n6311), .ZN(n6273) );
  OAI21_X1 U6988 ( .B1(n6388), .B2(n6315), .A(n6273), .ZN(U2835) );
  AOI21_X1 U6989 ( .B1(n6275), .B2(n6274), .A(n6243), .ZN(n7345) );
  INV_X1 U6990 ( .A(n7345), .ZN(n6279) );
  INV_X1 U6991 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6278) );
  OAI21_X1 U6992 ( .B1(n6282), .B2(n6277), .A(n6276), .ZN(n7153) );
  OAI222_X1 U6993 ( .A1(n6279), .A2(n6315), .B1(n6278), .B2(n6773), .C1(n7153), 
        .C2(n6320), .ZN(U2836) );
  OAI21_X1 U6994 ( .B1(n6280), .B2(n6281), .A(n6274), .ZN(n7131) );
  INV_X1 U6995 ( .A(n6282), .ZN(n6285) );
  NAND2_X1 U6996 ( .A1(n6566), .A2(n6283), .ZN(n6284) );
  NAND2_X1 U6997 ( .A1(n6285), .A2(n6284), .ZN(n7129) );
  OAI22_X1 U6998 ( .A1(n7129), .A2(n6320), .B1(n6286), .B2(n6773), .ZN(n6287)
         );
  INV_X1 U6999 ( .A(n6287), .ZN(n6288) );
  OAI21_X1 U7000 ( .B1(n7131), .B2(n6315), .A(n6288), .ZN(U2837) );
  NAND2_X1 U7001 ( .A1(n6758), .A2(n6289), .ZN(n6290) );
  AND2_X1 U7002 ( .A1(n6568), .A2(n6290), .ZN(n6582) );
  INV_X1 U7003 ( .A(n6582), .ZN(n7111) );
  INV_X1 U7004 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6296) );
  BUF_X1 U7005 ( .A(n6291), .Z(n6292) );
  NAND2_X1 U7006 ( .A1(n6293), .A2(n6294), .ZN(n6295) );
  NAND2_X1 U7007 ( .A1(n6292), .A2(n6295), .ZN(n7112) );
  OAI222_X1 U7008 ( .A1(n7111), .A2(n6320), .B1(n6773), .B2(n6296), .C1(n7112), 
        .C2(n6315), .ZN(U2839) );
  OAI21_X1 U7009 ( .B1(n6297), .B2(n6299), .A(n6298), .ZN(n7088) );
  NOR2_X1 U7010 ( .A1(n6310), .A2(n6300), .ZN(n6301) );
  OR2_X1 U7011 ( .A1(n6756), .A2(n6301), .ZN(n7087) );
  OAI22_X1 U7012 ( .A1(n7087), .A2(n6320), .B1(n7093), .B2(n6773), .ZN(n6302)
         );
  INV_X1 U7013 ( .A(n6302), .ZN(n6303) );
  OAI21_X1 U7014 ( .B1(n7088), .B2(n6315), .A(n6303), .ZN(U2841) );
  AND2_X1 U7015 ( .A1(n6305), .A2(n6306), .ZN(n6307) );
  OR2_X1 U7016 ( .A1(n6297), .A2(n6307), .ZN(n6813) );
  AND2_X1 U7017 ( .A1(n6319), .A2(n6308), .ZN(n6309) );
  NOR2_X1 U7018 ( .A1(n6310), .A2(n6309), .ZN(n7079) );
  AOI22_X1 U7019 ( .A1(n7079), .A2(n6769), .B1(EBX_REG_17__SCAN_IN), .B2(n6311), .ZN(n6312) );
  OAI21_X1 U7020 ( .B1(n6813), .B2(n6315), .A(n6312), .ZN(U2842) );
  NAND2_X1 U7021 ( .A1(n6256), .A2(n6313), .ZN(n6314) );
  AND2_X1 U7022 ( .A1(n6305), .A2(n6314), .ZN(n6437) );
  INV_X1 U7023 ( .A(n6315), .ZN(n6770) );
  NAND2_X1 U7024 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  NAND2_X1 U7025 ( .A1(n6319), .A2(n6318), .ZN(n7065) );
  OAI22_X1 U7026 ( .A1(n7065), .A2(n6320), .B1(n7071), .B2(n6773), .ZN(n6321)
         );
  AOI21_X1 U7027 ( .B1(n6437), .B2(n6770), .A(n6321), .ZN(n6322) );
  INV_X1 U7028 ( .A(n6322), .ZN(U2843) );
  AOI22_X1 U7029 ( .A1(n7434), .A2(DATAI_30_), .B1(n7437), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7030 ( .A1(n7438), .A2(DATAI_14_), .ZN(n6323) );
  OAI211_X1 U7031 ( .C1(n6356), .C2(n7335), .A(n6324), .B(n6323), .ZN(U2861)
         );
  AOI22_X1 U7032 ( .A1(n7434), .A2(DATAI_29_), .B1(n7437), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7033 ( .A1(n7438), .A2(DATAI_13_), .ZN(n6325) );
  OAI211_X1 U7034 ( .C1(n4716), .C2(n7335), .A(n6326), .B(n6325), .ZN(U2862)
         );
  AOI22_X1 U7035 ( .A1(n7434), .A2(DATAI_27_), .B1(n7437), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7036 ( .A1(n7438), .A2(DATAI_11_), .ZN(n6327) );
  OAI211_X1 U7037 ( .C1(n6329), .C2(n7335), .A(n6328), .B(n6327), .ZN(U2864)
         );
  AOI22_X1 U7038 ( .A1(n7434), .A2(DATAI_26_), .B1(n7437), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7039 ( .A1(n7438), .A2(DATAI_10_), .ZN(n6330) );
  OAI211_X1 U7040 ( .C1(n6368), .C2(n7335), .A(n6331), .B(n6330), .ZN(U2865)
         );
  AOI22_X1 U7041 ( .A1(n7434), .A2(DATAI_25_), .B1(n7437), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7042 ( .A1(n7438), .A2(DATAI_9_), .ZN(n6332) );
  OAI211_X1 U7043 ( .C1(n6334), .C2(n7335), .A(n6333), .B(n6332), .ZN(U2866)
         );
  AOI22_X1 U7044 ( .A1(n7434), .A2(DATAI_22_), .B1(n7437), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7045 ( .A1(n7438), .A2(DATAI_6_), .ZN(n6335) );
  OAI211_X1 U7046 ( .C1(n7131), .C2(n7335), .A(n6336), .B(n6335), .ZN(U2869)
         );
  AOI22_X1 U7047 ( .A1(n7434), .A2(DATAI_20_), .B1(n7437), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7048 ( .A1(n7438), .A2(DATAI_4_), .ZN(n6337) );
  OAI211_X1 U7049 ( .C1(n7112), .C2(n7335), .A(n6338), .B(n6337), .ZN(U2871)
         );
  AOI22_X1 U7050 ( .A1(n7434), .A2(DATAI_18_), .B1(n7437), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7051 ( .A1(n7438), .A2(DATAI_2_), .ZN(n6339) );
  OAI211_X1 U7052 ( .C1(n7088), .C2(n7335), .A(n6340), .B(n6339), .ZN(U2873)
         );
  INV_X1 U7053 ( .A(n6437), .ZN(n7066) );
  AOI22_X1 U7054 ( .A1(n7434), .A2(DATAI_16_), .B1(n7437), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7055 ( .A1(n7438), .A2(DATAI_0_), .ZN(n6341) );
  OAI211_X1 U7056 ( .C1(n7066), .C2(n7335), .A(n6342), .B(n6341), .ZN(U2875)
         );
  INV_X1 U7057 ( .A(DATAI_15_), .ZN(n6344) );
  INV_X1 U7058 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7334) );
  OAI222_X1 U7059 ( .A1(n6345), .A2(n7335), .B1(n6344), .B2(n6343), .C1(n6142), 
        .C2(n7334), .ZN(U2876) );
  NAND2_X1 U7060 ( .A1(n6908), .A2(REIP_REG_30__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U7061 ( .B1(n6448), .B2(n6346), .A(n6487), .ZN(n6347) );
  AOI21_X1 U7062 ( .B1(n6348), .B2(n6801), .A(n6347), .ZN(n6355) );
  NAND2_X1 U7063 ( .A1(n6349), .A2(n6426), .ZN(n6352) );
  NAND2_X1 U7064 ( .A1(n6350), .A2(n3633), .ZN(n6351) );
  NAND2_X1 U7065 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  NAND2_X1 U7066 ( .A1(n6486), .A2(n6819), .ZN(n6354) );
  OAI211_X1 U7067 ( .C1(n6356), .C2(n6791), .A(n6355), .B(n6354), .ZN(U2956)
         );
  XNOR2_X1 U7068 ( .A(n6360), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6523)
         );
  AND2_X1 U7069 ( .A1(n6908), .A2(REIP_REG_27__SCAN_IN), .ZN(n6517) );
  AOI21_X1 U7070 ( .B1(n4711), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6517), 
        .ZN(n6361) );
  OAI21_X1 U7071 ( .B1(n6822), .B2(n6362), .A(n6361), .ZN(n6363) );
  AOI21_X1 U7072 ( .B1(n6364), .B2(n6818), .A(n6363), .ZN(n6365) );
  OAI21_X1 U7073 ( .B1(n6804), .B2(n6523), .A(n6365), .ZN(U2959) );
  XNOR2_X1 U7074 ( .A(n3633), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6367)
         );
  XNOR2_X1 U7075 ( .A(n6366), .B(n6367), .ZN(n6533) );
  INV_X1 U7076 ( .A(n6368), .ZN(n6372) );
  AND2_X1 U7077 ( .A1(n6908), .A2(REIP_REG_26__SCAN_IN), .ZN(n6528) );
  AOI21_X1 U7078 ( .B1(n4711), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6528), 
        .ZN(n6369) );
  OAI21_X1 U7079 ( .B1(n6822), .B2(n6370), .A(n6369), .ZN(n6371) );
  AOI21_X1 U7080 ( .B1(n6372), .B2(n6818), .A(n6371), .ZN(n6373) );
  OAI21_X1 U7081 ( .B1(n6533), .B2(n6804), .A(n6373), .ZN(U2960) );
  XNOR2_X1 U7082 ( .A(n6374), .B(n6375), .ZN(n6541) );
  AND2_X1 U7083 ( .A1(n6908), .A2(REIP_REG_25__SCAN_IN), .ZN(n6534) );
  AOI21_X1 U7084 ( .B1(n4711), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6534), 
        .ZN(n6376) );
  OAI21_X1 U7085 ( .B1(n6822), .B2(n6377), .A(n6376), .ZN(n6378) );
  AOI21_X1 U7086 ( .B1(n6379), .B2(n6818), .A(n6378), .ZN(n6380) );
  OAI21_X1 U7087 ( .B1(n6804), .B2(n6541), .A(n6380), .ZN(U2961) );
  XNOR2_X1 U7088 ( .A(n3633), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6817)
         );
  INV_X1 U7089 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U7090 ( .A1(n3633), .A2(n6419), .ZN(n6383) );
  INV_X1 U7091 ( .A(n6578), .ZN(n6463) );
  NAND2_X1 U7092 ( .A1(n3633), .A2(n6463), .ZN(n6382) );
  INV_X1 U7093 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6575) );
  XNOR2_X1 U7094 ( .A(n3633), .B(n6575), .ZN(n6410) );
  NAND3_X1 U7095 ( .A1(n3633), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6386) );
  INV_X1 U7096 ( .A(n6816), .ZN(n6385) );
  NAND4_X1 U7097 ( .A1(n6385), .A2(n6426), .A3(n6384), .A4(n6419), .ZN(n6396)
         );
  XNOR2_X1 U7098 ( .A(n6387), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6549)
         );
  INV_X1 U7099 ( .A(n6388), .ZN(n7436) );
  NAND2_X1 U7100 ( .A1(n6908), .A2(REIP_REG_24__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7101 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6389)
         );
  OAI211_X1 U7102 ( .C1(n6822), .C2(n6390), .A(n6543), .B(n6389), .ZN(n6391)
         );
  AOI21_X1 U7103 ( .B1(n7436), .B2(n6818), .A(n6391), .ZN(n6392) );
  OAI21_X1 U7104 ( .B1(n6549), .B2(n6804), .A(n6392), .ZN(U2962) );
  OR3_X1 U7105 ( .A1(n6394), .A2(n6426), .A3(n6393), .ZN(n6395) );
  NAND2_X1 U7106 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  XNOR2_X1 U7107 ( .A(n6397), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6556)
         );
  NAND2_X1 U7108 ( .A1(n6908), .A2(REIP_REG_23__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7109 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6398)
         );
  OAI211_X1 U7110 ( .C1(n6822), .C2(n7158), .A(n6550), .B(n6398), .ZN(n6399)
         );
  AOI21_X1 U7111 ( .B1(n7345), .B2(n6818), .A(n6399), .ZN(n6400) );
  OAI21_X1 U7112 ( .B1(n6556), .B2(n6804), .A(n6400), .ZN(U2963) );
  XNOR2_X1 U7113 ( .A(n3633), .B(n6401), .ZN(n6402) );
  XNOR2_X1 U7114 ( .A(n6403), .B(n6402), .ZN(n6563) );
  NAND2_X1 U7115 ( .A1(n6908), .A2(REIP_REG_22__SCAN_IN), .ZN(n6557) );
  OAI21_X1 U7116 ( .B1(n6448), .B2(n6404), .A(n6557), .ZN(n6406) );
  NOR2_X1 U7117 ( .A1(n7131), .A2(n6791), .ZN(n6405) );
  AOI211_X1 U7118 ( .C1(n6801), .C2(n7134), .A(n6406), .B(n6405), .ZN(n6407)
         );
  OAI21_X1 U7119 ( .B1(n6563), .B2(n6804), .A(n6407), .ZN(U2964) );
  AOI21_X1 U7120 ( .B1(n6408), .B2(n6292), .A(n6280), .ZN(n7342) );
  INV_X1 U7121 ( .A(n7342), .ZN(n6417) );
  INV_X1 U7122 ( .A(n6409), .ZN(n6565) );
  NAND2_X1 U7123 ( .A1(n6411), .A2(n6410), .ZN(n6564) );
  NAND3_X1 U7124 ( .A1(n6565), .A2(n6819), .A3(n6564), .ZN(n6416) );
  INV_X1 U7125 ( .A(n7128), .ZN(n6414) );
  NAND2_X1 U7126 ( .A1(n6908), .A2(REIP_REG_21__SCAN_IN), .ZN(n6570) );
  OAI21_X1 U7127 ( .B1(n6448), .B2(n6412), .A(n6570), .ZN(n6413) );
  AOI21_X1 U7128 ( .B1(n6801), .B2(n6414), .A(n6413), .ZN(n6415) );
  OAI211_X1 U7129 ( .C1(n6791), .C2(n6417), .A(n6416), .B(n6415), .ZN(U2965)
         );
  NAND2_X1 U7130 ( .A1(n3633), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6418) );
  MUX2_X1 U7131 ( .A(n3633), .B(n6418), .S(n6816), .Z(n6420) );
  XNOR2_X1 U7132 ( .A(n6420), .B(n6419), .ZN(n6585) );
  NAND2_X1 U7133 ( .A1(n6908), .A2(REIP_REG_20__SCAN_IN), .ZN(n6577) );
  OAI21_X1 U7134 ( .B1(n6448), .B2(n7117), .A(n6577), .ZN(n6422) );
  NOR2_X1 U7135 ( .A1(n7112), .A2(n6791), .ZN(n6421) );
  AOI211_X1 U7136 ( .C1(n6801), .C2(n7114), .A(n6422), .B(n6421), .ZN(n6423)
         );
  OAI21_X1 U7137 ( .B1(n6585), .B2(n6804), .A(n6423), .ZN(U2966) );
  NAND2_X1 U7138 ( .A1(n3633), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6809) );
  INV_X1 U7139 ( .A(n6424), .ZN(n6425) );
  AOI21_X1 U7140 ( .B1(n6426), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6425), 
        .ZN(n6808) );
  NOR2_X1 U7141 ( .A1(n3633), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6806)
         );
  NAND2_X1 U7142 ( .A1(n6808), .A2(n6806), .ZN(n6811) );
  OAI21_X1 U7143 ( .B1(n6424), .B2(n6809), .A(n6811), .ZN(n6427) );
  XNOR2_X1 U7144 ( .A(n6427), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6602)
         );
  NAND2_X1 U7145 ( .A1(n6908), .A2(REIP_REG_18__SCAN_IN), .ZN(n6598) );
  OAI21_X1 U7146 ( .B1(n6448), .B2(n3701), .A(n6598), .ZN(n6429) );
  NOR2_X1 U7147 ( .A1(n7088), .A2(n6791), .ZN(n6428) );
  AOI211_X1 U7148 ( .C1(n6801), .C2(n7090), .A(n6429), .B(n6428), .ZN(n6430)
         );
  OAI21_X1 U7149 ( .B1(n6602), .B2(n6804), .A(n6430), .ZN(U2968) );
  XNOR2_X1 U7150 ( .A(n3633), .B(n6606), .ZN(n6432) );
  XNOR2_X1 U7151 ( .A(n6433), .B(n6432), .ZN(n6610) );
  NAND2_X1 U7152 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6434)
         );
  NAND2_X1 U7153 ( .A1(n6908), .A2(REIP_REG_16__SCAN_IN), .ZN(n6604) );
  OAI211_X1 U7154 ( .C1(n6822), .C2(n6435), .A(n6434), .B(n6604), .ZN(n6436)
         );
  AOI21_X1 U7155 ( .B1(n6437), .B2(n6818), .A(n6436), .ZN(n6438) );
  OAI21_X1 U7156 ( .B1(n6610), .B2(n6804), .A(n6438), .ZN(U2970) );
  INV_X1 U7157 ( .A(n6440), .ZN(n6441) );
  NOR2_X1 U7158 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  XNOR2_X1 U7159 ( .A(n6439), .B(n6443), .ZN(n6620) );
  NAND2_X1 U7160 ( .A1(n6908), .A2(REIP_REG_15__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U7161 ( .A1(n4711), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6444)
         );
  OAI211_X1 U7162 ( .C1(n6822), .C2(n6445), .A(n6614), .B(n6444), .ZN(n6446)
         );
  AOI21_X1 U7163 ( .B1(n6763), .B2(n6818), .A(n6446), .ZN(n6447) );
  OAI21_X1 U7164 ( .B1(n6620), .B2(n6804), .A(n6447), .ZN(U2971) );
  OAI22_X1 U7165 ( .A1(n6448), .A2(n4338), .B1(n6924), .B2(n6689), .ZN(n6450)
         );
  NOR2_X1 U7166 ( .A1(n7053), .A2(n6791), .ZN(n6449) );
  AOI211_X1 U7167 ( .C1(n6801), .C2(n7055), .A(n6450), .B(n6449), .ZN(n6451)
         );
  OAI21_X1 U7168 ( .B1(n6804), .B2(n6452), .A(n6451), .ZN(U2972) );
  INV_X1 U7169 ( .A(n6506), .ZN(n6496) );
  AND2_X1 U7170 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U7171 ( .A1(n6473), .A2(n6471), .ZN(n6466) );
  INV_X1 U7172 ( .A(n6453), .ZN(n6456) );
  INV_X1 U7173 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6455) );
  NOR2_X1 U7174 ( .A1(n6455), .A2(n6454), .ZN(n6605) );
  NAND3_X1 U7175 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6605), .ZN(n6586) );
  NOR2_X1 U7176 ( .A1(n6456), .A2(n6586), .ZN(n6588) );
  INV_X1 U7177 ( .A(n6457), .ZN(n6458) );
  AND2_X1 U7178 ( .A1(n6588), .A2(n6458), .ZN(n6469) );
  OR2_X1 U7179 ( .A1(n6589), .A2(n6469), .ZN(n6459) );
  AND2_X1 U7180 ( .A1(n6459), .A2(n6587), .ZN(n6462) );
  INV_X1 U7181 ( .A(n6462), .ZN(n6465) );
  NOR2_X1 U7182 ( .A1(n6912), .A2(n6586), .ZN(n6594) );
  NAND2_X1 U7183 ( .A1(n6594), .A2(n6460), .ZN(n6591) );
  OR2_X1 U7184 ( .A1(n6596), .A2(n6591), .ZN(n6470) );
  NAND2_X1 U7185 ( .A1(n6870), .A2(n6470), .ZN(n6461) );
  NAND2_X1 U7186 ( .A1(n6462), .A2(n6461), .ZN(n6842) );
  OR2_X1 U7187 ( .A1(n6842), .A2(n6463), .ZN(n6464) );
  OAI21_X1 U7188 ( .B1(n6465), .B2(n6467), .A(n6464), .ZN(n6576) );
  OAI21_X1 U7189 ( .B1(n6475), .B2(n6603), .A(n6576), .ZN(n6554) );
  AOI21_X1 U7190 ( .B1(n6477), .B2(n6466), .A(n6554), .ZN(n6545) );
  OAI21_X1 U7191 ( .B1(n6603), .B2(n6525), .A(n6545), .ZN(n6518) );
  AOI21_X1 U7192 ( .B1(n6496), .B2(n6467), .A(n6518), .ZN(n6495) );
  OAI21_X1 U7193 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6603), .A(n6495), 
        .ZN(n6491) );
  INV_X1 U7194 ( .A(n6491), .ZN(n6468) );
  OAI21_X1 U7195 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6603), .A(n6468), 
        .ZN(n6481) );
  INV_X1 U7196 ( .A(n6469), .ZN(n6472) );
  OAI22_X1 U7197 ( .A1(n6473), .A2(n6472), .B1(n6471), .B2(n6470), .ZN(n6474)
         );
  NAND2_X1 U7198 ( .A1(n6474), .A2(n6578), .ZN(n6571) );
  INV_X1 U7199 ( .A(n6475), .ZN(n6476) );
  NOR2_X1 U7200 ( .A1(n6551), .A2(n6477), .ZN(n6535) );
  NAND2_X1 U7201 ( .A1(n6535), .A2(n6525), .ZN(n6515) );
  INV_X1 U7202 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6478) );
  NOR4_X1 U7203 ( .A1(n6515), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6488), 
        .A4(n6478), .ZN(n6479) );
  AOI211_X1 U7204 ( .C1(n6481), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n6480), .B(n6479), .ZN(n6484) );
  NAND2_X1 U7205 ( .A1(n6482), .A2(n6917), .ZN(n6483) );
  OAI211_X1 U7206 ( .C1(n6485), .C2(n6619), .A(n6484), .B(n6483), .ZN(U2987)
         );
  NAND2_X1 U7207 ( .A1(n6486), .A2(n6915), .ZN(n6493) );
  INV_X1 U7208 ( .A(n6487), .ZN(n6490) );
  NOR3_X1 U7209 ( .A1(n6515), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n6488), 
        .ZN(n6489) );
  AOI211_X1 U7210 ( .C1(n6491), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6490), .B(n6489), .ZN(n6492) );
  OAI211_X1 U7211 ( .C1(n6494), .C2(n6884), .A(n6493), .B(n6492), .ZN(U2988)
         );
  INV_X1 U7212 ( .A(n6495), .ZN(n6499) );
  NOR3_X1 U7213 ( .A1(n6515), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n6496), 
        .ZN(n6497) );
  AOI211_X1 U7214 ( .C1(n6499), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n6498), .B(n6497), .ZN(n6503) );
  INV_X1 U7215 ( .A(n6500), .ZN(n6501) );
  NAND2_X1 U7216 ( .A1(n6501), .A2(n6917), .ZN(n6502) );
  OAI211_X1 U7217 ( .C1(n6504), .C2(n6619), .A(n6503), .B(n6502), .ZN(U2989)
         );
  INV_X1 U7218 ( .A(n6505), .ZN(n6510) );
  AOI211_X1 U7219 ( .C1(n6508), .C2(n6507), .A(n6506), .B(n6515), .ZN(n6509)
         );
  AOI211_X1 U7220 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n6518), .A(n6510), .B(n6509), .ZN(n6513) );
  NAND2_X1 U7221 ( .A1(n6511), .A2(n6917), .ZN(n6512) );
  OAI211_X1 U7222 ( .C1(n6514), .C2(n6619), .A(n6513), .B(n6512), .ZN(U2990)
         );
  NOR2_X1 U7223 ( .A1(n6515), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6516)
         );
  AOI211_X1 U7224 ( .C1(n6518), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6517), .B(n6516), .ZN(n6522) );
  INV_X1 U7225 ( .A(n6519), .ZN(n6520) );
  NAND2_X1 U7226 ( .A1(n6520), .A2(n6917), .ZN(n6521) );
  OAI211_X1 U7227 ( .C1(n6523), .C2(n6619), .A(n6522), .B(n6521), .ZN(U2991)
         );
  INV_X1 U7228 ( .A(n6545), .ZN(n6529) );
  INV_X1 U7229 ( .A(n6535), .ZN(n6524) );
  AOI211_X1 U7230 ( .C1(n6537), .C2(n6526), .A(n6525), .B(n6524), .ZN(n6527)
         );
  AOI211_X1 U7231 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n6529), .A(n6528), .B(n6527), .ZN(n6532) );
  NAND2_X1 U7232 ( .A1(n6530), .A2(n6917), .ZN(n6531) );
  OAI211_X1 U7233 ( .C1(n6533), .C2(n6619), .A(n6532), .B(n6531), .ZN(U2992)
         );
  AOI21_X1 U7234 ( .B1(n6535), .B2(n6537), .A(n6534), .ZN(n6536) );
  OAI21_X1 U7235 ( .B1(n6545), .B2(n6537), .A(n6536), .ZN(n6538) );
  AOI21_X1 U7236 ( .B1(n6539), .B2(n6917), .A(n6538), .ZN(n6540) );
  OAI21_X1 U7237 ( .B1(n6541), .B2(n6619), .A(n6540), .ZN(U2993) );
  INV_X1 U7238 ( .A(n6551), .ZN(n6542) );
  AOI21_X1 U7239 ( .B1(n6542), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6544) );
  OAI21_X1 U7240 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6546) );
  AOI21_X1 U7241 ( .B1(n6547), .B2(n6917), .A(n6546), .ZN(n6548) );
  OAI21_X1 U7242 ( .B1(n6549), .B2(n6619), .A(n6548), .ZN(U2994) );
  OAI21_X1 U7243 ( .B1(n6551), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6550), 
        .ZN(n6553) );
  NOR2_X1 U7244 ( .A1(n7153), .A2(n6884), .ZN(n6552) );
  AOI211_X1 U7245 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n6554), .A(n6553), .B(n6552), .ZN(n6555) );
  OAI21_X1 U7246 ( .B1(n6556), .B2(n6619), .A(n6555), .ZN(U2995) );
  INV_X1 U7247 ( .A(n6576), .ZN(n6561) );
  XNOR2_X1 U7248 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U7249 ( .B1(n6571), .B2(n6558), .A(n6557), .ZN(n6560) );
  NOR2_X1 U7250 ( .A1(n7129), .A2(n6884), .ZN(n6559) );
  AOI211_X1 U7251 ( .C1(n6561), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n6560), .B(n6559), .ZN(n6562) );
  OAI21_X1 U7252 ( .B1(n6563), .B2(n6619), .A(n6562), .ZN(U2996) );
  NAND3_X1 U7253 ( .A1(n6565), .A2(n6915), .A3(n6564), .ZN(n6574) );
  INV_X1 U7254 ( .A(n6566), .ZN(n6567) );
  AOI21_X1 U7255 ( .B1(n6569), .B2(n6568), .A(n6567), .ZN(n7124) );
  OAI21_X1 U7256 ( .B1(n6571), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6570), 
        .ZN(n6572) );
  AOI21_X1 U7257 ( .B1(n7124), .B2(n6917), .A(n6572), .ZN(n6573) );
  OAI211_X1 U7258 ( .C1(n6576), .C2(n6575), .A(n6574), .B(n6573), .ZN(U2997)
         );
  INV_X1 U7259 ( .A(n6577), .ZN(n6581) );
  NAND3_X1 U7260 ( .A1(n6594), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6906), .ZN(n6846) );
  NOR3_X1 U7261 ( .A1(n6846), .A2(n6579), .A3(n6578), .ZN(n6580) );
  AOI211_X1 U7262 ( .C1(n6842), .C2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6581), .B(n6580), .ZN(n6584) );
  NAND2_X1 U7263 ( .A1(n6582), .A2(n6917), .ZN(n6583) );
  OAI211_X1 U7264 ( .C1(n6585), .C2(n6619), .A(n6584), .B(n6583), .ZN(U2998)
         );
  NOR2_X1 U7265 ( .A1(n6586), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6907)
         );
  INV_X1 U7266 ( .A(n6907), .ZN(n6592) );
  OAI21_X1 U7267 ( .B1(n6589), .B2(n6588), .A(n6587), .ZN(n6590) );
  AOI21_X1 U7268 ( .B1(n6870), .B2(n6591), .A(n6590), .ZN(n6913) );
  OAI21_X1 U7269 ( .B1(n6593), .B2(n6592), .A(n6913), .ZN(n6600) );
  AND2_X1 U7270 ( .A1(n6906), .A2(n6594), .ZN(n6595) );
  NAND2_X1 U7271 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  OAI211_X1 U7272 ( .C1(n7087), .C2(n6884), .A(n6598), .B(n6597), .ZN(n6599)
         );
  AOI21_X1 U7273 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6600), .A(n6599), 
        .ZN(n6601) );
  OAI21_X1 U7274 ( .B1(n6602), .B2(n6619), .A(n6601), .ZN(U3000) );
  OAI21_X1 U7275 ( .B1(n6603), .B2(n6605), .A(n6905), .ZN(n6617) );
  OAI21_X1 U7276 ( .B1(n7065), .B2(n6884), .A(n6604), .ZN(n6608) );
  NAND2_X1 U7277 ( .A1(n6605), .A2(n6906), .ZN(n6611) );
  AOI221_X1 U7278 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n6606), .C2(n6612), .A(n6611), 
        .ZN(n6607) );
  AOI211_X1 U7279 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n6617), .A(n6608), .B(n6607), .ZN(n6609) );
  OAI21_X1 U7280 ( .B1(n6610), .B2(n6619), .A(n6609), .ZN(U3002) );
  INV_X1 U7281 ( .A(n6611), .ZN(n6613) );
  NAND2_X1 U7282 ( .A1(n6613), .A2(n6612), .ZN(n6615) );
  OAI211_X1 U7283 ( .C1(n6884), .C2(n6761), .A(n6615), .B(n6614), .ZN(n6616)
         );
  AOI21_X1 U7284 ( .B1(n6617), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6616), 
        .ZN(n6618) );
  OAI21_X1 U7285 ( .B1(n6620), .B2(n6619), .A(n6618), .ZN(U3003) );
  INV_X1 U7286 ( .A(n7174), .ZN(n6622) );
  OAI22_X1 U7287 ( .A1(n6622), .A2(n7169), .B1(n6621), .B2(n7217), .ZN(n6623)
         );
  MUX2_X1 U7288 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6623), .S(n7171), 
        .Z(U3456) );
  INV_X1 U7289 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6625) );
  INV_X1 U7290 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6830) );
  AOI21_X1 U7291 ( .B1(n6830), .B2(STATE_REG_1__SCAN_IN), .A(n7240), .ZN(n6651) );
  INV_X1 U7292 ( .A(n7229), .ZN(n6646) );
  NAND2_X1 U7293 ( .A1(n6830), .A2(n7240), .ZN(n6827) );
  AOI21_X1 U7294 ( .B1(n6624), .B2(n6827), .A(n6646), .ZN(n7226) );
  AOI21_X1 U7295 ( .B1(n6625), .B2(n6646), .A(n7226), .ZN(U3451) );
  NOR2_X1 U7296 ( .A1(n7229), .A2(n6626), .ZN(U3180) );
  NOR2_X1 U7297 ( .A1(n7229), .A2(n6627), .ZN(U3179) );
  INV_X1 U7298 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U7299 ( .A1(n7229), .A2(n6628), .ZN(U3178) );
  INV_X1 U7300 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U7301 ( .A1(n7229), .A2(n6629), .ZN(U3177) );
  NOR2_X1 U7302 ( .A1(n7229), .A2(n6630), .ZN(U3176) );
  INV_X1 U7303 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6631) );
  NOR2_X1 U7304 ( .A1(n7229), .A2(n6631), .ZN(U3175) );
  AND2_X1 U7305 ( .A1(n6646), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  NOR2_X1 U7306 ( .A1(n7229), .A2(n6632), .ZN(U3173) );
  AND2_X1 U7307 ( .A1(n6646), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  NOR2_X1 U7308 ( .A1(n7229), .A2(n6633), .ZN(U3171) );
  INV_X1 U7309 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6634) );
  NOR2_X1 U7310 ( .A1(n7229), .A2(n6634), .ZN(U3170) );
  INV_X1 U7311 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U7312 ( .A1(n7229), .A2(n6635), .ZN(U3169) );
  INV_X1 U7313 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U7314 ( .A1(n7229), .A2(n6636), .ZN(U3168) );
  INV_X1 U7315 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U7316 ( .A1(n7229), .A2(n6637), .ZN(U3167) );
  NOR2_X1 U7317 ( .A1(n7229), .A2(n6638), .ZN(U3166) );
  NOR2_X1 U7318 ( .A1(n7229), .A2(n6639), .ZN(U3165) );
  NOR2_X1 U7319 ( .A1(n7229), .A2(n6640), .ZN(U3164) );
  INV_X1 U7320 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6641) );
  NOR2_X1 U7321 ( .A1(n7229), .A2(n6641), .ZN(U3163) );
  INV_X1 U7322 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U7323 ( .A1(n7229), .A2(n6642), .ZN(U3162) );
  NOR2_X1 U7324 ( .A1(n7229), .A2(n6643), .ZN(U3161) );
  INV_X1 U7325 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6644) );
  NOR2_X1 U7326 ( .A1(n7229), .A2(n6644), .ZN(U3160) );
  NOR2_X1 U7327 ( .A1(n7229), .A2(n6645), .ZN(U3159) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6646), .ZN(U3158) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6646), .ZN(U3157) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6646), .ZN(U3156) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6646), .ZN(U3155) );
  AND2_X1 U7332 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6646), .ZN(U3154) );
  AND2_X1 U7333 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6646), .ZN(U3153) );
  AND2_X1 U7334 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6646), .ZN(U3152) );
  AND2_X1 U7335 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6646), .ZN(U3151) );
  INV_X1 U7336 ( .A(n6647), .ZN(n6648) );
  AND2_X1 U7337 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6648), .ZN(U3019)
         );
  AND2_X1 U7338 ( .A1(n6649), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7339 ( .B1(n6651), .B2(n6650), .A(n6829), .ZN(U2789) );
  AOI22_X1 U7340 ( .A1(n6668), .A2(LWORD_REG_0__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6653) );
  OAI21_X1 U7341 ( .B1(n7256), .B2(n6670), .A(n6653), .ZN(U2923) );
  AOI22_X1 U7342 ( .A1(n6668), .A2(LWORD_REG_1__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U7343 ( .B1(n7261), .B2(n6670), .A(n6654), .ZN(U2922) );
  AOI22_X1 U7344 ( .A1(n6668), .A2(LWORD_REG_2__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U7345 ( .B1(n7266), .B2(n6670), .A(n6655), .ZN(U2921) );
  AOI22_X1 U7346 ( .A1(n6668), .A2(LWORD_REG_3__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6656) );
  OAI21_X1 U7347 ( .B1(n7271), .B2(n6670), .A(n6656), .ZN(U2920) );
  AOI22_X1 U7348 ( .A1(n6668), .A2(LWORD_REG_4__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6657) );
  OAI21_X1 U7349 ( .B1(n7277), .B2(n6670), .A(n6657), .ZN(U2919) );
  AOI22_X1 U7350 ( .A1(n6668), .A2(LWORD_REG_5__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U7351 ( .B1(n4202), .B2(n6670), .A(n6658), .ZN(U2918) );
  AOI22_X1 U7352 ( .A1(n6668), .A2(LWORD_REG_6__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6659) );
  OAI21_X1 U7353 ( .B1(n4230), .B2(n6670), .A(n6659), .ZN(U2917) );
  AOI22_X1 U7354 ( .A1(n6668), .A2(LWORD_REG_7__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U7355 ( .B1(n7290), .B2(n6670), .A(n6660), .ZN(U2916) );
  AOI22_X1 U7356 ( .A1(n6668), .A2(LWORD_REG_8__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U7357 ( .B1(n7295), .B2(n6670), .A(n6661), .ZN(U2915) );
  AOI22_X1 U7358 ( .A1(n6668), .A2(LWORD_REG_9__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U7359 ( .B1(n7301), .B2(n6670), .A(n6662), .ZN(U2914) );
  AOI22_X1 U7360 ( .A1(n6668), .A2(LWORD_REG_10__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6663) );
  OAI21_X1 U7361 ( .B1(n7307), .B2(n6670), .A(n6663), .ZN(U2913) );
  AOI22_X1 U7362 ( .A1(n6668), .A2(LWORD_REG_11__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U7363 ( .B1(n7313), .B2(n6670), .A(n6664), .ZN(U2912) );
  AOI22_X1 U7364 ( .A1(n6668), .A2(LWORD_REG_12__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6665) );
  OAI21_X1 U7365 ( .B1(n4304), .B2(n6670), .A(n6665), .ZN(U2911) );
  AOI22_X1 U7366 ( .A1(n6668), .A2(LWORD_REG_13__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6666) );
  OAI21_X1 U7367 ( .B1(n7324), .B2(n6670), .A(n6666), .ZN(U2910) );
  AOI22_X1 U7368 ( .A1(n6668), .A2(LWORD_REG_14__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7369 ( .B1(n4341), .B2(n6670), .A(n6667), .ZN(U2909) );
  AOI22_X1 U7370 ( .A1(n6668), .A2(LWORD_REG_15__SCAN_IN), .B1(n6649), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6669) );
  OAI21_X1 U7371 ( .B1(n7334), .B2(n6670), .A(n6669), .ZN(U2908) );
  INV_X1 U7372 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6871) );
  INV_X1 U7373 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U7374 ( .A1(n6719), .A2(n6871), .B1(n6671), .B2(n6829), .C1(n5305), 
        .C2(n6713), .ZN(U3184) );
  INV_X1 U7375 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6673) );
  INV_X1 U7376 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6672) );
  OAI222_X1 U7377 ( .A1(n6719), .A2(n6673), .B1(n6672), .B2(n6829), .C1(n6871), 
        .C2(n6713), .ZN(U3185) );
  INV_X1 U7378 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6954) );
  INV_X1 U7379 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6674) );
  OAI222_X1 U7380 ( .A1(n6719), .A2(n6954), .B1(n6674), .B2(n6829), .C1(n6673), 
        .C2(n6713), .ZN(U3186) );
  OAI222_X1 U7381 ( .A1(n6719), .A2(n5242), .B1(n6675), .B2(n6829), .C1(n6954), 
        .C2(n6713), .ZN(U3187) );
  OAI222_X1 U7382 ( .A1(n6719), .A2(n5388), .B1(n6676), .B2(n6829), .C1(n5242), 
        .C2(n6713), .ZN(U3188) );
  INV_X1 U7383 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7002) );
  INV_X1 U7384 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U7385 ( .A1(n6719), .A2(n7002), .B1(n6677), .B2(n6829), .C1(n5388), 
        .C2(n6713), .ZN(U3189) );
  INV_X1 U7386 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6679) );
  INV_X1 U7387 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U7388 ( .A1(n6719), .A2(n6679), .B1(n6678), .B2(n6829), .C1(n7002), 
        .C2(n6713), .ZN(U3190) );
  OAI222_X1 U7389 ( .A1(n6719), .A2(n6681), .B1(n6680), .B2(n6829), .C1(n6679), 
        .C2(n6713), .ZN(U3191) );
  OAI222_X1 U7390 ( .A1(n6719), .A2(n6683), .B1(n6682), .B2(n6829), .C1(n6681), 
        .C2(n6713), .ZN(U3192) );
  INV_X1 U7391 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U7392 ( .A1(n6719), .A2(n7029), .B1(n6684), .B2(n6829), .C1(n6683), 
        .C2(n6713), .ZN(U3193) );
  INV_X1 U7393 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U7394 ( .A1(n6719), .A2(n6687), .B1(n6685), .B2(n6829), .C1(n7029), 
        .C2(n6713), .ZN(U3194) );
  INV_X1 U7395 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U7396 ( .A1(n6713), .A2(n6687), .B1(n6686), .B2(n6829), .C1(n6084), 
        .C2(n6719), .ZN(U3195) );
  INV_X1 U7397 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6688) );
  OAI222_X1 U7398 ( .A1(n6719), .A2(n6689), .B1(n6688), .B2(n6829), .C1(n6084), 
        .C2(n6713), .ZN(U3196) );
  INV_X1 U7399 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U7400 ( .A1(n6719), .A2(n7059), .B1(n6690), .B2(n6829), .C1(n6689), 
        .C2(n6713), .ZN(U3197) );
  INV_X1 U7401 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6691) );
  OAI222_X1 U7402 ( .A1(n6713), .A2(n7059), .B1(n6691), .B2(n6829), .C1(n7061), 
        .C2(n6719), .ZN(U3198) );
  INV_X1 U7403 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6693) );
  INV_X1 U7404 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6692) );
  OAI222_X1 U7405 ( .A1(n6719), .A2(n6693), .B1(n6692), .B2(n6829), .C1(n7061), 
        .C2(n6713), .ZN(U3199) );
  INV_X1 U7406 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7096) );
  INV_X1 U7407 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6694) );
  OAI222_X1 U7408 ( .A1(n6719), .A2(n7096), .B1(n6694), .B2(n6829), .C1(n6693), 
        .C2(n6713), .ZN(U3200) );
  INV_X1 U7409 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7097) );
  INV_X1 U7410 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7411 ( .A1(n6719), .A2(n7097), .B1(n6695), .B2(n6829), .C1(n7096), 
        .C2(n6713), .ZN(U3201) );
  INV_X1 U7412 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6696) );
  INV_X1 U7413 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7108) );
  OAI222_X1 U7414 ( .A1(n6713), .A2(n7097), .B1(n6696), .B2(n6829), .C1(n7108), 
        .C2(n6719), .ZN(U3202) );
  OAI222_X1 U7415 ( .A1(n6713), .A2(n7108), .B1(n6697), .B2(n6829), .C1(n6699), 
        .C2(n6719), .ZN(U3203) );
  INV_X1 U7416 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7137) );
  OAI222_X1 U7417 ( .A1(n6713), .A2(n6699), .B1(n6698), .B2(n6829), .C1(n7137), 
        .C2(n6719), .ZN(U3204) );
  OAI222_X1 U7418 ( .A1(n6719), .A2(n6702), .B1(n6700), .B2(n6829), .C1(n7137), 
        .C2(n6713), .ZN(U3205) );
  OAI222_X1 U7419 ( .A1(n6713), .A2(n6702), .B1(n6701), .B2(n6829), .C1(n6703), 
        .C2(n6719), .ZN(U3206) );
  OAI222_X1 U7420 ( .A1(n6719), .A2(n6706), .B1(n6704), .B2(n6829), .C1(n6703), 
        .C2(n6713), .ZN(U3207) );
  INV_X1 U7421 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6705) );
  INV_X1 U7422 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6708) );
  OAI222_X1 U7423 ( .A1(n6713), .A2(n6706), .B1(n6705), .B2(n6829), .C1(n6708), 
        .C2(n6719), .ZN(U3208) );
  OAI222_X1 U7424 ( .A1(n6713), .A2(n6708), .B1(n6707), .B2(n6829), .C1(n6710), 
        .C2(n6719), .ZN(U3209) );
  INV_X1 U7425 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6709) );
  OAI222_X1 U7426 ( .A1(n6713), .A2(n6710), .B1(n6709), .B2(n6829), .C1(n6712), 
        .C2(n6719), .ZN(U3210) );
  INV_X1 U7427 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6711) );
  OAI222_X1 U7428 ( .A1(n6713), .A2(n6712), .B1(n6711), .B2(n6829), .C1(n6715), 
        .C2(n6719), .ZN(U3211) );
  INV_X1 U7429 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6714) );
  OAI222_X1 U7430 ( .A1(n6713), .A2(n6715), .B1(n6714), .B2(n6829), .C1(n6716), 
        .C2(n6719), .ZN(U3212) );
  INV_X1 U7431 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6717) );
  OAI222_X1 U7432 ( .A1(n6719), .A2(n6718), .B1(n6717), .B2(n6829), .C1(n6716), 
        .C2(n6713), .ZN(U3213) );
  AOI22_X1 U7433 ( .A1(n6829), .A2(n6721), .B1(n6720), .B2(n7246), .ZN(U3445)
         );
  AOI221_X1 U7434 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6732) );
  NOR4_X1 U7435 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6725) );
  NOR4_X1 U7436 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6724) );
  NOR4_X1 U7437 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6723)
         );
  NOR4_X1 U7438 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6722) );
  NAND4_X1 U7439 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6731)
         );
  NOR4_X1 U7440 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6729)
         );
  AOI211_X1 U7441 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_21__SCAN_IN), .B(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6728) );
  NOR4_X1 U7442 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6727) );
  NOR4_X1 U7443 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6726) );
  NAND4_X1 U7444 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6730)
         );
  NOR2_X1 U7445 ( .A1(n6731), .A2(n6730), .ZN(n6744) );
  MUX2_X1 U7446 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6732), .S(n6744), .Z(
        U2795) );
  INV_X1 U7447 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7448 ( .A1(n6829), .A2(n6736), .B1(n6733), .B2(n7246), .ZN(U3446)
         );
  AOI21_X1 U7449 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6734) );
  OAI221_X1 U7450 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6734), .C1(n5305), .C2(
        REIP_REG_0__SCAN_IN), .A(n6744), .ZN(n6735) );
  OAI21_X1 U7451 ( .B1(n6744), .B2(n6736), .A(n6735), .ZN(U3468) );
  INV_X1 U7452 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6740) );
  INV_X1 U7453 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6737) );
  AOI22_X1 U7454 ( .A1(n6829), .A2(n6740), .B1(n6737), .B2(n7246), .ZN(U3447)
         );
  NOR3_X1 U7455 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n6738) );
  OAI21_X1 U7456 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6738), .A(n6744), .ZN(n6739)
         );
  OAI21_X1 U7457 ( .B1(n6744), .B2(n6740), .A(n6739), .ZN(U2794) );
  INV_X1 U7458 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6743) );
  INV_X1 U7459 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6741) );
  AOI22_X1 U7460 ( .A1(n6829), .A2(n6743), .B1(n6741), .B2(n7246), .ZN(U3448)
         );
  OAI21_X1 U7461 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6744), .ZN(n6742) );
  OAI21_X1 U7462 ( .B1(n6744), .B2(n6743), .A(n6742), .ZN(U3469) );
  INV_X1 U7463 ( .A(n6745), .ZN(n7021) );
  INV_X1 U7464 ( .A(n6746), .ZN(n6747) );
  AOI21_X1 U7465 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(n7016) );
  AOI22_X1 U7466 ( .A1(n7021), .A2(n6770), .B1(n6769), .B2(n7016), .ZN(n6750)
         );
  OAI21_X1 U7467 ( .B1(n6773), .B2(n6751), .A(n6750), .ZN(U2850) );
  AOI22_X1 U7468 ( .A1(n7342), .A2(n6770), .B1(n6769), .B2(n7124), .ZN(n6752)
         );
  OAI21_X1 U7469 ( .B1(n6773), .B2(n7121), .A(n6752), .ZN(U2838) );
  NAND2_X1 U7470 ( .A1(n6298), .A2(n6753), .ZN(n6754) );
  AND2_X1 U7471 ( .A1(n6293), .A2(n6754), .ZN(n7339) );
  OR2_X1 U7472 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  AND2_X1 U7473 ( .A1(n6758), .A2(n6757), .ZN(n7101) );
  AOI22_X1 U7474 ( .A1(n7339), .A2(n6770), .B1(n6769), .B2(n7101), .ZN(n6759)
         );
  OAI21_X1 U7475 ( .B1(n6773), .B2(n6760), .A(n6759), .ZN(U2840) );
  INV_X1 U7476 ( .A(n6761), .ZN(n6762) );
  AOI22_X1 U7477 ( .A1(n6763), .A2(n6770), .B1(n6769), .B2(n6762), .ZN(n6764)
         );
  OAI21_X1 U7478 ( .B1(n6773), .B2(n6765), .A(n6764), .ZN(U2844) );
  INV_X1 U7479 ( .A(n6766), .ZN(n6767) );
  XNOR2_X1 U7480 ( .A(n6768), .B(n6767), .ZN(n6957) );
  AOI22_X1 U7481 ( .A1(n6964), .A2(n6770), .B1(n6769), .B2(n6957), .ZN(n6771)
         );
  OAI21_X1 U7482 ( .B1(n6773), .B2(n6772), .A(n6771), .ZN(U2855) );
  AOI22_X1 U7483 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6779) );
  INV_X1 U7484 ( .A(n6931), .ZN(n6777) );
  XNOR2_X1 U7485 ( .A(n6775), .B(n6878), .ZN(n6776) );
  XNOR2_X1 U7486 ( .A(n6774), .B(n6776), .ZN(n6875) );
  AOI22_X1 U7487 ( .A1(n6777), .A2(n6818), .B1(n6875), .B2(n6819), .ZN(n6778)
         );
  OAI211_X1 U7488 ( .C1(n6822), .C2(n6938), .A(n6779), .B(n6778), .ZN(U2984)
         );
  AOI22_X1 U7489 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n6784) );
  XNOR2_X1 U7490 ( .A(n6781), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6782)
         );
  XNOR2_X1 U7491 ( .A(n6780), .B(n6782), .ZN(n6861) );
  AOI22_X1 U7492 ( .A1(n6861), .A2(n6819), .B1(n6818), .B2(n6944), .ZN(n6783)
         );
  OAI211_X1 U7493 ( .C1(n6822), .C2(n6951), .A(n6784), .B(n6783), .ZN(U2983)
         );
  AOI22_X1 U7494 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6790) );
  INV_X1 U7495 ( .A(n6787), .ZN(n6788) );
  AOI21_X1 U7496 ( .B1(n6785), .B2(n6786), .A(n6788), .ZN(n6856) );
  AOI22_X1 U7497 ( .A1(n6856), .A2(n6819), .B1(n6818), .B2(n6964), .ZN(n6789)
         );
  OAI211_X1 U7498 ( .C1(n6822), .C2(n6966), .A(n6790), .B(n6789), .ZN(U2982)
         );
  AOI22_X1 U7499 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n6795) );
  OAI22_X1 U7500 ( .A1(n6792), .A2(n6804), .B1(n6971), .B2(n6791), .ZN(n6793)
         );
  INV_X1 U7501 ( .A(n6793), .ZN(n6794) );
  OAI211_X1 U7502 ( .C1(n6822), .C2(n6972), .A(n6795), .B(n6794), .ZN(U2981)
         );
  AOI22_X1 U7503 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U7504 ( .A1(n6797), .A2(n6819), .B1(n6818), .B2(n6796), .ZN(n6798)
         );
  OAI211_X1 U7505 ( .C1(n6822), .C2(n6985), .A(n6799), .B(n6798), .ZN(U2980)
         );
  AOI22_X1 U7506 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6803) );
  INV_X1 U7507 ( .A(n6800), .ZN(n7043) );
  AOI22_X1 U7508 ( .A1(n7043), .A2(n6818), .B1(n7042), .B2(n6801), .ZN(n6802)
         );
  OAI211_X1 U7509 ( .C1(n6805), .C2(n6804), .A(n6803), .B(n6802), .ZN(U2974)
         );
  AOI22_X1 U7510 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6815) );
  INV_X1 U7511 ( .A(n6806), .ZN(n6807) );
  NAND2_X1 U7512 ( .A1(n6807), .A2(n6809), .ZN(n6810) );
  MUX2_X1 U7513 ( .A(n6810), .B(n6809), .S(n6808), .Z(n6812) );
  NAND2_X1 U7514 ( .A1(n6812), .A2(n6811), .ZN(n6909) );
  AOI22_X1 U7515 ( .A1(n6909), .A2(n6819), .B1(n6818), .B2(n7336), .ZN(n6814)
         );
  OAI211_X1 U7516 ( .C1(n6822), .C2(n7082), .A(n6815), .B(n6814), .ZN(U2969)
         );
  AOI22_X1 U7517 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4711), .B1(n6908), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U7518 ( .B1(n6381), .B2(n6817), .A(n6816), .ZN(n6843) );
  AOI22_X1 U7519 ( .A1(n6843), .A2(n6819), .B1(n6818), .B2(n7339), .ZN(n6820)
         );
  OAI211_X1 U7520 ( .C1(n6822), .C2(n7104), .A(n6821), .B(n6820), .ZN(U2967)
         );
  AND2_X1 U7521 ( .A1(n6823), .A2(n7221), .ZN(n6825) );
  OAI22_X1 U7522 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7207), .B1(n6825), .B2(
        n6824), .ZN(U2790) );
  OAI222_X1 U7523 ( .A1(n6829), .A2(n6827), .B1(n6829), .B2(n6826), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n7246), .ZN(U2791) );
  INV_X1 U7524 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6828) );
  AOI22_X1 U7525 ( .A1(n6829), .A2(READREQUEST_REG_SCAN_IN), .B1(n6828), .B2(
        n7246), .ZN(U3470) );
  INV_X1 U7526 ( .A(HOLD), .ZN(n7231) );
  NOR2_X1 U7527 ( .A1(n6830), .A2(n7231), .ZN(n7230) );
  INV_X1 U7528 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7233) );
  NOR2_X1 U7529 ( .A1(n7240), .A2(n7233), .ZN(n7239) );
  AOI21_X1 U7530 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7239), .ZN(n6832)
         );
  NAND2_X1 U7531 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7244) );
  OAI211_X1 U7532 ( .C1(n7230), .C2(n6832), .A(n6831), .B(n7244), .ZN(U3182)
         );
  NAND2_X1 U7533 ( .A1(READY_N), .A2(n3887), .ZN(n7204) );
  OAI211_X1 U7534 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(n7204), .B(n7216), .ZN(n6834) );
  OAI21_X1 U7535 ( .B1(n6835), .B2(n6834), .A(n6833), .ZN(U3150) );
  AOI211_X1 U7536 ( .C1(n4570), .C2(n7413), .A(n3887), .B(n6836), .ZN(n6837)
         );
  OAI21_X1 U7537 ( .B1(n6837), .B2(n7224), .A(n7216), .ZN(n6841) );
  AOI211_X1 U7538 ( .C1(n6668), .C2(n7250), .A(n6839), .B(n6838), .ZN(n6840)
         );
  MUX2_X1 U7539 ( .A(n6841), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6840), .Z(
        U3472) );
  AOI22_X1 U7540 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6842), .B1(n6908), .B2(REIP_REG_19__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7541 ( .A1(n6843), .A2(n6915), .B1(n6917), .B2(n7101), .ZN(n6844)
         );
  OAI211_X1 U7542 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6846), .A(n6845), .B(n6844), .ZN(U2999) );
  INV_X1 U7543 ( .A(n6847), .ZN(n6849) );
  AOI21_X1 U7544 ( .B1(n6849), .B2(n6917), .A(n6848), .ZN(n6853) );
  AOI22_X1 U7545 ( .A1(n6851), .A2(n6915), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6850), .ZN(n6852) );
  OAI211_X1 U7546 ( .C1(n6855), .C2(n6854), .A(n6853), .B(n6852), .ZN(U3005)
         );
  AOI22_X1 U7547 ( .A1(n6917), .A2(n6957), .B1(n6908), .B2(REIP_REG_4__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7548 ( .A1(n6856), .A2(n6915), .B1(INSTADDRPOINTER_REG_4__SCAN_IN), 
        .B2(n6862), .ZN(n6859) );
  OAI211_X1 U7549 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6880), .B(n6857), .ZN(n6858) );
  NAND3_X1 U7550 ( .A1(n6860), .A2(n6859), .A3(n6858), .ZN(U3014) );
  AOI22_X1 U7551 ( .A1(n6917), .A2(n6939), .B1(n6908), .B2(REIP_REG_3__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U7552 ( .A1(n6862), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6915), 
        .B2(n6861), .ZN(n6863) );
  OAI211_X1 U7553 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6865), .A(n6864), 
        .B(n6863), .ZN(U3015) );
  NAND2_X1 U7554 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6866), .ZN(n6879)
         );
  NAND2_X1 U7555 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6868) );
  OAI21_X1 U7556 ( .B1(n6878), .B2(n6868), .A(n6867), .ZN(n6869) );
  AND2_X1 U7557 ( .A1(n6870), .A2(n6869), .ZN(n6874) );
  INV_X1 U7558 ( .A(n6935), .ZN(n6872) );
  OAI22_X1 U7559 ( .A1(n6884), .A2(n6872), .B1(n6871), .B2(n6924), .ZN(n6873)
         );
  AOI211_X1 U7560 ( .C1(n6875), .C2(n6915), .A(n6874), .B(n6873), .ZN(n6876)
         );
  OAI221_X1 U7561 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6879), .C1(n6878), .C2(n6877), .A(n6876), .ZN(U3016) );
  NAND2_X1 U7562 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  NOR2_X1 U7563 ( .A1(n6882), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6886)
         );
  OAI21_X1 U7564 ( .B1(n6884), .B2(n6991), .A(n6883), .ZN(n6885) );
  AOI211_X1 U7565 ( .C1(n6887), .C2(n6915), .A(n6886), .B(n6885), .ZN(n6888)
         );
  OAI21_X1 U7566 ( .B1(n6890), .B2(n6889), .A(n6888), .ZN(U3011) );
  AOI21_X1 U7567 ( .B1(n6917), .B2(n7016), .A(n6891), .ZN(n6895) );
  AOI22_X1 U7568 ( .A1(n6893), .A2(n6915), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6892), .ZN(n6894) );
  OAI211_X1 U7569 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6896), .A(n6895), 
        .B(n6894), .ZN(U3009) );
  INV_X1 U7570 ( .A(n6897), .ZN(n7026) );
  INV_X1 U7571 ( .A(n6898), .ZN(n6899) );
  AOI21_X1 U7572 ( .B1(n6917), .B2(n7026), .A(n6899), .ZN(n6903) );
  INV_X1 U7573 ( .A(n6900), .ZN(n6901) );
  AOI22_X1 U7574 ( .A1(n6901), .A2(n6915), .B1(n6906), .B2(n6904), .ZN(n6902)
         );
  OAI211_X1 U7575 ( .C1(n6905), .C2(n6904), .A(n6903), .B(n6902), .ZN(U3007)
         );
  AOI22_X1 U7576 ( .A1(n6908), .A2(REIP_REG_17__SCAN_IN), .B1(n6907), .B2(
        n6906), .ZN(n6911) );
  AOI22_X1 U7577 ( .A1(n6909), .A2(n6915), .B1(n6917), .B2(n7079), .ZN(n6910)
         );
  OAI211_X1 U7578 ( .C1(n6913), .C2(n6912), .A(n6911), .B(n6910), .ZN(U3001)
         );
  INV_X1 U7579 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U7580 ( .A1(n6917), .A2(n6916), .B1(n6915), .B2(n6914), .ZN(n6923)
         );
  INV_X1 U7581 ( .A(n6918), .ZN(n6920) );
  OAI22_X1 U7582 ( .A1(n6921), .A2(n6920), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6919), .ZN(n6922) );
  OAI211_X1 U7583 ( .C1(n6925), .C2(n6924), .A(n6923), .B(n6922), .ZN(U3018)
         );
  AOI211_X1 U7584 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6941), .A(n6871), .B(n7106), 
        .ZN(n6928) );
  OAI22_X1 U7585 ( .A1(n7120), .A2(n6926), .B1(n5066), .B2(n6961), .ZN(n6927)
         );
  NOR2_X1 U7586 ( .A1(n6928), .A2(n6927), .ZN(n6937) );
  NAND3_X1 U7587 ( .A1(n7139), .A2(n6871), .A3(REIP_REG_1__SCAN_IN), .ZN(n6929) );
  OAI21_X1 U7588 ( .B1(n6930), .B2(n7122), .A(n6929), .ZN(n6934) );
  NOR2_X1 U7589 ( .A1(n6932), .A2(n6931), .ZN(n6933) );
  AOI211_X1 U7590 ( .C1(n6935), .C2(n7125), .A(n6934), .B(n6933), .ZN(n6936)
         );
  OAI211_X1 U7591 ( .C1(n6938), .C2(n7157), .A(n6937), .B(n6936), .ZN(U2825)
         );
  AOI22_X1 U7592 ( .A1(n7145), .A2(EBX_REG_3__SCAN_IN), .B1(n7125), .B2(n6939), 
        .ZN(n6950) );
  OR2_X1 U7593 ( .A1(n6953), .A2(n7075), .ZN(n6967) );
  NAND2_X1 U7594 ( .A1(n7074), .A2(n6967), .ZN(n6952) );
  AND2_X1 U7595 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6940) );
  AOI21_X1 U7596 ( .B1(n6941), .B2(n6940), .A(REIP_REG_3__SCAN_IN), .ZN(n6947)
         );
  OAI22_X1 U7597 ( .A1(n6942), .A2(n6961), .B1(n7122), .B2(n4152), .ZN(n6943)
         );
  INV_X1 U7598 ( .A(n6943), .ZN(n6946) );
  NAND2_X1 U7599 ( .A1(n6974), .A2(n6944), .ZN(n6945) );
  OAI211_X1 U7600 ( .C1(n6952), .C2(n6947), .A(n6946), .B(n6945), .ZN(n6948)
         );
  INV_X1 U7601 ( .A(n6948), .ZN(n6949) );
  OAI211_X1 U7602 ( .C1(n6951), .C2(n7157), .A(n6950), .B(n6949), .ZN(U2824)
         );
  NOR2_X1 U7603 ( .A1(n6952), .A2(n6954), .ZN(n6963) );
  NOR2_X1 U7604 ( .A1(n7147), .A2(n6953), .ZN(n6982) );
  AOI22_X1 U7605 ( .A1(EBX_REG_4__SCAN_IN), .A2(n7145), .B1(n6982), .B2(n6954), 
        .ZN(n6959) );
  NAND2_X1 U7606 ( .A1(n7144), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6955)
         );
  NAND2_X1 U7607 ( .A1(n6955), .A2(n7094), .ZN(n6956) );
  AOI21_X1 U7608 ( .B1(n7125), .B2(n6957), .A(n6956), .ZN(n6958) );
  OAI211_X1 U7609 ( .C1(n6961), .C2(n6960), .A(n6959), .B(n6958), .ZN(n6962)
         );
  AOI211_X1 U7610 ( .C1(n6964), .C2(n6974), .A(n6963), .B(n6962), .ZN(n6965)
         );
  OAI21_X1 U7611 ( .B1(n6966), .B2(n7157), .A(n6965), .ZN(U2823) );
  AOI21_X1 U7612 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6982), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6978) );
  OAI21_X1 U7613 ( .B1(n6983), .B2(n6967), .A(n7074), .ZN(n7003) );
  OAI22_X1 U7614 ( .A1(n7120), .A2(n6969), .B1(n7152), .B2(n6968), .ZN(n6970)
         );
  AOI211_X1 U7615 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n7086), 
        .B(n6970), .ZN(n6977) );
  INV_X1 U7616 ( .A(n6971), .ZN(n6975) );
  INV_X1 U7617 ( .A(n6972), .ZN(n6973) );
  AOI22_X1 U7618 ( .A1(n6975), .A2(n6974), .B1(n7133), .B2(n6973), .ZN(n6976)
         );
  OAI211_X1 U7619 ( .C1(n6978), .C2(n7003), .A(n6977), .B(n6976), .ZN(U2822)
         );
  OAI22_X1 U7620 ( .A1(n7120), .A2(n6980), .B1(n7152), .B2(n6979), .ZN(n6981)
         );
  AOI211_X1 U7621 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n7086), 
        .B(n6981), .ZN(n6990) );
  INV_X1 U7622 ( .A(n7003), .ZN(n6988) );
  INV_X1 U7623 ( .A(n6982), .ZN(n6984) );
  NOR2_X1 U7624 ( .A1(n6984), .A2(n6983), .ZN(n6999) );
  OAI22_X1 U7625 ( .A1(n6986), .A2(n7130), .B1(n6985), .B2(n7157), .ZN(n6987)
         );
  AOI221_X1 U7626 ( .B1(n6988), .B2(REIP_REG_6__SCAN_IN), .C1(n6999), .C2(
        n5388), .A(n6987), .ZN(n6989) );
  NAND2_X1 U7627 ( .A1(n6990), .A2(n6989), .ZN(U2821) );
  INV_X1 U7628 ( .A(n6991), .ZN(n6992) );
  AOI22_X1 U7629 ( .A1(n7145), .A2(EBX_REG_7__SCAN_IN), .B1(n7125), .B2(n6992), 
        .ZN(n6993) );
  NAND2_X1 U7630 ( .A1(n6993), .A2(n7094), .ZN(n6997) );
  OAI22_X1 U7631 ( .A1(n6995), .A2(n7130), .B1(n6994), .B2(n7157), .ZN(n6996)
         );
  AOI211_X1 U7632 ( .C1(PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n7144), .A(n6997), 
        .B(n6996), .ZN(n7001) );
  OAI211_X1 U7633 ( .C1(REIP_REG_6__SCAN_IN), .C2(REIP_REG_7__SCAN_IN), .A(
        n6999), .B(n6998), .ZN(n7000) );
  OAI211_X1 U7634 ( .C1(n7003), .C2(n7002), .A(n7001), .B(n7000), .ZN(U2820)
         );
  AOI21_X1 U7635 ( .B1(n7139), .B2(n7004), .A(REIP_REG_8__SCAN_IN), .ZN(n7013)
         );
  OAI22_X1 U7636 ( .A1(n7120), .A2(n7006), .B1(n7152), .B2(n7005), .ZN(n7007)
         );
  AOI211_X1 U7637 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n7086), 
        .B(n7007), .ZN(n7012) );
  INV_X1 U7638 ( .A(n7008), .ZN(n7010) );
  AOI22_X1 U7639 ( .A1(n7010), .A2(n7155), .B1(n7133), .B2(n7009), .ZN(n7011)
         );
  OAI211_X1 U7640 ( .C1(n7013), .C2(n7017), .A(n7012), .B(n7011), .ZN(U2819)
         );
  NOR3_X1 U7641 ( .A1(n7147), .A2(REIP_REG_9__SCAN_IN), .A3(n7014), .ZN(n7015)
         );
  AOI21_X1 U7642 ( .B1(n7016), .B2(n7125), .A(n7015), .ZN(n7025) );
  AOI22_X1 U7643 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n7144), .B1(
        EBX_REG_9__SCAN_IN), .B2(n7145), .ZN(n7024) );
  INV_X1 U7644 ( .A(n7017), .ZN(n7018) );
  AOI21_X1 U7645 ( .B1(REIP_REG_9__SCAN_IN), .B2(n7018), .A(n7086), .ZN(n7023)
         );
  INV_X1 U7646 ( .A(n7019), .ZN(n7020) );
  AOI22_X1 U7647 ( .A1(n7021), .A2(n7155), .B1(n7020), .B2(n7133), .ZN(n7022)
         );
  NAND4_X1 U7648 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(U2818)
         );
  AOI22_X1 U7649 ( .A1(n7125), .A2(n7026), .B1(PHYADDRPOINTER_REG_11__SCAN_IN), 
        .B2(n7144), .ZN(n7037) );
  INV_X1 U7650 ( .A(n7039), .ZN(n7030) );
  OR3_X1 U7651 ( .A1(n7147), .A2(REIP_REG_11__SCAN_IN), .A3(n7027), .ZN(n7028)
         );
  OAI21_X1 U7652 ( .B1(n7030), .B2(n7029), .A(n7028), .ZN(n7031) );
  AOI21_X1 U7653 ( .B1(EBX_REG_11__SCAN_IN), .B2(n7145), .A(n7031), .ZN(n7036)
         );
  INV_X1 U7654 ( .A(n7032), .ZN(n7033) );
  AOI22_X1 U7655 ( .A1(n7034), .A2(n7155), .B1(n7033), .B2(n7133), .ZN(n7035)
         );
  NAND4_X1 U7656 ( .A1(n7037), .A2(n7036), .A3(n7035), .A4(n7094), .ZN(U2816)
         );
  AOI22_X1 U7657 ( .A1(n7039), .A2(REIP_REG_12__SCAN_IN), .B1(n7125), .B2(
        n7038), .ZN(n7046) );
  OAI22_X1 U7658 ( .A1(REIP_REG_12__SCAN_IN), .A2(n7047), .B1(n7040), .B2(
        n7122), .ZN(n7041) );
  AOI211_X1 U7659 ( .C1(n7145), .C2(EBX_REG_12__SCAN_IN), .A(n7086), .B(n7041), 
        .ZN(n7045) );
  AOI22_X1 U7660 ( .A1(n7043), .A2(n7155), .B1(n7042), .B2(n7133), .ZN(n7044)
         );
  NAND3_X1 U7661 ( .A1(n7046), .A2(n7045), .A3(n7044), .ZN(U2815) );
  NOR2_X1 U7662 ( .A1(n7048), .A2(n7047), .ZN(n7050) );
  INV_X1 U7663 ( .A(n7060), .ZN(n7049) );
  MUX2_X1 U7664 ( .A(n7050), .B(n7049), .S(REIP_REG_14__SCAN_IN), .Z(n7051) );
  AOI211_X1 U7665 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7086), 
        .B(n7051), .ZN(n7057) );
  OAI22_X1 U7666 ( .A1(n7053), .A2(n7130), .B1(n7152), .B2(n7052), .ZN(n7054)
         );
  AOI21_X1 U7667 ( .B1(n7055), .B2(n7133), .A(n7054), .ZN(n7056) );
  OAI211_X1 U7668 ( .C1(n7058), .C2(n7120), .A(n7057), .B(n7056), .ZN(U2813)
         );
  XNOR2_X1 U7669 ( .A(n7061), .B(n7059), .ZN(n7062) );
  OAI22_X1 U7670 ( .A1(n7063), .A2(n7062), .B1(n7061), .B2(n7060), .ZN(n7064)
         );
  AOI211_X1 U7671 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7086), 
        .B(n7064), .ZN(n7070) );
  OAI22_X1 U7672 ( .A1(n7066), .A2(n7130), .B1(n7152), .B2(n7065), .ZN(n7067)
         );
  AOI21_X1 U7673 ( .B1(n7068), .B2(n7133), .A(n7067), .ZN(n7069) );
  OAI211_X1 U7674 ( .C1(n7071), .C2(n7120), .A(n7070), .B(n7069), .ZN(U2811)
         );
  AOI21_X1 U7675 ( .B1(n7073), .B2(n7072), .A(REIP_REG_17__SCAN_IN), .ZN(n7077) );
  OAI21_X1 U7676 ( .B1(n7075), .B2(n7083), .A(n7074), .ZN(n7105) );
  INV_X1 U7677 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7076) );
  OAI22_X1 U7678 ( .A1(n7077), .A2(n7105), .B1(n7076), .B2(n7122), .ZN(n7078)
         );
  AOI211_X1 U7679 ( .C1(n7145), .C2(EBX_REG_17__SCAN_IN), .A(n7086), .B(n7078), 
        .ZN(n7081) );
  AOI22_X1 U7680 ( .A1(n7336), .A2(n7155), .B1(n7125), .B2(n7079), .ZN(n7080)
         );
  OAI211_X1 U7681 ( .C1(n7082), .C2(n7157), .A(n7081), .B(n7080), .ZN(U2810)
         );
  INV_X1 U7682 ( .A(n7083), .ZN(n7084) );
  NAND2_X1 U7683 ( .A1(n7139), .A2(n7084), .ZN(n7118) );
  AOI22_X1 U7684 ( .A1(REIP_REG_18__SCAN_IN), .A2(n7105), .B1(n7118), .B2(
        n7096), .ZN(n7085) );
  AOI211_X1 U7685 ( .C1(n7144), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n7086), 
        .B(n7085), .ZN(n7092) );
  OAI22_X1 U7686 ( .A1(n7088), .A2(n7130), .B1(n7152), .B2(n7087), .ZN(n7089)
         );
  AOI21_X1 U7687 ( .B1(n7090), .B2(n7133), .A(n7089), .ZN(n7091) );
  OAI211_X1 U7688 ( .C1(n7093), .C2(n7120), .A(n7092), .B(n7091), .ZN(U2809)
         );
  INV_X1 U7689 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7095) );
  OAI21_X1 U7690 ( .B1(n7122), .B2(n7095), .A(n7094), .ZN(n7100) );
  XNOR2_X1 U7691 ( .A(n7097), .B(n7096), .ZN(n7098) );
  OAI22_X1 U7692 ( .A1(n7118), .A2(n7098), .B1(n7097), .B2(n7105), .ZN(n7099)
         );
  AOI211_X1 U7693 ( .C1(EBX_REG_19__SCAN_IN), .C2(n7145), .A(n7100), .B(n7099), 
        .ZN(n7103) );
  AOI22_X1 U7694 ( .A1(n7339), .A2(n7155), .B1(n7125), .B2(n7101), .ZN(n7102)
         );
  OAI211_X1 U7695 ( .C1(n7104), .C2(n7157), .A(n7103), .B(n7102), .ZN(U2808)
         );
  INV_X1 U7696 ( .A(n7119), .ZN(n7107) );
  OAI21_X1 U7697 ( .B1(n7107), .B2(n7106), .A(n7105), .ZN(n7135) );
  NAND2_X1 U7698 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n7109) );
  OAI21_X1 U7699 ( .B1(n7109), .B2(n7118), .A(n7108), .ZN(n7110) );
  AOI22_X1 U7700 ( .A1(EBX_REG_20__SCAN_IN), .A2(n7145), .B1(n7135), .B2(n7110), .ZN(n7116) );
  OAI22_X1 U7701 ( .A1(n7112), .A2(n7130), .B1(n7152), .B2(n7111), .ZN(n7113)
         );
  AOI21_X1 U7702 ( .B1(n7114), .B2(n7133), .A(n7113), .ZN(n7115) );
  OAI211_X1 U7703 ( .C1(n7117), .C2(n7122), .A(n7116), .B(n7115), .ZN(U2807)
         );
  NOR3_X1 U7704 ( .A1(REIP_REG_21__SCAN_IN), .A2(n7119), .A3(n7118), .ZN(n7136) );
  OAI22_X1 U7705 ( .A1(n6412), .A2(n7122), .B1(n7121), .B2(n7120), .ZN(n7123)
         );
  AOI211_X1 U7706 ( .C1(REIP_REG_21__SCAN_IN), .C2(n7135), .A(n7136), .B(n7123), .ZN(n7127) );
  AOI22_X1 U7707 ( .A1(n7342), .A2(n7155), .B1(n7125), .B2(n7124), .ZN(n7126)
         );
  OAI211_X1 U7708 ( .C1(n7128), .C2(n7157), .A(n7127), .B(n7126), .ZN(U2806)
         );
  AOI22_X1 U7709 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n7144), .B1(
        EBX_REG_22__SCAN_IN), .B2(n7145), .ZN(n7143) );
  OAI22_X1 U7710 ( .A1(n7131), .A2(n7130), .B1(n7152), .B2(n7129), .ZN(n7132)
         );
  AOI21_X1 U7711 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7142) );
  OAI21_X1 U7712 ( .B1(n7136), .B2(n7135), .A(REIP_REG_22__SCAN_IN), .ZN(n7141) );
  NAND3_X1 U7713 ( .A1(n7139), .A2(n7138), .A3(n7137), .ZN(n7140) );
  NAND4_X1 U7714 ( .A1(n7143), .A2(n7142), .A3(n7141), .A4(n7140), .ZN(U2805)
         );
  AOI22_X1 U7715 ( .A1(n7145), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n7144), .ZN(n7151) );
  NOR2_X1 U7716 ( .A1(n7147), .A2(n7146), .ZN(n7149) );
  OAI21_X1 U7717 ( .B1(REIP_REG_23__SCAN_IN), .B2(n7149), .A(n7148), .ZN(n7150) );
  OAI211_X1 U7718 ( .C1(n7153), .C2(n7152), .A(n7151), .B(n7150), .ZN(n7154)
         );
  AOI21_X1 U7719 ( .B1(n7345), .B2(n7155), .A(n7154), .ZN(n7156) );
  OAI21_X1 U7720 ( .B1(n7158), .B2(n7157), .A(n7156), .ZN(U2804) );
  NAND2_X1 U7721 ( .A1(n7159), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7177) );
  OR2_X1 U7722 ( .A1(n5092), .A2(n7160), .ZN(n7163) );
  NAND2_X1 U7723 ( .A1(n7161), .A2(n3650), .ZN(n7162) );
  NAND2_X1 U7724 ( .A1(n7163), .A2(n7162), .ZN(n7179) );
  INV_X1 U7725 ( .A(n7179), .ZN(n7165) );
  OAI22_X1 U7726 ( .A1(n7165), .A2(n7169), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n7164), .ZN(n7167) );
  OAI22_X1 U7727 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n7171), .B1(n7167), .B2(n7166), .ZN(n7168) );
  OAI21_X1 U7728 ( .B1(n7177), .B2(n7169), .A(n7168), .ZN(U3461) );
  NAND2_X1 U7729 ( .A1(n7170), .A2(n7214), .ZN(n7172) );
  OAI22_X1 U7730 ( .A1(n7173), .A2(n7172), .B1(n4175), .B2(n7171), .ZN(U3455)
         );
  AND2_X1 U7731 ( .A1(n7175), .A2(n7174), .ZN(n7189) );
  INV_X1 U7732 ( .A(n7175), .ZN(n7183) );
  NAND2_X1 U7733 ( .A1(n7175), .A2(n7176), .ZN(n7187) );
  NAND2_X1 U7734 ( .A1(n7177), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7178) );
  NOR2_X1 U7735 ( .A1(n7179), .A2(n7178), .ZN(n7181) );
  INV_X1 U7736 ( .A(n7181), .ZN(n7185) );
  INV_X1 U7737 ( .A(n7180), .ZN(n7182) );
  OAI22_X1 U7738 ( .A1(n7183), .A2(n7182), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7181), .ZN(n7184) );
  OAI21_X1 U7739 ( .B1(n7185), .B2(n7412), .A(n7184), .ZN(n7186) );
  AOI222_X1 U7740 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7187), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7186), .C1(n7187), .C2(n7186), 
        .ZN(n7188) );
  AOI222_X1 U7741 ( .A1(n7189), .A2(n7188), .B1(n7189), .B2(n7361), .C1(n7188), 
        .C2(n7361), .ZN(n7199) );
  INV_X1 U7742 ( .A(MORE_REG_SCAN_IN), .ZN(n7191) );
  AOI21_X1 U7743 ( .B1(n7192), .B2(n7191), .A(n7190), .ZN(n7195) );
  NOR4_X1 U7744 ( .A1(n7196), .A2(n7195), .A3(n7194), .A4(n7193), .ZN(n7197)
         );
  OAI211_X1 U7745 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7199), .A(n7198), .B(n7197), .ZN(n7220) );
  OAI22_X1 U7746 ( .A1(n7220), .A2(n7206), .B1(n7200), .B2(n7250), .ZN(n7201)
         );
  OAI21_X1 U7747 ( .B1(n7203), .B2(n7202), .A(n7201), .ZN(n7215) );
  AOI21_X1 U7748 ( .B1(n7215), .B2(n7204), .A(n7224), .ZN(n7218) );
  AOI21_X1 U7749 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7218), .A(n7205), .ZN(
        n7210) );
  OAI21_X1 U7750 ( .B1(READY_N), .B2(n7207), .A(n7206), .ZN(n7208) );
  NAND2_X1 U7751 ( .A1(n7215), .A2(n7208), .ZN(n7209) );
  OAI211_X1 U7752 ( .C1(n7211), .C2(n7215), .A(n7210), .B(n7209), .ZN(U3149)
         );
  OAI211_X1 U7753 ( .C1(n7214), .C2(n7215), .A(n7213), .B(n7212), .ZN(U3453)
         );
  OAI21_X1 U7754 ( .B1(n7217), .B2(n7216), .A(n7215), .ZN(n7225) );
  AOI211_X1 U7755 ( .C1(n7221), .C2(n7220), .A(n7219), .B(n7218), .ZN(n7222)
         );
  OAI221_X1 U7756 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n7225), .C1(n7224), .C2(
        n7223), .A(n7222), .ZN(U3148) );
  INV_X1 U7757 ( .A(n7226), .ZN(n7227) );
  OAI21_X1 U7758 ( .B1(n7229), .B2(n7413), .A(n7227), .ZN(U2792) );
  OAI21_X1 U7759 ( .B1(n7229), .B2(n7228), .A(n7227), .ZN(U3452) );
  INV_X1 U7760 ( .A(n7230), .ZN(n7236) );
  INV_X1 U7761 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7232) );
  NOR2_X1 U7762 ( .A1(n7232), .A2(n7231), .ZN(n7234) );
  INV_X1 U7763 ( .A(NA_N), .ZN(n7238) );
  AOI221_X1 U7764 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7238), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7242) );
  AOI221_X1 U7765 ( .B1(n7234), .B2(n7246), .C1(n7233), .C2(n7246), .A(n7242), 
        .ZN(n7235) );
  OAI221_X1 U7766 ( .B1(n7237), .B2(n7236), .C1(n7237), .C2(n7244), .A(n7235), 
        .ZN(U3181) );
  AOI21_X1 U7767 ( .B1(n7239), .B2(n7238), .A(STATE_REG_2__SCAN_IN), .ZN(n7245) );
  AOI221_X1 U7768 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7250), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7241) );
  AOI221_X1 U7769 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7241), .C2(HOLD), .A(n7240), .ZN(n7243) );
  OAI22_X1 U7770 ( .A1(n7245), .A2(n7244), .B1(n7243), .B2(n7242), .ZN(U3183)
         );
  AOI22_X1 U7771 ( .A1(n6829), .A2(n7248), .B1(n7247), .B2(n7246), .ZN(U3473)
         );
  OAI21_X1 U7772 ( .B1(n4570), .B2(n7250), .A(n7249), .ZN(n7327) );
  NOR2_X1 U7773 ( .A1(n7329), .A2(n7251), .ZN(n7254) );
  AOI21_X1 U7774 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n7330), .A(n7254), .ZN(n7252) );
  OAI21_X1 U7775 ( .B1(n7253), .B2(n7333), .A(n7252), .ZN(U2924) );
  AOI21_X1 U7776 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n7327), .A(n7254), .ZN(n7255) );
  OAI21_X1 U7777 ( .B1(n7256), .B2(n7333), .A(n7255), .ZN(U2939) );
  NOR2_X1 U7778 ( .A1(n7329), .A2(n7257), .ZN(n7259) );
  AOI21_X1 U7779 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n7330), .A(n7259), .ZN(n7258) );
  OAI21_X1 U7780 ( .B1(n4403), .B2(n7333), .A(n7258), .ZN(U2925) );
  AOI21_X1 U7781 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n7330), .A(n7259), .ZN(n7260) );
  OAI21_X1 U7782 ( .B1(n7261), .B2(n7333), .A(n7260), .ZN(U2940) );
  NOR2_X1 U7783 ( .A1(n7329), .A2(n5367), .ZN(n7264) );
  AOI21_X1 U7784 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n7330), .A(n7264), .ZN(n7262) );
  OAI21_X1 U7785 ( .B1(n7263), .B2(n7333), .A(n7262), .ZN(U2926) );
  AOI21_X1 U7786 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n7330), .A(n7264), .ZN(n7265) );
  OAI21_X1 U7787 ( .B1(n7266), .B2(n7333), .A(n7265), .ZN(U2941) );
  NOR2_X1 U7788 ( .A1(n7329), .A2(n7267), .ZN(n7269) );
  AOI21_X1 U7789 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n7330), .A(n7269), .ZN(n7268) );
  OAI21_X1 U7790 ( .B1(n4438), .B2(n7333), .A(n7268), .ZN(U2927) );
  AOI21_X1 U7791 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n7330), .A(n7269), .ZN(n7270) );
  OAI21_X1 U7792 ( .B1(n7271), .B2(n7333), .A(n7270), .ZN(U2942) );
  NOR2_X1 U7793 ( .A1(n7329), .A2(n7272), .ZN(n7275) );
  AOI21_X1 U7794 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n7330), .A(n7275), .ZN(n7273) );
  OAI21_X1 U7795 ( .B1(n7274), .B2(n7333), .A(n7273), .ZN(U2928) );
  AOI21_X1 U7796 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n7330), .A(n7275), .ZN(n7276) );
  OAI21_X1 U7797 ( .B1(n7277), .B2(n7333), .A(n7276), .ZN(U2943) );
  NOR2_X1 U7798 ( .A1(n7329), .A2(n5382), .ZN(n7280) );
  AOI21_X1 U7799 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n7330), .A(n7280), .ZN(n7278) );
  OAI21_X1 U7800 ( .B1(n7279), .B2(n7333), .A(n7278), .ZN(U2929) );
  AOI21_X1 U7801 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n7330), .A(n7280), .ZN(n7281) );
  OAI21_X1 U7802 ( .B1(n4202), .B2(n7333), .A(n7281), .ZN(U2944) );
  INV_X1 U7803 ( .A(DATAI_6_), .ZN(n7282) );
  NOR2_X1 U7804 ( .A1(n7329), .A2(n7282), .ZN(n7285) );
  AOI21_X1 U7805 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n7330), .A(n7285), .ZN(n7283) );
  OAI21_X1 U7806 ( .B1(n7284), .B2(n7333), .A(n7283), .ZN(U2930) );
  AOI21_X1 U7807 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n7330), .A(n7285), .ZN(n7286) );
  OAI21_X1 U7808 ( .B1(n4230), .B2(n7333), .A(n7286), .ZN(U2945) );
  NOR2_X1 U7809 ( .A1(n7329), .A2(n5849), .ZN(n7288) );
  AOI21_X1 U7810 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n7330), .A(n7288), .ZN(n7287) );
  OAI21_X1 U7811 ( .B1(n4506), .B2(n7333), .A(n7287), .ZN(U2931) );
  AOI21_X1 U7812 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n7330), .A(n7288), .ZN(n7289) );
  OAI21_X1 U7813 ( .B1(n7290), .B2(n7333), .A(n7289), .ZN(U2946) );
  NOR2_X1 U7814 ( .A1(n7329), .A2(n5851), .ZN(n7293) );
  AOI21_X1 U7815 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n7330), .A(n7293), .ZN(n7291) );
  OAI21_X1 U7816 ( .B1(n7292), .B2(n7333), .A(n7291), .ZN(U2932) );
  AOI21_X1 U7817 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n7330), .A(n7293), .ZN(n7294) );
  OAI21_X1 U7818 ( .B1(n7295), .B2(n7333), .A(n7294), .ZN(U2947) );
  NOR2_X1 U7819 ( .A1(n7329), .A2(n7296), .ZN(n7299) );
  AOI21_X1 U7820 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n7330), .A(n7299), .ZN(n7297) );
  OAI21_X1 U7821 ( .B1(n7298), .B2(n7333), .A(n7297), .ZN(U2933) );
  AOI21_X1 U7822 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n7330), .A(n7299), .ZN(n7300) );
  OAI21_X1 U7823 ( .B1(n7301), .B2(n7333), .A(n7300), .ZN(U2948) );
  NOR2_X1 U7824 ( .A1(n7329), .A2(n7302), .ZN(n7305) );
  AOI21_X1 U7825 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n7330), .A(n7305), .ZN(
        n7303) );
  OAI21_X1 U7826 ( .B1(n7304), .B2(n7333), .A(n7303), .ZN(U2934) );
  AOI21_X1 U7827 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n7330), .A(n7305), .ZN(
        n7306) );
  OAI21_X1 U7828 ( .B1(n7307), .B2(n7333), .A(n7306), .ZN(U2949) );
  NOR2_X1 U7829 ( .A1(n7329), .A2(n7308), .ZN(n7311) );
  AOI21_X1 U7830 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n7330), .A(n7311), .ZN(
        n7309) );
  OAI21_X1 U7831 ( .B1(n7310), .B2(n7333), .A(n7309), .ZN(U2935) );
  AOI21_X1 U7832 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n7330), .A(n7311), .ZN(
        n7312) );
  OAI21_X1 U7833 ( .B1(n7313), .B2(n7333), .A(n7312), .ZN(U2950) );
  NOR2_X1 U7834 ( .A1(n7329), .A2(n7314), .ZN(n7317) );
  AOI21_X1 U7835 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n7330), .A(n7317), .ZN(
        n7315) );
  OAI21_X1 U7836 ( .B1(n7316), .B2(n7333), .A(n7315), .ZN(U2936) );
  AOI21_X1 U7837 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n7330), .A(n7317), .ZN(
        n7318) );
  OAI21_X1 U7838 ( .B1(n4304), .B2(n7333), .A(n7318), .ZN(U2951) );
  NOR2_X1 U7839 ( .A1(n7329), .A2(n7319), .ZN(n7322) );
  AOI21_X1 U7840 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n7327), .A(n7322), .ZN(
        n7320) );
  OAI21_X1 U7841 ( .B1(n7321), .B2(n7333), .A(n7320), .ZN(U2937) );
  AOI21_X1 U7842 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n7327), .A(n7322), .ZN(
        n7323) );
  OAI21_X1 U7843 ( .B1(n7324), .B2(n7333), .A(n7323), .ZN(U2952) );
  NOR2_X1 U7844 ( .A1(n7329), .A2(n6080), .ZN(n7326) );
  AOI21_X1 U7845 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n7327), .A(n7326), .ZN(
        n7325) );
  OAI21_X1 U7846 ( .B1(n4740), .B2(n7333), .A(n7325), .ZN(U2938) );
  AOI21_X1 U7847 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n7327), .A(n7326), .ZN(
        n7328) );
  OAI21_X1 U7848 ( .B1(n4341), .B2(n7333), .A(n7328), .ZN(U2953) );
  INV_X1 U7849 ( .A(n7329), .ZN(n7331) );
  AOI22_X1 U7850 ( .A1(n7331), .A2(DATAI_15_), .B1(n7330), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n7332) );
  OAI21_X1 U7851 ( .B1(n7334), .B2(n7333), .A(n7332), .ZN(U2954) );
  INV_X1 U7852 ( .A(n7335), .ZN(n7435) );
  AOI22_X1 U7853 ( .A1(n7336), .A2(n7435), .B1(n7434), .B2(DATAI_17_), .ZN(
        n7338) );
  AOI22_X1 U7854 ( .A1(n7438), .A2(DATAI_1_), .B1(n7437), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U7855 ( .A1(n7338), .A2(n7337), .ZN(U2874) );
  AOI22_X1 U7856 ( .A1(n7339), .A2(n7435), .B1(n7434), .B2(DATAI_19_), .ZN(
        n7341) );
  AOI22_X1 U7857 ( .A1(n7438), .A2(DATAI_3_), .B1(n7437), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U7858 ( .A1(n7341), .A2(n7340), .ZN(U2872) );
  AOI22_X1 U7859 ( .A1(n7342), .A2(n7435), .B1(n7434), .B2(DATAI_21_), .ZN(
        n7344) );
  AOI22_X1 U7860 ( .A1(n7438), .A2(DATAI_5_), .B1(n7437), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U7861 ( .A1(n7344), .A2(n7343), .ZN(U2870) );
  AOI22_X1 U7862 ( .A1(n7345), .A2(n7435), .B1(n7434), .B2(DATAI_23_), .ZN(
        n7347) );
  AOI22_X1 U7863 ( .A1(n7438), .A2(DATAI_7_), .B1(n7437), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U7864 ( .A1(n7347), .A2(n7346), .ZN(U2868) );
  OAI21_X1 U7865 ( .B1(n7348), .B2(n7426), .A(n7400), .ZN(n7352) );
  INV_X1 U7866 ( .A(n7349), .ZN(n7399) );
  NOR2_X1 U7867 ( .A1(n7417), .A2(n7350), .ZN(n7537) );
  AOI21_X1 U7868 ( .B1(n7388), .B2(n7399), .A(n7537), .ZN(n7353) );
  INV_X1 U7869 ( .A(n7353), .ZN(n7351) );
  AOI22_X1 U7870 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7355), .B1(n7352), .B2(
        n7351), .ZN(n7543) );
  AOI22_X1 U7871 ( .A1(n7422), .A2(n7538), .B1(n7421), .B2(n7537), .ZN(n7357)
         );
  AOI21_X1 U7872 ( .B1(n7353), .B2(n7352), .A(n7424), .ZN(n7354) );
  OAI21_X1 U7873 ( .B1(n7415), .B2(n7355), .A(n7354), .ZN(n7540) );
  AOI22_X1 U7874 ( .A1(n7540), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n7430), 
        .B2(n7539), .ZN(n7356) );
  OAI211_X1 U7875 ( .C1(n7543), .C2(n7433), .A(n7357), .B(n7356), .ZN(U3124)
         );
  INV_X1 U7876 ( .A(n7368), .ZN(n7358) );
  OAI21_X1 U7877 ( .B1(n7358), .B2(n7426), .A(n7400), .ZN(n7366) );
  AND2_X1 U7878 ( .A1(n7360), .A2(n7359), .ZN(n7384) );
  NOR3_X1 U7879 ( .A1(n7412), .A2(n7361), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n7378) );
  INV_X1 U7880 ( .A(n7378), .ZN(n7362) );
  NOR2_X1 U7881 ( .A1(n7417), .A2(n7362), .ZN(n7544) );
  AOI21_X1 U7882 ( .B1(n7384), .B2(n7363), .A(n7544), .ZN(n7365) );
  INV_X1 U7883 ( .A(n7365), .ZN(n7364) );
  AOI22_X1 U7884 ( .A1(n7366), .A2(n7364), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7378), .ZN(n7549) );
  AOI22_X1 U7885 ( .A1(n7545), .A2(n7430), .B1(n7421), .B2(n7544), .ZN(n7370)
         );
  NAND2_X1 U7886 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  OAI211_X1 U7887 ( .C1(n7415), .C2(n7378), .A(n7408), .B(n7367), .ZN(n7546)
         );
  AOI22_X1 U7888 ( .A1(n7546), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7422), 
        .B2(n7551), .ZN(n7369) );
  OAI211_X1 U7889 ( .C1(n7549), .C2(n7433), .A(n7370), .B(n7369), .ZN(U3108)
         );
  NOR2_X1 U7890 ( .A1(n7556), .A2(n7426), .ZN(n7374) );
  AOI21_X1 U7891 ( .B1(n7374), .B2(n7373), .A(n7372), .ZN(n7383) );
  INV_X1 U7892 ( .A(n7383), .ZN(n7377) );
  NAND2_X1 U7893 ( .A1(n7417), .A2(n7378), .ZN(n7381) );
  INV_X1 U7894 ( .A(n7381), .ZN(n7550) );
  AOI22_X1 U7895 ( .A1(n7421), .A2(n7550), .B1(n7556), .B2(n7422), .ZN(n7386)
         );
  AOI211_X1 U7896 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7381), .A(n7380), .B(
        n7379), .ZN(n7382) );
  OAI21_X1 U7897 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7552) );
  AOI22_X1 U7898 ( .A1(n7552), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7430), 
        .B2(n7551), .ZN(n7385) );
  OAI211_X1 U7899 ( .C1(n7555), .C2(n7433), .A(n7386), .B(n7385), .ZN(U3100)
         );
  AOI21_X1 U7900 ( .B1(n7387), .B2(STATEBS16_REG_SCAN_IN), .A(n7426), .ZN(
        n7392) );
  NAND2_X1 U7901 ( .A1(n7388), .A2(n7418), .ZN(n7390) );
  NOR2_X1 U7902 ( .A1(n7417), .A2(n7393), .ZN(n7557) );
  INV_X1 U7903 ( .A(n7557), .ZN(n7389) );
  NAND2_X1 U7904 ( .A1(n7390), .A2(n7389), .ZN(n7396) );
  AOI22_X1 U7905 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7391), .B1(n7392), .B2(
        n7396), .ZN(n7562) );
  AOI22_X1 U7906 ( .A1(n7421), .A2(n7557), .B1(n7556), .B2(n7430), .ZN(n7398)
         );
  INV_X1 U7907 ( .A(n7392), .ZN(n7395) );
  AOI21_X1 U7908 ( .B1(n7426), .B2(n7393), .A(n7424), .ZN(n7394) );
  OAI21_X1 U7909 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7559) );
  AOI22_X1 U7910 ( .A1(n7559), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7422), 
        .B2(n7558), .ZN(n7397) );
  OAI211_X1 U7911 ( .C1(n7562), .C2(n7433), .A(n7398), .B(n7397), .ZN(U3092)
         );
  NOR2_X1 U7912 ( .A1(n7417), .A2(n7404), .ZN(n7563) );
  AOI21_X1 U7913 ( .B1(n7419), .B2(n7399), .A(n7563), .ZN(n7406) );
  INV_X1 U7914 ( .A(n7406), .ZN(n7402) );
  OAI21_X1 U7915 ( .B1(n7401), .B2(n7426), .A(n7400), .ZN(n7405) );
  AOI22_X1 U7916 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7403), .B1(n7402), .B2(
        n7405), .ZN(n7569) );
  AOI22_X1 U7917 ( .A1(n7430), .A2(n7565), .B1(n7421), .B2(n7563), .ZN(n7410)
         );
  AOI22_X1 U7918 ( .A1(n7406), .A2(n7405), .B1(n7426), .B2(n7404), .ZN(n7407)
         );
  NAND2_X1 U7919 ( .A1(n7408), .A2(n7407), .ZN(n7566) );
  AOI22_X1 U7920 ( .A1(n7566), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n7422), 
        .B2(n7564), .ZN(n7409) );
  OAI211_X1 U7921 ( .C1(n7569), .C2(n7433), .A(n7410), .B(n7409), .ZN(U3060)
         );
  NAND2_X1 U7922 ( .A1(n7412), .A2(n7411), .ZN(n7425) );
  OR2_X1 U7923 ( .A1(n7414), .A2(n7413), .ZN(n7416) );
  NAND2_X1 U7924 ( .A1(n7416), .A2(n7415), .ZN(n7429) );
  NOR2_X1 U7925 ( .A1(n7417), .A2(n7425), .ZN(n7570) );
  AOI21_X1 U7926 ( .B1(n7419), .B2(n7418), .A(n7570), .ZN(n7423) );
  OAI22_X1 U7927 ( .A1(n3887), .A2(n7425), .B1(n7429), .B2(n7423), .ZN(n7420)
         );
  AOI22_X1 U7928 ( .A1(n7422), .A2(n7573), .B1(n7421), .B2(n7570), .ZN(n7432)
         );
  INV_X1 U7929 ( .A(n7423), .ZN(n7428) );
  AOI21_X1 U7930 ( .B1(n7426), .B2(n7425), .A(n7424), .ZN(n7427) );
  OAI21_X1 U7931 ( .B1(n7429), .B2(n7428), .A(n7427), .ZN(n7575) );
  AOI22_X1 U7932 ( .A1(n7575), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n7430), 
        .B2(n3642), .ZN(n7431) );
  OAI211_X1 U7933 ( .C1(n7579), .C2(n7433), .A(n7432), .B(n7431), .ZN(U3028)
         );
  AOI22_X1 U7934 ( .A1(n7436), .A2(n7435), .B1(n7434), .B2(DATAI_24_), .ZN(
        n7440) );
  AOI22_X1 U7935 ( .A1(n7438), .A2(DATAI_8_), .B1(n7437), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U7936 ( .A1(n7440), .A2(n7439), .ZN(U2867) );
  AOI22_X1 U7937 ( .A1(n7452), .A2(n7539), .B1(n7451), .B2(n7537), .ZN(n7442)
         );
  AOI22_X1 U7938 ( .A1(n7540), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n7453), 
        .B2(n7538), .ZN(n7441) );
  OAI211_X1 U7939 ( .C1(n7543), .C2(n7456), .A(n7442), .B(n7441), .ZN(U3125)
         );
  AOI22_X1 U7940 ( .A1(n7545), .A2(n7452), .B1(n7451), .B2(n7544), .ZN(n7444)
         );
  AOI22_X1 U7941 ( .A1(n7546), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7453), 
        .B2(n7551), .ZN(n7443) );
  OAI211_X1 U7942 ( .C1(n7549), .C2(n7456), .A(n7444), .B(n7443), .ZN(U3109)
         );
  AOI22_X1 U7943 ( .A1(n7451), .A2(n7550), .B1(n7556), .B2(n7453), .ZN(n7446)
         );
  AOI22_X1 U7944 ( .A1(n7552), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7452), 
        .B2(n7551), .ZN(n7445) );
  OAI211_X1 U7945 ( .C1(n7555), .C2(n7456), .A(n7446), .B(n7445), .ZN(U3101)
         );
  AOI22_X1 U7946 ( .A1(n7451), .A2(n7557), .B1(n7556), .B2(n7452), .ZN(n7448)
         );
  AOI22_X1 U7947 ( .A1(n7559), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7453), 
        .B2(n7558), .ZN(n7447) );
  OAI211_X1 U7948 ( .C1(n7562), .C2(n7456), .A(n7448), .B(n7447), .ZN(U3093)
         );
  AOI22_X1 U7949 ( .A1(n7452), .A2(n7565), .B1(n7451), .B2(n7563), .ZN(n7450)
         );
  AOI22_X1 U7950 ( .A1(n7566), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n7453), 
        .B2(n7564), .ZN(n7449) );
  OAI211_X1 U7951 ( .C1(n7569), .C2(n7456), .A(n7450), .B(n7449), .ZN(U3061)
         );
  AOI22_X1 U7952 ( .A1(n7452), .A2(n3642), .B1(n7451), .B2(n7570), .ZN(n7455)
         );
  AOI22_X1 U7953 ( .A1(n7575), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n7453), 
        .B2(n7573), .ZN(n7454) );
  OAI211_X1 U7954 ( .C1(n7579), .C2(n7456), .A(n7455), .B(n7454), .ZN(U3029)
         );
  AOI22_X1 U7955 ( .A1(n7468), .A2(n7538), .B1(n7467), .B2(n7537), .ZN(n7458)
         );
  AOI22_X1 U7956 ( .A1(n7540), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n7469), 
        .B2(n7539), .ZN(n7457) );
  OAI211_X1 U7957 ( .C1(n7543), .C2(n7472), .A(n7458), .B(n7457), .ZN(U3126)
         );
  AOI22_X1 U7958 ( .A1(n7551), .A2(n7468), .B1(n7467), .B2(n7544), .ZN(n7460)
         );
  AOI22_X1 U7959 ( .A1(n7546), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7469), 
        .B2(n7545), .ZN(n7459) );
  OAI211_X1 U7960 ( .C1(n7549), .C2(n7472), .A(n7460), .B(n7459), .ZN(U3110)
         );
  AOI22_X1 U7961 ( .A1(n7467), .A2(n7550), .B1(n7556), .B2(n7468), .ZN(n7462)
         );
  AOI22_X1 U7962 ( .A1(n7552), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7469), 
        .B2(n7551), .ZN(n7461) );
  OAI211_X1 U7963 ( .C1(n7555), .C2(n7472), .A(n7462), .B(n7461), .ZN(U3102)
         );
  AOI22_X1 U7964 ( .A1(n7467), .A2(n7557), .B1(n7556), .B2(n7469), .ZN(n7464)
         );
  AOI22_X1 U7965 ( .A1(n7559), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7468), 
        .B2(n7558), .ZN(n7463) );
  OAI211_X1 U7966 ( .C1(n7562), .C2(n7472), .A(n7464), .B(n7463), .ZN(U3094)
         );
  AOI22_X1 U7967 ( .A1(n7469), .A2(n7565), .B1(n7467), .B2(n7563), .ZN(n7466)
         );
  AOI22_X1 U7968 ( .A1(n7566), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n7468), 
        .B2(n7564), .ZN(n7465) );
  OAI211_X1 U7969 ( .C1(n7569), .C2(n7472), .A(n7466), .B(n7465), .ZN(U3062)
         );
  AOI22_X1 U7970 ( .A1(n7468), .A2(n7573), .B1(n7467), .B2(n7570), .ZN(n7471)
         );
  AOI22_X1 U7971 ( .A1(n7575), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n7469), 
        .B2(n3642), .ZN(n7470) );
  OAI211_X1 U7972 ( .C1(n7579), .C2(n7472), .A(n7471), .B(n7470), .ZN(U3030)
         );
  AOI22_X1 U7973 ( .A1(n7485), .A2(n7539), .B1(n7483), .B2(n7537), .ZN(n7474)
         );
  AOI22_X1 U7974 ( .A1(n7540), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n7484), 
        .B2(n7538), .ZN(n7473) );
  OAI211_X1 U7975 ( .C1(n7543), .C2(n7488), .A(n7474), .B(n7473), .ZN(U3127)
         );
  AOI22_X1 U7976 ( .A1(n7545), .A2(n7485), .B1(n7483), .B2(n7544), .ZN(n7476)
         );
  AOI22_X1 U7977 ( .A1(n7546), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7484), 
        .B2(n7551), .ZN(n7475) );
  OAI211_X1 U7978 ( .C1(n7549), .C2(n7488), .A(n7476), .B(n7475), .ZN(U3111)
         );
  AOI22_X1 U7979 ( .A1(n7483), .A2(n7550), .B1(n7556), .B2(n7484), .ZN(n7478)
         );
  AOI22_X1 U7980 ( .A1(n7552), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7485), 
        .B2(n7551), .ZN(n7477) );
  OAI211_X1 U7981 ( .C1(n7555), .C2(n7488), .A(n7478), .B(n7477), .ZN(U3103)
         );
  AOI22_X1 U7982 ( .A1(n7483), .A2(n7557), .B1(n7556), .B2(n7485), .ZN(n7480)
         );
  AOI22_X1 U7983 ( .A1(n7559), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n7484), 
        .B2(n7558), .ZN(n7479) );
  OAI211_X1 U7984 ( .C1(n7562), .C2(n7488), .A(n7480), .B(n7479), .ZN(U3095)
         );
  AOI22_X1 U7985 ( .A1(n7484), .A2(n7564), .B1(n7483), .B2(n7563), .ZN(n7482)
         );
  AOI22_X1 U7986 ( .A1(n7566), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n7485), 
        .B2(n7565), .ZN(n7481) );
  OAI211_X1 U7987 ( .C1(n7569), .C2(n7488), .A(n7482), .B(n7481), .ZN(U3063)
         );
  AOI22_X1 U7988 ( .A1(n7484), .A2(n7573), .B1(n7483), .B2(n7570), .ZN(n7487)
         );
  AOI22_X1 U7989 ( .A1(n7575), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n7485), 
        .B2(n3642), .ZN(n7486) );
  OAI211_X1 U7990 ( .C1(n7579), .C2(n7488), .A(n7487), .B(n7486), .ZN(U3031)
         );
  AOI22_X1 U7991 ( .A1(n7501), .A2(n7539), .B1(n7499), .B2(n7537), .ZN(n7490)
         );
  AOI22_X1 U7992 ( .A1(n7540), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n7500), 
        .B2(n7538), .ZN(n7489) );
  OAI211_X1 U7993 ( .C1(n7543), .C2(n7504), .A(n7490), .B(n7489), .ZN(U3128)
         );
  AOI22_X1 U7994 ( .A1(n7545), .A2(n7501), .B1(n7499), .B2(n7544), .ZN(n7492)
         );
  AOI22_X1 U7995 ( .A1(n7546), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7500), 
        .B2(n7551), .ZN(n7491) );
  OAI211_X1 U7996 ( .C1(n7549), .C2(n7504), .A(n7492), .B(n7491), .ZN(U3112)
         );
  AOI22_X1 U7997 ( .A1(n7499), .A2(n7550), .B1(n7556), .B2(n7500), .ZN(n7494)
         );
  AOI22_X1 U7998 ( .A1(n7552), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7501), 
        .B2(n7551), .ZN(n7493) );
  OAI211_X1 U7999 ( .C1(n7555), .C2(n7504), .A(n7494), .B(n7493), .ZN(U3104)
         );
  AOI22_X1 U8000 ( .A1(n7499), .A2(n7557), .B1(n7556), .B2(n7501), .ZN(n7496)
         );
  AOI22_X1 U8001 ( .A1(n7559), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7500), 
        .B2(n7558), .ZN(n7495) );
  OAI211_X1 U8002 ( .C1(n7562), .C2(n7504), .A(n7496), .B(n7495), .ZN(U3096)
         );
  AOI22_X1 U8003 ( .A1(n7500), .A2(n7564), .B1(n7499), .B2(n7563), .ZN(n7498)
         );
  AOI22_X1 U8004 ( .A1(n7566), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n7501), 
        .B2(n7565), .ZN(n7497) );
  OAI211_X1 U8005 ( .C1(n7569), .C2(n7504), .A(n7498), .B(n7497), .ZN(U3064)
         );
  AOI22_X1 U8006 ( .A1(n7500), .A2(n7573), .B1(n7499), .B2(n7570), .ZN(n7503)
         );
  AOI22_X1 U8007 ( .A1(n7575), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n7501), 
        .B2(n3642), .ZN(n7502) );
  OAI211_X1 U8008 ( .C1(n7579), .C2(n7504), .A(n7503), .B(n7502), .ZN(U3032)
         );
  AOI22_X1 U8009 ( .A1(n7516), .A2(n7539), .B1(n7515), .B2(n7537), .ZN(n7506)
         );
  AOI22_X1 U8010 ( .A1(n7540), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n7517), 
        .B2(n7538), .ZN(n7505) );
  OAI211_X1 U8011 ( .C1(n7543), .C2(n7520), .A(n7506), .B(n7505), .ZN(U3129)
         );
  AOI22_X1 U8012 ( .A1(n7551), .A2(n7517), .B1(n7515), .B2(n7544), .ZN(n7508)
         );
  AOI22_X1 U8013 ( .A1(n7546), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7516), 
        .B2(n7545), .ZN(n7507) );
  OAI211_X1 U8014 ( .C1(n7549), .C2(n7520), .A(n7508), .B(n7507), .ZN(U3113)
         );
  AOI22_X1 U8015 ( .A1(n7515), .A2(n7550), .B1(n7556), .B2(n7517), .ZN(n7510)
         );
  AOI22_X1 U8016 ( .A1(n7552), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7516), 
        .B2(n7551), .ZN(n7509) );
  OAI211_X1 U8017 ( .C1(n7555), .C2(n7520), .A(n7510), .B(n7509), .ZN(U3105)
         );
  AOI22_X1 U8018 ( .A1(n7515), .A2(n7557), .B1(n7556), .B2(n7516), .ZN(n7512)
         );
  AOI22_X1 U8019 ( .A1(n7559), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n7517), 
        .B2(n7558), .ZN(n7511) );
  OAI211_X1 U8020 ( .C1(n7562), .C2(n7520), .A(n7512), .B(n7511), .ZN(U3097)
         );
  AOI22_X1 U8021 ( .A1(n7517), .A2(n7564), .B1(n7515), .B2(n7563), .ZN(n7514)
         );
  AOI22_X1 U8022 ( .A1(n7566), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n7516), 
        .B2(n7565), .ZN(n7513) );
  OAI211_X1 U8023 ( .C1(n7569), .C2(n7520), .A(n7514), .B(n7513), .ZN(U3065)
         );
  AOI22_X1 U8024 ( .A1(n7516), .A2(n3642), .B1(n7515), .B2(n7570), .ZN(n7519)
         );
  AOI22_X1 U8025 ( .A1(n7575), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n7517), 
        .B2(n7573), .ZN(n7518) );
  OAI211_X1 U8026 ( .C1(n7579), .C2(n7520), .A(n7519), .B(n7518), .ZN(U3033)
         );
  AOI22_X1 U8027 ( .A1(n7532), .A2(n7538), .B1(n7531), .B2(n7537), .ZN(n7522)
         );
  AOI22_X1 U8028 ( .A1(n7540), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n7533), 
        .B2(n7539), .ZN(n7521) );
  OAI211_X1 U8029 ( .C1(n7543), .C2(n7536), .A(n7522), .B(n7521), .ZN(U3130)
         );
  AOI22_X1 U8030 ( .A1(n7545), .A2(n7533), .B1(n7531), .B2(n7544), .ZN(n7524)
         );
  AOI22_X1 U8031 ( .A1(n7546), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7532), 
        .B2(n7551), .ZN(n7523) );
  OAI211_X1 U8032 ( .C1(n7549), .C2(n7536), .A(n7524), .B(n7523), .ZN(U3114)
         );
  AOI22_X1 U8033 ( .A1(n7531), .A2(n7550), .B1(n7556), .B2(n7532), .ZN(n7526)
         );
  AOI22_X1 U8034 ( .A1(n7552), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7533), 
        .B2(n7551), .ZN(n7525) );
  OAI211_X1 U8035 ( .C1(n7555), .C2(n7536), .A(n7526), .B(n7525), .ZN(U3106)
         );
  AOI22_X1 U8036 ( .A1(n7558), .A2(n7532), .B1(n7531), .B2(n7557), .ZN(n7528)
         );
  AOI22_X1 U8037 ( .A1(n7559), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7533), 
        .B2(n7556), .ZN(n7527) );
  OAI211_X1 U8038 ( .C1(n7562), .C2(n7536), .A(n7528), .B(n7527), .ZN(U3098)
         );
  AOI22_X1 U8039 ( .A1(n7533), .A2(n7565), .B1(n7531), .B2(n7563), .ZN(n7530)
         );
  AOI22_X1 U8040 ( .A1(n7566), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n7532), 
        .B2(n7564), .ZN(n7529) );
  OAI211_X1 U8041 ( .C1(n7569), .C2(n7536), .A(n7530), .B(n7529), .ZN(U3066)
         );
  AOI22_X1 U8042 ( .A1(n7532), .A2(n7573), .B1(n7531), .B2(n7570), .ZN(n7535)
         );
  AOI22_X1 U8043 ( .A1(n7575), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n7533), 
        .B2(n3642), .ZN(n7534) );
  OAI211_X1 U8044 ( .C1(n7579), .C2(n7536), .A(n7535), .B(n7534), .ZN(U3034)
         );
  AOI22_X1 U8045 ( .A1(n7574), .A2(n7538), .B1(n7571), .B2(n7537), .ZN(n7542)
         );
  AOI22_X1 U8046 ( .A1(n7540), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n7572), 
        .B2(n7539), .ZN(n7541) );
  OAI211_X1 U8047 ( .C1(n7543), .C2(n7578), .A(n7542), .B(n7541), .ZN(U3131)
         );
  AOI22_X1 U8048 ( .A1(n7545), .A2(n7572), .B1(n7571), .B2(n7544), .ZN(n7548)
         );
  AOI22_X1 U8049 ( .A1(n7546), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7574), 
        .B2(n7551), .ZN(n7547) );
  OAI211_X1 U8050 ( .C1(n7549), .C2(n7578), .A(n7548), .B(n7547), .ZN(U3115)
         );
  AOI22_X1 U8051 ( .A1(n7571), .A2(n7550), .B1(n7556), .B2(n7574), .ZN(n7554)
         );
  AOI22_X1 U8052 ( .A1(n7552), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7572), 
        .B2(n7551), .ZN(n7553) );
  OAI211_X1 U8053 ( .C1(n7555), .C2(n7578), .A(n7554), .B(n7553), .ZN(U3107)
         );
  AOI22_X1 U8054 ( .A1(n7571), .A2(n7557), .B1(n7556), .B2(n7572), .ZN(n7561)
         );
  AOI22_X1 U8055 ( .A1(n7559), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7574), 
        .B2(n7558), .ZN(n7560) );
  OAI211_X1 U8056 ( .C1(n7562), .C2(n7578), .A(n7561), .B(n7560), .ZN(U3099)
         );
  AOI22_X1 U8057 ( .A1(n7574), .A2(n7564), .B1(n7571), .B2(n7563), .ZN(n7568)
         );
  AOI22_X1 U8058 ( .A1(n7566), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7572), 
        .B2(n7565), .ZN(n7567) );
  OAI211_X1 U8059 ( .C1(n7569), .C2(n7578), .A(n7568), .B(n7567), .ZN(U3067)
         );
  AOI22_X1 U8060 ( .A1(n7572), .A2(n3642), .B1(n7571), .B2(n7570), .ZN(n7577)
         );
  AOI22_X1 U8061 ( .A1(n7575), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n7574), 
        .B2(n7573), .ZN(n7576) );
  OAI211_X1 U8062 ( .C1(n7579), .C2(n7578), .A(n7577), .B(n7576), .ZN(U3035)
         );
  INV_X1 U3833 ( .A(n3964), .ZN(n3687) );
  XNOR2_X1 U4568 ( .A(n4083), .B(n4084), .ZN(n4087) );
  NAND2_X1 U3693 ( .A1(n4222), .A2(n4221), .ZN(n4616) );
  NAND2_X1 U3699 ( .A1(n4100), .A2(n4101), .ZN(n5031) );
  CLKBUF_X1 U3671 ( .A(n3962), .Z(n4015) );
  CLKBUF_X1 U3697 ( .A(n4093), .Z(n4094) );
  AND4_X1 U3834 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3850)
         );
  NAND2_X1 U4014 ( .A1(n4613), .A2(n4612), .ZN(n4614) );
  CLKBUF_X1 U4019 ( .A(n4070), .Z(n5092) );
  XNOR2_X1 U4406 ( .A(n4087), .B(n4056), .ZN(n5083) );
  CLKBUF_X1 U4593 ( .A(n6209), .Z(n6210) );
  NOR2_X2 U4602 ( .A1(n6209), .A2(n3644), .ZN(n4746) );
endmodule

