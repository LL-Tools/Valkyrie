

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9583, n9584, n9585, n9586, n9587, n9588, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477;

  INV_X2 U11027 ( .A(n20924), .ZN(n20856) );
  OAI21_X1 U11028 ( .B1(n20504), .B2(n20519), .A(n20731), .ZN(n20521) );
  INV_X1 U11029 ( .A(n21013), .ZN(n14888) );
  NOR2_X1 U11030 ( .A1(n19390), .A2(n19175), .ZN(n19226) );
  INV_X2 U11031 ( .A(n16495), .ZN(n20133) );
  INV_X1 U11032 ( .A(n20970), .ZN(n21002) );
  AND2_X1 U11033 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11287), .ZN(
        n16951) );
  AND2_X1 U11034 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9663) );
  OR2_X1 U11035 ( .A1(n12571), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17571) );
  AND2_X1 U11036 ( .A1(n12211), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12246) );
  AND2_X1 U11037 ( .A1(n10127), .A2(n9605), .ZN(n20560) );
  NOR2_X2 U11038 ( .A1(n9605), .A2(n10678), .ZN(n10817) );
  CLKBUF_X2 U11039 ( .A(n11185), .Z(n9585) );
  XNOR2_X1 U11040 ( .A(n10685), .B(n10684), .ZN(n13244) );
  BUF_X1 U11041 ( .A(n10659), .Z(n10146) );
  OAI21_X1 U11042 ( .B1(n9804), .B2(n9803), .A(n10663), .ZN(n9802) );
  INV_X1 U11043 ( .A(n18476), .ZN(n19449) );
  NAND2_X2 U11044 ( .A1(n11809), .A2(n11810), .ZN(n12405) );
  CLKBUF_X2 U11045 ( .A(n10658), .Z(n11185) );
  CLKBUF_X2 U11046 ( .A(n10652), .Z(n11173) );
  INV_X1 U11047 ( .A(n21477), .ZN(n9591) );
  INV_X1 U11048 ( .A(n11733), .ZN(n11835) );
  BUF_X1 U11049 ( .A(n12324), .Z(n12256) );
  CLKBUF_X1 U11050 ( .A(n12321), .Z(n12263) );
  CLKBUF_X2 U11051 ( .A(n11728), .Z(n12334) );
  INV_X1 U11052 ( .A(n11192), .ZN(n12775) );
  INV_X1 U11055 ( .A(n14317), .ZN(n14569) );
  CLKBUF_X3 U11056 ( .A(n13867), .Z(n9597) );
  INV_X1 U11057 ( .A(n9583), .ZN(n9588) );
  INV_X1 U11058 ( .A(n14041), .ZN(n13389) );
  INV_X1 U11060 ( .A(n21477), .ZN(n9592) );
  NAND2_X1 U11061 ( .A1(n9899), .A2(n14568), .ZN(n10169) );
  OR2_X1 U11062 ( .A1(n11600), .A2(n11599), .ZN(n14299) );
  INV_X1 U11063 ( .A(n21477), .ZN(n9590) );
  NAND2_X1 U11064 ( .A1(n10926), .A2(n10947), .ZN(n13320) );
  NAND2_X1 U11065 ( .A1(n10947), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13324) );
  INV_X1 U11066 ( .A(n9583), .ZN(n9587) );
  INV_X1 U11067 ( .A(n21477), .ZN(n9593) );
  NAND2_X2 U11069 ( .A1(n14132), .A2(n14518), .ZN(n17438) );
  AND2_X1 U11070 ( .A1(n11694), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11573) );
  AND2_X1 U11071 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14216) );
  AND2_X1 U11072 ( .A1(n10179), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11574) );
  NOR2_X2 U11073 ( .A1(n17192), .A2(n20636), .ZN(n20743) );
  INV_X1 U11074 ( .A(n20731), .ZN(n20636) );
  AND3_X1 U11075 ( .A1(n10496), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13569) );
  CLKBUF_X2 U11076 ( .A(n12117), .Z(n12284) );
  AND2_X1 U11077 ( .A1(n11220), .A2(n17205), .ZN(n10603) );
  INV_X1 U11078 ( .A(n13320), .ZN(n13391) );
  NOR2_X1 U11079 ( .A1(n11054), .A2(n10378), .ZN(n11035) );
  OR2_X1 U11080 ( .A1(n10965), .A2(n10371), .ZN(n11028) );
  OR2_X1 U11081 ( .A1(n16814), .A2(n16815), .ZN(n16789) );
  CLKBUF_X3 U11082 ( .A(n10698), .Z(n9624) );
  INV_X1 U11083 ( .A(n13092), .ZN(n9594) );
  NAND2_X1 U11084 ( .A1(n12609), .A2(n14299), .ZN(n11665) );
  INV_X1 U11085 ( .A(n11660), .ZN(n9602) );
  AND2_X2 U11086 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14214) );
  NAND2_X1 U11087 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  INV_X1 U11088 ( .A(n16297), .ZN(n16250) );
  INV_X1 U11090 ( .A(n20319), .ZN(n20316) );
  AND2_X1 U11091 ( .A1(n10679), .A2(n14039), .ZN(n20726) );
  BUF_X1 U11092 ( .A(n13867), .Z(n9599) );
  NOR2_X1 U11094 ( .A1(n11665), .A2(n14569), .ZN(n10295) );
  INV_X2 U11095 ( .A(n21018), .ZN(n20983) );
  NAND2_X1 U11096 ( .A1(n13189), .A2(n11095), .ZN(n11543) );
  INV_X1 U11097 ( .A(n16282), .ZN(n16288) );
  INV_X1 U11098 ( .A(n12490), .ZN(n11342) );
  NAND2_X1 U11099 ( .A1(n10617), .A2(n10618), .ZN(n10664) );
  OAI21_X1 U11100 ( .B1(n10143), .B2(n10027), .A(n10026), .ZN(n11551) );
  AOI21_X1 U11101 ( .B1(n16758), .B2(n16699), .A(n16698), .ZN(n16732) );
  AND2_X1 U11102 ( .A1(n11238), .A2(n11212), .ZN(n17266) );
  OR2_X1 U11103 ( .A1(n14062), .A2(n17814), .ZN(n13147) );
  INV_X1 U11104 ( .A(n18167), .ZN(n18179) );
  INV_X1 U11105 ( .A(n19089), .ZN(n19080) );
  INV_X1 U11106 ( .A(n19304), .ZN(n19269) );
  INV_X1 U11107 ( .A(n21006), .ZN(n21014) );
  NAND2_X1 U11108 ( .A1(n14686), .A2(n14688), .ZN(n14687) );
  INV_X1 U11109 ( .A(n15029), .ZN(n15022) );
  INV_X1 U11110 ( .A(n14304), .ZN(n14541) );
  AOI21_X1 U11111 ( .B1(n14666), .B2(n14665), .A(n14664), .ZN(n15093) );
  AOI21_X1 U11112 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(n15221) );
  AOI21_X1 U11113 ( .B1(n13701), .B2(n13702), .A(n13251), .ZN(n13717) );
  CLKBUF_X3 U11114 ( .A(n10620), .Z(n11297) );
  INV_X1 U11115 ( .A(n20409), .ZN(n20457) );
  INV_X1 U11116 ( .A(n10457), .ZN(n18518) );
  AOI211_X1 U11117 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14641), .A(n14632), 
        .B(n14631), .ZN(n14633) );
  XNOR2_X1 U11118 ( .A(n13718), .B(n13717), .ZN(n20889) );
  INV_X1 U11119 ( .A(n19088), .ZN(n19100) );
  NAND2_X1 U11120 ( .A1(n13042), .A2(n13044), .ZN(n9583) );
  INV_X1 U11121 ( .A(n9583), .ZN(n9586) );
  NAND2_X1 U11122 ( .A1(n13036), .A2(n14518), .ZN(n9584) );
  INV_X4 U11124 ( .A(n17438), .ZN(n17465) );
  XNOR2_X2 U11125 ( .A(n9921), .B(n14392), .ZN(n14213) );
  NAND2_X2 U11126 ( .A1(n11705), .A2(n11706), .ZN(n9921) );
  NOR2_X4 U11127 ( .A1(n14858), .A2(n14956), .ZN(n14846) );
  AOI21_X2 U11128 ( .B1(n14004), .B2(n9998), .A(n9683), .ZN(n9997) );
  NAND2_X2 U11129 ( .A1(n10648), .A2(n10647), .ZN(n10658) );
  AND2_X4 U11130 ( .A1(n9624), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11395) );
  AOI21_X4 U11131 ( .B1(n16528), .B2(n20912), .A(n10306), .ZN(n16273) );
  XNOR2_X2 U11132 ( .A(n12778), .B(n12777), .ZN(n16528) );
  NAND2_X2 U11133 ( .A1(n17646), .A2(n10797), .ZN(n17060) );
  AND2_X4 U11135 ( .A1(n13031), .A2(n14131), .ZN(n13076) );
  XNOR2_X2 U11136 ( .A(n17299), .B(n17297), .ZN(n17296) );
  NAND2_X2 U11137 ( .A1(n9991), .A2(n14022), .ZN(n17299) );
  AND2_X1 U11138 ( .A1(n13043), .A2(n14132), .ZN(n13860) );
  CLKBUF_X3 U11139 ( .A(n13860), .Z(n17466) );
  AND2_X4 U11141 ( .A1(n14131), .A2(n14518), .ZN(n13057) );
  NOR2_X4 U11142 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14131) );
  AND2_X4 U11143 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14518) );
  NOR2_X2 U11144 ( .A1(n19094), .A2(n19396), .ZN(n19093) );
  INV_X4 U11145 ( .A(n9594), .ZN(n9595) );
  INV_X2 U11146 ( .A(n9594), .ZN(n9596) );
  NOR2_X2 U11147 ( .A1(n13141), .A2(n13965), .ZN(n17814) );
  AND2_X1 U11148 ( .A1(n13036), .A2(n13031), .ZN(n13867) );
  NOR2_X2 U11149 ( .A1(n19104), .A2(n17689), .ZN(n17693) );
  AND2_X1 U11150 ( .A1(n10327), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9932) );
  INV_X1 U11151 ( .A(n14484), .ZN(n9600) );
  INV_X2 U11153 ( .A(n19009), .ZN(n18970) );
  CLKBUF_X2 U11154 ( .A(n12583), .Z(n15245) );
  INV_X1 U11155 ( .A(n20704), .ZN(n20765) );
  AND2_X1 U11156 ( .A1(n17331), .A2(n17330), .ZN(n19857) );
  INV_X1 U11157 ( .A(n20257), .ZN(n9601) );
  NOR2_X1 U11159 ( .A1(n20143), .A2(n20636), .ZN(n20755) );
  INV_X1 U11160 ( .A(n11350), .ZN(n14348) );
  NOR2_X1 U11161 ( .A1(n20271), .A2(n20636), .ZN(n20767) );
  CLKBUF_X2 U11162 ( .A(n13244), .Z(n20214) );
  NAND2_X2 U11163 ( .A1(n19375), .A2(n19398), .ZN(n19304) );
  CLKBUF_X2 U11164 ( .A(n13245), .Z(n13666) );
  AND2_X1 U11166 ( .A1(n10637), .A2(n10633), .ZN(n9941) );
  NAND2_X1 U11167 ( .A1(n9799), .A2(n11297), .ZN(n10659) );
  CLKBUF_X2 U11168 ( .A(n11098), .Z(n11186) );
  OR2_X1 U11169 ( .A1(n10639), .A2(n11309), .ZN(n10647) );
  INV_X1 U11171 ( .A(n11488), .ZN(n11305) );
  NAND2_X1 U11172 ( .A1(n19426), .A2(n18518), .ZN(n13135) );
  NAND2_X1 U11173 ( .A1(n10323), .A2(n12621), .ZN(n13843) );
  CLKBUF_X2 U11174 ( .A(n10604), .Z(n11192) );
  CLKBUF_X2 U11175 ( .A(n11323), .Z(n12489) );
  INV_X4 U11176 ( .A(n19430), .ZN(n14057) );
  INV_X2 U11177 ( .A(n13829), .ZN(n14579) );
  INV_X2 U11179 ( .A(n12626), .ZN(n10323) );
  NAND2_X2 U11180 ( .A1(n10134), .A2(n10133), .ZN(n17183) );
  INV_X2 U11181 ( .A(n13322), .ZN(n13392) );
  INV_X1 U11182 ( .A(n13324), .ZN(n13390) );
  AND2_X2 U11183 ( .A1(n13413), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10773) );
  CLKBUF_X2 U11185 ( .A(n10699), .Z(n13413) );
  BUF_X2 U11186 ( .A(n12201), .Z(n12017) );
  CLKBUF_X2 U11187 ( .A(n11625), .Z(n12176) );
  CLKBUF_X2 U11188 ( .A(n12257), .Z(n12322) );
  INV_X1 U11189 ( .A(n13069), .ZN(n9608) );
  BUF_X2 U11190 ( .A(n12332), .Z(n9607) );
  CLKBUF_X2 U11191 ( .A(n11746), .Z(n12255) );
  CLKBUF_X3 U11192 ( .A(n13569), .Z(n9609) );
  CLKBUF_X2 U11193 ( .A(n13569), .Z(n9617) );
  CLKBUF_X2 U11194 ( .A(n13569), .Z(n9616) );
  AND2_X1 U11195 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14221) );
  NOR2_X1 U11196 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11575) );
  AND2_X1 U11197 ( .A1(n13211), .A2(n10484), .ZN(n13212) );
  AND2_X1 U11198 ( .A1(n10092), .A2(n10091), .ZN(n16921) );
  NOR2_X1 U11199 ( .A1(n9699), .A2(n16918), .ZN(n16933) );
  AND2_X1 U11200 ( .A1(n10136), .A2(n10135), .ZN(n16886) );
  NAND2_X1 U11201 ( .A1(n9919), .A2(n9918), .ZN(n16691) );
  OR2_X1 U11202 ( .A1(n16580), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9862) );
  NOR2_X1 U11203 ( .A1(n16583), .A2(n12449), .ZN(n16918) );
  NOR2_X1 U11204 ( .A1(n10475), .A2(n13201), .ZN(n16788) );
  XNOR2_X1 U11205 ( .A(n12355), .B(n12354), .ZN(n15042) );
  NAND2_X1 U11206 ( .A1(n16579), .A2(n9785), .ZN(n16571) );
  NOR3_X1 U11207 ( .A1(n10236), .A2(n10235), .A3(n15861), .ZN(n10234) );
  NAND2_X1 U11208 ( .A1(n16579), .A2(n10914), .ZN(n16543) );
  INV_X1 U11209 ( .A(n16583), .ZN(n9603) );
  NAND2_X1 U11210 ( .A1(n13505), .A2(n13504), .ZN(n16310) );
  OR2_X1 U11211 ( .A1(n13505), .A2(n13504), .ZN(n10149) );
  OAI21_X1 U11212 ( .B1(n16641), .B2(n10424), .A(n10421), .ZN(n16600) );
  XNOR2_X1 U11213 ( .A(n14597), .B(n13214), .ZN(n14531) );
  NAND2_X1 U11214 ( .A1(n16547), .A2(n16805), .ZN(n16800) );
  OAI21_X1 U11215 ( .B1(n13193), .B2(n10363), .A(n10361), .ZN(n10475) );
  AND2_X1 U11216 ( .A1(n12852), .A2(n12851), .ZN(n12853) );
  AND2_X1 U11217 ( .A1(n15863), .A2(n15862), .ZN(n10235) );
  AND2_X1 U11218 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  NOR2_X1 U11219 ( .A1(n18751), .A2(n19006), .ZN(n17491) );
  NAND2_X1 U11220 ( .A1(n13481), .A2(n13480), .ZN(n13505) );
  NAND2_X1 U11221 ( .A1(n10125), .A2(n10123), .ZN(n16641) );
  NAND2_X1 U11222 ( .A1(n13193), .A2(n10362), .ZN(n10361) );
  CLKBUF_X1 U11223 ( .A(n14686), .Z(n14701) );
  NOR2_X1 U11224 ( .A1(n13196), .A2(n16544), .ZN(n13193) );
  NAND2_X1 U11225 ( .A1(n10031), .A2(n9637), .ZN(n10125) );
  CLKBUF_X1 U11226 ( .A(n16321), .Z(n16334) );
  NAND2_X1 U11227 ( .A1(n9831), .A2(n10069), .ZN(n9791) );
  OR2_X1 U11228 ( .A1(n16322), .A2(n16325), .ZN(n13481) );
  AND2_X1 U11229 ( .A1(n11551), .A2(n11550), .ZN(n13196) );
  AOI211_X1 U11230 ( .C1(n21014), .C2(P1_EBX_REG_3__SCAN_IN), .A(n14892), .B(
        n14891), .ZN(n14893) );
  NAND2_X1 U11231 ( .A1(n15848), .A2(n11538), .ZN(n12492) );
  AND2_X1 U11232 ( .A1(n16831), .A2(n11290), .ZN(n16806) );
  AND2_X1 U11233 ( .A1(n15897), .A2(n10356), .ZN(n15848) );
  NOR2_X1 U11234 ( .A1(n16749), .A2(n9780), .ZN(n10383) );
  AOI21_X1 U11235 ( .B1(n16768), .B2(n16696), .A(n16695), .ZN(n16758) );
  NAND2_X1 U11236 ( .A1(n10126), .A2(n9700), .ZN(n10420) );
  AND2_X1 U11237 ( .A1(n16842), .A2(n16844), .ZN(n16831) );
  AND2_X1 U11238 ( .A1(n10304), .A2(n10303), .ZN(n10302) );
  NAND2_X1 U11239 ( .A1(n10906), .A2(n10908), .ZN(n16749) );
  AND2_X1 U11240 ( .A1(n10069), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9935) );
  AND2_X1 U11241 ( .A1(n17841), .A2(n10198), .ZN(n17834) );
  INV_X1 U11242 ( .A(n16533), .ZN(n10218) );
  AND2_X1 U11243 ( .A1(n12276), .A2(n10305), .ZN(n10304) );
  AOI21_X1 U11244 ( .B1(n10423), .B2(n9717), .A(n10422), .ZN(n10421) );
  NAND2_X1 U11245 ( .A1(n10045), .A2(n17040), .ZN(n10069) );
  XNOR2_X1 U11246 ( .A(n12501), .B(n11558), .ZN(n12850) );
  AND3_X1 U11247 ( .A1(n11549), .A2(n11548), .A3(n16554), .ZN(n11550) );
  AOI21_X1 U11248 ( .B1(n20492), .B2(n9869), .A(n20493), .ZN(n20500) );
  OR2_X1 U11249 ( .A1(n17069), .A2(n11005), .ZN(n11007) );
  NAND2_X1 U11250 ( .A1(n9793), .A2(n17071), .ZN(n10852) );
  CLKBUF_X1 U11251 ( .A(n17060), .Z(n17061) );
  INV_X1 U11252 ( .A(n10366), .ZN(n11557) );
  OR2_X1 U11253 ( .A1(n12984), .A2(n12252), .ZN(n12986) );
  NAND2_X1 U11254 ( .A1(n17105), .A2(n17104), .ZN(n17646) );
  NAND2_X1 U11255 ( .A1(n13277), .A2(n10155), .ZN(n16353) );
  NOR2_X1 U11256 ( .A1(n15206), .A2(n15208), .ZN(n12585) );
  NAND2_X1 U11257 ( .A1(n17184), .A2(n17219), .ZN(n20468) );
  AND2_X1 U11258 ( .A1(n11090), .A2(n11095), .ZN(n15917) );
  INV_X1 U11259 ( .A(n10848), .ZN(n9604) );
  AND2_X1 U11260 ( .A1(n9846), .A2(n10847), .ZN(n10849) );
  AND2_X1 U11261 ( .A1(n9845), .A2(n10879), .ZN(n10883) );
  INV_X1 U11262 ( .A(n20876), .ZN(n17184) );
  AND2_X1 U11263 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18924), .ZN(
        n19157) );
  AND2_X1 U11264 ( .A1(n11038), .A2(n11037), .ZN(n15997) );
  AND2_X1 U11265 ( .A1(n11077), .A2(n10367), .ZN(n15899) );
  NAND2_X1 U11266 ( .A1(n10010), .A2(n10013), .ZN(n18891) );
  NAND2_X1 U11267 ( .A1(n17340), .A2(n19007), .ZN(n19289) );
  NOR2_X1 U11268 ( .A1(n18969), .A2(n19236), .ZN(n18924) );
  OR2_X1 U11269 ( .A1(n14666), .A2(n12854), .ZN(n12984) );
  AND2_X1 U11270 ( .A1(n10822), .A2(n10827), .ZN(n10018) );
  AND2_X1 U11271 ( .A1(n11047), .A2(n11046), .ZN(n16072) );
  OAI21_X1 U11272 ( .B1(n10720), .B2(n10721), .A(n10116), .ZN(n10115) );
  AND4_X1 U11273 ( .A1(n10162), .A2(n10163), .A3(n10160), .A4(n10161), .ZN(
        n10070) );
  NAND2_X1 U11274 ( .A1(n12246), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12250) );
  AND2_X1 U11275 ( .A1(n10118), .A2(n10117), .ZN(n10116) );
  OR2_X1 U11276 ( .A1(n20677), .A2(n10725), .ZN(n10160) );
  NOR2_X2 U11277 ( .A1(n19857), .A2(n19906), .ZN(n17816) );
  CLKBUF_X1 U11278 ( .A(n14570), .Z(n15008) );
  NAND2_X1 U11279 ( .A1(n14203), .A2(n10408), .ZN(n16163) );
  AND2_X1 U11280 ( .A1(n11035), .A2(n16360), .ZN(n11033) );
  INV_X1 U11281 ( .A(n11833), .ZN(n11834) );
  OR2_X1 U11282 ( .A1(n20217), .A2(n11281), .ZN(n11282) );
  OR2_X1 U11283 ( .A1(n16909), .A2(n20218), .ZN(n11283) );
  AOI22_X1 U11284 ( .A1(n10816), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n20726), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11285 ( .A1(n10819), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n20560), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10162) );
  OR2_X1 U11286 ( .A1(n18905), .A2(n10272), .ZN(n18992) );
  XNOR2_X1 U11287 ( .A(n18905), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19322) );
  OR2_X1 U11288 ( .A1(n13240), .A2(n13241), .ZN(n10148) );
  AND2_X1 U11289 ( .A1(n10674), .A2(n14039), .ZN(n10818) );
  AND2_X1 U11290 ( .A1(n14039), .A2(n10671), .ZN(n20629) );
  NOR2_X2 U11291 ( .A1(n14039), .A2(n10670), .ZN(n10816) );
  NAND2_X1 U11292 ( .A1(n13228), .A2(n13227), .ZN(n13256) );
  INV_X1 U11293 ( .A(n10691), .ZN(n10690) );
  NAND2_X1 U11294 ( .A1(n10686), .A2(n17649), .ZN(n20257) );
  NAND2_X1 U11295 ( .A1(n11563), .A2(n17267), .ZN(n20217) );
  NAND2_X1 U11296 ( .A1(n11563), .A2(n11263), .ZN(n16909) );
  OR2_X1 U11297 ( .A1(n19875), .A2(n17329), .ZN(n17330) );
  INV_X1 U11298 ( .A(n20871), .ZN(n20251) );
  INV_X1 U11299 ( .A(n11056), .ZN(n9976) );
  NAND2_X1 U11300 ( .A1(n17296), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10274) );
  AND2_X1 U11301 ( .A1(n10689), .A2(n20243), .ZN(n10687) );
  NAND2_X1 U11302 ( .A1(n11822), .A2(n11821), .ZN(n14336) );
  NAND2_X2 U11303 ( .A1(n21035), .A2(n14317), .ZN(n14963) );
  NOR2_X1 U11304 ( .A1(n10688), .A2(n20214), .ZN(n10686) );
  NAND2_X1 U11305 ( .A1(n9977), .A2(n9761), .ZN(n11056) );
  INV_X2 U11306 ( .A(n20112), .ZN(n16418) );
  NAND2_X1 U11307 ( .A1(n12530), .A2(n11780), .ZN(n11802) );
  NOR2_X2 U11308 ( .A1(n19874), .A2(n18679), .ZN(n20042) );
  BUF_X2 U11309 ( .A(n9618), .Z(n9605) );
  NAND2_X1 U11310 ( .A1(n12535), .A2(n12534), .ZN(n13808) );
  NAND2_X1 U11311 ( .A1(n9802), .A2(n9800), .ZN(n10242) );
  NAND2_X2 U11312 ( .A1(n17117), .A2(n17116), .ZN(n20731) );
  CLKBUF_X1 U11313 ( .A(n14900), .Z(n21206) );
  OAI21_X1 U11314 ( .B1(n14900), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11741), 
        .ZN(n12530) );
  OR2_X1 U11315 ( .A1(n13676), .A2(n11240), .ZN(n10064) );
  CLKBUF_X1 U11316 ( .A(n21169), .Z(n21309) );
  OAI21_X1 U11317 ( .B1(n13245), .B2(n17114), .A(n13248), .ZN(n13663) );
  OR2_X1 U11318 ( .A1(n14098), .A2(n16226), .ZN(n10407) );
  AND2_X1 U11319 ( .A1(n14175), .A2(n9724), .ZN(n16204) );
  NAND2_X1 U11320 ( .A1(n9992), .A2(n14015), .ZN(n19029) );
  AND2_X1 U11321 ( .A1(n10656), .A2(n10657), .ZN(n10244) );
  NAND2_X1 U11322 ( .A1(n13620), .A2(n17287), .ZN(n20077) );
  CLKBUF_X1 U11323 ( .A(n11790), .Z(n14290) );
  NAND2_X1 U11324 ( .A1(n10650), .A2(n10649), .ZN(n10667) );
  NAND2_X1 U11325 ( .A1(n10050), .A2(n10049), .ZN(n11238) );
  AOI21_X1 U11326 ( .B1(n10662), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10643), .ZN(n10644) );
  NAND2_X1 U11327 ( .A1(n10435), .A2(n10651), .ZN(n10655) );
  OR2_X1 U11328 ( .A1(n12824), .A2(n11164), .ZN(n12825) );
  AOI22_X1 U11329 ( .A1(n10662), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n10130), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U11330 ( .A1(n10662), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10435) );
  AND2_X1 U11331 ( .A1(n10645), .A2(n10464), .ZN(n10650) );
  NAND2_X2 U11332 ( .A1(n14026), .A2(n14025), .ZN(n19006) );
  NAND2_X1 U11333 ( .A1(n10637), .A2(n9990), .ZN(n10662) );
  INV_X1 U11334 ( .A(n10659), .ZN(n11175) );
  CLKBUF_X1 U11335 ( .A(n12418), .Z(n13849) );
  AND2_X1 U11336 ( .A1(n13133), .A2(n19430), .ZN(n9962) );
  NAND2_X1 U11337 ( .A1(n11954), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12030) );
  INV_X1 U11338 ( .A(n10639), .ZN(n9799) );
  AND2_X1 U11339 ( .A1(n11242), .A2(n10065), .ZN(n11259) );
  OAI21_X1 U11340 ( .B1(n11674), .B2(n12599), .A(n12727), .ZN(n11676) );
  NAND2_X1 U11341 ( .A1(n10619), .A2(n13680), .ZN(n10639) );
  NOR2_X1 U11342 ( .A1(n13007), .A2(n18776), .ZN(n18764) );
  AND2_X1 U11343 ( .A1(n12809), .A2(n10285), .ZN(n12813) );
  NOR2_X1 U11344 ( .A1(n13135), .A2(n14083), .ZN(n13133) );
  NOR3_X1 U11345 ( .A1(n18518), .A2(n13129), .A3(n14083), .ZN(n14084) );
  NAND2_X1 U11346 ( .A1(n12410), .A2(n10492), .ZN(n12615) );
  AND2_X1 U11347 ( .A1(n10623), .A2(n10622), .ZN(n11226) );
  AND2_X1 U11348 ( .A1(n10771), .A2(n10770), .ZN(n10952) );
  AND3_X1 U11349 ( .A1(n10589), .A2(n10590), .A3(n10606), .ZN(n10621) );
  OR2_X1 U11350 ( .A1(n10878), .A2(n10877), .ZN(n11347) );
  INV_X2 U11351 ( .A(n11223), .ZN(n10599) );
  NAND2_X1 U11352 ( .A1(n19449), .A2(n18479), .ZN(n9975) );
  NAND2_X1 U11353 ( .A1(n15500), .A2(n14541), .ZN(n12411) );
  AND2_X1 U11354 ( .A1(n10753), .A2(n10752), .ZN(n11303) );
  INV_X2 U11355 ( .A(n11309), .ZN(n16324) );
  AND4_X1 U11356 ( .A1(n10704), .A2(n10703), .A3(n10702), .A4(n10701), .ZN(
        n10716) );
  XNOR2_X2 U11357 ( .A(n13996), .B(n18611), .ZN(n13999) );
  INV_X2 U11358 ( .A(U212), .ZN(n17753) );
  NAND2_X1 U11359 ( .A1(n9602), .A2(n14568), .ZN(n11662) );
  NAND2_X1 U11360 ( .A1(n9632), .A2(n9681), .ZN(n13996) );
  NAND2_X1 U11361 ( .A1(n10463), .A2(n10467), .ZN(n18479) );
  CLKBUF_X1 U11362 ( .A(n10595), .Z(n17239) );
  OR2_X1 U11363 ( .A1(n13109), .A2(n13108), .ZN(n18476) );
  BUF_X2 U11364 ( .A(n10620), .Z(n11309) );
  INV_X1 U11365 ( .A(n10620), .ZN(n10601) );
  OR2_X1 U11366 ( .A1(n13087), .A2(n13086), .ZN(n13985) );
  NOR2_X1 U11367 ( .A1(n18896), .A2(n13006), .ZN(n18878) );
  AND4_X2 U11368 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13049), .ZN(
        n19430) );
  OR2_X2 U11369 ( .A1(n17764), .A2(n17708), .ZN(n17766) );
  NAND2_X2 U11370 ( .A1(n10563), .A2(n10562), .ZN(n10625) );
  NAND2_X1 U11371 ( .A1(n10551), .A2(n10550), .ZN(n17224) );
  NAND2_X1 U11372 ( .A1(n10539), .A2(n10538), .ZN(n10595) );
  NAND2_X1 U11373 ( .A1(n9994), .A2(n9993), .ZN(n10593) );
  NAND2_X1 U11374 ( .A1(n10433), .A2(n10431), .ZN(n10620) );
  INV_X2 U11375 ( .A(n11663), .ZN(n9899) );
  INV_X1 U11377 ( .A(n14568), .ZN(n11659) );
  CLKBUF_X1 U11378 ( .A(n11663), .Z(n14294) );
  AND2_X1 U11379 ( .A1(n10488), .A2(n10491), .ZN(n12609) );
  NAND2_X1 U11380 ( .A1(n10489), .A2(n11609), .ZN(n11663) );
  AND4_X1 U11381 ( .A1(n10769), .A2(n10768), .A3(n10767), .A4(n10766), .ZN(
        n10770) );
  OR2_X2 U11382 ( .A1(n11642), .A2(n11641), .ZN(n14304) );
  NAND2_X1 U11383 ( .A1(n11580), .A2(n10490), .ZN(n11660) );
  OR2_X1 U11384 ( .A1(n12794), .A2(n12790), .ZN(n12792) );
  OR2_X2 U11385 ( .A1(n11618), .A2(n11619), .ZN(n14317) );
  AND3_X1 U11386 ( .A1(n10509), .A2(n14056), .A3(n10508), .ZN(n10416) );
  AND2_X1 U11387 ( .A1(n10511), .A2(n10510), .ZN(n10415) );
  AND2_X1 U11388 ( .A1(n10515), .A2(n9687), .ZN(n9995) );
  AND2_X1 U11389 ( .A1(n10498), .A2(n10497), .ZN(n9911) );
  AND3_X1 U11390 ( .A1(n10541), .A2(n14056), .A3(n10540), .ZN(n10544) );
  AND2_X1 U11391 ( .A1(n10506), .A2(n10504), .ZN(n9913) );
  INV_X2 U11392 ( .A(n17799), .ZN(U215) );
  INV_X1 U11393 ( .A(n9584), .ZN(n9619) );
  AND4_X1 U11394 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11580) );
  BUF_X2 U11395 ( .A(n13859), .Z(n18420) );
  INV_X2 U11396 ( .A(n21466), .ZN(n21067) );
  BUF_X2 U11397 ( .A(n11734), .Z(n12333) );
  BUF_X2 U11398 ( .A(n11745), .Z(n12331) );
  AND2_X2 U11399 ( .A1(n10705), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10802) );
  AND2_X2 U11400 ( .A1(n10576), .A2(n14056), .ZN(n13397) );
  CLKBUF_X3 U11401 ( .A(n13859), .Z(n18395) );
  CLKBUF_X3 U11402 ( .A(n13110), .Z(n18421) );
  NAND2_X2 U11403 ( .A1(n20018), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19996) );
  NAND2_X2 U11404 ( .A1(n20018), .A2(n19934), .ZN(n19982) );
  NAND2_X2 U11405 ( .A1(n13366), .A2(n14056), .ZN(n14041) );
  AND2_X1 U11406 ( .A1(n13042), .A2(n13043), .ZN(n13110) );
  CLKBUF_X3 U11407 ( .A(n13103), .Z(n18342) );
  AND2_X1 U11408 ( .A1(n13036), .A2(n13044), .ZN(n13092) );
  AND2_X2 U11409 ( .A1(n14245), .A2(n14224), .ZN(n12330) );
  NOR2_X1 U11410 ( .A1(n19039), .A2(n19038), .ZN(n18963) );
  INV_X2 U11411 ( .A(n17802), .ZN(n17804) );
  AND2_X1 U11412 ( .A1(n14131), .A2(n13044), .ZN(n13081) );
  NOR2_X1 U11413 ( .A1(n9850), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13036) );
  AND2_X1 U11414 ( .A1(n14130), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13043) );
  AND2_X1 U11415 ( .A1(n14119), .A2(n13037), .ZN(n13103) );
  AND2_X1 U11416 ( .A1(n10164), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17158) );
  NAND2_X1 U11417 ( .A1(n18133), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19039) );
  INV_X1 U11418 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14143) );
  AND2_X1 U11419 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14119) );
  INV_X1 U11420 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14077) );
  INV_X1 U11421 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10496) );
  NOR2_X2 U11422 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13044) );
  AND2_X2 U11423 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14132) );
  INV_X2 U11424 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n11308) );
  NOR2_X2 U11425 ( .A1(n11871), .A2(n14877), .ZN(n11891) );
  NAND3_X2 U11426 ( .A1(n10207), .A2(n11064), .A3(n9821), .ZN(n10143) );
  AND2_X4 U11427 ( .A1(n13042), .A2(n14518), .ZN(n13868) );
  NOR2_X2 U11428 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17939), .ZN(n17921) );
  NAND2_X1 U11429 ( .A1(n10689), .A2(n20214), .ZN(n10691) );
  NOR2_X2 U11430 ( .A1(n16113), .A2(n10390), .ZN(n16075) );
  OR2_X1 U11431 ( .A1(n13719), .A2(n16300), .ZN(n10688) );
  INV_X1 U11432 ( .A(n13223), .ZN(n9611) );
  CLKBUF_X1 U11433 ( .A(n9605), .Z(n9614) );
  BUF_X4 U11434 ( .A(n13223), .Z(n14039) );
  CLKBUF_X1 U11435 ( .A(n9605), .Z(n9613) );
  XNOR2_X1 U11437 ( .A(n11101), .B(n10242), .ZN(n9618) );
  INV_X2 U11438 ( .A(n19096), .ZN(n19083) );
  OAI21_X1 U11439 ( .B1(n11307), .B2(n10602), .A(n9873), .ZN(n9872) );
  NAND2_X2 U11440 ( .A1(n9914), .A2(n13229), .ZN(n11307) );
  INV_X2 U11441 ( .A(n9584), .ZN(n9620) );
  NOR2_X2 U11442 ( .A1(n12030), .A2(n11981), .ZN(n12053) );
  NOR2_X2 U11443 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17866), .ZN(n17851) );
  INV_X2 U11445 ( .A(n17183), .ZN(n11244) );
  AND2_X2 U11446 ( .A1(n14712), .A2(n10305), .ZN(n14686) );
  NOR2_X4 U11447 ( .A1(n14740), .A2(n14728), .ZN(n14712) );
  AND2_X1 U11448 ( .A1(n14245), .A2(n14224), .ZN(n9623) );
  NOR2_X4 U11449 ( .A1(n19003), .A2(n19210), .ZN(n18902) );
  AOI22_X4 U11450 ( .A1(n19088), .A2(n19289), .B1(n18970), .B2(n19291), .ZN(
        n19003) );
  NOR2_X2 U11451 ( .A1(n17644), .A2(n12799), .ZN(n12802) );
  NOR2_X2 U11452 ( .A1(n16227), .A2(n10407), .ZN(n14096) );
  NOR4_X2 U11453 ( .A1(n18389), .A2(n18017), .A3(n18034), .A4(n18377), .ZN(
        n18362) );
  NOR2_X2 U11454 ( .A1(n17916), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17887) );
  NOR2_X2 U11455 ( .A1(n11900), .A2(n20981), .ZN(n11931) );
  AND2_X1 U11456 ( .A1(n15040), .A2(n14561), .ZN(n9627) );
  AND2_X4 U11457 ( .A1(n15040), .A2(n14561), .ZN(n21018) );
  INV_X2 U11458 ( .A(n16273), .ZN(n20080) );
  AND2_X2 U11459 ( .A1(n20080), .A2(n20083), .ZN(n16282) );
  NAND2_X1 U11460 ( .A1(n10332), .A2(n9703), .ZN(n12595) );
  NAND2_X1 U11461 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  NAND2_X1 U11462 ( .A1(n10638), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10642) );
  OR2_X1 U11463 ( .A1(n14294), .A2(n21369), .ZN(n11809) );
  OR2_X1 U11464 ( .A1(n10659), .A2(n20808), .ZN(n10464) );
  AND2_X1 U11465 ( .A1(n17224), .A2(n10596), .ZN(n10622) );
  AND4_X1 U11466 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10813) );
  AND2_X1 U11467 ( .A1(n13148), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13974) );
  AOI21_X1 U11468 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19861), .A(
        n13153), .ZN(n13977) );
  NAND3_X1 U11469 ( .A1(n10101), .A2(n15157), .A3(n9932), .ZN(n10337) );
  NAND2_X1 U11470 ( .A1(n10951), .A2(n11555), .ZN(n9811) );
  AND2_X1 U11471 ( .A1(n10456), .A2(n13144), .ZN(n13961) );
  AND2_X1 U11472 ( .A1(n20912), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13679) );
  NAND2_X1 U11473 ( .A1(n16669), .A2(n10041), .ZN(n16604) );
  AND2_X1 U11474 ( .A1(n10042), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10041) );
  NAND2_X1 U11475 ( .A1(n10950), .A2(n13643), .ZN(n13617) );
  NAND3_X1 U11476 ( .A1(n9723), .A2(n10248), .A3(n14222), .ZN(n11658) );
  BUF_X1 U11477 ( .A(n12335), .Z(n12279) );
  AND2_X1 U11478 ( .A1(n11890), .A2(n11889), .ZN(n11895) );
  AND2_X2 U11479 ( .A1(n11572), .A2(n11573), .ZN(n11745) );
  AND2_X2 U11480 ( .A1(n14216), .A2(n14214), .ZN(n12117) );
  OR2_X1 U11481 ( .A1(n14304), .A2(n21369), .ZN(n11810) );
  AND3_X2 U11482 ( .A1(n14304), .A2(n14294), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12397) );
  NAND2_X1 U11483 ( .A1(n10564), .A2(n10625), .ZN(n10602) );
  AND2_X1 U11484 ( .A1(n11553), .A2(n16553), .ZN(n13194) );
  AND2_X1 U11485 ( .A1(n10622), .A2(n10597), .ZN(n10598) );
  AOI21_X1 U11486 ( .B1(n20074), .B2(n11559), .A(n16692), .ZN(n10022) );
  NAND2_X1 U11487 ( .A1(n10612), .A2(n10611), .ZN(n11241) );
  NAND2_X1 U11488 ( .A1(n10132), .A2(n10667), .ZN(n10247) );
  NAND2_X1 U11489 ( .A1(n11207), .A2(n11206), .ZN(n10052) );
  NAND2_X1 U11490 ( .A1(n13942), .A2(n14006), .ZN(n10255) );
  OR2_X1 U11491 ( .A1(n15500), .A2(n21369), .ZN(n12310) );
  NOR2_X1 U11492 ( .A1(n15028), .A2(n10293), .ZN(n10292) );
  INV_X1 U11493 ( .A(n10481), .ZN(n10293) );
  OAI211_X1 U11494 ( .C1(n10327), .C2(n9782), .A(n10102), .B(n10334), .ZN(
        n10338) );
  INV_X1 U11495 ( .A(n10329), .ZN(n10100) );
  NOR2_X1 U11496 ( .A1(n10329), .A2(n10099), .ZN(n10103) );
  AND2_X1 U11497 ( .A1(n9729), .A2(n11659), .ZN(n10294) );
  AND2_X1 U11498 ( .A1(n14568), .A2(n14542), .ZN(n12562) );
  NAND2_X1 U11499 ( .A1(n9908), .A2(n9906), .ZN(n12610) );
  NAND2_X1 U11500 ( .A1(n11770), .A2(n11769), .ZN(n11788) );
  INV_X1 U11501 ( .A(n12397), .ZN(n12387) );
  NAND2_X1 U11502 ( .A1(n15916), .A2(n10400), .ZN(n10399) );
  INV_X1 U11503 ( .A(n11160), .ZN(n10400) );
  NOR2_X2 U11504 ( .A1(n11297), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11304) );
  NAND2_X1 U11505 ( .A1(n10447), .A2(n10446), .ZN(n10450) );
  NOR2_X1 U11506 ( .A1(n13409), .A2(n13435), .ZN(n10447) );
  INV_X1 U11507 ( .A(n16350), .ZN(n10443) );
  NOR2_X1 U11508 ( .A1(n10453), .A2(n10156), .ZN(n10155) );
  NAND2_X1 U11509 ( .A1(n13276), .A2(n16359), .ZN(n10156) );
  NOR2_X1 U11510 ( .A1(n10625), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11323) );
  INV_X1 U11511 ( .A(n13197), .ZN(n16544) );
  NAND2_X1 U11512 ( .A1(n9714), .A2(n9984), .ZN(n9790) );
  INV_X1 U11513 ( .A(n10912), .ZN(n10382) );
  INV_X1 U11514 ( .A(n14351), .ZN(n10354) );
  INV_X1 U11515 ( .A(n14282), .ZN(n11475) );
  AND2_X1 U11516 ( .A1(n10237), .A2(n10139), .ZN(n10138) );
  NOR2_X1 U11517 ( .A1(n10238), .A2(n11338), .ZN(n10237) );
  NOR2_X1 U11518 ( .A1(n9989), .A2(n9914), .ZN(n10066) );
  NOR2_X1 U11519 ( .A1(n13006), .A2(n10194), .ZN(n10193) );
  INV_X1 U11520 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10194) );
  NOR2_X1 U11521 ( .A1(n17308), .A2(n10014), .ZN(n10013) );
  AND2_X1 U11522 ( .A1(n19006), .A2(n9774), .ZN(n10014) );
  NAND2_X1 U11523 ( .A1(n14019), .A2(n14018), .ZN(n14023) );
  NAND2_X1 U11524 ( .A1(n13977), .A2(n13165), .ZN(n13971) );
  NAND2_X1 U11525 ( .A1(n13146), .A2(n13964), .ZN(n14059) );
  INV_X2 U11526 ( .A(n14542), .ZN(n14546) );
  INV_X2 U11527 ( .A(n12346), .ZN(n12352) );
  INV_X1 U11528 ( .A(n14613), .ZN(n10303) );
  NOR2_X1 U11529 ( .A1(n15027), .A2(n15028), .ZN(n14493) );
  OR2_X1 U11530 ( .A1(n17532), .A2(n20927), .ZN(n13724) );
  NAND2_X1 U11531 ( .A1(n15077), .A2(n15069), .ZN(n15068) );
  INV_X1 U11532 ( .A(n12995), .ZN(n10170) );
  NAND2_X1 U11533 ( .A1(n17271), .A2(n13611), .ZN(n13616) );
  NOR2_X1 U11534 ( .A1(n15872), .A2(n15873), .ZN(n15855) );
  AND2_X1 U11535 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  INV_X1 U11536 ( .A(n16014), .ZN(n10340) );
  INV_X1 U11537 ( .A(n10068), .ZN(n9880) );
  AOI21_X1 U11538 ( .B1(n16629), .B2(n20213), .A(n16628), .ZN(n10068) );
  INV_X1 U11539 ( .A(n10216), .ZN(n9917) );
  AND2_X1 U11540 ( .A1(n10357), .A2(n11536), .ZN(n10356) );
  XNOR2_X1 U11541 ( .A(n13192), .B(n10389), .ZN(n13198) );
  NAND2_X1 U11542 ( .A1(n10208), .A2(n16767), .ZN(n10207) );
  AND2_X1 U11543 ( .A1(n16596), .A2(n10466), .ZN(n11064) );
  AOI21_X1 U11544 ( .B1(n9811), .B2(n9808), .A(n9718), .ZN(n9821) );
  NAND2_X1 U11545 ( .A1(n9984), .A2(n10383), .ZN(n9822) );
  NAND2_X1 U11546 ( .A1(n16748), .A2(n10908), .ZN(n16728) );
  AND2_X1 U11547 ( .A1(n10343), .A2(n11337), .ZN(n10342) );
  INV_X1 U11548 ( .A(n16225), .ZN(n10343) );
  NOR2_X1 U11549 ( .A1(n13663), .A2(n13250), .ZN(n13251) );
  INV_X1 U11550 ( .A(n13679), .ZN(n17114) );
  NOR2_X1 U11551 ( .A1(n20876), .A2(n17219), .ZN(n20315) );
  INV_X1 U11552 ( .A(n20881), .ZN(n20906) );
  AND2_X1 U11553 ( .A1(n20876), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20735) );
  OR2_X1 U11554 ( .A1(n20889), .A2(n20251), .ZN(n20673) );
  NAND2_X1 U11555 ( .A1(n20876), .A2(n17219), .ZN(n20627) );
  INV_X1 U11556 ( .A(n13971), .ZN(n19876) );
  NAND2_X1 U11557 ( .A1(n10199), .A2(n18756), .ZN(n10195) );
  NAND2_X1 U11558 ( .A1(n10269), .A2(n10267), .ZN(n10008) );
  NAND2_X1 U11559 ( .A1(n10271), .A2(n10268), .ZN(n10267) );
  AND2_X1 U11560 ( .A1(n10271), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10270) );
  NAND2_X1 U11561 ( .A1(n17317), .A2(n18890), .ZN(n18780) );
  AND4_X1 U11562 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13038), .ZN(
        n13050) );
  AND4_X1 U11563 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        n13049) );
  AND4_X1 U11564 ( .A1(n13030), .A2(n13029), .A3(n13028), .A4(n13027), .ZN(
        n13052) );
  OR2_X2 U11565 ( .A1(n13724), .A2(n17514), .ZN(n20932) );
  OR2_X1 U11566 ( .A1(n13616), .A2(n17677), .ZN(n20908) );
  INV_X1 U11567 ( .A(n20073), .ZN(n16290) );
  AOI21_X1 U11568 ( .B1(n12484), .B2(n20213), .A(n12483), .ZN(n12485) );
  NAND2_X1 U11569 ( .A1(n10047), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9886) );
  NOR2_X1 U11570 ( .A1(n20039), .A2(n19910), .ZN(n20026) );
  INV_X1 U11571 ( .A(n18486), .ZN(n18480) );
  OAI211_X1 U11572 ( .C1(n19116), .C2(n9859), .A(n19397), .B(n9858), .ZN(n9857) );
  NAND2_X1 U11573 ( .A1(n9860), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9859) );
  OR2_X1 U11574 ( .A1(n19111), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9858) );
  NAND2_X1 U11575 ( .A1(n19224), .A2(n19110), .ZN(n9860) );
  NAND2_X1 U11576 ( .A1(n12405), .A2(n12359), .ZN(n9898) );
  AND3_X1 U11577 ( .A1(n10324), .A2(n10322), .A3(n13843), .ZN(n11683) );
  AND2_X1 U11578 ( .A1(n12730), .A2(n12731), .ZN(n10322) );
  AND2_X1 U11579 ( .A1(n13719), .A2(n13666), .ZN(n10689) );
  NAND3_X1 U11580 ( .A1(n10788), .A2(n10787), .A3(n10474), .ZN(n10932) );
  NOR2_X1 U11581 ( .A1(n12385), .A2(n12384), .ZN(n12391) );
  AND2_X1 U11582 ( .A1(n14336), .A2(n11858), .ZN(n10249) );
  OR2_X1 U11583 ( .A1(n11868), .A2(n11867), .ZN(n12565) );
  AND2_X1 U11584 ( .A1(n11620), .A2(n11682), .ZN(n10248) );
  INV_X1 U11585 ( .A(n11686), .ZN(n12410) );
  INV_X1 U11586 ( .A(n11662), .ZN(n12612) );
  AND2_X1 U11587 ( .A1(n11744), .A2(n11742), .ZN(n11725) );
  AOI21_X1 U11588 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17510), .A(
        n12391), .ZN(n12401) );
  NAND2_X1 U11589 ( .A1(n10636), .A2(n12775), .ZN(n9990) );
  NOR2_X1 U11590 ( .A1(n10419), .A2(n10210), .ZN(n10209) );
  INV_X1 U11591 ( .A(n16699), .ZN(n10210) );
  NAND2_X1 U11592 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10161) );
  AND2_X1 U11593 ( .A1(n17176), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10044) );
  AOI21_X1 U11594 ( .B1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n10819), .A(n9688), .ZN(n10028) );
  OAI22_X1 U11595 ( .A1(n20503), .A2(n13303), .B1(n17230), .B2(n17245), .ZN(
        n10038) );
  OAI211_X1 U11596 ( .C1(n13456), .C2(n20378), .A(n10040), .B(n10718), .ZN(
        n10039) );
  NAND2_X1 U11597 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10040) );
  NAND2_X1 U11598 ( .A1(n10130), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10129) );
  AND2_X1 U11599 ( .A1(n10596), .A2(n11297), .ZN(n10574) );
  NAND2_X1 U11600 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10182) );
  OAI211_X1 U11601 ( .C1(n13967), .C2(n13143), .A(n13137), .B(n13136), .ZN(
        n13138) );
  INV_X1 U11602 ( .A(n10255), .ZN(n13940) );
  AND2_X1 U11603 ( .A1(n13158), .A2(n13157), .ZN(n13979) );
  INV_X1 U11604 ( .A(n12240), .ZN(n12211) );
  NAND2_X1 U11605 ( .A1(n12085), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12103) );
  INV_X1 U11606 ( .A(n12084), .ZN(n12085) );
  NOR2_X1 U11607 ( .A1(n12038), .A2(n10085), .ZN(n10084) );
  INV_X1 U11608 ( .A(n14849), .ZN(n10085) );
  XNOR2_X1 U11609 ( .A(n10330), .B(n11877), .ZN(n12508) );
  NAND2_X1 U11610 ( .A1(n14109), .A2(n12538), .ZN(n12546) );
  NOR2_X1 U11611 ( .A1(n14317), .A2(n11775), .ZN(n11791) );
  OR2_X1 U11612 ( .A1(n13818), .A2(n11795), .ZN(n11796) );
  INV_X1 U11613 ( .A(n14837), .ZN(n10317) );
  INV_X1 U11614 ( .A(n14947), .ZN(n12672) );
  INV_X1 U11615 ( .A(n10328), .ZN(n10327) );
  OAI21_X1 U11616 ( .B1(n10329), .B2(n17571), .A(n12580), .ZN(n10328) );
  NAND2_X1 U11617 ( .A1(n17577), .A2(n12560), .ZN(n10104) );
  NAND2_X1 U11618 ( .A1(n11834), .A2(n9933), .ZN(n12554) );
  AND2_X1 U11619 ( .A1(n14336), .A2(n9934), .ZN(n9933) );
  AND2_X1 U11620 ( .A1(n9735), .A2(n11858), .ZN(n9934) );
  AND2_X1 U11622 ( .A1(n14546), .A2(n14304), .ZN(n11685) );
  AND2_X1 U11623 ( .A1(n10248), .A2(n9723), .ZN(n11680) );
  NAND2_X1 U11624 ( .A1(n11664), .A2(n14304), .ZN(n12637) );
  OAI21_X1 U11625 ( .B1(n12620), .B2(n20927), .A(n9892), .ZN(n9896) );
  INV_X1 U11626 ( .A(n9893), .ZN(n9892) );
  OAI21_X1 U11627 ( .B1(n12619), .B2(n20927), .A(n15176), .ZN(n9893) );
  OR2_X1 U11628 ( .A1(n11766), .A2(n11765), .ZN(n12531) );
  OR2_X1 U11629 ( .A1(n11756), .A2(n11755), .ZN(n12572) );
  OR3_X1 U11630 ( .A1(n11788), .A2(n11774), .A3(n11773), .ZN(n11780) );
  OAI211_X1 U11631 ( .C1(n17525), .C2(n21203), .A(n11704), .B(n11703), .ZN(
        n11706) );
  NAND2_X1 U11632 ( .A1(n11663), .A2(n14317), .ZN(n11657) );
  INV_X1 U11633 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14233) );
  AOI221_X1 U11634 ( .B1(n21468), .B2(n15520), .C1(n17632), .C2(n15520), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n15533) );
  INV_X1 U11635 ( .A(n10169), .ZN(n12621) );
  INV_X1 U11636 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21203) );
  NOR2_X1 U11637 ( .A1(n17205), .A2(n10595), .ZN(n10565) );
  AND2_X1 U11638 ( .A1(n10369), .A2(n11088), .ZN(n10368) );
  NOR2_X1 U11639 ( .A1(n11082), .A2(n10370), .ZN(n10369) );
  NAND2_X1 U11640 ( .A1(n16687), .A2(n10232), .ZN(n10231) );
  NAND2_X1 U11641 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  INV_X1 U11642 ( .A(n10966), .ZN(n10377) );
  NOR2_X1 U11643 ( .A1(n16061), .A2(n16042), .ZN(n10413) );
  NOR2_X1 U11644 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13367) );
  NOR2_X1 U11645 ( .A1(n10707), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10803) );
  AOI211_X1 U11646 ( .C1(n13506), .C2(n13503), .A(n14094), .B(n13544), .ZN(
        n13504) );
  NAND2_X1 U11647 ( .A1(n10452), .A2(n16338), .ZN(n10449) );
  NAND2_X1 U11648 ( .A1(n10454), .A2(n16363), .ZN(n10453) );
  NOR2_X1 U11649 ( .A1(n16372), .A2(n16367), .ZN(n10454) );
  NAND2_X1 U11650 ( .A1(n10624), .A2(n10625), .ZN(n9989) );
  NOR2_X1 U11651 ( .A1(n16576), .A2(n12814), .ZN(n10297) );
  NOR2_X1 U11652 ( .A1(n16760), .A2(n10301), .ZN(n10300) );
  NAND2_X1 U11653 ( .A1(n10243), .A2(n10657), .ZN(n11101) );
  NAND2_X1 U11654 ( .A1(n13192), .A2(n9781), .ZN(n9982) );
  OR2_X1 U11655 ( .A1(n15894), .A2(n11555), .ZN(n13197) );
  AOI21_X1 U11656 ( .B1(n11550), .B2(n11551), .A(n13195), .ZN(n16545) );
  NAND2_X1 U11657 ( .A1(n10349), .A2(n10348), .ZN(n10347) );
  INV_X1 U11658 ( .A(n15963), .ZN(n10348) );
  INV_X1 U11659 ( .A(n15983), .ZN(n10349) );
  NOR2_X1 U11660 ( .A1(n11277), .A2(n10056), .ZN(n10055) );
  INV_X1 U11661 ( .A(n11276), .ZN(n10056) );
  OR2_X1 U11662 ( .A1(n16094), .A2(n11555), .ZN(n11072) );
  NAND2_X1 U11663 ( .A1(n10394), .A2(n11125), .ZN(n10393) );
  INV_X1 U11664 ( .A(n16101), .ZN(n10394) );
  INV_X1 U11665 ( .A(n14260), .ZN(n11416) );
  AND2_X1 U11666 ( .A1(n11115), .A2(n16190), .ZN(n10410) );
  NAND2_X1 U11667 ( .A1(n9943), .A2(n9942), .ZN(n10908) );
  NOR2_X1 U11668 ( .A1(n11555), .A2(n17024), .ZN(n9942) );
  NAND2_X1 U11669 ( .A1(n10850), .A2(n9604), .ZN(n10851) );
  NAND2_X1 U11670 ( .A1(n9980), .A2(n9979), .ZN(n9978) );
  NAND2_X1 U11671 ( .A1(n20273), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U11672 ( .A1(n10960), .A2(n9914), .ZN(n9980) );
  OAI21_X1 U11673 ( .B1(n11342), .B2(n20808), .A(n11313), .ZN(n11317) );
  CLKBUF_X1 U11674 ( .A(n10624), .Z(n13254) );
  NAND2_X1 U11675 ( .A1(n10665), .A2(n10664), .ZN(n10414) );
  CLKBUF_X1 U11676 ( .A(n10708), .Z(n10709) );
  NAND2_X1 U11677 ( .A1(n20912), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U11678 ( .A1(n10051), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U11679 ( .A1(n10052), .A2(n11210), .ZN(n10051) );
  CLKBUF_X1 U11680 ( .A(n11242), .Z(n11243) );
  NOR2_X2 U11681 ( .A1(n10691), .A2(n14039), .ZN(n20436) );
  AOI22_X1 U11682 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10519) );
  INV_X1 U11683 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n17256) );
  NAND2_X1 U11684 ( .A1(n9911), .A2(n10499), .ZN(n9910) );
  XNOR2_X1 U11685 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10928) );
  NOR2_X1 U11686 ( .A1(n13135), .A2(n13132), .ZN(n13145) );
  NOR2_X1 U11687 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  AND2_X1 U11688 ( .A1(n13043), .A2(n14131), .ZN(n13859) );
  NOR2_X1 U11689 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13037) );
  INV_X1 U11690 ( .A(n10261), .ZN(n10260) );
  INV_X1 U11691 ( .A(n19438), .ZN(n13130) );
  NAND2_X1 U11692 ( .A1(n9855), .A2(n17338), .ZN(n19008) );
  XNOR2_X1 U11693 ( .A(n17335), .B(n17339), .ZN(n9855) );
  NAND2_X1 U11694 ( .A1(n19036), .A2(n13952), .ZN(n13954) );
  OR2_X1 U11695 ( .A1(n19346), .A2(n13939), .ZN(n13952) );
  INV_X1 U11696 ( .A(n14011), .ZN(n14019) );
  INV_X1 U11697 ( .A(n19066), .ZN(n9998) );
  INV_X1 U11698 ( .A(n14004), .ZN(n9999) );
  NAND2_X1 U11699 ( .A1(n19063), .A2(n13948), .ZN(n13949) );
  AOI21_X1 U11700 ( .B1(n14059), .B2(n14058), .A(n14064), .ZN(n14087) );
  NOR2_X1 U11701 ( .A1(n14060), .A2(n19879), .ZN(n14085) );
  NOR2_X1 U11702 ( .A1(n14304), .A2(n14542), .ZN(n14235) );
  OR2_X1 U11703 ( .A1(n14209), .A2(n14208), .ZN(n14429) );
  AND2_X1 U11704 ( .A1(n11684), .A2(n11659), .ZN(n12856) );
  AND2_X1 U11705 ( .A1(n14304), .A2(n14542), .ZN(n13829) );
  OAI21_X1 U11706 ( .B1(n9891), .B2(n9890), .A(n11784), .ZN(n14079) );
  AND2_X1 U11707 ( .A1(n12856), .A2(n9625), .ZN(n13842) );
  OR4_X1 U11708 ( .A1(n17532), .A2(n14546), .A3(n11674), .A4(n21467), .ZN(
        n12408) );
  NOR2_X1 U11709 ( .A1(n14687), .A2(n12984), .ZN(n14664) );
  NOR2_X1 U11710 ( .A1(n14687), .A2(n12854), .ZN(n14663) );
  OR2_X1 U11711 ( .A1(n15142), .A2(n12295), .ZN(n12109) );
  NAND2_X1 U11712 ( .A1(n14846), .A2(n9757), .ZN(n14740) );
  NAND2_X1 U11713 ( .A1(n12053), .A2(n12052), .ZN(n12067) );
  AND2_X1 U11714 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12052) );
  OR2_X1 U11715 ( .A1(n14936), .A2(n14935), .ZN(n14938) );
  NAND2_X1 U11716 ( .A1(n11852), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11871) );
  AND2_X1 U11717 ( .A1(n14608), .A2(n14609), .ZN(n14611) );
  AND2_X1 U11718 ( .A1(n14640), .A2(n14629), .ZN(n14608) );
  NAND2_X1 U11719 ( .A1(n9923), .A2(n12765), .ZN(n9922) );
  NAND2_X1 U11720 ( .A1(n14696), .A2(n9765), .ZN(n14653) );
  INV_X1 U11721 ( .A(n14651), .ZN(n10319) );
  NOR2_X1 U11722 ( .A1(n14653), .A2(n14638), .ZN(n14640) );
  NAND2_X1 U11723 ( .A1(n12991), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10178) );
  NOR2_X1 U11724 ( .A1(n15334), .A2(n9904), .ZN(n15321) );
  AND2_X1 U11725 ( .A1(n21127), .A2(n15323), .ZN(n9904) );
  NAND2_X1 U11726 ( .A1(n15471), .A2(n9905), .ZN(n15339) );
  OR2_X1 U11727 ( .A1(n15376), .A2(n15353), .ZN(n9905) );
  NAND2_X1 U11728 ( .A1(n14773), .A2(n9702), .ZN(n14716) );
  INV_X1 U11729 ( .A(n14714), .ZN(n10321) );
  INV_X1 U11730 ( .A(n21130), .ZN(n15468) );
  AND2_X1 U11731 ( .A1(n17612), .A2(n10312), .ZN(n14957) );
  AND2_X1 U11732 ( .A1(n10314), .A2(n10313), .ZN(n10312) );
  INV_X1 U11733 ( .A(n14959), .ZN(n10313) );
  NOR2_X1 U11734 ( .A1(n13847), .A2(n12744), .ZN(n14220) );
  NAND2_X1 U11735 ( .A1(n12418), .A2(n11675), .ZN(n12624) );
  NAND2_X1 U11736 ( .A1(n9894), .A2(n13624), .ZN(n12749) );
  BUF_X1 U11737 ( .A(n12512), .Z(n15526) );
  OR2_X1 U11738 ( .A1(n21170), .A2(n15805), .ZN(n15540) );
  OR2_X2 U11739 ( .A1(n11590), .A2(n11589), .ZN(n14568) );
  NOR2_X1 U11741 ( .A1(n15560), .A2(n15527), .ZN(n21199) );
  NOR2_X2 U11742 ( .A1(n14974), .A2(n15264), .ZN(n14329) );
  NOR2_X1 U11743 ( .A1(n15560), .A2(n15559), .ZN(n15802) );
  INV_X1 U11744 ( .A(n15533), .ZN(n15642) );
  AND2_X1 U11745 ( .A1(n15560), .A2(n15527), .ZN(n15597) );
  INV_X1 U11746 ( .A(n15562), .ZN(n14400) );
  NAND2_X1 U11747 ( .A1(n11557), .A2(n11556), .ZN(n12501) );
  NAND2_X1 U11748 ( .A1(n15899), .A2(n16330), .ZN(n13189) );
  AND2_X1 U11749 ( .A1(n16005), .A2(n15999), .ZN(n15970) );
  INV_X1 U11750 ( .A(n16020), .ZN(n16017) );
  NOR2_X1 U11751 ( .A1(n16136), .A2(n10229), .ZN(n16090) );
  AND2_X1 U11752 ( .A1(n20273), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10966) );
  OR2_X1 U11753 ( .A1(n10965), .A2(n10966), .ZN(n11015) );
  AND2_X1 U11754 ( .A1(n10398), .A2(n15933), .ZN(n10395) );
  NOR2_X1 U11755 ( .A1(n15885), .A2(n10399), .ZN(n10398) );
  NAND2_X1 U11756 ( .A1(n14092), .A2(n10150), .ZN(n16375) );
  AND2_X1 U11757 ( .A1(n10151), .A2(n16383), .ZN(n10150) );
  AND2_X1 U11758 ( .A1(n13263), .A2(n10152), .ZN(n10151) );
  INV_X1 U11759 ( .A(n16387), .ZN(n10152) );
  OR2_X1 U11760 ( .A1(n13432), .A2(n9760), .ZN(n10440) );
  NAND2_X1 U11761 ( .A1(n9760), .A2(n13432), .ZN(n10441) );
  NOR2_X1 U11762 ( .A1(n17266), .A2(n16324), .ZN(n13676) );
  INV_X1 U11763 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16576) );
  NOR2_X1 U11764 ( .A1(n10290), .A2(n10287), .ZN(n10285) );
  INV_X1 U11765 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U11766 ( .A1(n11123), .A2(n9666), .ZN(n11124) );
  OR2_X1 U11767 ( .A1(n12493), .A2(n10048), .ZN(n10047) );
  AND2_X1 U11768 ( .A1(n20236), .A2(n12494), .ZN(n10048) );
  OAI21_X1 U11769 ( .B1(n15848), .B2(n11538), .A(n12492), .ZN(n13583) );
  NOR2_X1 U11770 ( .A1(n10384), .A2(n9864), .ZN(n9863) );
  INV_X1 U11771 ( .A(n10914), .ZN(n9864) );
  INV_X1 U11772 ( .A(n13198), .ZN(n10362) );
  NAND2_X1 U11773 ( .A1(n9987), .A2(n10389), .ZN(n9986) );
  NAND2_X1 U11774 ( .A1(n15897), .A2(n10359), .ZN(n15865) );
  XNOR2_X1 U11775 ( .A(n11552), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11549) );
  AND2_X1 U11776 ( .A1(n11513), .A2(n11512), .ZN(n16047) );
  NAND2_X1 U11777 ( .A1(n12495), .A2(n10090), .ZN(n10089) );
  INV_X1 U11778 ( .A(n12449), .ZN(n10090) );
  NOR2_X1 U11779 ( .A1(n10353), .A2(n10351), .ZN(n10350) );
  INV_X1 U11780 ( .A(n16059), .ZN(n10351) );
  NOR2_X1 U11781 ( .A1(n10089), .A2(n16961), .ZN(n9938) );
  AND3_X1 U11782 ( .A1(n11491), .A2(n11490), .A3(n11489), .ZN(n14351) );
  INV_X1 U11783 ( .A(n9960), .ZN(n9959) );
  OAI21_X1 U11784 ( .B1(n10418), .B2(n9961), .A(n16671), .ZN(n9960) );
  INV_X1 U11785 ( .A(n12451), .ZN(n9961) );
  NAND2_X1 U11786 ( .A1(n9811), .A2(n9809), .ZN(n9806) );
  NOR2_X1 U11787 ( .A1(n16720), .A2(n11274), .ZN(n9918) );
  INV_X1 U11788 ( .A(n16727), .ZN(n9919) );
  NOR2_X2 U11789 ( .A1(n16163), .A2(n16145), .ZN(n16147) );
  NOR2_X1 U11790 ( .A1(n17087), .A2(n10057), .ZN(n17015) );
  NAND2_X1 U11791 ( .A1(n9719), .A2(n10061), .ZN(n10057) );
  NAND2_X1 U11792 ( .A1(n11116), .A2(n9671), .ZN(n11117) );
  NAND2_X1 U11793 ( .A1(n9883), .A2(n9935), .ZN(n9792) );
  NAND2_X1 U11794 ( .A1(n9870), .A2(n9705), .ZN(n9831) );
  OAI21_X1 U11795 ( .B1(n17105), .B2(n10214), .A(n10212), .ZN(n10999) );
  AND3_X1 U11796 ( .A1(n11336), .A2(n11335), .A3(n11334), .ZN(n16245) );
  INV_X1 U11797 ( .A(n20315), .ZN(n20433) );
  NOR2_X1 U11798 ( .A1(n20673), .A2(n20433), .ZN(n20437) );
  NOR2_X1 U11799 ( .A1(n20520), .A2(n20881), .ZN(n9869) );
  CLKBUF_X1 U11800 ( .A(n13229), .Z(n13230) );
  NAND2_X1 U11801 ( .A1(n20916), .A2(n17115), .ZN(n17116) );
  NAND2_X1 U11802 ( .A1(n17668), .A2(n20912), .ZN(n17117) );
  AND2_X1 U11803 ( .A1(n17264), .A2(n10945), .ZN(n13611) );
  NAND2_X1 U11804 ( .A1(n13129), .A2(n9975), .ZN(n9972) );
  NAND2_X1 U11805 ( .A1(n9974), .A2(n19442), .ZN(n9973) );
  NAND2_X1 U11806 ( .A1(n18620), .A2(n9975), .ZN(n9974) );
  NAND2_X1 U11807 ( .A1(n13985), .A2(n13145), .ZN(n17806) );
  INV_X1 U11808 ( .A(n19922), .ZN(n20027) );
  INV_X1 U11809 ( .A(n17328), .ZN(n19879) );
  NAND2_X1 U11810 ( .A1(n13026), .A2(n13025), .ZN(n17841) );
  INV_X1 U11811 ( .A(n10197), .ZN(n10196) );
  OAI21_X1 U11812 ( .B1(n10198), .B2(n17862), .A(n10198), .ZN(n10197) );
  NAND2_X1 U11813 ( .A1(n13021), .A2(n13020), .ZN(n17872) );
  INV_X1 U11814 ( .A(n18768), .ZN(n13020) );
  NAND2_X1 U11815 ( .A1(n10202), .A2(n9708), .ZN(n17934) );
  NAND2_X1 U11816 ( .A1(n9656), .A2(n17936), .ZN(n10203) );
  NAND2_X1 U11817 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  INV_X1 U11818 ( .A(n18846), .ZN(n10204) );
  INV_X1 U11819 ( .A(n17945), .ZN(n10205) );
  OR2_X1 U11820 ( .A1(n13936), .A2(n13935), .ZN(n14024) );
  OR2_X1 U11821 ( .A1(n13926), .A2(n13925), .ZN(n14017) );
  NOR2_X1 U11822 ( .A1(n18812), .A2(n18822), .ZN(n18797) );
  INV_X1 U11823 ( .A(n18855), .ZN(n10192) );
  NAND2_X1 U11824 ( .A1(n10005), .A2(n10004), .ZN(n17319) );
  AND2_X1 U11825 ( .A1(n18780), .A2(n10006), .ZN(n10005) );
  NAND2_X1 U11826 ( .A1(n18890), .A2(n10007), .ZN(n10006) );
  OAI211_X1 U11827 ( .C1(n18952), .C2(n10012), .A(n17312), .B(n10011), .ZN(
        n17315) );
  NAND2_X1 U11828 ( .A1(n18952), .A2(n19006), .ZN(n10010) );
  NAND2_X1 U11829 ( .A1(n10256), .A2(n10261), .ZN(n18918) );
  INV_X1 U11830 ( .A(n13147), .ZN(n13960) );
  NAND2_X1 U11831 ( .A1(n19006), .A2(n10273), .ZN(n10272) );
  XNOR2_X1 U11832 ( .A(n14003), .B(n19367), .ZN(n19067) );
  AND2_X1 U11833 ( .A1(n19876), .A2(n13984), .ZN(n19873) );
  OAI21_X1 U11834 ( .B1(n12862), .B2(n14960), .A(n12863), .ZN(n12864) );
  CLKBUF_X1 U11835 ( .A(n12433), .Z(n15006) );
  OAI21_X1 U11836 ( .B1(n15310), .B2(n20932), .A(n10080), .ZN(n10079) );
  INV_X1 U11837 ( .A(n15083), .ZN(n10080) );
  OR2_X1 U11838 ( .A1(n14634), .A2(n14637), .ZN(n10077) );
  OR2_X1 U11839 ( .A1(n15320), .A2(n20932), .ZN(n13003) );
  OAI21_X1 U11840 ( .B1(n14831), .B2(n14811), .A(n14936), .ZN(n15209) );
  AND2_X2 U11841 ( .A1(n20932), .A2(n12997), .ZN(n21094) );
  INV_X1 U11842 ( .A(n15264), .ZN(n21101) );
  AND2_X1 U11843 ( .A1(n10114), .A2(n10113), .ZN(n12598) );
  NAND2_X1 U11844 ( .A1(n15034), .A2(n12596), .ZN(n10113) );
  AND2_X1 U11845 ( .A1(n15434), .A2(n15342), .ZN(n21130) );
  NAND2_X1 U11846 ( .A1(n15423), .A2(n17600), .ZN(n17591) );
  OR2_X1 U11847 ( .A1(n21134), .A2(n15467), .ZN(n15423) );
  AND2_X1 U11848 ( .A1(n15803), .A2(n15802), .ZN(n21363) );
  INV_X1 U11849 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21400) );
  AND2_X1 U11850 ( .A1(n15860), .A2(n16290), .ZN(n15861) );
  NOR2_X1 U11851 ( .A1(n15859), .A2(n16538), .ZN(n10236) );
  AND2_X1 U11852 ( .A1(n12843), .A2(n12842), .ZN(n20072) );
  OAI21_X1 U11853 ( .B1(n16267), .B2(n20200), .A(n10309), .ZN(n10308) );
  AOI21_X1 U11854 ( .B1(n17168), .B2(n16301), .A(n10310), .ZN(n10309) );
  OAI21_X1 U11855 ( .B1(n20887), .B2(n20077), .A(n10311), .ZN(n10310) );
  XNOR2_X1 U11856 ( .A(n12492), .B(n12491), .ZN(n16424) );
  NAND2_X1 U11857 ( .A1(n20178), .A2(n20909), .ZN(n20145) );
  OAI21_X1 U11858 ( .B1(n16543), .B2(n9843), .A(n9842), .ZN(n9834) );
  NAND2_X1 U11859 ( .A1(n11188), .A2(n9775), .ZN(n11189) );
  XNOR2_X1 U11860 ( .A(n9866), .B(n12494), .ZN(n12445) );
  NAND2_X1 U11861 ( .A1(n9987), .A2(n9795), .ZN(n16809) );
  NAND2_X1 U11862 ( .A1(n16543), .A2(n16805), .ZN(n9795) );
  INV_X1 U11863 ( .A(n16318), .ZN(n16808) );
  NAND2_X1 U11864 ( .A1(n16627), .A2(n16615), .ZN(n9820) );
  NOR2_X1 U11865 ( .A1(n16614), .A2(n16773), .ZN(n9819) );
  NOR2_X1 U11866 ( .A1(n9880), .A2(n10403), .ZN(n9879) );
  NOR2_X1 U11867 ( .A1(n9880), .A2(n9778), .ZN(n9876) );
  AND2_X1 U11868 ( .A1(n10094), .A2(n16626), .ZN(n9882) );
  NOR2_X1 U11869 ( .A1(n9880), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9877) );
  NAND2_X1 U11870 ( .A1(n13617), .A2(n11161), .ZN(n17654) );
  AND2_X1 U11871 ( .A1(n17654), .A2(n17120), .ZN(n20213) );
  INV_X1 U11872 ( .A(n20213), .ZN(n20194) );
  INV_X1 U11873 ( .A(n17654), .ZN(n20204) );
  XNOR2_X1 U11874 ( .A(n9817), .B(n12505), .ZN(n16531) );
  NOR2_X1 U11875 ( .A1(n15845), .A2(n11555), .ZN(n12504) );
  NAND2_X1 U11876 ( .A1(n9841), .A2(n9835), .ZN(n9844) );
  NAND2_X1 U11877 ( .A1(n16543), .A2(n9833), .ZN(n9841) );
  INV_X1 U11878 ( .A(n9836), .ZN(n9835) );
  NOR2_X1 U11879 ( .A1(n20219), .A2(n12779), .ZN(n9833) );
  INV_X1 U11880 ( .A(n16424), .ZN(n10016) );
  XNOR2_X1 U11881 ( .A(n9916), .B(n11561), .ZN(n12444) );
  OAI21_X1 U11882 ( .B1(n11087), .B2(n10217), .A(n9917), .ZN(n9916) );
  INV_X1 U11883 ( .A(n12445), .ZN(n9865) );
  INV_X1 U11884 ( .A(n16809), .ZN(n9789) );
  NAND2_X1 U11885 ( .A1(n11087), .A2(n11086), .ZN(n16566) );
  NAND2_X1 U11886 ( .A1(n9862), .A2(n16571), .ZN(n16852) );
  OAI21_X1 U11887 ( .B1(n10143), .B2(n10142), .A(n10140), .ZN(n16575) );
  NAND2_X1 U11888 ( .A1(n9945), .A2(n16581), .ZN(n16864) );
  NAND2_X1 U11889 ( .A1(n9946), .A2(n11279), .ZN(n9945) );
  NAND2_X1 U11890 ( .A1(n16604), .A2(n16603), .ZN(n10135) );
  INV_X1 U11891 ( .A(n16602), .ZN(n10136) );
  OAI211_X1 U11892 ( .C1(n9952), .C2(n9739), .A(n9949), .B(n9947), .ZN(n16898)
         );
  OR2_X1 U11893 ( .A1(n9950), .A2(n9739), .ZN(n9949) );
  NAND2_X1 U11894 ( .A1(n9952), .A2(n9948), .ZN(n9947) );
  NAND2_X1 U11895 ( .A1(n16641), .A2(n9953), .ZN(n9952) );
  NAND2_X1 U11896 ( .A1(n9603), .A2(n10402), .ZN(n16627) );
  OAI21_X1 U11897 ( .B1(n16913), .B2(n10094), .A(n16626), .ZN(n9881) );
  NAND2_X1 U11898 ( .A1(n10088), .A2(n10087), .ZN(n10092) );
  AOI21_X1 U11899 ( .B1(n9652), .B2(n10089), .A(n10093), .ZN(n10087) );
  NAND2_X1 U11900 ( .A1(n16583), .A2(n9652), .ZN(n10088) );
  NAND2_X1 U11901 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10094), .ZN(
        n10093) );
  NAND2_X1 U11902 ( .A1(n16691), .A2(n16978), .ZN(n16973) );
  AND2_X1 U11903 ( .A1(n11563), .A2(n11262), .ZN(n17090) );
  INV_X1 U11904 ( .A(n17090), .ZN(n20242) );
  AND2_X1 U11905 ( .A1(n11563), .A2(n20902), .ZN(n17661) );
  AND2_X1 U11906 ( .A1(n10148), .A2(n13252), .ZN(n13718) );
  AND2_X2 U11907 ( .A1(n14033), .A2(n14037), .ZN(n20876) );
  INV_X1 U11908 ( .A(n14034), .ZN(n14036) );
  AND2_X1 U11909 ( .A1(n20462), .A2(n20461), .ZN(n20501) );
  NAND2_X1 U11910 ( .A1(n17833), .A2(n18170), .ZN(n17845) );
  AND2_X1 U11911 ( .A1(n9825), .A2(n17848), .ZN(n9824) );
  OR2_X1 U11912 ( .A1(n17849), .A2(n19991), .ZN(n9825) );
  NAND2_X1 U11913 ( .A1(n17847), .A2(n19991), .ZN(n9826) );
  NAND2_X1 U11914 ( .A1(n17870), .A2(n17867), .ZN(n17866) );
  INV_X1 U11915 ( .A(n18185), .ZN(n18170) );
  NAND2_X1 U11916 ( .A1(n18480), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n18482) );
  NAND2_X1 U11917 ( .A1(n18500), .A2(n9649), .ZN(n18486) );
  INV_X1 U11918 ( .A(n18576), .ZN(n18615) );
  AND2_X1 U11919 ( .A1(n14103), .A2(n9967), .ZN(n18612) );
  INV_X1 U11920 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19895) );
  XNOR2_X1 U11921 ( .A(n10279), .B(n17679), .ZN(n17684) );
  NAND2_X1 U11922 ( .A1(n17537), .A2(n17536), .ZN(n10279) );
  NAND2_X1 U11923 ( .A1(n17496), .A2(n17696), .ZN(n10263) );
  AND2_X1 U11924 ( .A1(n10262), .A2(n17703), .ZN(n10002) );
  OR2_X1 U11925 ( .A1(n17497), .A2(n17538), .ZN(n10262) );
  OR2_X1 U11926 ( .A1(n17541), .A2(n17696), .ZN(n10264) );
  AOI21_X1 U11927 ( .B1(n19105), .B2(n19878), .A(n9851), .ZN(n19108) );
  INV_X1 U11928 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20039) );
  NAND2_X1 U11929 ( .A1(n19390), .A2(n19400), .ZN(n19384) );
  INV_X1 U11930 ( .A(n19384), .ZN(n19392) );
  OR2_X1 U11931 ( .A1(n19875), .A2(n19390), .ZN(n19404) );
  AND2_X1 U11932 ( .A1(n9897), .A2(n12360), .ZN(n12366) );
  NAND2_X1 U11933 ( .A1(n12377), .A2(n10167), .ZN(n12360) );
  INV_X1 U11934 ( .A(n10168), .ZN(n10167) );
  INV_X1 U11935 ( .A(n11259), .ZN(n10638) );
  OAI21_X1 U11936 ( .B1(n17246), .B2(n17256), .A(n10639), .ZN(n10640) );
  CLKBUF_X1 U11937 ( .A(n12323), .Z(n12300) );
  AND2_X1 U11938 ( .A1(n11658), .A2(n11721), .ZN(n11656) );
  AOI22_X1 U11939 ( .A1(n20726), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10819), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10820) );
  OAI22_X1 U11940 ( .A1(n11437), .A2(n13323), .B1(n10804), .B2(n9981), .ZN(
        n10805) );
  INV_X1 U11941 ( .A(n10803), .ZN(n9981) );
  NAND2_X1 U11942 ( .A1(n9799), .A2(n9798), .ZN(n10436) );
  NOR2_X1 U11943 ( .A1(n16324), .A2(n20809), .ZN(n9798) );
  AND2_X1 U11944 ( .A1(n16300), .A2(n10685), .ZN(n10668) );
  NAND2_X1 U11945 ( .A1(n12383), .A2(n12382), .ZN(n12385) );
  XNOR2_X1 U11946 ( .A(n11823), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12384) );
  CLKBUF_X1 U11947 ( .A(n12330), .Z(n12262) );
  INV_X1 U11949 ( .A(n12581), .ZN(n10325) );
  INV_X1 U11950 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U11951 ( .A1(n11630), .A2(n12609), .ZN(n11631) );
  AND2_X1 U11952 ( .A1(n9907), .A2(n12406), .ZN(n9906) );
  INV_X1 U11953 ( .A(n11809), .ZN(n11767) );
  INV_X1 U11954 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11694) );
  OR2_X1 U11955 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  NAND2_X1 U11956 ( .A1(n11803), .A2(n10097), .ZN(n11833) );
  CLKBUF_X1 U11957 ( .A(n11698), .Z(n11699) );
  INV_X1 U11958 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11567) );
  OR2_X1 U11959 ( .A1(n11820), .A2(n11819), .ZN(n12518) );
  NOR2_X1 U11960 ( .A1(n12363), .A2(n12405), .ZN(n12396) );
  NAND2_X1 U11961 ( .A1(n10699), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10512) );
  NAND2_X1 U11962 ( .A1(n10601), .A2(n11244), .ZN(n11194) );
  INV_X1 U11963 ( .A(n10882), .ZN(n9814) );
  NOR2_X1 U11964 ( .A1(n9940), .A2(n11555), .ZN(n9939) );
  INV_X1 U11965 ( .A(n10883), .ZN(n9940) );
  AOI21_X1 U11966 ( .B1(n10816), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(n9685), .ZN(n10858) );
  NAND2_X1 U11967 ( .A1(n20273), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U11968 ( .A1(n10955), .A2(n9914), .ZN(n10957) );
  INV_X1 U11969 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13233) );
  INV_X1 U11970 ( .A(n10932), .ZN(n11320) );
  NAND2_X1 U11971 ( .A1(n9697), .A2(n10632), .ZN(n10241) );
  OAI21_X1 U11972 ( .B1(n10652), .B2(n10628), .A(n10487), .ZN(n10629) );
  AND2_X1 U11973 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14044) );
  AND2_X1 U11974 ( .A1(n10694), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10947) );
  AOI22_X1 U11975 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10573) );
  AND2_X1 U11976 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10501) );
  AOI21_X1 U11977 ( .B1(n10706), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10500) );
  AND2_X1 U11978 ( .A1(n20679), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10925) );
  INV_X2 U11979 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10926) );
  OAI21_X1 U11980 ( .B1(n10932), .B2(n11192), .A(n10931), .ZN(n10955) );
  NAND2_X1 U11981 ( .A1(n11192), .A2(n11201), .ZN(n10931) );
  NAND2_X1 U11982 ( .A1(n14090), .A2(n9854), .ZN(n13942) );
  NOR2_X1 U11983 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12392), .ZN(
        n12415) );
  AND2_X1 U11984 ( .A1(n14700), .A2(n12128), .ZN(n10305) );
  NOR2_X1 U11985 ( .A1(n10083), .A2(n9766), .ZN(n10082) );
  INV_X1 U11986 ( .A(n10084), .ZN(n10083) );
  NOR2_X1 U11987 ( .A1(n14848), .A2(n14807), .ZN(n14808) );
  OAI21_X1 U11988 ( .B1(n12530), .B2(n14546), .A(n12529), .ZN(n12537) );
  AOI21_X1 U11989 ( .B1(n15116), .B2(n10334), .A(n10251), .ZN(n10250) );
  INV_X1 U11990 ( .A(n10252), .ZN(n10251) );
  AOI21_X1 U11991 ( .B1(n10334), .B2(n9647), .A(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10252) );
  INV_X1 U11992 ( .A(n14676), .ZN(n10320) );
  NAND2_X1 U11993 ( .A1(n12585), .A2(n9660), .ZN(n15168) );
  INV_X1 U11994 ( .A(n14948), .ZN(n10318) );
  INV_X1 U11995 ( .A(n12714), .ZN(n12711) );
  AND2_X1 U11996 ( .A1(n10473), .A2(n17611), .ZN(n10314) );
  AND2_X1 U11997 ( .A1(n13829), .A2(n12626), .ZN(n12714) );
  NAND2_X1 U11998 ( .A1(n10175), .A2(n12746), .ZN(n10174) );
  AND2_X1 U11999 ( .A1(n12523), .A2(n12747), .ZN(n10173) );
  AOI21_X1 U12000 ( .B1(n12548), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12550) );
  NAND2_X1 U12001 ( .A1(n10105), .A2(n12511), .ZN(n12551) );
  NAND2_X1 U12002 ( .A1(n12508), .A2(n12562), .ZN(n10105) );
  NAND2_X1 U12003 ( .A1(n11664), .A2(n12609), .ZN(n14222) );
  AND2_X1 U12004 ( .A1(n12410), .A2(n12409), .ZN(n12737) );
  AND4_X1 U12005 ( .A1(n11608), .A2(n11607), .A3(n11606), .A4(n11605), .ZN(
        n11609) );
  NAND2_X1 U12006 ( .A1(n11727), .A2(n11726), .ZN(n21169) );
  INV_X1 U12007 ( .A(n11725), .ZN(n11726) );
  INV_X1 U12008 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U12009 ( .A1(n10620), .A2(n17183), .ZN(n10604) );
  NAND2_X1 U12010 ( .A1(n9643), .A2(n10379), .ZN(n10378) );
  INV_X1 U12011 ( .A(n11040), .ZN(n10379) );
  NOR2_X1 U12012 ( .A1(n11045), .A2(n9758), .ZN(n10381) );
  NAND2_X1 U12013 ( .A1(n10230), .A2(n16678), .ZN(n10229) );
  INV_X1 U12014 ( .A(n10231), .ZN(n10230) );
  INV_X1 U12015 ( .A(n11051), .ZN(n9977) );
  NAND2_X1 U12016 ( .A1(n10372), .A2(n16404), .ZN(n10371) );
  INV_X1 U12017 ( .A(n10373), .ZN(n10372) );
  INV_X1 U12018 ( .A(n11347), .ZN(n10962) );
  NOR2_X1 U12019 ( .A1(n16208), .A2(n17638), .ZN(n20079) );
  NAND2_X1 U12020 ( .A1(n11138), .A2(n9667), .ZN(n11139) );
  NAND3_X1 U12021 ( .A1(n13230), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11309), 
        .ZN(n14094) );
  INV_X1 U12022 ( .A(n10707), .ZN(n13570) );
  CLKBUF_X1 U12023 ( .A(n13413), .Z(n13571) );
  INV_X1 U12024 ( .A(n14094), .ZN(n13473) );
  INV_X1 U12025 ( .A(n16370), .ZN(n10455) );
  NOR2_X1 U12026 ( .A1(n16805), .A2(n12494), .ZN(n10387) );
  AND2_X1 U12027 ( .A1(n12830), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12832) );
  AND2_X1 U12028 ( .A1(n12828), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12830) );
  NAND2_X1 U12029 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12813), .ZN(
        n12478) );
  NOR2_X1 U12030 ( .A1(n16635), .A2(n10289), .ZN(n10288) );
  INV_X1 U12031 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10289) );
  INV_X1 U12032 ( .A(n10245), .ZN(n9804) );
  INV_X1 U12033 ( .A(n9843), .ZN(n9840) );
  NOR2_X1 U12034 ( .A1(n16775), .A2(n10389), .ZN(n10388) );
  AND2_X1 U12035 ( .A1(n15883), .A2(n11532), .ZN(n10359) );
  AND2_X1 U12036 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  INV_X1 U12037 ( .A(n15866), .ZN(n10358) );
  AOI21_X1 U12038 ( .B1(n10141), .B2(n16573), .A(n10430), .ZN(n10026) );
  INV_X1 U12039 ( .A(n11019), .ZN(n9807) );
  AND2_X1 U12040 ( .A1(n10418), .A2(n9809), .ZN(n9808) );
  NAND2_X1 U12041 ( .A1(n10209), .A2(n10020), .ZN(n10019) );
  NAND2_X1 U12042 ( .A1(n10209), .A2(n20074), .ZN(n10021) );
  INV_X1 U12043 ( .A(n10022), .ZN(n10020) );
  AOI21_X1 U12044 ( .B1(n10123), .B2(n10122), .A(n9717), .ZN(n10121) );
  INV_X1 U12045 ( .A(n16650), .ZN(n10122) );
  NOR2_X1 U12046 ( .A1(n10401), .A2(n16961), .ZN(n10042) );
  NAND2_X1 U12047 ( .A1(n10402), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10401) );
  NOR2_X1 U12048 ( .A1(n10412), .A2(n16029), .ZN(n10411) );
  INV_X1 U12049 ( .A(n10413), .ZN(n10412) );
  OR3_X1 U12050 ( .A1(n16016), .A2(n11555), .A3(n16615), .ZN(n16612) );
  AND2_X1 U12051 ( .A1(n11514), .A2(n11518), .ZN(n10341) );
  NAND2_X1 U12052 ( .A1(n9958), .A2(n9956), .ZN(n10031) );
  AOI21_X1 U12053 ( .B1(n9959), .B2(n9961), .A(n9957), .ZN(n9956) );
  NAND2_X1 U12054 ( .A1(n10420), .A2(n9959), .ZN(n9958) );
  INV_X1 U12055 ( .A(n16661), .ZN(n9957) );
  NOR2_X1 U12056 ( .A1(n10000), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U12057 ( .A1(n16699), .A2(n16692), .ZN(n10000) );
  AND3_X1 U12058 ( .A1(n11415), .A2(n11414), .A3(n11413), .ZN(n14260) );
  NAND2_X1 U12059 ( .A1(n9814), .A2(n10883), .ZN(n10905) );
  OAI21_X1 U12060 ( .B1(n10951), .B2(n9810), .A(n10022), .ZN(n16694) );
  INV_X1 U12061 ( .A(n10951), .ZN(n9848) );
  INV_X1 U12062 ( .A(n10478), .ZN(n9793) );
  AND2_X1 U12063 ( .A1(n10993), .A2(n10213), .ZN(n10212) );
  NAND2_X1 U12064 ( .A1(n16248), .A2(n11559), .ZN(n10213) );
  INV_X1 U12065 ( .A(n16248), .ZN(n10214) );
  NAND2_X1 U12066 ( .A1(n10718), .A2(n10601), .ZN(n10139) );
  NOR2_X1 U12067 ( .A1(n10115), .A2(n10044), .ZN(n10043) );
  NOR2_X1 U12068 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  AND3_X1 U12069 ( .A1(n10682), .A2(n10029), .A3(n10028), .ZN(n10036) );
  OR2_X1 U12070 ( .A1(n11307), .A2(n11312), .ZN(n11321) );
  OR2_X1 U12071 ( .A1(n16324), .A2(n17125), .ZN(n11298) );
  NAND2_X1 U12072 ( .A1(n10062), .A2(n13643), .ZN(n11268) );
  AND4_X1 U12073 ( .A1(n13636), .A2(n17276), .A3(n11256), .A4(n11255), .ZN(
        n11257) );
  NAND2_X1 U12074 ( .A1(n13676), .A2(n9753), .ZN(n10063) );
  NAND2_X1 U12075 ( .A1(n13473), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13249) );
  AND4_X1 U12076 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10714) );
  NAND2_X1 U12077 ( .A1(n10247), .A2(n10246), .ZN(n9868) );
  INV_X1 U12078 ( .A(n10244), .ZN(n9794) );
  AND2_X1 U12079 ( .A1(n10941), .A2(n10940), .ZN(n11211) );
  OR2_X1 U12080 ( .A1(n10939), .A2(n10938), .ZN(n10941) );
  NAND2_X1 U12081 ( .A1(n10532), .A2(n14056), .ZN(n10539) );
  NAND2_X1 U12082 ( .A1(n10537), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10538) );
  NOR2_X1 U12083 ( .A1(n20636), .A2(n20868), .ZN(n17187) );
  XNOR2_X1 U12084 ( .A(n14056), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10919) );
  NAND2_X1 U12085 ( .A1(n10918), .A2(n10917), .ZN(n10921) );
  NAND2_X1 U12086 ( .A1(n11251), .A2(n10575), .ZN(n11214) );
  INV_X1 U12087 ( .A(n13014), .ZN(n10201) );
  INV_X1 U12088 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9850) );
  AND2_X1 U12089 ( .A1(n10181), .A2(n10180), .ZN(n18026) );
  INV_X1 U12090 ( .A(n19012), .ZN(n10180) );
  NOR2_X1 U12091 ( .A1(n13005), .A2(n10182), .ZN(n10181) );
  INV_X1 U12092 ( .A(n19102), .ZN(n10007) );
  INV_X1 U12093 ( .A(n17319), .ZN(n17321) );
  NAND2_X1 U12094 ( .A1(n18890), .A2(n10268), .ZN(n10271) );
  NOR2_X1 U12095 ( .A1(n18939), .A2(n18927), .ZN(n10261) );
  AND2_X1 U12096 ( .A1(n10281), .A2(n17303), .ZN(n10280) );
  NOR2_X1 U12097 ( .A1(n17334), .A2(n17333), .ZN(n17335) );
  NAND2_X1 U12098 ( .A1(n19008), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19007) );
  OAI21_X1 U12099 ( .B1(n13942), .B2(n14006), .A(n10255), .ZN(n13941) );
  AND4_X1 U12100 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n13032), .ZN(
        n13051) );
  OAI221_X1 U12101 ( .B1(n19895), .B2(P3_STATE2_REG_2__SCAN_IN), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n20039), .A(n14526), .ZN(n19424) );
  AOI21_X1 U12102 ( .B1(n13979), .B2(n13978), .A(n13983), .ZN(n17328) );
  CLKBUF_X1 U12103 ( .A(n12613), .Z(n12614) );
  NAND2_X1 U12104 ( .A1(n10294), .A2(n12526), .ZN(n13654) );
  AND2_X1 U12105 ( .A1(n12664), .A2(n12663), .ZN(n14959) );
  AND3_X1 U12106 ( .A1(n11935), .A2(n11934), .A3(n11933), .ZN(n14956) );
  CLKBUF_X1 U12107 ( .A(n12730), .Z(n14885) );
  NAND2_X1 U12108 ( .A1(n14884), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14886) );
  AND2_X1 U12109 ( .A1(n12708), .A2(n12707), .ZN(n14651) );
  NAND2_X1 U12110 ( .A1(n14317), .A2(n11660), .ZN(n12432) );
  AND2_X1 U12111 ( .A1(n13817), .A2(n11798), .ZN(n14078) );
  AND2_X1 U12112 ( .A1(n12212), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12213) );
  NAND2_X1 U12113 ( .A1(n12213), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12312) );
  NOR2_X1 U12114 ( .A1(n12254), .A2(n12210), .ZN(n12236) );
  AOI22_X1 U12115 ( .A1(n15106), .A2(n14538), .B1(n12274), .B2(n12273), .ZN(
        n14688) );
  OR2_X1 U12116 ( .A1(n12129), .A2(n15130), .ZN(n12131) );
  AND2_X1 U12117 ( .A1(n12104), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12105) );
  NAND2_X1 U12118 ( .A1(n12105), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12129) );
  AND2_X1 U12119 ( .A1(n14846), .A2(n10082), .ZN(n14756) );
  AND2_X1 U12120 ( .A1(n14770), .A2(n12056), .ZN(n14771) );
  NAND2_X1 U12121 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n11947), .ZN(
        n11952) );
  INV_X1 U12122 ( .A(n11946), .ZN(n11947) );
  NAND2_X1 U12123 ( .A1(n14846), .A2(n14849), .ZN(n14848) );
  CLKBUF_X1 U12124 ( .A(n14846), .Z(n14847) );
  CLKBUF_X1 U12125 ( .A(n14858), .Z(n14955) );
  NAND2_X1 U12126 ( .A1(n11907), .A2(n11906), .ZN(n14492) );
  AOI21_X1 U12127 ( .B1(n12553), .B2(n12027), .A(n11894), .ZN(n15028) );
  INV_X1 U12128 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U12129 ( .A1(n11856), .A2(n11855), .ZN(n14484) );
  INV_X1 U12130 ( .A(n14387), .ZN(n11855) );
  AND2_X1 U12131 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11824), .ZN(
        n11852) );
  NAND2_X1 U12132 ( .A1(n11832), .A2(n11831), .ZN(n10074) );
  XNOR2_X1 U12133 ( .A(n12546), .B(n21123), .ZN(n14195) );
  AOI21_X1 U12134 ( .B1(n11779), .B2(n9890), .A(n10284), .ZN(n10283) );
  INV_X1 U12135 ( .A(n11801), .ZN(n10284) );
  NAND2_X1 U12136 ( .A1(n14078), .A2(n14079), .ZN(n14198) );
  NOR2_X1 U12137 ( .A1(n9931), .A2(n12597), .ZN(n9926) );
  AND2_X1 U12138 ( .A1(n9645), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9929) );
  NOR2_X1 U12139 ( .A1(n15044), .A2(n12757), .ZN(n10112) );
  NAND2_X1 U12140 ( .A1(n14696), .A2(n9744), .ZN(n14673) );
  NAND2_X1 U12141 ( .A1(n14696), .A2(n9743), .ZN(n14675) );
  OR2_X1 U12142 ( .A1(n10336), .A2(n10334), .ZN(n10331) );
  AND2_X1 U12143 ( .A1(n15146), .A2(n9783), .ZN(n10336) );
  NAND3_X1 U12144 ( .A1(n10337), .A2(n10333), .A3(n10338), .ZN(n10332) );
  NOR2_X1 U12145 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  NAND2_X1 U12146 ( .A1(n10096), .A2(n10334), .ZN(n15103) );
  NOR2_X1 U12147 ( .A1(n10335), .A2(n9647), .ZN(n10171) );
  AND2_X1 U12148 ( .A1(n12700), .A2(n12699), .ZN(n14709) );
  NOR3_X1 U12149 ( .A1(n15118), .A2(n15117), .A3(n15136), .ZN(n15119) );
  NAND2_X1 U12150 ( .A1(n14773), .A2(n9636), .ZN(n14725) );
  AND2_X1 U12151 ( .A1(n14773), .A2(n9677), .ZN(n14750) );
  XNOR2_X1 U12152 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15146) );
  AND2_X1 U12153 ( .A1(n12691), .A2(n12690), .ZN(n14767) );
  OR2_X1 U12154 ( .A1(n12592), .A2(n15169), .ZN(n15158) );
  AND2_X1 U12155 ( .A1(n14773), .A2(n12687), .ZN(n14776) );
  XNOR2_X1 U12156 ( .A(n15227), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15173) );
  NAND2_X1 U12157 ( .A1(n15227), .A2(n15408), .ZN(n15171) );
  AND2_X1 U12158 ( .A1(n12685), .A2(n12684), .ZN(n14800) );
  NAND2_X1 U12159 ( .A1(n9662), .A2(n10316), .ZN(n10315) );
  INV_X1 U12160 ( .A(n14812), .ZN(n10316) );
  AND2_X1 U12161 ( .A1(n12585), .A2(n10172), .ZN(n15195) );
  INV_X1 U12162 ( .A(n15204), .ZN(n10172) );
  NAND2_X1 U12163 ( .A1(n10318), .A2(n9662), .ZN(n14839) );
  AND2_X1 U12164 ( .A1(n12671), .A2(n12670), .ZN(n14947) );
  NAND2_X1 U12165 ( .A1(n10318), .A2(n12672), .ZN(n14950) );
  NAND2_X1 U12166 ( .A1(n17573), .A2(n17571), .ZN(n10326) );
  NAND2_X1 U12167 ( .A1(n17612), .A2(n10314), .ZN(n14958) );
  NAND2_X1 U12168 ( .A1(n10104), .A2(n12561), .ZN(n17573) );
  NAND2_X1 U12169 ( .A1(n12559), .A2(n12558), .ZN(n17578) );
  NAND2_X1 U12170 ( .A1(n15504), .A2(n21369), .ZN(n12996) );
  NOR2_X2 U12171 ( .A1(n14429), .A2(n12646), .ZN(n14487) );
  XNOR2_X1 U12172 ( .A(n12551), .B(n17627), .ZN(n17585) );
  OR2_X1 U12173 ( .A1(n12749), .A2(n15501), .ZN(n15434) );
  XNOR2_X1 U12174 ( .A(n11788), .B(n11787), .ZN(n12532) );
  OR2_X1 U12175 ( .A1(n12530), .A2(n11780), .ZN(n11781) );
  INV_X1 U12176 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11823) );
  INV_X1 U12177 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10111) );
  INV_X1 U12178 ( .A(n17532), .ZN(n13851) );
  OR2_X1 U12179 ( .A1(n21175), .A2(n15561), .ZN(n15564) );
  INV_X1 U12180 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17510) );
  INV_X1 U12181 ( .A(n12609), .ZN(n14309) );
  AND2_X1 U12182 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15533), .ZN(n14324) );
  AND2_X1 U12183 ( .A1(n15762), .A2(n21285), .ZN(n15768) );
  NAND2_X1 U12184 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21389) );
  CLKBUF_X1 U12185 ( .A(n11220), .Z(n11221) );
  NOR2_X1 U12186 ( .A1(n11544), .A2(n10365), .ZN(n10364) );
  NOR2_X1 U12187 ( .A1(n15901), .A2(n15904), .ZN(n15888) );
  NAND2_X1 U12188 ( .A1(n11099), .A2(n9746), .ZN(n11100) );
  AND2_X1 U12189 ( .A1(n10368), .A2(n11155), .ZN(n10367) );
  NAND2_X1 U12190 ( .A1(n11077), .A2(n10368), .ZN(n11094) );
  INV_X1 U12191 ( .A(n15970), .ZN(n15952) );
  NAND2_X1 U12192 ( .A1(n11077), .A2(n11078), .ZN(n11083) );
  AND2_X1 U12193 ( .A1(n16625), .A2(n10226), .ZN(n10225) );
  NOR2_X1 U12194 ( .A1(n16638), .A2(n10227), .ZN(n10226) );
  NAND2_X1 U12195 ( .A1(n10380), .A2(n10381), .ZN(n11060) );
  NAND2_X1 U12196 ( .A1(n16065), .A2(n16645), .ZN(n16048) );
  NOR3_X1 U12197 ( .A1(n16136), .A2(n10233), .A3(n10229), .ZN(n16077) );
  INV_X1 U12198 ( .A(n16664), .ZN(n10233) );
  NOR2_X1 U12199 ( .A1(n16136), .A2(n10231), .ZN(n16105) );
  NOR2_X1 U12200 ( .A1(n16136), .A2(n16709), .ZN(n16118) );
  NAND2_X1 U12201 ( .A1(n10374), .A2(n20107), .ZN(n10373) );
  INV_X1 U12202 ( .A(n10375), .ZN(n10374) );
  NAND2_X1 U12203 ( .A1(n16182), .A2(n16745), .ZN(n16167) );
  NOR2_X1 U12204 ( .A1(n16196), .A2(n16762), .ZN(n16182) );
  NAND2_X1 U12205 ( .A1(n20079), .A2(n20081), .ZN(n16196) );
  AND2_X1 U12206 ( .A1(n14033), .A2(n13255), .ZN(n16218) );
  NAND2_X1 U12207 ( .A1(n16290), .A2(n20187), .ZN(n10311) );
  AND2_X1 U12208 ( .A1(n12779), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12209 ( .A1(n11181), .A2(n9752), .ZN(n11182) );
  NAND2_X1 U12210 ( .A1(n11169), .A2(n9747), .ZN(n11170) );
  INV_X1 U12211 ( .A(n10399), .ZN(n10397) );
  NAND2_X1 U12212 ( .A1(n11136), .A2(n9674), .ZN(n11137) );
  NAND2_X1 U12213 ( .A1(n11135), .A2(n10413), .ZN(n16043) );
  NOR2_X1 U12214 ( .A1(n9661), .A2(n10445), .ZN(n10444) );
  INV_X1 U12215 ( .A(n13255), .ZN(n10445) );
  NAND2_X1 U12216 ( .A1(n11113), .A2(n9670), .ZN(n11114) );
  CLKBUF_X1 U12217 ( .A(n14092), .Z(n14095) );
  AND2_X1 U12218 ( .A1(n10449), .A2(n10451), .ZN(n10448) );
  NOR2_X1 U12219 ( .A1(n13364), .A2(n13363), .ZN(n16350) );
  INV_X1 U12220 ( .A(n16353), .ZN(n10442) );
  AND2_X1 U12221 ( .A1(n11520), .A2(n11519), .ZN(n16014) );
  NOR2_X1 U12222 ( .A1(n10453), .A2(n16377), .ZN(n10154) );
  AND2_X2 U12223 ( .A1(n13593), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n17185)
         );
  NAND2_X1 U12224 ( .A1(n10385), .A2(n12779), .ZN(n9843) );
  NAND2_X1 U12225 ( .A1(n10386), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9842) );
  NOR2_X1 U12226 ( .A1(n12825), .A2(n12953), .ZN(n12828) );
  AND2_X1 U12227 ( .A1(n9646), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10296) );
  NAND2_X1 U12228 ( .A1(n12820), .A2(n9646), .ZN(n12822) );
  NAND2_X1 U12229 ( .A1(n12820), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12816) );
  INV_X1 U12230 ( .A(n12478), .ZN(n12818) );
  AND2_X1 U12231 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12818), .ZN(
        n12820) );
  NAND2_X1 U12232 ( .A1(n12809), .A2(n10288), .ZN(n12784) );
  NAND2_X1 U12233 ( .A1(n12809), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12811) );
  NOR2_X1 U12234 ( .A1(n12449), .A2(n10406), .ZN(n10405) );
  NAND2_X1 U12235 ( .A1(n11132), .A2(n9673), .ZN(n11133) );
  NOR2_X1 U12236 ( .A1(n12806), .A2(n16093), .ZN(n12807) );
  AND2_X1 U12237 ( .A1(n12807), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12809) );
  NAND2_X1 U12238 ( .A1(n10391), .A2(n16088), .ZN(n10390) );
  INV_X1 U12239 ( .A(n10393), .ZN(n10391) );
  INV_X1 U12240 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12803) );
  OR2_X1 U12241 ( .A1(n12804), .A2(n12803), .ZN(n12806) );
  NAND2_X1 U12242 ( .A1(n12789), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12804) );
  NOR2_X1 U12243 ( .A1(n12792), .A2(n16707), .ZN(n12789) );
  INV_X1 U12244 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16707) );
  AND2_X1 U12245 ( .A1(n9634), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U12246 ( .A1(n12802), .A2(n9634), .ZN(n12796) );
  NAND2_X1 U12247 ( .A1(n12802), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12801) );
  AND2_X1 U12248 ( .A1(n12802), .A2(n10300), .ZN(n12797) );
  INV_X1 U12249 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16760) );
  NAND2_X1 U12250 ( .A1(n11106), .A2(n9669), .ZN(n11107) );
  NAND2_X1 U12251 ( .A1(n10245), .A2(n10661), .ZN(n9805) );
  NAND2_X1 U12252 ( .A1(n11103), .A2(n9693), .ZN(n11105) );
  NOR2_X1 U12253 ( .A1(n12798), .A2(n17655), .ZN(n12800) );
  NAND2_X1 U12254 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U12256 ( .A1(n16530), .A2(n17090), .ZN(n10046) );
  NAND2_X1 U12257 ( .A1(n12495), .A2(n9838), .ZN(n9837) );
  NAND2_X1 U12258 ( .A1(n12495), .A2(n9840), .ZN(n9839) );
  INV_X1 U12259 ( .A(n9842), .ZN(n9838) );
  NAND2_X1 U12260 ( .A1(n16806), .A2(n11291), .ZN(n12493) );
  NOR2_X1 U12261 ( .A1(n10221), .A2(n10430), .ZN(n10220) );
  NAND2_X1 U12262 ( .A1(n9983), .A2(n10222), .ZN(n10219) );
  NAND2_X1 U12263 ( .A1(n11554), .A2(n11550), .ZN(n9983) );
  AND2_X1 U12264 ( .A1(n11529), .A2(n11528), .ZN(n15914) );
  AND2_X1 U12265 ( .A1(n16979), .A2(n10053), .ZN(n16844) );
  NOR2_X1 U12266 ( .A1(n10054), .A2(n11280), .ZN(n10053) );
  INV_X1 U12267 ( .A(n10055), .ZN(n10054) );
  INV_X1 U12268 ( .A(n10023), .ZN(n11087) );
  AOI21_X1 U12269 ( .B1(n10143), .B2(n10140), .A(n10024), .ZN(n10023) );
  NAND2_X1 U12270 ( .A1(n10025), .A2(n16573), .ZN(n10024) );
  NAND2_X1 U12271 ( .A1(n10140), .A2(n10142), .ZN(n10025) );
  NAND2_X1 U12272 ( .A1(n11150), .A2(n9749), .ZN(n11151) );
  NAND2_X1 U12273 ( .A1(n10346), .A2(n15946), .ZN(n10345) );
  INV_X1 U12274 ( .A(n10347), .ZN(n10346) );
  AND2_X1 U12275 ( .A1(n16579), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16580) );
  NAND2_X1 U12276 ( .A1(n11148), .A2(n9748), .ZN(n11149) );
  CLKBUF_X1 U12277 ( .A(n15966), .Z(n15987) );
  AND2_X1 U12278 ( .A1(n11525), .A2(n11524), .ZN(n15963) );
  NOR2_X1 U12279 ( .A1(n16584), .A2(n10073), .ZN(n10071) );
  NAND2_X1 U12280 ( .A1(n16979), .A2(n10055), .ZN(n16878) );
  INV_X1 U12281 ( .A(n16598), .ZN(n10422) );
  OR2_X1 U12282 ( .A1(n12455), .A2(n16632), .ZN(n10425) );
  NAND2_X1 U12283 ( .A1(n10121), .A2(n10124), .ZN(n10119) );
  INV_X1 U12284 ( .A(n12450), .ZN(n10404) );
  AND2_X1 U12285 ( .A1(n11135), .A2(n10411), .ZN(n16028) );
  CLKBUF_X1 U12286 ( .A(n12458), .Z(n12459) );
  NOR2_X1 U12287 ( .A1(n16611), .A2(n10426), .ZN(n9953) );
  AND2_X1 U12288 ( .A1(n9950), .A2(n9739), .ZN(n9948) );
  AOI21_X1 U12289 ( .B1(n16620), .B2(n9954), .A(n9951), .ZN(n9950) );
  INV_X1 U12290 ( .A(n16621), .ZN(n9951) );
  INV_X1 U12291 ( .A(n16631), .ZN(n10429) );
  INV_X1 U12292 ( .A(n12452), .ZN(n10428) );
  INV_X1 U12293 ( .A(n16632), .ZN(n9954) );
  NAND2_X1 U12294 ( .A1(n10354), .A2(n11475), .ZN(n10352) );
  NAND2_X1 U12295 ( .A1(n11126), .A2(n9672), .ZN(n11127) );
  INV_X1 U12296 ( .A(n16113), .ZN(n10392) );
  OR2_X1 U12297 ( .A1(n11071), .A2(n16961), .ZN(n16671) );
  AND3_X1 U12298 ( .A1(n11435), .A2(n11434), .A3(n11433), .ZN(n14268) );
  NAND2_X1 U12299 ( .A1(n11118), .A2(n9665), .ZN(n11119) );
  INV_X1 U12300 ( .A(n14276), .ZN(n11393) );
  AND2_X1 U12301 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  INV_X1 U12302 ( .A(n16161), .ZN(n10409) );
  INV_X1 U12303 ( .A(n16749), .ZN(n10907) );
  AND3_X1 U12304 ( .A1(n11372), .A2(n11371), .A3(n11370), .ZN(n14273) );
  CLKBUF_X1 U12305 ( .A(n14271), .Z(n14277) );
  INV_X1 U12306 ( .A(n10045), .ZN(n16754) );
  NAND2_X1 U12307 ( .A1(n9811), .A2(n20074), .ZN(n16693) );
  AND3_X1 U12308 ( .A1(n11341), .A2(n11340), .A3(n11339), .ZN(n16225) );
  NAND2_X1 U12309 ( .A1(n10973), .A2(n9978), .ZN(n10991) );
  NAND2_X1 U12310 ( .A1(n17105), .A2(n11555), .ZN(n10211) );
  NAND2_X1 U12311 ( .A1(n10059), .A2(n20235), .ZN(n17087) );
  AND2_X1 U12312 ( .A1(n11270), .A2(n11271), .ZN(n10059) );
  NOR2_X1 U12313 ( .A1(n10058), .A2(n10060), .ZN(n17098) );
  INV_X1 U12314 ( .A(n20235), .ZN(n10058) );
  NAND2_X1 U12315 ( .A1(n13224), .A2(n11308), .ZN(n13247) );
  AND2_X1 U12316 ( .A1(n11231), .A2(n11230), .ZN(n17127) );
  NAND2_X1 U12317 ( .A1(n9713), .A2(n10591), .ZN(n11229) );
  INV_X1 U12318 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17138) );
  INV_X1 U12319 ( .A(n17677), .ZN(n13643) );
  NAND2_X1 U12320 ( .A1(n10127), .A2(n9611), .ZN(n20319) );
  INV_X1 U12321 ( .A(n10819), .ZN(n20348) );
  INV_X1 U12322 ( .A(n10854), .ZN(n20528) );
  INV_X1 U12323 ( .A(n20870), .ZN(n20346) );
  NAND2_X2 U12324 ( .A1(n10527), .A2(n10526), .ZN(n17205) );
  NAND2_X1 U12325 ( .A1(n10525), .A2(n14056), .ZN(n10526) );
  NAND2_X1 U12326 ( .A1(n20876), .A2(n17220), .ZN(n20674) );
  INV_X1 U12327 ( .A(n20680), .ZN(n20687) );
  OR2_X1 U12328 ( .A1(n20674), .A2(n20673), .ZN(n20682) );
  NAND2_X1 U12329 ( .A1(n17185), .A2(n17187), .ZN(n20290) );
  NAND2_X1 U12330 ( .A1(n17187), .A2(n17186), .ZN(n20289) );
  NAND2_X1 U12331 ( .A1(n10556), .A2(n14056), .ZN(n10563) );
  INV_X1 U12332 ( .A(n20280), .ZN(n20287) );
  OR2_X1 U12333 ( .A1(n10939), .A2(n10940), .ZN(n11208) );
  XNOR2_X1 U12334 ( .A(n10921), .B(n10919), .ZN(n11204) );
  OR2_X1 U12335 ( .A1(n12834), .A2(n12833), .ZN(n16274) );
  NAND2_X1 U12336 ( .A1(n17887), .A2(n17892), .ZN(n17871) );
  NOR2_X1 U12337 ( .A1(n9628), .A2(n13014), .ZN(n17945) );
  NOR2_X1 U12338 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18030), .ZN(n18014) );
  NAND2_X1 U12339 ( .A1(n18041), .A2(n18034), .ZN(n18030) );
  INV_X1 U12340 ( .A(n18052), .ZN(n18013) );
  NOR2_X1 U12341 ( .A1(n18126), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n18110) );
  INV_X1 U12342 ( .A(n13173), .ZN(n13181) );
  NOR2_X1 U12343 ( .A1(n18624), .A2(n18626), .ZN(n9963) );
  OR2_X1 U12344 ( .A1(n13878), .A2(n13877), .ZN(n14016) );
  OR2_X1 U12345 ( .A1(n18597), .A2(n18474), .ZN(n18590) );
  NOR3_X1 U12346 ( .A1(n14057), .A2(n18620), .A3(n14497), .ZN(n14086) );
  INV_X1 U12347 ( .A(n9975), .ZN(n14103) );
  OAI21_X1 U12348 ( .B1(n14062), .B2(n14061), .A(n20027), .ZN(n18619) );
  NAND2_X1 U12349 ( .A1(n18764), .A2(n9644), .ZN(n13023) );
  AND2_X1 U12350 ( .A1(n18764), .A2(n9772), .ZN(n13022) );
  NOR2_X1 U12351 ( .A1(n9740), .A2(n13016), .ZN(n10191) );
  NAND2_X1 U12352 ( .A1(n10190), .A2(n10193), .ZN(n18854) );
  NAND2_X1 U12353 ( .A1(n18052), .A2(n18026), .ZN(n18941) );
  AND2_X1 U12354 ( .A1(n17376), .A2(n10259), .ZN(n10257) );
  NOR2_X1 U12355 ( .A1(n9852), .A2(n19290), .ZN(n9851) );
  INV_X1 U12356 ( .A(n19104), .ZN(n9852) );
  NAND2_X1 U12357 ( .A1(n19158), .A2(n18744), .ZN(n19105) );
  NAND2_X1 U12358 ( .A1(n9754), .A2(n18794), .ZN(n18793) );
  CLKBUF_X1 U12359 ( .A(n18804), .Z(n18848) );
  AND2_X1 U12360 ( .A1(n17301), .A2(n10282), .ZN(n10281) );
  NAND2_X1 U12361 ( .A1(n17302), .A2(n10280), .ZN(n18973) );
  NOR2_X1 U12362 ( .A1(n13985), .A2(n13130), .ZN(n14069) );
  NOR2_X1 U12363 ( .A1(n19322), .A2(n18890), .ZN(n17351) );
  AND2_X1 U12364 ( .A1(n14024), .A2(n17386), .ZN(n14025) );
  INV_X1 U12365 ( .A(n14023), .ZN(n14026) );
  NAND2_X1 U12366 ( .A1(n19025), .A2(n13955), .ZN(n17336) );
  NOR2_X1 U12367 ( .A1(n17336), .A2(n17337), .ZN(n17334) );
  XNOR2_X1 U12368 ( .A(n13954), .B(n10254), .ZN(n19026) );
  INV_X1 U12369 ( .A(n13953), .ZN(n10254) );
  NAND2_X1 U12370 ( .A1(n19026), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19025) );
  NAND2_X1 U12371 ( .A1(n19049), .A2(n13951), .ZN(n9847) );
  OAI21_X1 U12372 ( .B1(n19067), .B2(n9999), .A(n9997), .ZN(n14010) );
  XNOR2_X1 U12373 ( .A(n13949), .B(n10253), .ZN(n19050) );
  INV_X1 U12374 ( .A(n13950), .ZN(n10253) );
  NAND2_X1 U12375 ( .A1(n19050), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19049) );
  AND2_X1 U12376 ( .A1(n19227), .A2(n19430), .ZN(n19878) );
  INV_X1 U12377 ( .A(n13905), .ZN(n19094) );
  NAND3_X1 U12378 ( .A1(n20039), .A2(n20009), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19756) );
  INV_X1 U12379 ( .A(n13985), .ZN(n19434) );
  NOR2_X2 U12380 ( .A1(n13098), .A2(n13097), .ZN(n19438) );
  INV_X1 U12381 ( .A(n18479), .ZN(n19446) );
  NAND2_X1 U12382 ( .A1(n20030), .A2(n19424), .ZN(n19523) );
  NOR2_X1 U12383 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n13166) );
  OAI211_X1 U12384 ( .C1(n14057), .C2(n20027), .A(n20023), .B(n17812), .ZN(
        n19898) );
  NAND2_X1 U12385 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20023) );
  OR3_X1 U12386 ( .A1(n17532), .A2(n11674), .A3(n20927), .ZN(n14536) );
  NAND2_X1 U12387 ( .A1(n14536), .A2(n14535), .ZN(n21462) );
  INV_X1 U12388 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20981) );
  INV_X1 U12389 ( .A(n21016), .ZN(n20980) );
  AND2_X1 U12390 ( .A1(n14884), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21016) );
  INV_X1 U12391 ( .A(n20974), .ZN(n20989) );
  OR2_X1 U12392 ( .A1(n14611), .A2(n14610), .ZN(n15287) );
  AND2_X1 U12393 ( .A1(n12859), .A2(n13624), .ZN(n21035) );
  INV_X1 U12394 ( .A(n14567), .ZN(n15005) );
  NOR2_X1 U12395 ( .A1(n15022), .A2(n14082), .ZN(n15023) );
  OR2_X1 U12396 ( .A1(n12419), .A2(n13836), .ZN(n12420) );
  INV_X1 U12397 ( .A(n15023), .ZN(n15033) );
  INV_X1 U12398 ( .A(n21069), .ZN(n21044) );
  OR2_X1 U12399 ( .A1(n21090), .A2(n14542), .ZN(n14443) );
  AOI21_X1 U12400 ( .B1(n14599), .B2(n14598), .A(n14597), .ZN(n15051) );
  NAND2_X1 U12401 ( .A1(n12988), .A2(n12987), .ZN(n14650) );
  OR2_X1 U12402 ( .A1(n14664), .A2(n12985), .ZN(n12988) );
  INV_X1 U12403 ( .A(n14663), .ZN(n14665) );
  AND2_X1 U12404 ( .A1(n14712), .A2(n12128), .ZN(n10480) );
  INV_X1 U12405 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15130) );
  INV_X1 U12406 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15177) );
  AND2_X1 U12407 ( .A1(n14938), .A2(n14937), .ZN(n17556) );
  INV_X1 U12408 ( .A(n20932), .ZN(n21102) );
  AND2_X1 U12409 ( .A1(n15271), .A2(n21142), .ZN(n9902) );
  XNOR2_X1 U12410 ( .A(n12725), .B(n14581), .ZN(n14573) );
  NAND2_X1 U12411 ( .A1(n15036), .A2(n15037), .ZN(n15047) );
  INV_X1 U12412 ( .A(n12993), .ZN(n10177) );
  NAND2_X1 U12413 ( .A1(n15339), .A2(n12755), .ZN(n15334) );
  AND3_X1 U12414 ( .A1(n15386), .A2(n21129), .A3(n15385), .ZN(n15428) );
  INV_X1 U12415 ( .A(n15482), .ZN(n21145) );
  OR2_X1 U12416 ( .A1(n12749), .A2(n12745), .ZN(n17600) );
  NAND2_X1 U12417 ( .A1(n9894), .A2(n9759), .ZN(n15342) );
  OR2_X1 U12418 ( .A1(n12749), .A2(n12625), .ZN(n15482) );
  NAND2_X1 U12419 ( .A1(n13653), .A2(n9776), .ZN(n12623) );
  INV_X1 U12420 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21307) );
  CLKBUF_X1 U12422 ( .A(n12539), .Z(n14285) );
  AND2_X1 U12423 ( .A1(n15560), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15603) );
  INV_X1 U12424 ( .A(n21285), .ZN(n21311) );
  CLKBUF_X1 U12425 ( .A(n14213), .Z(n15531) );
  OAI21_X1 U12426 ( .B1(n14251), .B2(n17635), .A(n15642), .ZN(n21153) );
  NOR2_X1 U12427 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15504) );
  OAI22_X1 U12428 ( .A1(n15541), .A2(n15540), .B1(n15539), .B2(n21201), .ZN(
        n21165) );
  AOI22_X1 U12429 ( .A1(n15568), .A2(n15565), .B1(n15723), .B2(n15640), .ZN(
        n15596) );
  OAI21_X1 U12430 ( .B1(n21209), .B2(n21239), .A(n21208), .ZN(n21243) );
  OAI21_X1 U12431 ( .B1(n21202), .B2(n21201), .A(n21200), .ZN(n21240) );
  AOI22_X1 U12432 ( .A1(n15646), .A2(n15643), .B1(n15640), .B2(n15798), .ZN(
        n15675) );
  INV_X1 U12433 ( .A(n15672), .ZN(n14424) );
  OAI211_X1 U12434 ( .C1(n15680), .C2(n17636), .A(n15679), .B(n15678), .ZN(
        n15711) );
  AOI22_X1 U12435 ( .A1(n15731), .A2(n15726), .B1(n15723), .B2(n15799), .ZN(
        n15760) );
  AOI22_X1 U12436 ( .A1(n15768), .A2(n15764), .B1(n15765), .B2(n15798), .ZN(
        n15797) );
  INV_X1 U12437 ( .A(n21314), .ZN(n15812) );
  INV_X1 U12438 ( .A(n21323), .ZN(n15815) );
  INV_X1 U12439 ( .A(n21329), .ZN(n15818) );
  INV_X1 U12440 ( .A(n21341), .ZN(n15824) );
  INV_X1 U12441 ( .A(n21347), .ZN(n15827) );
  INV_X1 U12442 ( .A(n21353), .ZN(n15830) );
  INV_X1 U12443 ( .A(n21361), .ZN(n15837) );
  OAI211_X1 U12444 ( .C1(n15832), .C2(n15809), .A(n21208), .B(n15808), .ZN(
        n15831) );
  NOR2_X1 U12445 ( .A1(n15642), .A2(n14303), .ZN(n21314) );
  INV_X1 U12446 ( .A(n15683), .ZN(n21313) );
  NOR2_X1 U12447 ( .A1(n15642), .A2(n14313), .ZN(n21323) );
  INV_X1 U12448 ( .A(n15687), .ZN(n21322) );
  NOR2_X1 U12449 ( .A1(n15642), .A2(n14308), .ZN(n21329) );
  NOR2_X1 U12450 ( .A1(n15642), .A2(n14298), .ZN(n21335) );
  INV_X1 U12451 ( .A(n15695), .ZN(n21334) );
  NOR2_X1 U12452 ( .A1(n15642), .A2(n14390), .ZN(n21341) );
  INV_X1 U12453 ( .A(n15699), .ZN(n21340) );
  NOR2_X1 U12454 ( .A1(n15642), .A2(n14490), .ZN(n21347) );
  NOR2_X1 U12455 ( .A1(n15642), .A2(n15032), .ZN(n21353) );
  INV_X1 U12456 ( .A(n15707), .ZN(n21352) );
  INV_X1 U12457 ( .A(n15712), .ZN(n21359) );
  AND2_X1 U12458 ( .A1(n15803), .A2(n15597), .ZN(n21164) );
  AND2_X1 U12459 ( .A1(n15803), .A2(n14400), .ZN(n15833) );
  NAND2_X1 U12460 ( .A1(n13625), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17527) );
  NOR2_X1 U12461 ( .A1(n13625), .A2(n11775), .ZN(n17632) );
  NOR2_X1 U12462 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21468) );
  AND2_X1 U12463 ( .A1(n17531), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n17637) );
  NOR2_X1 U12464 ( .A1(n21377), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21461) );
  NAND2_X1 U12465 ( .A1(n17114), .A2(n17113), .ZN(n20916) );
  AND2_X1 U12466 ( .A1(n15970), .A2(n10224), .ZN(n15936) );
  NOR2_X1 U12467 ( .A1(n15951), .A2(n9737), .ZN(n10224) );
  AND2_X1 U12468 ( .A1(n11017), .A2(n9654), .ZN(n16173) );
  INV_X1 U12469 ( .A(n20072), .ZN(n16292) );
  OR2_X1 U12470 ( .A1(n20908), .A2(n12776), .ZN(n20073) );
  INV_X1 U12471 ( .A(n20077), .ZN(n16294) );
  INV_X1 U12472 ( .A(n13666), .ZN(n16300) );
  OR2_X1 U12473 ( .A1(n13202), .A2(n13206), .ZN(n16794) );
  INV_X1 U12474 ( .A(n13203), .ZN(n13205) );
  CLKBUF_X1 U12475 ( .A(n16375), .Z(n16376) );
  NOR2_X1 U12476 ( .A1(n11487), .A2(n11486), .ZN(n16387) );
  NAND2_X1 U12477 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n16414) );
  AND2_X1 U12478 ( .A1(n20112), .A2(n10625), .ZN(n20108) );
  INV_X1 U12479 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n16255) );
  INV_X1 U12480 ( .A(n20108), .ZN(n20101) );
  CLKBUF_X1 U12481 ( .A(n16344), .Z(n16345) );
  INV_X1 U12482 ( .A(n20115), .ZN(n16513) );
  AND2_X1 U12483 ( .A1(n14165), .A2(n17186), .ZN(n20115) );
  AND2_X1 U12484 ( .A1(n14165), .A2(n17185), .ZN(n20116) );
  OR2_X1 U12485 ( .A1(n14165), .A2(n20114), .ZN(n16522) );
  NOR2_X1 U12486 ( .A1(n13663), .A2(n13665), .ZN(n17219) );
  AND4_X1 U12487 ( .A1(n13664), .A2(n13230), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n11308), .ZN(n13665) );
  INV_X1 U12488 ( .A(n16517), .ZN(n20134) );
  NAND2_X1 U12489 ( .A1(n13677), .A2(n13762), .ZN(n13678) );
  INV_X1 U12490 ( .A(n20145), .ZN(n20176) );
  CLKBUF_X1 U12491 ( .A(n13794), .Z(n13791) );
  NOR2_X2 U12492 ( .A1(n13670), .A2(n16324), .ZN(n13783) );
  INV_X1 U12493 ( .A(n16794), .ZN(n15879) );
  NAND2_X1 U12494 ( .A1(n13210), .A2(n9985), .ZN(n10484) );
  INV_X1 U12495 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16635) );
  INV_X1 U12496 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17644) );
  INV_X1 U12497 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17655) );
  INV_X1 U12498 ( .A(n9866), .ZN(n16537) );
  NAND2_X1 U12499 ( .A1(n13198), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U12500 ( .A1(n13210), .A2(n9986), .ZN(n16799) );
  AND2_X1 U12501 ( .A1(n9655), .A2(n15867), .ZN(n16796) );
  NAND2_X1 U12502 ( .A1(n10143), .A2(n11076), .ZN(n16588) );
  OAI21_X1 U12503 ( .B1(n16583), .B2(n10403), .A(n16615), .ZN(n9920) );
  NAND2_X1 U12504 ( .A1(n16641), .A2(n10032), .ZN(n16924) );
  NAND2_X1 U12505 ( .A1(n10034), .A2(n10033), .ZN(n10032) );
  INV_X1 U12506 ( .A(n16642), .ZN(n10033) );
  NAND2_X1 U12507 ( .A1(n10125), .A2(n16651), .ZN(n10034) );
  NAND2_X1 U12508 ( .A1(n9936), .A2(n9706), .ZN(n16928) );
  NAND2_X1 U12509 ( .A1(n16669), .A2(n9937), .ZN(n9936) );
  AND2_X1 U12510 ( .A1(n9938), .A2(n10406), .ZN(n9937) );
  NAND2_X1 U12511 ( .A1(n16979), .A2(n11276), .ZN(n16942) );
  OAI21_X1 U12512 ( .B1(n10420), .B2(n9961), .A(n9959), .ZN(n16663) );
  OAI21_X1 U12513 ( .B1(n16669), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16583), .ZN(n16971) );
  INV_X1 U12514 ( .A(n9984), .ZN(n16750) );
  OR2_X1 U12515 ( .A1(n11272), .A2(n17087), .ZN(n17049) );
  NAND2_X1 U12516 ( .A1(n16909), .A2(n20217), .ZN(n20236) );
  INV_X1 U12517 ( .A(n17219), .ZN(n17220) );
  OR2_X1 U12518 ( .A1(n20881), .A2(n20050), .ZN(n20868) );
  INV_X1 U12519 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20894) );
  NAND2_X1 U12520 ( .A1(n20559), .A2(n11308), .ZN(n20881) );
  NAND2_X1 U12521 ( .A1(n14175), .A2(n11330), .ZN(n16246) );
  NOR2_X1 U12522 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17288) );
  NOR2_X1 U12523 ( .A1(n17266), .A2(n11308), .ZN(n17668) );
  NAND2_X1 U12524 ( .A1(n17179), .A2(n17178), .ZN(n20311) );
  NOR2_X1 U12525 ( .A1(n20383), .A2(n20382), .ZN(n20405) );
  OAI21_X1 U12526 ( .B1(n10465), .B2(n11308), .A(n20441), .ZN(n20458) );
  NOR2_X1 U12527 ( .A1(n20500), .A2(n20501), .ZN(n20502) );
  INV_X1 U12528 ( .A(n20492), .ZN(n20550) );
  OAI21_X1 U12529 ( .B1(n20558), .B2(n20557), .A(n20556), .ZN(n20580) );
  INV_X1 U12530 ( .A(n20592), .ZN(n20607) );
  NOR2_X2 U12531 ( .A1(n20627), .A2(n20346), .ZN(n20622) );
  AOI21_X1 U12532 ( .B1(n20559), .B2(n17237), .A(n17236), .ZN(n20621) );
  OAI21_X1 U12533 ( .B1(n20639), .B2(n20638), .A(n20637), .ZN(n20670) );
  OAI22_X1 U12534 ( .A1(n17729), .A2(n20290), .B1(n16505), .B2(n20289), .ZN(
        n20696) );
  OAI22_X1 U12535 ( .A1(n17727), .A2(n20290), .B1(n16497), .B2(n20289), .ZN(
        n20700) );
  OAI22_X1 U12536 ( .A1(n20275), .A2(n20290), .B1(n20274), .B2(n20289), .ZN(
        n20708) );
  OAI22_X1 U12537 ( .A1(n20291), .A2(n20290), .B1(n16469), .B2(n20289), .ZN(
        n20717) );
  INV_X1 U12538 ( .A(n20691), .ZN(n20730) );
  INV_X1 U12539 ( .A(n20683), .ZN(n20741) );
  AND2_X1 U12540 ( .A1(n11297), .A2(n20287), .ZN(n20742) );
  INV_X1 U12541 ( .A(n20692), .ZN(n20747) );
  AND2_X1 U12542 ( .A1(n17239), .A2(n20287), .ZN(n20748) );
  AND2_X1 U12543 ( .A1(n20731), .A2(n17238), .ZN(n20749) );
  INV_X1 U12544 ( .A(n20696), .ZN(n20753) );
  INV_X1 U12545 ( .A(n20654), .ZN(n20760) );
  AND2_X1 U12546 ( .A1(n20731), .A2(n17210), .ZN(n20761) );
  INV_X1 U12547 ( .A(n20708), .ZN(n20771) );
  AND2_X1 U12548 ( .A1(n20731), .A2(n20278), .ZN(n20773) );
  INV_X1 U12549 ( .A(n20712), .ZN(n20777) );
  INV_X1 U12550 ( .A(n20682), .ZN(n20783) );
  NOR2_X1 U12551 ( .A1(n20733), .A2(n20727), .ZN(n20781) );
  AND2_X1 U12552 ( .A1(n20731), .A2(n20284), .ZN(n20780) );
  INV_X1 U12553 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17290) );
  NAND2_X1 U12554 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20917) );
  INV_X1 U12555 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20861) );
  NAND2_X1 U12556 ( .A1(n20026), .A2(n19876), .ZN(n18679) );
  INV_X1 U12557 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20030) );
  XNOR2_X1 U12558 ( .A(n17834), .B(n10188), .ZN(n10187) );
  INV_X1 U12559 ( .A(n17835), .ZN(n10188) );
  INV_X1 U12560 ( .A(n17840), .ZN(n10184) );
  INV_X1 U12561 ( .A(n10200), .ZN(n17853) );
  OAI21_X1 U12562 ( .B1(n17872), .B2(n17862), .A(n10196), .ZN(n10200) );
  NOR2_X1 U12563 ( .A1(n17871), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17870) );
  NOR2_X1 U12564 ( .A1(n17861), .A2(n17862), .ZN(n17860) );
  AND2_X1 U12565 ( .A1(n17872), .A2(n10198), .ZN(n17861) );
  AND2_X1 U12566 ( .A1(n10206), .A2(n10198), .ZN(n17935) );
  NOR2_X1 U12567 ( .A1(n17962), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17946) );
  NAND2_X1 U12568 ( .A1(n17946), .A2(n18279), .ZN(n17939) );
  NAND2_X1 U12569 ( .A1(n17969), .A2(n18306), .ZN(n17962) );
  NOR2_X1 U12570 ( .A1(n17983), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17969) );
  NOR2_X1 U12571 ( .A1(n18056), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n18041) );
  NAND2_X1 U12572 ( .A1(n18063), .A2(n18062), .ZN(n18056) );
  NOR2_X1 U12573 ( .A1(n18077), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n18063) );
  NOR2_X1 U12574 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18100), .ZN(n18084) );
  NAND2_X1 U12575 ( .A1(n18110), .A2(n18102), .ZN(n18100) );
  NOR2_X1 U12576 ( .A1(n18154), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n18129) );
  NAND2_X1 U12577 ( .A1(n18129), .A2(n18442), .ZN(n18126) );
  INV_X1 U12578 ( .A(n18176), .ZN(n18157) );
  AND3_X1 U12579 ( .A1(n9830), .A2(n9829), .A3(n9828), .ZN(n18168) );
  INV_X1 U12580 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n9828) );
  NOR2_X2 U12581 ( .A1(n20009), .A2(n18189), .ZN(n18176) );
  NOR2_X1 U12582 ( .A1(n18240), .A2(n17392), .ZN(n18246) );
  AND2_X1 U12583 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18307), .ZN(n18294) );
  NOR2_X1 U12584 ( .A1(n18320), .A2(n18335), .ZN(n18307) );
  INV_X1 U12585 ( .A(n18361), .ZN(n18337) );
  NOR2_X2 U12586 ( .A1(n13075), .A2(n13074), .ZN(n10457) );
  NOR3_X1 U12587 ( .A1(n19430), .A2(n19426), .A3(n14497), .ZN(n18468) );
  NOR2_X1 U12588 ( .A1(n18470), .A2(n10457), .ZN(n18471) );
  NAND2_X1 U12589 ( .A1(n18500), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n18495) );
  NOR2_X1 U12590 ( .A1(n18628), .A2(n18504), .ZN(n18500) );
  INV_X1 U12591 ( .A(n18511), .ZN(n18505) );
  NAND2_X1 U12592 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18505), .ZN(n18504) );
  NOR2_X1 U12593 ( .A1(n18526), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U12594 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .ZN(n9970) );
  NAND2_X1 U12595 ( .A1(n18556), .A2(n9968), .ZN(n18514) );
  AND2_X1 U12596 ( .A1(n9969), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n9968) );
  NOR2_X1 U12597 ( .A1(n18518), .A2(n18552), .ZN(n18546) );
  NAND2_X1 U12598 ( .A1(n18556), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18552) );
  NOR2_X1 U12599 ( .A1(n18560), .A2(n18730), .ZN(n18556) );
  NAND2_X1 U12600 ( .A1(n9965), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n9964) );
  INV_X1 U12601 ( .A(n18564), .ZN(n9965) );
  NAND2_X1 U12602 ( .A1(n9678), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n18560) );
  NAND2_X1 U12603 ( .A1(n18593), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n18585) );
  AND2_X1 U12604 ( .A1(n9967), .A2(n9966), .ZN(n18593) );
  NOR3_X1 U12605 ( .A1(n18590), .A2(n18660), .A3(n18663), .ZN(n9966) );
  INV_X1 U12606 ( .A(n14024), .ZN(n18594) );
  INV_X1 U12607 ( .A(n14016), .ZN(n18598) );
  NOR2_X1 U12608 ( .A1(n18679), .A2(n18619), .ZN(n18672) );
  INV_X1 U12609 ( .A(n18729), .ZN(n18718) );
  NOR2_X1 U12610 ( .A1(n18726), .A2(n19430), .ZN(n18727) );
  NOR2_X1 U12611 ( .A1(n18896), .A2(n9740), .ZN(n18842) );
  INV_X1 U12612 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18967) );
  INV_X1 U12613 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18984) );
  OR2_X1 U12614 ( .A1(n19099), .A2(n18591), .ZN(n18991) );
  INV_X2 U12615 ( .A(n18991), .ZN(n19011) );
  INV_X1 U12616 ( .A(n19479), .ZN(n19801) );
  AND2_X1 U12617 ( .A1(n17816), .A2(n19430), .ZN(n19088) );
  INV_X1 U12618 ( .A(n17816), .ZN(n17342) );
  NAND2_X1 U12619 ( .A1(n20030), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19095) );
  AND2_X1 U12620 ( .A1(n10009), .A2(n10008), .ZN(n18769) );
  INV_X1 U12621 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19217) );
  AND2_X2 U12622 ( .A1(n19269), .A2(n19314), .ZN(n19227) );
  NOR2_X1 U12623 ( .A1(n19266), .A2(n18939), .ZN(n18919) );
  NAND2_X1 U12624 ( .A1(n17302), .A2(n17301), .ZN(n18979) );
  NAND2_X1 U12625 ( .A1(n9996), .A2(n14004), .ZN(n19055) );
  NAND2_X1 U12626 ( .A1(n19067), .A2(n19066), .ZN(n9996) );
  INV_X1 U12627 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19367) );
  NAND2_X1 U12628 ( .A1(n13990), .A2(n20026), .ZN(n19390) );
  INV_X1 U12629 ( .A(n19880), .ZN(n19375) );
  INV_X1 U12630 ( .A(n19878), .ZN(n19379) );
  INV_X1 U12631 ( .A(n19389), .ZN(n19406) );
  INV_X1 U12632 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19861) );
  INV_X1 U12633 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14104) );
  INV_X1 U12634 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14130) );
  AOI211_X1 U12635 ( .C1(n20026), .C2(n19884), .A(n19425), .B(n14066), .ZN(
        n14523) );
  OR2_X1 U12636 ( .A1(n19918), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n20037) );
  AND2_X1 U12637 ( .A1(n12431), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14974)
         );
  AOI21_X1 U12639 ( .B1(n15100), .B2(n21031), .A(n12864), .ZN(n12983) );
  AOI21_X1 U12640 ( .B1(n15042), .B2(n21101), .A(n15041), .ZN(n15043) );
  NOR2_X1 U12641 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  INV_X1 U12642 ( .A(n10079), .ZN(n10078) );
  NOR2_X1 U12643 ( .A1(n14635), .A2(n15264), .ZN(n10076) );
  OAI21_X1 U12644 ( .B1(n15209), .B2(n15264), .A(n9716), .ZN(P1_U2986) );
  INV_X1 U12645 ( .A(n15213), .ZN(n9888) );
  OR2_X1 U12646 ( .A1(n15446), .A2(n20932), .ZN(n9889) );
  OAI21_X1 U12647 ( .B1(n15272), .B2(n15482), .A(n9900), .ZN(P1_U3000) );
  AOI211_X1 U12648 ( .C1(n15267), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9900)
         );
  AND2_X1 U12649 ( .A1(n15266), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9903) );
  OAI21_X1 U12650 ( .B1(n15270), .B2(n15269), .A(n15268), .ZN(n9901) );
  AND2_X1 U12651 ( .A1(n15858), .A2(n10234), .ZN(n15864) );
  AND2_X1 U12652 ( .A1(n16266), .A2(n10307), .ZN(n16268) );
  INV_X1 U12653 ( .A(n10308), .ZN(n10307) );
  NAND2_X1 U12654 ( .A1(n10159), .A2(n10157), .ZN(P2_U2857) );
  INV_X1 U12655 ( .A(n10158), .ZN(n10157) );
  NAND2_X1 U12656 ( .A1(n13601), .A2(n20108), .ZN(n10159) );
  OAI21_X1 U12657 ( .B1(n13602), .B2(n16418), .A(n13603), .ZN(n10158) );
  NAND2_X1 U12658 ( .A1(n16531), .A2(n20196), .ZN(n9816) );
  INV_X1 U12659 ( .A(n12443), .ZN(n12448) );
  NAND2_X1 U12660 ( .A1(n12444), .A2(n20196), .ZN(n12447) );
  OAI21_X1 U12661 ( .B1(n16826), .B2(n20211), .A(n11166), .ZN(n11167) );
  OAI21_X1 U12662 ( .B1(n16852), .B2(n16773), .A(n9861), .ZN(P2_U2990) );
  AOI21_X1 U12663 ( .B1(n16850), .B2(n20196), .A(n16572), .ZN(n9861) );
  OAI21_X1 U12664 ( .B1(n16864), .B2(n16773), .A(n9944), .ZN(P2_U2991) );
  AOI21_X1 U12665 ( .B1(n16862), .B2(n20196), .A(n16582), .ZN(n9944) );
  INV_X1 U12666 ( .A(n12487), .ZN(n12488) );
  NAND2_X1 U12667 ( .A1(n9820), .A2(n9819), .ZN(n9818) );
  NAND2_X1 U12668 ( .A1(n9878), .A2(n9875), .ZN(n16630) );
  AOI21_X1 U12669 ( .B1(n16913), .B2(n9877), .A(n9876), .ZN(n9875) );
  NAND2_X1 U12670 ( .A1(n9603), .A2(n9879), .ZN(n9878) );
  NAND2_X1 U12671 ( .A1(n10016), .A2(n20238), .ZN(n10015) );
  NOR2_X1 U12672 ( .A1(n9884), .A2(n9844), .ZN(n10344) );
  NAND2_X1 U12673 ( .A1(n16531), .A2(n17661), .ZN(n10017) );
  NAND2_X1 U12674 ( .A1(n9865), .A2(n12495), .ZN(n11564) );
  NAND2_X1 U12675 ( .A1(n12444), .A2(n17661), .ZN(n11565) );
  NAND2_X1 U12676 ( .A1(n9789), .A2(n12495), .ZN(n9788) );
  OAI211_X1 U12677 ( .C1(n16887), .C2(n20241), .A(n10166), .B(n10165), .ZN(
        P2_U3025) );
  NOR2_X1 U12678 ( .A1(n16884), .A2(n16885), .ZN(n10166) );
  NAND2_X1 U12679 ( .A1(n16886), .A2(n12495), .ZN(n10165) );
  OAI211_X1 U12680 ( .C1(n16908), .C2(n20241), .A(n10265), .B(n9853), .ZN(
        P2_U3028) );
  NOR2_X1 U12681 ( .A1(n16906), .A2(n10266), .ZN(n10265) );
  AND2_X1 U12682 ( .A1(n16907), .A2(n20238), .ZN(n10266) );
  AOI21_X1 U12683 ( .B1(n16920), .B2(n20238), .A(n16919), .ZN(n10091) );
  NAND2_X1 U12684 ( .A1(n16973), .A2(n9679), .ZN(n16983) );
  NAND2_X1 U12685 ( .A1(n10186), .A2(n10183), .ZN(P3_U2641) );
  NOR4_X1 U12686 ( .A1(n10185), .A2(n17838), .A3(n17837), .A4(n10184), .ZN(
        n10183) );
  NAND2_X1 U12687 ( .A1(n10187), .A2(n18097), .ZN(n10186) );
  NOR2_X1 U12688 ( .A1(n17845), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10185) );
  OAI21_X1 U12689 ( .B1(n17845), .B2(n9827), .A(n9707), .ZN(P3_U2642) );
  NOR2_X1 U12690 ( .A1(n17851), .A2(n14514), .ZN(n9827) );
  NAND2_X1 U12691 ( .A1(n9826), .A2(n9824), .ZN(n9823) );
  OR2_X1 U12692 ( .A1(n18480), .A2(n10472), .ZN(n18481) );
  AOI21_X1 U12693 ( .B1(n10277), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10276), .ZN(n10275) );
  NAND2_X1 U12694 ( .A1(n17684), .A2(n19326), .ZN(n10278) );
  OR2_X1 U12695 ( .A1(n17540), .A2(n17683), .ZN(n10276) );
  NAND2_X1 U12696 ( .A1(n10003), .A2(n10001), .ZN(P3_U2833) );
  AND2_X1 U12697 ( .A1(n10264), .A2(n9732), .ZN(n10001) );
  NAND2_X1 U12698 ( .A1(n17700), .A2(n19326), .ZN(n10003) );
  NAND2_X1 U12699 ( .A1(n19392), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9856) );
  XOR2_X2 U12700 ( .A(n13013), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n9628) );
  INV_X4 U12701 ( .A(n11312), .ZN(n11324) );
  NAND2_X1 U12702 ( .A1(n10455), .A2(n13290), .ZN(n16366) );
  NAND4_X1 U12703 ( .A1(n10609), .A2(n10592), .A3(n10624), .A4(n10593), .ZN(
        n11223) );
  NAND2_X1 U12704 ( .A1(n12554), .A2(n12507), .ZN(n12583) );
  INV_X2 U12705 ( .A(n15227), .ZN(n10334) );
  AND2_X1 U12706 ( .A1(n13277), .A2(n9770), .ZN(n13408) );
  AND3_X1 U12707 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9629) );
  INV_X2 U12708 ( .A(n10652), .ZN(n11098) );
  AND4_X1 U12709 ( .A1(n13894), .A2(n13893), .A3(n13892), .A4(n13891), .ZN(
        n9630) );
  NAND2_X1 U12710 ( .A1(n15915), .A2(n15916), .ZN(n11159) );
  NAND2_X1 U12711 ( .A1(n14712), .A2(n10304), .ZN(n14612) );
  NOR2_X1 U12712 ( .A1(n10355), .A2(n10352), .ZN(n14350) );
  OR2_X1 U12713 ( .A1(n12462), .A2(n15983), .ZN(n15962) );
  AND2_X1 U12714 ( .A1(n10338), .A2(n10476), .ZN(n9631) );
  AND4_X1 U12715 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n9632) );
  NOR2_X1 U12716 ( .A1(n10355), .A2(n10353), .ZN(n14475) );
  INV_X2 U12717 ( .A(n10593), .ZN(n9914) );
  AND2_X1 U12718 ( .A1(n12809), .A2(n10286), .ZN(n9633) );
  AND2_X1 U12719 ( .A1(n10300), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9634) );
  AND2_X1 U12720 ( .A1(n10031), .A2(n10035), .ZN(n16649) );
  OR2_X1 U12721 ( .A1(n10908), .A2(n9780), .ZN(n9635) );
  AND2_X1 U12722 ( .A1(n9677), .A2(n14726), .ZN(n9636) );
  NAND2_X1 U12723 ( .A1(n10392), .A2(n11125), .ZN(n16100) );
  NOR2_X1 U12724 ( .A1(n16344), .A2(n13409), .ZN(n16337) );
  INV_X1 U12725 ( .A(n10153), .ZN(n16358) );
  AND2_X1 U12726 ( .A1(n10035), .A2(n16650), .ZN(n9637) );
  INV_X1 U12727 ( .A(n16614), .ZN(n9955) );
  INV_X1 U12728 ( .A(n10141), .ZN(n10140) );
  AND2_X1 U12729 ( .A1(n10425), .A2(n12454), .ZN(n9638) );
  AND3_X1 U12730 ( .A1(n10856), .A2(n10855), .A3(n10857), .ZN(n9639) );
  NOR2_X1 U12731 ( .A1(n16619), .A2(n16618), .ZN(n9640) );
  NAND2_X1 U12732 ( .A1(n10442), .A2(n13352), .ZN(n16349) );
  OR2_X1 U12733 ( .A1(n10883), .A2(n11559), .ZN(n9641) );
  NAND2_X1 U12734 ( .A1(n20912), .A2(n17290), .ZN(n17246) );
  INV_X1 U12735 ( .A(n17246), .ZN(n10130) );
  NAND2_X1 U12736 ( .A1(n14095), .A2(n13263), .ZN(n16386) );
  NAND2_X1 U12737 ( .A1(n9767), .A2(n14175), .ZN(n16224) );
  AND2_X1 U12738 ( .A1(n10455), .A2(n10454), .ZN(n9642) );
  AND2_X1 U12739 ( .A1(n10381), .A2(n9764), .ZN(n9643) );
  AND2_X1 U12740 ( .A1(n9629), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9644) );
  NOR2_X1 U12741 ( .A1(n15045), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9645) );
  AND2_X1 U12742 ( .A1(n10297), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9646) );
  NAND4_X1 U12743 ( .A1(n15120), .A2(n15366), .A3(n15361), .A4(n15113), .ZN(
        n9647) );
  AND2_X1 U12744 ( .A1(n10914), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9648) );
  AND2_X1 U12745 ( .A1(n9963), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9649) );
  NOR2_X2 U12746 ( .A1(n20468), .A2(n20346), .ZN(n9650) );
  AND2_X2 U12747 ( .A1(n13554), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10765) );
  INV_X1 U12748 ( .A(n9608), .ZN(n18410) );
  AND2_X2 U12749 ( .A1(n10700), .A2(n13367), .ZN(n10758) );
  AND2_X2 U12750 ( .A1(n13568), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10743) );
  AND4_X1 U12751 ( .A1(n13890), .A2(n13889), .A3(n13888), .A4(n13887), .ZN(
        n9651) );
  NAND2_X1 U12752 ( .A1(n16937), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9652) );
  AND2_X1 U12754 ( .A1(n10067), .A2(n10139), .ZN(n9653) );
  OR2_X1 U12755 ( .A1(n10965), .A2(n10375), .ZN(n9654) );
  NOR2_X1 U12756 ( .A1(n12462), .A2(n10347), .ZN(n15945) );
  NAND2_X1 U12757 ( .A1(n14493), .A2(n14492), .ZN(n14491) );
  NOR2_X1 U12758 ( .A1(n16113), .A2(n10393), .ZN(n16087) );
  AND2_X1 U12759 ( .A1(n10990), .A2(n11000), .ZN(n10964) );
  NAND2_X1 U12760 ( .A1(n10101), .A2(n10327), .ZN(n15154) );
  NAND2_X1 U12761 ( .A1(n15897), .A2(n10357), .ZN(n9655) );
  OR2_X1 U12762 ( .A1(n17936), .A2(n18846), .ZN(n9656) );
  AND2_X1 U12763 ( .A1(n11135), .A2(n11134), .ZN(n9657) );
  AND2_X1 U12764 ( .A1(n18500), .A2(n9963), .ZN(n9658) );
  OR2_X1 U12765 ( .A1(n17064), .A2(n10883), .ZN(n9659) );
  NAND2_X1 U12766 ( .A1(n15227), .A2(n12584), .ZN(n9660) );
  NAND2_X1 U12767 ( .A1(n11025), .A2(n16681), .ZN(n10419) );
  AND2_X1 U12768 ( .A1(n10295), .A2(n10294), .ZN(n12603) );
  AND2_X1 U12769 ( .A1(n18905), .A2(n17305), .ZN(n17308) );
  AND2_X1 U12770 ( .A1(n13256), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9661) );
  NOR2_X1 U12771 ( .A1(n13203), .A2(n11178), .ZN(n13202) );
  AND2_X1 U12772 ( .A1(n12672), .A2(n10317), .ZN(n9662) );
  AND2_X1 U12773 ( .A1(n11515), .A2(n10339), .ZN(n12463) );
  NAND2_X1 U12774 ( .A1(n11515), .A2(n10341), .ZN(n16013) );
  NAND2_X1 U12775 ( .A1(n10420), .A2(n11025), .ZN(n16683) );
  OR2_X1 U12776 ( .A1(n10146), .A2(n20815), .ZN(n9664) );
  OR2_X1 U12777 ( .A1(n10146), .A2(n16721), .ZN(n9665) );
  OR2_X1 U12778 ( .A1(n10146), .A2(n16685), .ZN(n9666) );
  OR2_X1 U12779 ( .A1(n10146), .A2(n20834), .ZN(n9667) );
  OR2_X1 U12780 ( .A1(n10146), .A2(n20829), .ZN(n9668) );
  OR2_X1 U12781 ( .A1(n10146), .A2(n11346), .ZN(n9669) );
  OR2_X1 U12782 ( .A1(n10146), .A2(n20819), .ZN(n9670) );
  OR2_X1 U12783 ( .A1(n10146), .A2(n20821), .ZN(n9671) );
  OR2_X1 U12784 ( .A1(n10146), .A2(n16675), .ZN(n9672) );
  OR2_X1 U12785 ( .A1(n10146), .A2(n16643), .ZN(n9673) );
  OR2_X1 U12786 ( .A1(n10146), .A2(n20832), .ZN(n9674) );
  OR2_X1 U12787 ( .A1(n10146), .A2(n20827), .ZN(n9675) );
  OR2_X1 U12788 ( .A1(n10146), .A2(n20836), .ZN(n9676) );
  NOR2_X2 U12789 ( .A1(n13128), .A2(n13127), .ZN(n19442) );
  INV_X1 U12790 ( .A(n19442), .ZN(n13129) );
  AND2_X1 U12791 ( .A1(n12693), .A2(n12687), .ZN(n9677) );
  INV_X1 U12792 ( .A(n10419), .ZN(n10418) );
  NAND2_X1 U12793 ( .A1(n10326), .A2(n17570), .ZN(n15223) );
  NOR2_X1 U12794 ( .A1(n18585), .A2(n9964), .ZN(n9678) );
  NAND2_X1 U12795 ( .A1(n19289), .A2(n19251), .ZN(n19266) );
  AND2_X1 U12796 ( .A1(n16972), .A2(n12495), .ZN(n9679) );
  AND2_X1 U12797 ( .A1(n12820), .A2(n10297), .ZN(n9680) );
  AND4_X1 U12798 ( .A1(n13886), .A2(n13885), .A3(n13884), .A4(n13883), .ZN(
        n9681) );
  NAND2_X1 U12799 ( .A1(n10211), .A2(n16248), .ZN(n17081) );
  NOR2_X1 U12800 ( .A1(n12592), .A2(n15155), .ZN(n10476) );
  INV_X1 U12801 ( .A(n10476), .ZN(n10335) );
  NAND2_X1 U12802 ( .A1(n11077), .A2(n10369), .ZN(n9682) );
  AOI21_X1 U12803 ( .B1(n15168), .B2(n12590), .A(n12589), .ZN(n15157) );
  NOR2_X1 U12804 ( .A1(n13063), .A2(n13062), .ZN(n19426) );
  INV_X1 U12805 ( .A(n19426), .ZN(n18620) );
  NOR2_X1 U12806 ( .A1(n14687), .A2(n12986), .ZN(n14634) );
  NAND2_X1 U12807 ( .A1(n11515), .A2(n11514), .ZN(n16037) );
  INV_X2 U12808 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14056) );
  AND2_X1 U12809 ( .A1(n19053), .A2(n19354), .ZN(n9683) );
  AND2_X1 U12810 ( .A1(n16669), .A2(n10042), .ZN(n16614) );
  AND2_X1 U12811 ( .A1(n16310), .A2(n10149), .ZN(n16315) );
  NAND2_X1 U12812 ( .A1(n10652), .A2(n10926), .ZN(n10605) );
  NAND2_X1 U12813 ( .A1(n10420), .A2(n10418), .ZN(n16672) );
  AND4_X1 U12814 ( .A1(n10839), .A2(n10838), .A3(n10837), .A4(n10836), .ZN(
        n9684) );
  AND2_X1 U12815 ( .A1(n10819), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U12816 ( .A1(n14846), .A2(n10084), .ZN(n10086) );
  NOR2_X1 U12817 ( .A1(n16337), .A2(n16338), .ZN(n9686) );
  NAND2_X1 U12818 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n9687) );
  INV_X1 U12819 ( .A(n16061), .ZN(n11134) );
  AND3_X1 U12820 ( .A1(n10679), .A2(n9605), .A3(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n9688) );
  AND2_X1 U12821 ( .A1(n11108), .A2(n9664), .ZN(n9689) );
  AND2_X1 U12822 ( .A1(n11128), .A2(n9675), .ZN(n9690) );
  AND2_X1 U12823 ( .A1(n11130), .A2(n9668), .ZN(n9691) );
  AND2_X1 U12824 ( .A1(n11140), .A2(n9676), .ZN(n9692) );
  AND2_X1 U12825 ( .A1(n10332), .A2(n10331), .ZN(n15102) );
  OR2_X1 U12826 ( .A1(n10659), .A2(n11104), .ZN(n9693) );
  AND3_X1 U12827 ( .A1(n10692), .A2(n10680), .A3(n10681), .ZN(n9694) );
  AND2_X1 U12828 ( .A1(n10436), .A2(n10651), .ZN(n9695) );
  AOI21_X1 U12829 ( .B1(n13244), .B2(n13679), .A(n13243), .ZN(n13701) );
  AND3_X1 U12830 ( .A1(n10625), .A2(n10601), .A3(n17224), .ZN(n9696) );
  AND2_X1 U12831 ( .A1(n11244), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9697) );
  AND2_X1 U12832 ( .A1(n10100), .A2(n10098), .ZN(n9698) );
  AND2_X1 U12833 ( .A1(n16659), .A2(n16936), .ZN(n9699) );
  AND2_X1 U12834 ( .A1(n9806), .A2(n11019), .ZN(n9700) );
  OR2_X1 U12835 ( .A1(n13915), .A2(n13914), .ZN(n14006) );
  AND2_X1 U12836 ( .A1(n16543), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9701) );
  INV_X1 U12837 ( .A(n10223), .ZN(n15901) );
  NOR2_X1 U12838 ( .A1(n15918), .A2(n16560), .ZN(n10223) );
  AND2_X1 U12839 ( .A1(n9636), .A2(n10321), .ZN(n9702) );
  AND2_X1 U12840 ( .A1(n10331), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12841 ( .A1(n10512), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9704) );
  NAND2_X1 U12842 ( .A1(n16754), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9705) );
  INV_X1 U12843 ( .A(n10124), .ZN(n10123) );
  NAND2_X1 U12844 ( .A1(n16642), .A2(n16651), .ZN(n10124) );
  OR2_X1 U12845 ( .A1(n9652), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9706) );
  NOR2_X1 U12846 ( .A1(n17846), .A2(n9823), .ZN(n9707) );
  AND2_X1 U12847 ( .A1(n14622), .A2(n14621), .ZN(n14635) );
  OR2_X1 U12848 ( .A1(n9656), .A2(n10201), .ZN(n9708) );
  OR2_X1 U12849 ( .A1(n11054), .A2(n11045), .ZN(n9709) );
  OR2_X1 U12850 ( .A1(n9635), .A2(n10382), .ZN(n9710) );
  AND3_X1 U12851 ( .A1(n10820), .A2(n10828), .A3(n10821), .ZN(n9711) );
  OR2_X1 U12852 ( .A1(n10330), .A2(n11878), .ZN(n9712) );
  NOR2_X1 U12853 ( .A1(n10621), .A2(n17183), .ZN(n9713) );
  AND2_X1 U12854 ( .A1(n10383), .A2(n10912), .ZN(n9714) );
  NAND2_X1 U12855 ( .A1(n10380), .A2(n9643), .ZN(n9715) );
  AND2_X1 U12856 ( .A1(n9889), .A2(n9888), .ZN(n9716) );
  OR3_X1 U12857 ( .A1(n11067), .A2(n11555), .A3(n16626), .ZN(n16620) );
  INV_X1 U12858 ( .A(n10424), .ZN(n10423) );
  NAND2_X1 U12859 ( .A1(n9638), .A2(n16597), .ZN(n10424) );
  OR2_X1 U12860 ( .A1(n12455), .A2(n10426), .ZN(n9717) );
  AND2_X1 U12861 ( .A1(n14696), .A2(n14695), .ZN(n12860) );
  AND2_X1 U12862 ( .A1(n10418), .A2(n9807), .ZN(n9718) );
  AND2_X1 U12863 ( .A1(n11273), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9719) );
  AND2_X1 U12864 ( .A1(n14712), .A2(n10302), .ZN(n14596) );
  INV_X1 U12865 ( .A(n16579), .ZN(n9946) );
  NAND2_X1 U12866 ( .A1(n11086), .A2(n9741), .ZN(n10430) );
  OR2_X1 U12867 ( .A1(n16799), .A2(n20219), .ZN(n9720) );
  AND2_X1 U12868 ( .A1(n16641), .A2(n12452), .ZN(n9721) );
  INV_X1 U12869 ( .A(n9923), .ZN(n12991) );
  AND2_X1 U12870 ( .A1(n11373), .A2(n14347), .ZN(n9722) );
  AND2_X1 U12871 ( .A1(n11632), .A2(n11631), .ZN(n9723) );
  INV_X1 U12872 ( .A(n9895), .ZN(n21129) );
  OAI21_X1 U12873 ( .B1(n15342), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n9896), .ZN(n9895) );
  AND2_X1 U12874 ( .A1(n11330), .A2(n10342), .ZN(n9724) );
  AND2_X1 U12875 ( .A1(n16812), .A2(n16811), .ZN(n9725) );
  NAND2_X1 U12876 ( .A1(n17183), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20913) );
  INV_X1 U12877 ( .A(n20913), .ZN(n13680) );
  AND2_X1 U12878 ( .A1(n10863), .A2(n10862), .ZN(n9726) );
  AND2_X1 U12879 ( .A1(n10411), .A2(n16011), .ZN(n9727) );
  INV_X1 U12880 ( .A(n16586), .ZN(n10142) );
  AND2_X1 U12881 ( .A1(n9857), .A2(n9856), .ZN(n9728) );
  AND2_X1 U12882 ( .A1(n9602), .A2(n9899), .ZN(n9729) );
  AND2_X1 U12883 ( .A1(n10119), .A2(n9638), .ZN(n9730) );
  OR2_X1 U12884 ( .A1(n12540), .A2(n11809), .ZN(n9731) );
  AND2_X1 U12885 ( .A1(n10263), .A2(n10002), .ZN(n9732) );
  AND2_X1 U12886 ( .A1(n10131), .A2(n10129), .ZN(n9733) );
  AND2_X1 U12887 ( .A1(n9982), .A2(n13194), .ZN(n10222) );
  INV_X1 U12888 ( .A(n10222), .ZN(n10221) );
  OR2_X1 U12889 ( .A1(n10965), .A2(n10373), .ZN(n9734) );
  AND2_X1 U12890 ( .A1(n11877), .A2(n11896), .ZN(n9735) );
  NAND2_X1 U12891 ( .A1(n10147), .A2(n13252), .ZN(n14034) );
  AND2_X1 U12892 ( .A1(n10046), .A2(n16527), .ZN(n9736) );
  INV_X1 U12893 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16733) );
  INV_X1 U12894 ( .A(n20074), .ZN(n9810) );
  INV_X1 U12895 ( .A(n13365), .ZN(n13567) );
  INV_X1 U12896 ( .A(n10705), .ZN(n13365) );
  INV_X1 U12897 ( .A(n13432), .ZN(n10439) );
  AOI21_X1 U12898 ( .B1(n14087), .B2(n20026), .A(n14086), .ZN(n18475) );
  INV_X1 U12899 ( .A(n18475), .ZN(n9967) );
  NOR2_X1 U12900 ( .A1(n12780), .A2(n9680), .ZN(n9737) );
  NAND2_X1 U12901 ( .A1(n11563), .A2(n11562), .ZN(n20219) );
  NAND2_X1 U12902 ( .A1(n9745), .A2(n11475), .ZN(n14281) );
  NAND2_X1 U12903 ( .A1(n14348), .A2(n14347), .ZN(n14272) );
  NOR2_X2 U12904 ( .A1(n14325), .A2(n11775), .ZN(n12027) );
  INV_X1 U12905 ( .A(n12027), .ZN(n9890) );
  AND2_X1 U12906 ( .A1(n14092), .A2(n10151), .ZN(n16382) );
  INV_X1 U12907 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n9829) );
  AND2_X1 U12908 ( .A1(n16065), .A2(n10226), .ZN(n9738) );
  NAND2_X1 U12909 ( .A1(n12516), .A2(n12515), .ZN(n12548) );
  INV_X1 U12910 ( .A(n12548), .ZN(n10175) );
  NAND2_X1 U12911 ( .A1(n14203), .A2(n10410), .ZN(n16160) );
  NAND2_X1 U12912 ( .A1(n14203), .A2(n16190), .ZN(n16176) );
  AND2_X1 U12913 ( .A1(n16613), .A2(n16612), .ZN(n9739) );
  AND2_X1 U12914 ( .A1(n10676), .A2(n14039), .ZN(n10854) );
  NAND2_X1 U12915 ( .A1(n10193), .A2(n10192), .ZN(n9740) );
  OR2_X1 U12916 ( .A1(n16564), .A2(n16843), .ZN(n9741) );
  AND2_X1 U12917 ( .A1(n10334), .A2(n12594), .ZN(n9742) );
  AND2_X1 U12918 ( .A1(n14695), .A2(n12861), .ZN(n9743) );
  AND2_X1 U12919 ( .A1(n9743), .A2(n10320), .ZN(n9744) );
  NOR2_X1 U12920 ( .A1(n14258), .A2(n14268), .ZN(n14263) );
  NAND2_X1 U12921 ( .A1(n13277), .A2(n13276), .ZN(n16370) );
  INV_X1 U12922 ( .A(n16660), .ZN(n10035) );
  AND2_X1 U12923 ( .A1(n14263), .A2(n14264), .ZN(n9745) );
  INV_X1 U12924 ( .A(n9745), .ZN(n10355) );
  NAND2_X1 U12925 ( .A1(n17612), .A2(n17611), .ZN(n14494) );
  INV_X1 U12926 ( .A(n14485), .ZN(n9887) );
  OR2_X1 U12927 ( .A1(n10146), .A2(n20848), .ZN(n9746) );
  OR2_X1 U12928 ( .A1(n10146), .A2(n20851), .ZN(n9747) );
  OR2_X1 U12929 ( .A1(n10146), .A2(n16589), .ZN(n9748) );
  OR2_X1 U12930 ( .A1(n10146), .A2(n20842), .ZN(n9749) );
  OR2_X1 U12931 ( .A1(n10146), .A2(n20844), .ZN(n9750) );
  OR2_X1 U12932 ( .A1(n10146), .A2(n20853), .ZN(n9751) );
  OR2_X1 U12933 ( .A1(n10146), .A2(n12844), .ZN(n9752) );
  NAND2_X1 U12934 ( .A1(n16206), .A2(n11348), .ZN(n14344) );
  OR2_X1 U12935 ( .A1(n16227), .A2(n16226), .ZN(n14097) );
  NAND4_X1 U12936 ( .A1(n10814), .A2(n10813), .A3(n10812), .A4(n10811), .ZN(
        n10924) );
  NAND2_X1 U12937 ( .A1(n11563), .A2(n11540), .ZN(n20227) );
  INV_X1 U12938 ( .A(n13475), .ZN(n10451) );
  INV_X1 U12939 ( .A(n19006), .ZN(n18890) );
  INV_X1 U12940 ( .A(n11078), .ZN(n10370) );
  AND2_X1 U12941 ( .A1(n17239), .A2(n13640), .ZN(n9753) );
  NOR2_X1 U12942 ( .A1(n10429), .A2(n10428), .ZN(n10427) );
  INV_X1 U12943 ( .A(n10427), .ZN(n10426) );
  NOR2_X1 U12944 ( .A1(n18514), .A2(n18518), .ZN(n18510) );
  AND2_X1 U12945 ( .A1(n18804), .A2(n17316), .ZN(n9754) );
  AND2_X1 U12946 ( .A1(n11153), .A2(n9750), .ZN(n9755) );
  AND2_X1 U12947 ( .A1(n11179), .A2(n9751), .ZN(n9756) );
  AND2_X1 U12948 ( .A1(n10082), .A2(n14741), .ZN(n9757) );
  AND2_X1 U12949 ( .A1(n20273), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n9758) );
  NOR2_X1 U12950 ( .A1(n12743), .A2(n20927), .ZN(n9759) );
  NAND2_X1 U12951 ( .A1(n13277), .A2(n10154), .ZN(n10153) );
  INV_X2 U12952 ( .A(n12582), .ZN(n15227) );
  INV_X1 U12953 ( .A(n10789), .ZN(n10238) );
  AND2_X1 U12954 ( .A1(n10443), .A2(n13352), .ZN(n9760) );
  NAND2_X1 U12955 ( .A1(n20273), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n9761) );
  OR2_X1 U12956 ( .A1(n19875), .A2(n17386), .ZN(n19290) );
  NAND2_X1 U12957 ( .A1(n20273), .A2(n11032), .ZN(n9762) );
  AND2_X1 U12958 ( .A1(n18556), .A2(n9969), .ZN(n9763) );
  NAND2_X1 U12959 ( .A1(n20273), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n9764) );
  AND2_X1 U12960 ( .A1(n9744), .A2(n10319), .ZN(n9765) );
  INV_X1 U12961 ( .A(n13435), .ZN(n10452) );
  NOR3_X1 U12962 ( .A1(n10439), .A2(n13434), .A3(n16340), .ZN(n13435) );
  INV_X1 U12963 ( .A(n9891), .ZN(n15560) );
  NAND2_X1 U12964 ( .A1(n11781), .A2(n11802), .ZN(n9891) );
  INV_X1 U12965 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12781) );
  INV_X1 U12966 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20679) );
  NAND2_X1 U12967 ( .A1(n14755), .A2(n12056), .ZN(n9766) );
  AND2_X1 U12968 ( .A1(n11330), .A2(n11337), .ZN(n9767) );
  INV_X1 U12969 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20809) );
  INV_X1 U12970 ( .A(n10287), .ZN(n10286) );
  NAND2_X1 U12971 ( .A1(n10288), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U12972 ( .A1(n17302), .A2(n10281), .ZN(n9768) );
  INV_X1 U12973 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20912) );
  INV_X1 U12974 ( .A(n18735), .ZN(n10199) );
  NOR2_X1 U12975 ( .A1(n11488), .A2(n11555), .ZN(n9769) );
  AND2_X1 U12976 ( .A1(n10155), .A2(n9760), .ZN(n9770) );
  AND2_X1 U12977 ( .A1(n10789), .A2(n10139), .ZN(n9771) );
  AND2_X1 U12978 ( .A1(n9644), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9772) );
  INV_X1 U12979 ( .A(n11272), .ZN(n10061) );
  INV_X1 U12980 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17859) );
  NOR2_X2 U12981 ( .A1(n13668), .A2(n11309), .ZN(n13794) );
  INV_X1 U12982 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10189) );
  INV_X1 U12983 ( .A(n16709), .ZN(n10232) );
  INV_X1 U12984 ( .A(n10360), .ZN(n13594) );
  NAND2_X1 U12985 ( .A1(n10625), .A2(n10593), .ZN(n10360) );
  INV_X1 U12986 ( .A(n16773), .ZN(n20205) );
  OR2_X1 U12987 ( .A1(n13617), .A2(n11297), .ZN(n16773) );
  OR2_X1 U12988 ( .A1(n10146), .A2(n20858), .ZN(n9773) );
  NAND3_X1 U12989 ( .A1(n17304), .A2(n18939), .A3(n18927), .ZN(n9774) );
  NOR2_X1 U12990 ( .A1(n18941), .A2(n18943), .ZN(n17954) );
  INV_X1 U12991 ( .A(n16645), .ZN(n10227) );
  INV_X1 U12992 ( .A(n16625), .ZN(n10228) );
  NAND2_X1 U12993 ( .A1(n18764), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18731) );
  INV_X1 U12994 ( .A(n13188), .ZN(n10365) );
  INV_X1 U12995 ( .A(n11665), .ZN(n12526) );
  AND2_X1 U12996 ( .A1(n11187), .A2(n9773), .ZN(n9775) );
  OR2_X1 U12997 ( .A1(n12727), .A2(n9899), .ZN(n9776) );
  AND2_X1 U12998 ( .A1(n10280), .A2(n19287), .ZN(n9777) );
  INV_X1 U12999 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18723) );
  INV_X1 U13000 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13231) );
  NOR2_X1 U13001 ( .A1(n16773), .A2(n9882), .ZN(n9778) );
  AND2_X1 U13002 ( .A1(n11097), .A2(n11297), .ZN(n20196) );
  AND2_X1 U13003 ( .A1(n18764), .A2(n9629), .ZN(n9779) );
  INV_X1 U13004 ( .A(n20927), .ZN(n13624) );
  INV_X1 U13005 ( .A(n9628), .ZN(n10198) );
  INV_X1 U13006 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16557) );
  INV_X1 U13007 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21369) );
  NAND2_X1 U13008 ( .A1(n10388), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10384) );
  INV_X1 U13009 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10094) );
  INV_X1 U13010 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10273) );
  AND2_X1 U13011 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18133) );
  NAND4_X1 U13012 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9780) );
  NAND2_X1 U13013 ( .A1(n17954), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18896) );
  OR2_X1 U13014 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9781) );
  NAND3_X1 U13015 ( .A1(n15159), .A2(n15408), .A3(n15395), .ZN(n9782) );
  INV_X1 U13016 ( .A(n10386), .ZN(n10385) );
  NAND2_X1 U13017 ( .A1(n10388), .A2(n10387), .ZN(n10386) );
  AND2_X1 U13018 ( .A1(n12762), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9783) );
  AND2_X1 U13019 ( .A1(n18963), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18052) );
  INV_X1 U13020 ( .A(n10259), .ZN(n10258) );
  NOR2_X1 U13021 ( .A1(n10260), .A2(n17304), .ZN(n10259) );
  AND2_X1 U13022 ( .A1(n9648), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9784) );
  INV_X1 U13023 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10389) );
  INV_X1 U13024 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10282) );
  INV_X1 U13025 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n9830) );
  INV_X1 U13026 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10268) );
  INV_X1 U13027 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10376) );
  INV_X1 U13028 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10406) );
  AND2_X1 U13029 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9785) );
  INV_X1 U13030 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10301) );
  INV_X1 U13031 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10298) );
  INV_X1 U13032 ( .A(n10403), .ZN(n10402) );
  NAND2_X1 U13033 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  INV_X1 U13034 ( .A(n10073), .ZN(n10072) );
  NAND2_X1 U13035 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10073) );
  AND2_X1 U13036 ( .A1(n10405), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9786) );
  INV_X1 U13037 ( .A(n20128), .ZN(n20138) );
  OAI22_X1 U13038 ( .A1(n20681), .A2(n20716), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n20687), .ZN(n20723) );
  OAI21_X1 U13039 ( .B1(n10819), .B2(n20372), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20356) );
  NAND3_X1 U13040 ( .A1(n17290), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17677) );
  AOI211_X1 U13041 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16265), .B(n16264), .ZN(n16266) );
  INV_X1 U13042 ( .A(n16275), .ZN(n20092) );
  NOR4_X2 U13043 ( .A1(n14498), .A2(n18470), .A3(n18450), .A4(n18438), .ZN(
        n18436) );
  INV_X1 U13044 ( .A(n18468), .ZN(n18470) );
  NOR2_X4 U13045 ( .A1(n21476), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21439) );
  NOR2_X1 U13046 ( .A1(n20273), .A2(n20280), .ZN(n9787) );
  INV_X4 U13047 ( .A(n9914), .ZN(n20273) );
  NAND3_X1 U13048 ( .A1(n16813), .A2(n9788), .A3(n9725), .ZN(P2_U3019) );
  AND2_X2 U13049 ( .A1(n10815), .A2(n9604), .ZN(n10478) );
  AND3_X2 U13050 ( .A1(n9832), .A2(n10067), .A3(n10138), .ZN(n10848) );
  OAI21_X1 U13051 ( .B1(n11223), .B2(n11218), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9988) );
  NAND2_X1 U13052 ( .A1(n10594), .A2(n11223), .ZN(n10632) );
  NAND2_X2 U13053 ( .A1(n9790), .A2(n9710), .ZN(n16579) );
  NAND2_X2 U13054 ( .A1(n9792), .A2(n9791), .ZN(n9984) );
  NAND3_X1 U13055 ( .A1(n10636), .A2(n12775), .A3(n10605), .ZN(n10616) );
  NAND3_X1 U13056 ( .A1(n10605), .A2(n12775), .A3(n10614), .ZN(n10615) );
  XNOR2_X2 U13057 ( .A(n9868), .B(n9794), .ZN(n13719) );
  NAND3_X2 U13058 ( .A1(n9796), .A2(n9797), .A3(n9659), .ZN(n9883) );
  NAND2_X1 U13059 ( .A1(n10880), .A2(n9848), .ZN(n9796) );
  NAND3_X1 U13060 ( .A1(n17063), .A2(n10951), .A3(n17064), .ZN(n9797) );
  AND2_X1 U13061 ( .A1(n9986), .A2(n20205), .ZN(n9985) );
  NAND2_X1 U13062 ( .A1(n16579), .A2(n9648), .ZN(n9987) );
  NAND2_X1 U13063 ( .A1(n9801), .A2(n10245), .ZN(n9800) );
  NOR2_X1 U13064 ( .A1(n10663), .A2(n9803), .ZN(n9801) );
  INV_X1 U13065 ( .A(n10661), .ZN(n9803) );
  NAND2_X1 U13066 ( .A1(n11102), .A2(n9805), .ZN(n16227) );
  NAND3_X1 U13067 ( .A1(n16798), .A2(n16797), .A3(n9720), .ZN(P2_U3018) );
  NAND3_X1 U13068 ( .A1(n9813), .A2(n9641), .A3(n9812), .ZN(n10045) );
  NAND2_X1 U13069 ( .A1(n10882), .A2(n11555), .ZN(n9812) );
  NAND2_X1 U13070 ( .A1(n9939), .A2(n9814), .ZN(n9813) );
  OAI21_X1 U13071 ( .B1(n16561), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16543), .ZN(n16823) );
  NOR2_X2 U13072 ( .A1(n16571), .A2(n16830), .ZN(n16561) );
  OR2_X2 U13073 ( .A1(n16823), .A2(n20219), .ZN(n16824) );
  NAND3_X1 U13074 ( .A1(n9816), .A2(n16532), .A3(n9815), .ZN(P2_U2983) );
  OAI21_X1 U13075 ( .B1(n9834), .B2(n9701), .A(n20205), .ZN(n9815) );
  NAND3_X1 U13076 ( .A1(n12500), .A2(n16534), .A3(n12499), .ZN(n9817) );
  XNOR2_X2 U13077 ( .A(n10882), .B(n10883), .ZN(n10951) );
  NAND2_X2 U13078 ( .A1(n10848), .A2(n10849), .ZN(n10882) );
  OAI211_X1 U13079 ( .C1(n16898), .C2(n20211), .A(n9818), .B(n9640), .ZN(
        P2_U2995) );
  NAND2_X1 U13080 ( .A1(n16669), .A2(n9786), .ZN(n16913) );
  NAND2_X2 U13081 ( .A1(n9822), .A2(n9635), .ZN(n16669) );
  NAND2_X2 U13082 ( .A1(n16669), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16583) );
  NAND2_X1 U13083 ( .A1(n9849), .A2(n10951), .ZN(n9870) );
  NAND2_X1 U13084 ( .A1(n9832), .A2(n10789), .ZN(n9915) );
  NAND3_X1 U13085 ( .A1(n10067), .A2(n9832), .A3(n9771), .ZN(n10095) );
  NAND4_X1 U13086 ( .A1(n10043), .A2(n10070), .A3(n10128), .A4(n10731), .ZN(
        n9832) );
  OAI21_X1 U13087 ( .B1(n16543), .B2(n9839), .A(n9837), .ZN(n9836) );
  NAND4_X1 U13088 ( .A1(n9726), .A2(n9639), .A3(n10858), .A4(n10861), .ZN(
        n9845) );
  NAND4_X1 U13089 ( .A1(n9711), .A2(n10018), .A3(n10823), .A4(n10826), .ZN(
        n9846) );
  NAND3_X1 U13090 ( .A1(n9694), .A2(n10036), .A3(n10037), .ZN(n10067) );
  NAND2_X1 U13091 ( .A1(n9847), .A2(n19037), .ZN(n19036) );
  OAI21_X1 U13092 ( .B1(n19037), .B2(n9847), .A(n19036), .ZN(n19342) );
  NAND2_X1 U13093 ( .A1(n17063), .A2(n17064), .ZN(n9849) );
  NOR2_X2 U13094 ( .A1(n19266), .A2(n10258), .ZN(n19158) );
  NAND3_X1 U13095 ( .A1(n9881), .A2(n16627), .A3(n12495), .ZN(n9853) );
  NAND2_X1 U13096 ( .A1(n18611), .A2(n13905), .ZN(n9854) );
  OR2_X2 U13097 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  NAND2_X1 U13098 ( .A1(n16579), .A2(n9863), .ZN(n9866) );
  NAND4_X1 U13099 ( .A1(n9867), .A2(n10591), .A3(n11244), .A4(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10239) );
  INV_X1 U13100 ( .A(n10621), .ZN(n9867) );
  NAND2_X1 U13101 ( .A1(n13719), .A2(n13679), .ZN(n13239) );
  NAND2_X1 U13102 ( .A1(n10683), .A2(n10666), .ZN(n10246) );
  NAND2_X1 U13103 ( .A1(n10881), .A2(n9870), .ZN(n16753) );
  AND2_X2 U13104 ( .A1(n10603), .A2(n9872), .ZN(n11213) );
  NAND3_X1 U13105 ( .A1(n10622), .A2(n10603), .A3(n9871), .ZN(n10131) );
  AND2_X1 U13106 ( .A1(n9872), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9871) );
  NAND2_X1 U13107 ( .A1(n9696), .A2(n9874), .ZN(n9873) );
  INV_X1 U13108 ( .A(n10607), .ZN(n9874) );
  NAND2_X1 U13109 ( .A1(n9883), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10881) );
  XNOR2_X1 U13110 ( .A(n9883), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17059) );
  INV_X1 U13111 ( .A(n13229), .ZN(n10624) );
  NOR2_X2 U13112 ( .A1(n10593), .A2(n13229), .ZN(n10606) );
  NAND2_X1 U13113 ( .A1(n10593), .A2(n13229), .ZN(n10607) );
  NAND2_X2 U13114 ( .A1(n9910), .A2(n9912), .ZN(n13229) );
  INV_X1 U13115 ( .A(n11194), .ZN(n10623) );
  NAND3_X1 U13116 ( .A1(n9736), .A2(n9886), .A3(n9885), .ZN(n9884) );
  NAND4_X1 U13117 ( .A1(n16776), .A2(n12779), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9885) );
  NAND2_X2 U13118 ( .A1(n9600), .A2(n9887), .ZN(n15027) );
  NAND2_X1 U13119 ( .A1(n12620), .A2(n12619), .ZN(n9894) );
  NAND2_X1 U13120 ( .A1(n12402), .A2(n9898), .ZN(n9897) );
  AND2_X1 U13121 ( .A1(n11662), .A2(n9899), .ZN(n10492) );
  AND3_X1 U13122 ( .A1(n14569), .A2(n9899), .A3(n14325), .ZN(n12855) );
  NAND2_X1 U13123 ( .A1(n12612), .A2(n9899), .ZN(n12409) );
  AOI21_X1 U13124 ( .B1(n12572), .B2(n9899), .A(n21369), .ZN(n11786) );
  NAND2_X2 U13125 ( .A1(n9908), .A2(n12406), .ZN(n17532) );
  INV_X1 U13126 ( .A(n12608), .ZN(n9907) );
  NAND2_X1 U13127 ( .A1(n9909), .A2(n12404), .ZN(n9908) );
  NAND3_X1 U13128 ( .A1(n12400), .A2(n12398), .A3(n12399), .ZN(n9909) );
  NAND3_X1 U13129 ( .A1(n9913), .A2(n10505), .A3(n10507), .ZN(n9912) );
  XNOR2_X2 U13130 ( .A(n9653), .B(n9915), .ZN(n17105) );
  NAND2_X1 U13131 ( .A1(n16579), .A2(n9784), .ZN(n13210) );
  NAND2_X1 U13132 ( .A1(n9984), .A2(n10907), .ZN(n16748) );
  NOR2_X1 U13133 ( .A1(n16727), .A2(n16720), .ZN(n16719) );
  AND2_X1 U13134 ( .A1(n9955), .A2(n9920), .ZN(n16896) );
  NAND3_X1 U13135 ( .A1(n9921), .A2(n11709), .A3(n21369), .ZN(n10075) );
  OR2_X1 U13136 ( .A1(n9921), .A2(n14292), .ZN(n13838) );
  NAND2_X1 U13137 ( .A1(n9921), .A2(n11709), .ZN(n14232) );
  NAND3_X1 U13138 ( .A1(n15084), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n9922), .ZN(n15069) );
  NOR2_X2 U13139 ( .A1(n12992), .A2(n9742), .ZN(n15077) );
  AND2_X2 U13140 ( .A1(n9923), .A2(n10334), .ZN(n12992) );
  NAND2_X2 U13141 ( .A1(n12595), .A2(n15103), .ZN(n9923) );
  OAI21_X1 U13142 ( .B1(n15272), .B2(n20932), .A(n15043), .ZN(P1_U2968) );
  NAND3_X1 U13143 ( .A1(n9924), .A2(n9925), .A3(n9930), .ZN(n15272) );
  NAND3_X1 U13144 ( .A1(n9928), .A2(n9927), .A3(n9931), .ZN(n9924) );
  NAND2_X1 U13145 ( .A1(n15038), .A2(n9926), .ZN(n9925) );
  NAND3_X1 U13146 ( .A1(n15036), .A2(n15037), .A3(n9645), .ZN(n9927) );
  NAND2_X1 U13147 ( .A1(n15038), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9928) );
  NAND3_X1 U13148 ( .A1(n15036), .A2(n15037), .A3(n9929), .ZN(n9930) );
  INV_X1 U13149 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9931) );
  NAND3_X1 U13150 ( .A1(n10634), .A2(n9941), .A3(n10635), .ZN(n10665) );
  INV_X1 U13151 ( .A(n10905), .ZN(n9943) );
  AOI21_X1 U13152 ( .B1(n16641), .B2(n10427), .A(n9954), .ZN(n16622) );
  NOR2_X2 U13153 ( .A1(n13147), .A2(n9962), .ZN(n13964) );
  INV_X1 U13154 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n9971) );
  NAND3_X1 U13155 ( .A1(n13963), .A2(n9973), .A3(n9972), .ZN(n13965) );
  NAND2_X2 U13156 ( .A1(n9976), .A2(n9762), .ZN(n11054) );
  NOR2_X2 U13157 ( .A1(n10973), .A2(n9978), .ZN(n10990) );
  NOR2_X1 U13158 ( .A1(n10688), .A2(n20243), .ZN(n10127) );
  NOR2_X2 U13159 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10700) );
  AOI21_X2 U13160 ( .B1(n11241), .B2(n10613), .A(n9988), .ZN(n10636) );
  NOR2_X1 U13161 ( .A1(n20133), .A2(n9989), .ZN(n14165) );
  NAND2_X1 U13162 ( .A1(n10561), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10562) );
  NAND2_X2 U13163 ( .A1(n10337), .A2(n9631), .ZN(n15116) );
  NAND2_X1 U13164 ( .A1(n14213), .A2(n21369), .ZN(n11822) );
  NOR2_X1 U13165 ( .A1(n10099), .A2(n9782), .ZN(n10098) );
  NAND2_X1 U13166 ( .A1(n11685), .A2(n14294), .ZN(n10324) );
  NAND2_X1 U13167 ( .A1(n15068), .A2(n12766), .ZN(n15036) );
  NAND2_X1 U13168 ( .A1(n10075), .A2(n9731), .ZN(n11723) );
  NAND2_X2 U13169 ( .A1(n10599), .A2(n10598), .ZN(n10652) );
  AOI211_X1 U13170 ( .C1(n17661), .C2(n16930), .A(n16929), .B(n16928), .ZN(
        n16931) );
  NAND2_X1 U13171 ( .A1(n10066), .A2(n11226), .ZN(n10065) );
  NOR2_X1 U13172 ( .A1(n10604), .A2(n20912), .ZN(n10597) );
  NAND2_X1 U13173 ( .A1(n15068), .A2(n10112), .ZN(n10114) );
  NAND2_X1 U13174 ( .A1(n17584), .A2(n17585), .ZN(n17583) );
  NAND2_X1 U13175 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  AND2_X1 U13176 ( .A1(n10514), .A2(n10513), .ZN(n10417) );
  NAND3_X1 U13177 ( .A1(n9995), .A2(n10417), .A3(n9704), .ZN(n9993) );
  INV_X1 U13178 ( .A(n10114), .ZN(n15038) );
  NAND2_X1 U13179 ( .A1(n11724), .A2(n21169), .ZN(n14900) );
  NAND2_X1 U13180 ( .A1(n19029), .A2(n19028), .ZN(n9991) );
  NAND2_X1 U13181 ( .A1(n19042), .A2(n14013), .ZN(n9992) );
  NAND2_X1 U13182 ( .A1(n10416), .A2(n10415), .ZN(n9994) );
  NAND2_X1 U13183 ( .A1(n19078), .A2(n19077), .ZN(n14002) );
  NAND2_X1 U13184 ( .A1(n19085), .A2(n13998), .ZN(n19077) );
  NAND2_X1 U13185 ( .A1(n19093), .A2(n19086), .ZN(n19085) );
  XNOR2_X2 U13186 ( .A(n18611), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19086) );
  XNOR2_X1 U13187 ( .A(n13999), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19078) );
  NAND2_X4 U13188 ( .A1(n9651), .A2(n9630), .ZN(n18611) );
  INV_X1 U13189 ( .A(n18781), .ZN(n10009) );
  NAND3_X1 U13190 ( .A1(n10009), .A2(n10008), .A3(n19110), .ZN(n10004) );
  NAND2_X1 U13191 ( .A1(n10013), .A2(n18890), .ZN(n10011) );
  INV_X1 U13192 ( .A(n10013), .ZN(n10012) );
  OAI21_X2 U13193 ( .B1(n18952), .B2(n9774), .A(n19006), .ZN(n17309) );
  NAND3_X1 U13194 ( .A1(n10344), .A2(n10017), .A3(n10015), .ZN(P2_U3015) );
  OAI21_X1 U13195 ( .B1(n10951), .B2(n10021), .A(n10019), .ZN(n10208) );
  NAND2_X1 U13196 ( .A1(n16573), .A2(n16586), .ZN(n10027) );
  AOI22_X1 U13197 ( .A1(n10030), .A2(n10690), .B1(n20316), .B2(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10029) );
  AND2_X1 U13198 ( .A1(n9614), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10030) );
  INV_X1 U13199 ( .A(n20677), .ZN(n20684) );
  NAND2_X1 U13200 ( .A1(n10690), .A2(n14039), .ZN(n20677) );
  NAND3_X1 U13201 ( .A1(n16694), .A2(n16699), .A3(n16767), .ZN(n10126) );
  INV_X1 U13202 ( .A(n11270), .ZN(n10060) );
  INV_X2 U13203 ( .A(n11268), .ZN(n11563) );
  NAND3_X1 U13204 ( .A1(n10064), .A2(n10063), .A3(n11257), .ZN(n10062) );
  NAND2_X1 U13205 ( .A1(n11260), .A2(n11259), .ZN(n10646) );
  NAND2_X2 U13206 ( .A1(n11213), .A2(n10622), .ZN(n11260) );
  NAND2_X1 U13207 ( .A1(n16669), .A2(n10072), .ZN(n16659) );
  AND2_X1 U13208 ( .A1(n16669), .A2(n10071), .ZN(n16602) );
  NAND2_X1 U13209 ( .A1(n14255), .A2(n10074), .ZN(n14388) );
  XNOR2_X1 U13210 ( .A(n14255), .B(n10074), .ZN(n14898) );
  NAND2_X1 U13211 ( .A1(n10077), .A2(n14636), .ZN(n15079) );
  NAND2_X1 U13212 ( .A1(n10077), .A2(n10076), .ZN(n10081) );
  NAND2_X1 U13213 ( .A1(n10081), .A2(n10078), .ZN(P1_U2973) );
  INV_X1 U13214 ( .A(n10086), .ZN(n14770) );
  NAND2_X1 U13215 ( .A1(n10095), .A2(n11338), .ZN(n10815) );
  NOR2_X4 U13216 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14245) );
  NAND3_X1 U13217 ( .A1(n10338), .A2(n10337), .A3(n10171), .ZN(n10096) );
  XNOR2_X1 U13218 ( .A(n10097), .B(n11802), .ZN(n12539) );
  XNOR2_X2 U13219 ( .A(n11723), .B(n11722), .ZN(n10097) );
  INV_X1 U13220 ( .A(n12561), .ZN(n10099) );
  NAND2_X1 U13221 ( .A1(n10104), .A2(n10103), .ZN(n10101) );
  NAND2_X1 U13222 ( .A1(n10104), .A2(n9698), .ZN(n10102) );
  INV_X1 U13223 ( .A(n10107), .ZN(n21097) );
  NAND3_X1 U13224 ( .A1(n10109), .A2(n12549), .A3(n10106), .ZN(n17584) );
  NAND2_X1 U13225 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U13226 ( .A1(n12524), .A2(n12523), .ZN(n10107) );
  INV_X1 U13227 ( .A(n12550), .ZN(n10108) );
  NAND3_X1 U13228 ( .A1(n14479), .A2(n10174), .A3(n10110), .ZN(n10109) );
  NAND2_X1 U13229 ( .A1(n12524), .A2(n10173), .ZN(n10110) );
  AND2_X2 U13230 ( .A1(n14224), .A2(n11574), .ZN(n12201) );
  AND2_X2 U13231 ( .A1(n10111), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14224) );
  OR2_X2 U13232 ( .A1(n11657), .A2(n11662), .ZN(n15500) );
  NAND3_X1 U13233 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A3(
        n9613), .ZN(n10118) );
  NAND3_X1 U13234 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A3(
        n14039), .ZN(n10117) );
  NAND2_X1 U13235 ( .A1(n10120), .A2(n9730), .ZN(n16599) );
  NAND2_X1 U13236 ( .A1(n16649), .A2(n10121), .ZN(n10120) );
  NAND2_X2 U13237 ( .A1(n11007), .A2(n11006), .ZN(n16767) );
  INV_X1 U13238 ( .A(n10726), .ZN(n10128) );
  NAND2_X1 U13239 ( .A1(n10414), .A2(n10644), .ZN(n10132) );
  INV_X1 U13240 ( .A(n10414), .ZN(n10683) );
  NAND2_X1 U13241 ( .A1(n10144), .A2(n14056), .ZN(n10133) );
  NAND2_X1 U13242 ( .A1(n10145), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10134) );
  AND2_X4 U13243 ( .A1(n10708), .A2(n17248), .ZN(n10705) );
  AND2_X2 U13244 ( .A1(n10137), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10708) );
  INV_X1 U13245 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10137) );
  OAI21_X2 U13246 ( .B1(n11076), .B2(n10142), .A(n16585), .ZN(n10141) );
  NAND4_X1 U13247 ( .A1(n10579), .A2(n10580), .A3(n10578), .A4(n10577), .ZN(
        n10144) );
  NAND4_X1 U13248 ( .A1(n10583), .A2(n10584), .A3(n10582), .A4(n10581), .ZN(
        n10145) );
  NAND2_X1 U13249 ( .A1(n13717), .A2(n10148), .ZN(n10147) );
  NAND3_X1 U13250 ( .A1(n10149), .A2(n16310), .A3(n16317), .ZN(n16316) );
  AOI21_X2 U13251 ( .B1(n16316), .B2(n16310), .A(n13545), .ZN(n16305) );
  NAND2_X1 U13252 ( .A1(n14033), .A2(n10444), .ZN(n14092) );
  NOR2_X2 U13253 ( .A1(n14039), .A2(n10677), .ZN(n10819) );
  INV_X1 U13254 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10164) );
  AND2_X4 U13255 ( .A1(n17158), .A2(n10926), .ZN(n10699) );
  NAND2_X1 U13256 ( .A1(n14309), .A2(n10169), .ZN(n11632) );
  OAI21_X1 U13257 ( .B1(n14541), .B2(n10169), .A(n12359), .ZN(n10168) );
  AOI21_X1 U13258 ( .B1(n12733), .B2(n10169), .A(n12732), .ZN(n12735) );
  NAND2_X1 U13259 ( .A1(n10170), .A2(n12621), .ZN(n17514) );
  NAND2_X1 U13260 ( .A1(n12613), .A2(n14546), .ZN(n12418) );
  NOR2_X2 U13261 ( .A1(n11658), .A2(n12411), .ZN(n12613) );
  NAND2_X1 U13262 ( .A1(n10249), .A2(n11834), .ZN(n10330) );
  NAND2_X1 U13263 ( .A1(n14193), .A2(n12547), .ZN(n14479) );
  INV_X1 U13264 ( .A(n12992), .ZN(n15085) );
  NOR2_X1 U13265 ( .A1(n12992), .A2(n10176), .ZN(n12994) );
  NAND2_X1 U13266 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  INV_X1 U13267 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10179) );
  AND4_X2 U13268 ( .A1(n10179), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11625) );
  INV_X1 U13269 ( .A(n18896), .ZN(n10190) );
  NAND2_X1 U13270 ( .A1(n10190), .A2(n10191), .ZN(n18812) );
  OAI22_X1 U13271 ( .A1(n17872), .A2(n10195), .B1(n18735), .B2(n10196), .ZN(
        n17852) );
  NAND2_X1 U13272 ( .A1(n9628), .A2(n10203), .ZN(n10202) );
  INV_X1 U13273 ( .A(n10206), .ZN(n17944) );
  NAND2_X1 U13274 ( .A1(n10215), .A2(n10219), .ZN(n16535) );
  NAND2_X1 U13275 ( .A1(n11087), .A2(n10220), .ZN(n10215) );
  OAI21_X1 U13276 ( .B1(n10217), .B2(n10220), .A(n16534), .ZN(n10216) );
  OAI21_X2 U13277 ( .B1(n15888), .B2(n20080), .A(n16549), .ZN(n15872) );
  NAND2_X1 U13278 ( .A1(n16065), .A2(n10225), .ZN(n16020) );
  AND3_X2 U13279 ( .A1(n10241), .A2(n10240), .A3(n10239), .ZN(n10637) );
  NAND3_X1 U13280 ( .A1(n11251), .A2(n10575), .A3(n13680), .ZN(n10240) );
  XNOR2_X2 U13281 ( .A(n11101), .B(n10242), .ZN(n13223) );
  NAND3_X1 U13282 ( .A1(n10244), .A2(n10246), .A3(n10247), .ZN(n10243) );
  NAND2_X1 U13283 ( .A1(n11185), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10245) );
  NAND2_X1 U13284 ( .A1(n11834), .A2(n14336), .ZN(n11857) );
  NAND2_X1 U13285 ( .A1(n12595), .A2(n10250), .ZN(n15053) );
  INV_X1 U13286 ( .A(n19266), .ZN(n10256) );
  NAND2_X1 U13287 ( .A1(n10256), .A2(n10257), .ZN(n17697) );
  NAND3_X1 U13288 ( .A1(n18806), .A2(n18793), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17317) );
  NAND3_X1 U13289 ( .A1(n18806), .A2(n18793), .A3(n10270), .ZN(n10269) );
  NAND2_X2 U13290 ( .A1(n10274), .A2(n17300), .ZN(n18905) );
  NAND2_X1 U13291 ( .A1(n10278), .A2(n10275), .ZN(P3_U2832) );
  NAND2_X1 U13292 ( .A1(n17541), .A2(n17542), .ZN(n10277) );
  NAND2_X2 U13293 ( .A1(n17302), .A2(n9777), .ZN(n18952) );
  OAI21_X1 U13294 ( .B1(n12539), .B2(n11778), .A(n10283), .ZN(n14199) );
  INV_X1 U13295 ( .A(n15027), .ZN(n10291) );
  NAND3_X1 U13296 ( .A1(n14492), .A2(n10291), .A3(n10292), .ZN(n14858) );
  NAND3_X1 U13297 ( .A1(n10295), .A2(n10294), .A3(n14304), .ZN(n11674) );
  NAND2_X1 U13298 ( .A1(n12820), .A2(n10296), .ZN(n12824) );
  NAND2_X1 U13299 ( .A1(n12802), .A2(n10299), .ZN(n12794) );
  NAND2_X1 U13300 ( .A1(n16273), .A2(n20083), .ZN(n16297) );
  NOR2_X2 U13301 ( .A1(n14948), .A2(n10315), .ZN(n14940) );
  NAND2_X1 U13302 ( .A1(n14580), .A2(n11665), .ZN(n12734) );
  NAND2_X2 U13303 ( .A1(n12637), .A2(n12626), .ZN(n14580) );
  NAND3_X1 U13304 ( .A1(n11683), .A2(n12734), .A3(n11666), .ZN(n11667) );
  NAND2_X1 U13305 ( .A1(n14541), .A2(n14542), .ZN(n12730) );
  NAND2_X1 U13306 ( .A1(n10325), .A2(n17570), .ZN(n10329) );
  NAND2_X1 U13307 ( .A1(n15116), .A2(n15146), .ZN(n15115) );
  NAND2_X1 U13308 ( .A1(n14348), .A2(n9722), .ZN(n14271) );
  INV_X1 U13309 ( .A(n14271), .ZN(n11394) );
  NOR2_X2 U13310 ( .A1(n12462), .A2(n10345), .ZN(n15930) );
  NAND2_X1 U13311 ( .A1(n9745), .A2(n10350), .ZN(n16045) );
  NAND3_X1 U13312 ( .A1(n11475), .A2(n10354), .A3(n14476), .ZN(n10353) );
  AND2_X1 U13313 ( .A1(n15897), .A2(n11532), .ZN(n15882) );
  NAND2_X1 U13314 ( .A1(n11543), .A2(n13188), .ZN(n13191) );
  NAND2_X1 U13315 ( .A1(n11543), .A2(n10364), .ZN(n10366) );
  NAND2_X1 U13316 ( .A1(n11545), .A2(n10366), .ZN(n15877) );
  INV_X1 U13317 ( .A(n11054), .ZN(n10380) );
  OAI211_X2 U13318 ( .C1(n17060), .C2(n9663), .A(n10852), .B(n17062), .ZN(
        n17063) );
  AND2_X1 U13319 ( .A1(n15932), .A2(n15933), .ZN(n15915) );
  NAND2_X1 U13320 ( .A1(n15932), .A2(n10395), .ZN(n13203) );
  AND2_X1 U13321 ( .A1(n15932), .A2(n10396), .ZN(n11171) );
  AND2_X1 U13322 ( .A1(n10397), .A2(n15933), .ZN(n10396) );
  AND2_X2 U13323 ( .A1(n11135), .A2(n9727), .ZN(n12458) );
  OAI21_X1 U13324 ( .B1(n10664), .B2(n10665), .A(n10414), .ZN(n13245) );
  NAND2_X1 U13325 ( .A1(n10432), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10431) );
  NAND4_X1 U13326 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10432) );
  NAND2_X1 U13327 ( .A1(n10434), .A2(n14056), .ZN(n10433) );
  NAND4_X1 U13328 ( .A1(n10569), .A2(n10567), .A3(n10566), .A4(n10568), .ZN(
        n10434) );
  NAND3_X1 U13329 ( .A1(n10653), .A2(n10437), .A3(n10436), .ZN(n10654) );
  NAND4_X1 U13330 ( .A1(n10435), .A2(n10653), .A3(n9695), .A4(n10437), .ZN(
        n10657) );
  NAND2_X1 U13331 ( .A1(n10658), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U13332 ( .A1(n16353), .A2(n10439), .ZN(n10438) );
  OAI211_X1 U13333 ( .C1(n16353), .C2(n10441), .A(n10440), .B(n10438), .ZN(
        n16343) );
  INV_X1 U13334 ( .A(n16344), .ZN(n10446) );
  NAND2_X1 U13335 ( .A1(n10450), .A2(n10449), .ZN(n13476) );
  NAND2_X1 U13336 ( .A1(n10450), .A2(n10448), .ZN(n16322) );
  NAND2_X1 U13337 ( .A1(n17491), .A2(n17322), .ZN(n17537) );
  OR2_X1 U13338 ( .A1(n12583), .A2(n15435), .ZN(n12586) );
  INV_X1 U13339 ( .A(n12583), .ZN(n12582) );
  CLKBUF_X1 U13340 ( .A(n14479), .Z(n21096) );
  XNOR2_X1 U13341 ( .A(n13663), .B(n13249), .ZN(n13702) );
  NAND2_X1 U13342 ( .A1(n14196), .A2(n11801), .ZN(n14255) );
  AND2_X1 U13343 ( .A1(n14335), .A2(n15526), .ZN(n15719) );
  CLKBUF_X1 U13344 ( .A(n16748), .Z(n17033) );
  NAND2_X1 U13345 ( .A1(n11306), .A2(n11305), .ZN(n11311) );
  NAND2_X1 U13346 ( .A1(n11800), .A2(n11799), .ZN(n14196) );
  INV_X1 U13347 ( .A(n14198), .ZN(n11799) );
  INV_X1 U13348 ( .A(n14199), .ZN(n11800) );
  CLKBUF_X1 U13349 ( .A(n13719), .Z(n17168) );
  OR2_X1 U13350 ( .A1(n13719), .A2(n10673), .ZN(n10677) );
  OR2_X1 U13351 ( .A1(n13719), .A2(n10669), .ZN(n10675) );
  INV_X1 U13352 ( .A(n14336), .ZN(n14337) );
  AND2_X1 U13353 ( .A1(n14285), .A2(n14336), .ZN(n15803) );
  CLKBUF_X1 U13354 ( .A(n14258), .Z(n14267) );
  NAND2_X1 U13355 ( .A1(n11790), .A2(n21369), .ZN(n11770) );
  INV_X1 U13356 ( .A(n11171), .ZN(n15886) );
  XNOR2_X1 U13357 ( .A(n11744), .B(n11743), .ZN(n11790) );
  NAND2_X1 U13358 ( .A1(n11679), .A2(n11678), .ZN(n11744) );
  INV_X1 U13359 ( .A(n14773), .ZN(n14802) );
  XNOR2_X1 U13360 ( .A(n12598), .B(n12597), .ZN(n13222) );
  NOR2_X1 U13361 ( .A1(n14579), .A2(n14576), .ZN(n12641) );
  NAND2_X1 U13362 ( .A1(n10882), .A2(n10851), .ZN(n10853) );
  NOR2_X1 U13363 ( .A1(n11314), .A2(n10954), .ZN(n10981) );
  NAND2_X1 U13364 ( .A1(n12457), .A2(n15985), .ZN(n15966) );
  NAND2_X1 U13365 ( .A1(n10610), .A2(n17205), .ZN(n10611) );
  NOR2_X1 U13366 ( .A1(n17205), .A2(n10588), .ZN(n10589) );
  OR2_X1 U13367 ( .A1(n13583), .A2(n16517), .ZN(n13599) );
  OR2_X1 U13368 ( .A1(n13583), .A2(n20077), .ZN(n12852) );
  NOR2_X1 U13369 ( .A1(n11542), .A2(n11541), .ZN(n11566) );
  INV_X1 U13370 ( .A(n16781), .ZN(n15863) );
  NOR2_X1 U13371 ( .A1(n20273), .A2(n20280), .ZN(n20766) );
  AND2_X1 U13372 ( .A1(n20273), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13373 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10816), .B1(
        n17176), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10682) );
  NAND2_X1 U13374 ( .A1(n11237), .A2(n11236), .ZN(n13602) );
  INV_X1 U13375 ( .A(n14388), .ZN(n11856) );
  AOI21_X1 U13376 ( .B1(n16530), .B2(n20213), .A(n16529), .ZN(n16532) );
  NOR2_X1 U13377 ( .A1(n10606), .A2(n17239), .ZN(n10586) );
  AND3_X1 U13378 ( .A1(n10546), .A2(n10545), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13379 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10705), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13380 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U13381 ( .A1(n13139), .A2(n13138), .ZN(n10456) );
  INV_X1 U13382 ( .A(n17814), .ZN(n18680) );
  INV_X1 U13383 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20559) );
  OR2_X1 U13384 ( .A1(n16493), .A2(n20227), .ZN(n10458) );
  OR2_X1 U13385 ( .A1(n16942), .A2(n16911), .ZN(n10459) );
  AND3_X1 U13386 ( .A1(n12471), .A2(n12480), .A3(n12470), .ZN(n10460) );
  OR2_X1 U13387 ( .A1(n12477), .A2(n20219), .ZN(n10461) );
  NAND2_X2 U13388 ( .A1(n15029), .A2(n14082), .ZN(n15031) );
  INV_X1 U13389 ( .A(n20087), .ZN(n15862) );
  AND2_X1 U13390 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10462) );
  INV_X1 U13391 ( .A(n14960), .ZN(n21030) );
  NAND2_X1 U13392 ( .A1(n21035), .A2(n14569), .ZN(n14960) );
  AND4_X1 U13393 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n10463) );
  OR2_X1 U13394 ( .A1(n19523), .A2(n19756), .ZN(n19479) );
  INV_X1 U13395 ( .A(n9612), .ZN(n18880) );
  NOR2_X1 U13396 ( .A1(n19095), .A2(n19083), .ZN(n17343) );
  INV_X1 U13397 ( .A(n11251), .ZN(n11258) );
  NOR2_X1 U13398 ( .A1(n20555), .A2(n20435), .ZN(n10465) );
  INV_X1 U13399 ( .A(n9610), .ZN(n12720) );
  INV_X1 U13400 ( .A(n11555), .ZN(n11559) );
  AND2_X1 U13401 ( .A1(n16597), .A2(n11063), .ZN(n10466) );
  INV_X1 U13402 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n10937) );
  AND4_X1 U13403 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n13115), .ZN(
        n10467) );
  AND2_X1 U13404 ( .A1(n13003), .A2(n13002), .ZN(n10468) );
  OR2_X1 U13405 ( .A1(n13198), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10469) );
  OR2_X1 U13406 ( .A1(n13794), .A2(n13669), .ZN(n13743) );
  AND2_X1 U13407 ( .A1(n10543), .A2(n10542), .ZN(n10470) );
  INV_X2 U13408 ( .A(n18703), .ZN(n18726) );
  INV_X2 U13409 ( .A(n18471), .ZN(n18458) );
  AND2_X1 U13410 ( .A1(n13599), .A2(n13598), .ZN(n10471) );
  NAND2_X1 U13411 ( .A1(n12729), .A2(n12728), .ZN(n17622) );
  AND2_X1 U13412 ( .A1(n18615), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10472) );
  INV_X1 U13413 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18912) );
  INV_X1 U13414 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11088) );
  INV_X1 U13415 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18899) );
  INV_X1 U13416 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13625) );
  AND2_X1 U13417 ( .A1(n14861), .A2(n14862), .ZN(n10473) );
  AND3_X1 U13418 ( .A1(n10786), .A2(n10785), .A3(n10784), .ZN(n10474) );
  INV_X1 U13419 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20789) );
  INV_X1 U13420 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19882) );
  INV_X1 U13421 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13148) );
  NOR2_X2 U13422 ( .A1(n20627), .A2(n20534), .ZN(n10477) );
  OR2_X1 U13423 ( .A1(n20627), .A2(n20633), .ZN(n20675) );
  INV_X1 U13424 ( .A(n20256), .ZN(n20724) );
  OR2_X1 U13425 ( .A1(n20627), .A2(n20673), .ZN(n20256) );
  INV_X1 U13426 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n17636) );
  INV_X1 U13427 ( .A(n15176), .ZN(n21133) );
  INV_X1 U13428 ( .A(n17205), .ZN(n10609) );
  AND2_X1 U13429 ( .A1(n14791), .A2(n14811), .ZN(n10479) );
  OR2_X1 U13430 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12295) );
  INV_X1 U13431 ( .A(n14712), .ZN(n14727) );
  NAND3_X1 U13432 ( .A1(n11920), .A2(n11919), .A3(n11918), .ZN(n10481) );
  OR2_X1 U13433 ( .A1(n10795), .A2(n20234), .ZN(n10482) );
  INV_X1 U13434 ( .A(n15897), .ZN(n15913) );
  OR2_X1 U13435 ( .A1(n13602), .A2(n20087), .ZN(n10483) );
  OR2_X1 U13436 ( .A1(n12477), .A2(n16773), .ZN(n10485) );
  OR2_X1 U13437 ( .A1(n16823), .A2(n16773), .ZN(n10486) );
  AND2_X1 U13438 ( .A1(n17246), .A2(n10627), .ZN(n10487) );
  AND4_X1 U13439 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n10488) );
  AND4_X1 U13440 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n10489) );
  AND4_X1 U13441 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n10490) );
  AND4_X1 U13442 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n10491) );
  NAND2_X1 U13443 ( .A1(n11662), .A2(n14299), .ZN(n11682) );
  AOI22_X1 U13444 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10818), .B1(
        n10854), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10680) );
  OR2_X1 U13445 ( .A1(n11845), .A2(n11844), .ZN(n12520) );
  OR2_X1 U13446 ( .A1(n12381), .A2(n12380), .ZN(n12383) );
  INV_X1 U13447 ( .A(n10640), .ZN(n10641) );
  AOI22_X1 U13448 ( .A1(n10706), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10545) );
  AND2_X1 U13449 ( .A1(n21307), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12370) );
  INV_X1 U13450 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12210) );
  OR2_X1 U13451 ( .A1(n11888), .A2(n11887), .ZN(n12564) );
  OAI21_X1 U13452 ( .B1(n12996), .B2(n15722), .A(n11695), .ZN(n11671) );
  AND2_X1 U13453 ( .A1(n13369), .A2(n13368), .ZN(n13535) );
  AOI22_X1 U13454 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13455 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10580) );
  INV_X1 U13456 ( .A(n12250), .ZN(n12212) );
  INV_X1 U13457 ( .A(n14713), .ZN(n12128) );
  INV_X1 U13458 ( .A(n11952), .ZN(n11953) );
  OR2_X1 U13459 ( .A1(n11740), .A2(n11739), .ZN(n12525) );
  INV_X1 U13460 ( .A(n12572), .ZN(n12506) );
  OR2_X1 U13461 ( .A1(n11697), .A2(n11696), .ZN(n11707) );
  NAND2_X1 U13462 ( .A1(n12397), .A2(n12562), .ZN(n12402) );
  INV_X1 U13463 ( .A(n16115), .ZN(n11125) );
  INV_X1 U13464 ( .A(n13535), .ZN(n13558) );
  AND2_X1 U13465 ( .A1(n16333), .A2(n16323), .ZN(n13479) );
  AND2_X1 U13466 ( .A1(n13408), .A2(n13432), .ZN(n13409) );
  INV_X1 U13467 ( .A(n17224), .ZN(n11218) );
  NAND2_X1 U13468 ( .A1(n13143), .A2(n13131), .ZN(n13132) );
  AND2_X1 U13469 ( .A1(n14017), .A2(n14016), .ZN(n14018) );
  NAND2_X1 U13470 ( .A1(n12037), .A2(n10479), .ZN(n12038) );
  AND2_X1 U13471 ( .A1(n12313), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12314) );
  NAND2_X1 U13472 ( .A1(n12236), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12240) );
  AND2_X1 U13473 ( .A1(n11953), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11954) );
  INV_X1 U13474 ( .A(n11791), .ZN(n12346) );
  INV_X1 U13475 ( .A(n11720), .ZN(n12540) );
  NOR2_X1 U13476 ( .A1(n13807), .A2(n12506), .ZN(n12507) );
  INV_X1 U13477 ( .A(n16377), .ZN(n13276) );
  INV_X1 U13478 ( .A(n16354), .ZN(n13352) );
  INV_X1 U13479 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U13480 ( .A1(n10957), .A2(n10956), .ZN(n10979) );
  INV_X1 U13481 ( .A(n16047), .ZN(n11514) );
  OR2_X2 U13482 ( .A1(n10965), .A2(n20273), .ZN(n11095) );
  NAND2_X1 U13483 ( .A1(n10601), .A2(n11333), .ZN(n10718) );
  NOR2_X2 U13484 ( .A1(n10952), .A2(n20273), .ZN(n11314) );
  AOI21_X1 U13485 ( .B1(n13247), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13246), .ZN(n13248) );
  OR2_X1 U13486 ( .A1(n13976), .A2(n13164), .ZN(n13165) );
  INV_X1 U13487 ( .A(n14544), .ZN(n14550) );
  AND2_X1 U13488 ( .A1(n12275), .A2(n14688), .ZN(n12276) );
  AND2_X1 U13489 ( .A1(n11775), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12351) );
  OR2_X1 U13490 ( .A1(n12995), .A2(n14872), .ZN(n14218) );
  NAND2_X1 U13491 ( .A1(n12314), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14533) );
  OR2_X1 U13492 ( .A1(n12131), .A2(n12130), .ZN(n12254) );
  OR2_X1 U13493 ( .A1(n12067), .A2(n15177), .ZN(n12084) );
  INV_X1 U13494 ( .A(n14774), .ZN(n12687) );
  AND2_X1 U13495 ( .A1(n15605), .A2(n21285), .ZN(n15607) );
  NAND2_X1 U13496 ( .A1(n11808), .A2(n11807), .ZN(n14392) );
  XNOR2_X1 U13497 ( .A(n11833), .B(n14336), .ZN(n12512) );
  INV_X1 U13498 ( .A(n17527), .ZN(n17525) );
  AND2_X1 U13499 ( .A1(n20273), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11045) );
  AND2_X1 U13500 ( .A1(n13502), .A2(n13501), .ZN(n13544) );
  INV_X1 U13501 ( .A(n14273), .ZN(n11373) );
  NAND2_X1 U13502 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12449) );
  INV_X1 U13503 ( .A(n15849), .ZN(n11536) );
  AND2_X1 U13504 ( .A1(n11535), .A2(n11534), .ZN(n15866) );
  OR3_X1 U13505 ( .A1(n15958), .A2(n11555), .A3(n11279), .ZN(n11086) );
  AND2_X1 U13506 ( .A1(n16613), .A2(n16621), .ZN(n12454) );
  AND2_X1 U13507 ( .A1(n16910), .A2(n16936), .ZN(n16911) );
  AND3_X1 U13508 ( .A1(n11392), .A2(n11391), .A3(n11390), .ZN(n14276) );
  INV_X1 U13509 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17024) );
  NOR2_X1 U13510 ( .A1(n20876), .A2(n20050), .ZN(n20464) );
  INV_X1 U13511 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17248) );
  NOR2_X1 U13512 ( .A1(n10457), .A2(n19438), .ZN(n13963) );
  CLKBUF_X3 U13513 ( .A(n13081), .Z(n18271) );
  NOR2_X1 U13514 ( .A1(n13958), .A2(n17806), .ZN(n14062) );
  NOR2_X1 U13515 ( .A1(n18598), .A2(n13938), .ZN(n13937) );
  AND2_X1 U13516 ( .A1(n18873), .A2(n17311), .ZN(n18806) );
  NAND2_X1 U13517 ( .A1(n17814), .A2(n14057), .ZN(n14058) );
  OR2_X1 U13518 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  NAND2_X1 U13519 ( .A1(n14550), .A2(n14548), .ZN(n21006) );
  NAND2_X1 U13520 ( .A1(n14550), .A2(n14549), .ZN(n20970) );
  NAND2_X1 U13521 ( .A1(n14961), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12863) );
  AND2_X1 U13522 ( .A1(n12678), .A2(n12677), .ZN(n14812) );
  NAND2_X1 U13523 ( .A1(n11931), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11946) );
  OR2_X1 U13524 ( .A1(n15245), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15045) );
  AND2_X1 U13525 ( .A1(n15227), .A2(n15449), .ZN(n15206) );
  INV_X1 U13526 ( .A(n21148), .ZN(n17601) );
  INV_X1 U13527 ( .A(n17591), .ZN(n17592) );
  AND2_X1 U13528 ( .A1(n21172), .A2(n21171), .ZN(n21174) );
  OR2_X1 U13529 ( .A1(n21175), .A2(n15562), .ZN(n15635) );
  NAND2_X1 U13530 ( .A1(n21250), .A2(n14400), .ZN(n15672) );
  OR2_X1 U13531 ( .A1(n15677), .A2(n15682), .ZN(n15678) );
  AND2_X1 U13532 ( .A1(n11805), .A2(n14293), .ZN(n15681) );
  INV_X1 U13533 ( .A(n15559), .ZN(n15527) );
  AOI21_X1 U13534 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21307), .A(n15642), 
        .ZN(n21315) );
  AND2_X1 U13535 ( .A1(n11523), .A2(n11522), .ZN(n15983) );
  INV_X1 U13536 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16093) );
  NOR2_X2 U13537 ( .A1(n15966), .A2(n15967), .ZN(n15948) );
  INV_X1 U13538 ( .A(n13544), .ZN(n16309) );
  AND3_X1 U13539 ( .A1(n11474), .A2(n11473), .A3(n11472), .ZN(n14282) );
  INV_X1 U13540 ( .A(n13669), .ZN(n13670) );
  AOI21_X1 U13541 ( .B1(n16329), .B2(n20213), .A(n11165), .ZN(n11166) );
  NOR2_X1 U13542 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  AND2_X1 U13543 ( .A1(n11517), .A2(n11516), .ZN(n16039) );
  OR2_X1 U13544 ( .A1(n10935), .A2(n10936), .ZN(n17263) );
  NAND2_X1 U13545 ( .A1(n20889), .A2(n20251), .ZN(n20534) );
  OR2_X1 U13546 ( .A1(n20468), .A2(n20633), .ZN(n20409) );
  AND2_X1 U13547 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20462) );
  OR2_X1 U13548 ( .A1(n20674), .A2(n20534), .ZN(n20492) );
  OR2_X1 U13549 ( .A1(n20889), .A2(n20871), .ZN(n20633) );
  AND2_X1 U13550 ( .A1(n20676), .A2(n20873), .ZN(n20680) );
  NAND2_X1 U13551 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20731), .ZN(n20280) );
  NOR2_X1 U13552 ( .A1(n18157), .A2(n17346), .ZN(n13177) );
  NAND2_X1 U13553 ( .A1(n20042), .A2(n18620), .ZN(n13173) );
  OAI211_X2 U13554 ( .C1(P3_STATEBS16_REG_SCAN_IN), .C2(n20028), .A(n13181), 
        .B(n13180), .ZN(n18185) );
  NAND2_X1 U13555 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18294), .ZN(n18278) );
  INV_X1 U13556 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18034) );
  INV_X1 U13557 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18732) );
  NAND2_X1 U13558 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13006) );
  INV_X1 U13559 ( .A(n14059), .ZN(n14521) );
  INV_X1 U13560 ( .A(n19635), .ZN(n19681) );
  OR2_X1 U13561 ( .A1(n17527), .A2(n21369), .ZN(n20927) );
  OR2_X1 U13562 ( .A1(n20958), .A2(n14823), .ZN(n17565) );
  OR2_X1 U13563 ( .A1(n21462), .A2(n14540), .ZN(n14884) );
  INV_X1 U13564 ( .A(n21035), .ZN(n14961) );
  INV_X2 U13565 ( .A(n14443), .ZN(n21091) );
  NAND2_X1 U13566 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  AOI21_X1 U13567 ( .B1(n14687), .B2(n12854), .A(n14663), .ZN(n15100) );
  NAND2_X1 U13568 ( .A1(n11891), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11900) );
  NOR2_X2 U13569 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21285) );
  OAI21_X1 U13570 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12582), .A(
        n12586), .ZN(n15208) );
  NOR2_X1 U13571 ( .A1(n17592), .A2(n17597), .ZN(n21113) );
  INV_X1 U13572 ( .A(n17600), .ZN(n21127) );
  NAND2_X1 U13573 ( .A1(n13851), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15520) );
  INV_X1 U13574 ( .A(n21198), .ZN(n21155) );
  OR2_X1 U13575 ( .A1(n15526), .A2(n14285), .ZN(n21175) );
  INV_X1 U13576 ( .A(n15564), .ZN(n21194) );
  OAI22_X1 U13577 ( .A1(n15610), .A2(n15609), .B1(n11775), .B2(n15608), .ZN(
        n15632) );
  INV_X1 U13578 ( .A(n21210), .ZN(n21242) );
  AND2_X1 U13579 ( .A1(n14285), .A2(n14337), .ZN(n21250) );
  AND2_X1 U13580 ( .A1(n21250), .A2(n15802), .ZN(n21271) );
  AND2_X1 U13581 ( .A1(n21250), .A2(n15597), .ZN(n15716) );
  AND2_X1 U13582 ( .A1(n15719), .A2(n15802), .ZN(n21302) );
  OAI21_X1 U13583 ( .B1(n14360), .B2(n15724), .A(n21315), .ZN(n14384) );
  AND2_X1 U13584 ( .A1(n15719), .A2(n15597), .ZN(n15795) );
  OAI21_X1 U13585 ( .B1(n21317), .B2(n21316), .A(n21315), .ZN(n21364) );
  NOR2_X2 U13586 ( .A1(n15264), .A2(n14440), .ZN(n14328) );
  INV_X1 U13587 ( .A(n21206), .ZN(n15805) );
  INV_X1 U13588 ( .A(n15691), .ZN(n21328) );
  INV_X1 U13589 ( .A(n15703), .ZN(n21346) );
  NOR2_X1 U13590 ( .A1(n15642), .A2(n14496), .ZN(n21361) );
  INV_X1 U13591 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21390) );
  AOI21_X1 U13592 ( .B1(n12850), .B2(n16290), .A(n12849), .ZN(n12851) );
  AND2_X1 U13593 ( .A1(n16262), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16275) );
  NOR2_X1 U13594 ( .A1(n16414), .A2(n16391), .ZN(n16415) );
  AND2_X1 U13595 ( .A1(n14095), .A2(n16220), .ZN(n16217) );
  NOR2_X2 U13596 ( .A1(n20133), .A2(n10360), .ZN(n20114) );
  OR2_X1 U13597 ( .A1(n13639), .A2(n13581), .ZN(n13582) );
  INV_X1 U13598 ( .A(n20909), .ZN(n20175) );
  INV_X1 U13599 ( .A(n20132), .ZN(n17210) );
  AND2_X1 U13600 ( .A1(n17654), .A2(n13633), .ZN(n20209) );
  INV_X1 U13601 ( .A(n20227), .ZN(n20238) );
  XNOR2_X1 U13602 ( .A(n13701), .B(n13702), .ZN(n20871) );
  NOR2_X2 U13603 ( .A1(n20534), .A2(n20433), .ZN(n20310) );
  NOR2_X2 U13604 ( .A1(n20534), .A2(n20468), .ZN(n20342) );
  AND2_X1 U13605 ( .A1(n20889), .A2(n20871), .ZN(n20870) );
  NOR2_X1 U13606 ( .A1(n20433), .A2(n20633), .ZN(n20427) );
  OAI21_X1 U13607 ( .B1(n20501), .B2(n11308), .A(n20467), .ZN(n20488) );
  NOR2_X2 U13608 ( .A1(n20673), .A2(n20468), .ZN(n20520) );
  NOR2_X1 U13609 ( .A1(n20674), .A2(n20346), .ZN(n20592) );
  NOR2_X2 U13610 ( .A1(n20674), .A2(n20633), .ZN(n20669) );
  INV_X1 U13611 ( .A(n20675), .ZN(n20718) );
  OAI22_X1 U13612 ( .A1(n17725), .A2(n20290), .B1(n16488), .B2(n20289), .ZN(
        n20704) );
  AND2_X1 U13613 ( .A1(n10625), .A2(n20287), .ZN(n20778) );
  NAND2_X1 U13614 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17115) );
  INV_X1 U13615 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20806) );
  NOR2_X1 U13616 ( .A1(n14521), .A2(n13147), .ZN(n19874) );
  NOR2_X1 U13617 ( .A1(n20041), .A2(n14060), .ZN(n19880) );
  NOR2_X1 U13618 ( .A1(n18179), .A2(n13170), .ZN(n17881) );
  NOR2_X1 U13619 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18005), .ZN(n17992) );
  INV_X1 U13620 ( .A(n18186), .ZN(n18132) );
  NOR2_X2 U13621 ( .A1(n19898), .A2(n13173), .ZN(n18167) );
  INV_X1 U13622 ( .A(n18280), .ZN(n18240) );
  NOR2_X1 U13623 ( .A1(n18518), .A2(n18278), .ZN(n18280) );
  NAND2_X1 U13624 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18350), .ZN(n18335) );
  INV_X1 U13625 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18442) );
  OAI21_X1 U13626 ( .B1(n14085), .B2(n14084), .A(n20026), .ZN(n14497) );
  NOR2_X1 U13627 ( .A1(n18642), .A2(n18545), .ZN(n18540) );
  INV_X1 U13628 ( .A(n18531), .ZN(n18550) );
  INV_X1 U13629 ( .A(n18610), .ZN(n18613) );
  INV_X1 U13630 ( .A(n19095), .ZN(n18932) );
  OR2_X1 U13631 ( .A1(n13866), .A2(n13865), .ZN(n17386) );
  AND2_X1 U13632 ( .A1(n19027), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18935) );
  INV_X1 U13633 ( .A(n19291), .ZN(n18969) );
  INV_X1 U13634 ( .A(n17491), .ZN(n18754) );
  INV_X1 U13635 ( .A(n19164), .ZN(n19179) );
  INV_X1 U13636 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n19228) );
  NOR2_X2 U13637 ( .A1(n19404), .A2(n18591), .ZN(n19326) );
  INV_X1 U13638 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n19346) );
  INV_X1 U13639 ( .A(n19390), .ZN(n19397) );
  INV_X1 U13640 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19866) );
  NOR2_X1 U13641 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n20040) );
  INV_X1 U13642 ( .A(n19423), .ZN(n19455) );
  INV_X1 U13643 ( .A(n19516), .ZN(n19518) );
  INV_X1 U13644 ( .A(n19588), .ZN(n19575) );
  INV_X1 U13645 ( .A(n19653), .ZN(n19655) );
  INV_X1 U13646 ( .A(n19696), .ZN(n19702) );
  INV_X1 U13647 ( .A(n19830), .ZN(n19742) );
  INV_X1 U13648 ( .A(n19477), .ZN(n19790) );
  AND2_X1 U13649 ( .A1(n19759), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19807) );
  INV_X1 U13650 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19918) );
  INV_X1 U13651 ( .A(n17185), .ZN(n17186) );
  NOR2_X1 U13652 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13608), .ZN(n17787)
         );
  INV_X1 U13653 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21204) );
  OR2_X1 U13654 ( .A1(n15040), .A2(n14560), .ZN(n20974) );
  INV_X1 U13655 ( .A(n21024), .ZN(n14918) );
  INV_X1 U13656 ( .A(n15093), .ZN(n14979) );
  INV_X1 U13657 ( .A(n17556), .ZN(n15014) );
  AND2_X1 U13658 ( .A1(n12420), .A2(n13624), .ZN(n15029) );
  OR2_X1 U13659 ( .A1(n21069), .A2(n14541), .ZN(n14163) );
  OR2_X1 U13660 ( .A1(n13724), .A2(n13723), .ZN(n21069) );
  NOR2_X1 U13661 ( .A1(n14536), .A2(n14437), .ZN(n14444) );
  OR2_X2 U13662 ( .A1(n21094), .A2(n13824), .ZN(n21106) );
  NAND2_X1 U13663 ( .A1(n12989), .A2(n21285), .ZN(n15264) );
  AOI21_X1 U13664 ( .B1(n15536), .B2(n15540), .A(n15535), .ZN(n21158) );
  OR2_X1 U13665 ( .A1(n21175), .A2(n15528), .ZN(n21198) );
  NAND2_X1 U13666 ( .A1(n15598), .A2(n15597), .ZN(n21210) );
  NAND2_X1 U13667 ( .A1(n21250), .A2(n21199), .ZN(n21275) );
  AOI21_X1 U13668 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(n14428) );
  NAND2_X1 U13669 ( .A1(n15719), .A2(n21199), .ZN(n21306) );
  NAND2_X1 U13670 ( .A1(n15719), .A2(n14400), .ZN(n15757) );
  NAND2_X1 U13671 ( .A1(n15803), .A2(n21199), .ZN(n21367) );
  INV_X1 U13672 ( .A(n21335), .ZN(n15821) );
  NOR2_X1 U13673 ( .A1(n14288), .A2(n14287), .ZN(n14333) );
  INV_X1 U13674 ( .A(n21389), .ZN(n21467) );
  NOR2_X1 U13675 ( .A1(n21461), .A2(n21392), .ZN(n21450) );
  INV_X1 U13676 ( .A(n21439), .ZN(n21436) );
  OR3_X1 U13677 ( .A1(n12838), .A2(n17677), .A3(n17272), .ZN(n13668) );
  INV_X1 U13678 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20050) );
  INV_X1 U13679 ( .A(n16301), .ZN(n20087) );
  INV_X1 U13680 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n16404) );
  AND2_X1 U13681 ( .A1(n11232), .A2(n13643), .ZN(n20112) );
  NAND2_X1 U13682 ( .A1(n10588), .A2(n16495), .ZN(n16517) );
  AND2_X1 U13683 ( .A1(n13582), .A2(n13643), .ZN(n16495) );
  AND2_X1 U13684 ( .A1(n20138), .A2(n16517), .ZN(n16525) );
  INV_X1 U13685 ( .A(n16522), .ZN(n20142) );
  NAND2_X1 U13686 ( .A1(n13679), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20909) );
  NAND2_X1 U13687 ( .A1(n13678), .A2(n20911), .ZN(n20178) );
  INV_X1 U13688 ( .A(n13794), .ZN(n13762) );
  INV_X1 U13689 ( .A(n11167), .ZN(n11168) );
  INV_X1 U13690 ( .A(n20196), .ZN(n20211) );
  INV_X1 U13691 ( .A(n20209), .ZN(n20199) );
  INV_X1 U13692 ( .A(n12475), .ZN(n12476) );
  INV_X1 U13693 ( .A(n17661), .ZN(n20241) );
  INV_X1 U13694 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20885) );
  NAND2_X1 U13695 ( .A1(n13646), .A2(n13645), .ZN(n17149) );
  OAI22_X1 U13696 ( .A1(n20255), .A2(n20288), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n20259), .ZN(n20295) );
  INV_X1 U13697 ( .A(n20311), .ZN(n20307) );
  NAND2_X1 U13698 ( .A1(n20315), .A2(n20870), .ZN(n20377) );
  INV_X1 U13699 ( .A(n20427), .ZN(n20425) );
  INV_X1 U13700 ( .A(n20437), .ZN(n20491) );
  OAI22_X1 U13701 ( .A1(n20499), .A2(n20498), .B1(n20497), .B2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n20524) );
  INV_X1 U13702 ( .A(n20604), .ZN(n20595) );
  AOI21_X1 U13703 ( .B1(n17233), .B2(n17232), .A(n17231), .ZN(n20626) );
  INV_X1 U13704 ( .A(n20749), .ZN(n20699) );
  INV_X1 U13705 ( .A(n20773), .ZN(n20715) );
  INV_X1 U13706 ( .A(n20700), .ZN(n20759) );
  INV_X1 U13707 ( .A(n20717), .ZN(n20787) );
  INV_X1 U13708 ( .A(n20867), .ZN(n20788) );
  INV_X1 U13709 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U13710 ( .A1(n19895), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19910) );
  INV_X1 U13711 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19038) );
  INV_X1 U13712 ( .A(n18235), .ZN(n18239) );
  AND2_X1 U13713 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18337), .ZN(n18350) );
  INV_X1 U13714 ( .A(n18451), .ZN(n18473) );
  NAND2_X1 U13715 ( .A1(n18476), .A2(n18576), .ZN(n18531) );
  INV_X1 U13716 ( .A(n17386), .ZN(n18591) );
  INV_X1 U13717 ( .A(n18612), .ZN(n18607) );
  NAND2_X1 U13718 ( .A1(n18672), .A2(n18620), .ZN(n18645) );
  INV_X1 U13719 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18663) );
  INV_X1 U13720 ( .A(n18672), .ZN(n18677) );
  AOI211_X1 U13721 ( .C1(n20028), .C2(n14057), .A(n18680), .B(n18679), .ZN(
        n18703) );
  INV_X1 U13722 ( .A(n18727), .ZN(n18720) );
  OR3_X1 U13723 ( .A1(n14057), .A2(n18680), .A3(n18679), .ZN(n18729) );
  INV_X1 U13724 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19162) );
  INV_X1 U13725 ( .A(n18935), .ZN(n18962) );
  NAND2_X1 U13726 ( .A1(n17816), .A2(n14057), .ZN(n19099) );
  INV_X1 U13727 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19174) );
  INV_X2 U13728 ( .A(n19400), .ZN(n19402) );
  INV_X1 U13729 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19287) );
  INV_X1 U13730 ( .A(n19326), .ZN(n19310) );
  NAND2_X2 U13731 ( .A1(n20040), .A2(n13166), .ZN(n19400) );
  INV_X1 U13732 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19860) );
  INV_X1 U13733 ( .A(n19535), .ZN(n19544) );
  INV_X1 U13734 ( .A(n19621), .ZN(n19634) );
  INV_X1 U13735 ( .A(n19826), .ZN(n19745) );
  INV_X1 U13736 ( .A(n19797), .ZN(n19763) );
  INV_X1 U13737 ( .A(n19788), .ZN(n19781) );
  INV_X1 U13738 ( .A(n19764), .ZN(n19812) );
  INV_X1 U13739 ( .A(n18097), .ZN(n19913) );
  INV_X1 U13740 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20009) );
  INV_X1 U13741 ( .A(n20006), .ZN(n20003) );
  INV_X1 U13742 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19932) );
  INV_X1 U13743 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19958) );
  INV_X1 U13744 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20144) );
  INV_X1 U13745 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20812) );
  NAND2_X1 U13746 ( .A1(n13004), .A2(n10468), .ZN(P1_U2974) );
  INV_X1 U13747 ( .A(n11234), .ZN(P2_U2856) );
  NAND2_X1 U13748 ( .A1(n10486), .A2(n11168), .ZN(P2_U2988) );
  OR2_X1 U13749 ( .A1(n13187), .A2(n13186), .ZN(P3_U2640) );
  AND2_X2 U13750 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10694) );
  AND2_X4 U13751 ( .A1(n10694), .A2(n10926), .ZN(n10706) );
  AOI22_X1 U13752 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10495) );
  NAND2_X2 U13753 ( .A1(n10700), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10503) );
  INV_X4 U13754 ( .A(n10503), .ZN(n10576) );
  NOR2_X2 U13755 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10493) );
  AND2_X4 U13756 ( .A1(n10493), .A2(n17138), .ZN(n13554) );
  AOI22_X1 U13757 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10494) );
  AND3_X1 U13758 ( .A1(n10495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10494), .ZN(n10499) );
  AND2_X4 U13759 ( .A1(n10708), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10698) );
  AND2_X4 U13760 ( .A1(n10694), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13366) );
  AOI22_X1 U13761 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13762 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10497) );
  INV_X1 U13763 ( .A(n10500), .ZN(n10502) );
  NOR2_X1 U13764 ( .A1(n10502), .A2(n10501), .ZN(n10507) );
  AOI22_X1 U13765 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10506) );
  INV_X4 U13766 ( .A(n10503), .ZN(n13568) );
  AOI22_X1 U13767 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13768 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13769 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13770 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13771 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U13772 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13773 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13774 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13775 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13776 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13777 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13778 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10516) );
  NAND4_X1 U13779 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10520) );
  NAND2_X1 U13780 ( .A1(n10520), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10527) );
  AOI22_X1 U13781 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13782 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13783 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13784 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10521) );
  NAND4_X1 U13785 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  AOI22_X1 U13786 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13787 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13788 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13789 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10528) );
  NAND4_X1 U13790 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  AOI22_X1 U13791 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13792 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13793 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13794 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10533) );
  NAND4_X1 U13795 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10537) );
  AOI22_X1 U13796 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13797 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13798 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13799 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13800 ( .A1(n10544), .A2(n10470), .ZN(n10551) );
  AOI22_X1 U13801 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13802 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10705), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13803 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10547) );
  NAND3_X1 U13804 ( .A1(n10549), .A2(n10548), .A3(n10547), .ZN(n10550) );
  INV_X1 U13805 ( .A(n17224), .ZN(n10564) );
  AOI22_X1 U13806 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13807 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13808 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13809 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10552) );
  NAND4_X1 U13810 ( .A1(n10555), .A2(n10554), .A3(n10553), .A4(n10552), .ZN(
        n10556) );
  AOI22_X1 U13811 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13812 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13813 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13814 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10561) );
  INV_X2 U13815 ( .A(n10602), .ZN(n10613) );
  AND3_X2 U13816 ( .A1(n9874), .A2(n10565), .A3(n10613), .ZN(n10619) );
  INV_X1 U13817 ( .A(n10619), .ZN(n11251) );
  NAND3_X1 U13818 ( .A1(n10606), .A2(n10613), .A3(n10565), .ZN(n10935) );
  AOI22_X1 U13819 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13820 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13821 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13822 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13823 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13824 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U13825 ( .A1(n10935), .A2(n10574), .ZN(n10575) );
  AOI22_X1 U13826 ( .A1(n10576), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13827 ( .A1(n10706), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13828 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10699), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13829 ( .A1(n13568), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13830 ( .A1(n10705), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10706), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13831 ( .A1(n10698), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13366), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10581) );
  MUX2_X1 U13832 ( .A(n10624), .B(n10625), .S(n17205), .Z(n10587) );
  NAND2_X1 U13833 ( .A1(n11307), .A2(n11218), .ZN(n10585) );
  NAND3_X1 U13834 ( .A1(n10587), .A2(n10586), .A3(n10585), .ZN(n10591) );
  AND2_X1 U13835 ( .A1(n17224), .A2(n10595), .ZN(n10590) );
  INV_X1 U13836 ( .A(n10625), .ZN(n10588) );
  NAND2_X1 U13837 ( .A1(n11307), .A2(n10601), .ZN(n11222) );
  INV_X1 U13838 ( .A(n11222), .ZN(n10594) );
  INV_X1 U13839 ( .A(n10625), .ZN(n10592) );
  INV_X1 U13840 ( .A(n10637), .ZN(n10600) );
  INV_X1 U13841 ( .A(n10595), .ZN(n10596) );
  NAND2_X1 U13842 ( .A1(n10600), .A2(n10605), .ZN(n10618) );
  NAND2_X1 U13843 ( .A1(n11194), .A2(n10604), .ZN(n11220) );
  INV_X1 U13844 ( .A(n10606), .ZN(n10608) );
  NAND2_X1 U13845 ( .A1(n10608), .A2(n10607), .ZN(n11216) );
  NAND2_X1 U13846 ( .A1(n11216), .A2(n10609), .ZN(n10612) );
  INV_X1 U13847 ( .A(n11307), .ZN(n10610) );
  AND2_X1 U13848 ( .A1(n10622), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13850 ( .A1(n10621), .A2(n11244), .ZN(n11242) );
  NAND3_X1 U13851 ( .A1(n11260), .A2(n10647), .A3(n11259), .ZN(n10626) );
  NAND2_X1 U13852 ( .A1(n10626), .A2(n10462), .ZN(n10635) );
  INV_X1 U13853 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20063) );
  INV_X1 U13854 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13855 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10627) );
  INV_X1 U13856 ( .A(n10629), .ZN(n10630) );
  OAI21_X1 U13857 ( .B1(n10659), .B2(n20063), .A(n10630), .ZN(n10631) );
  INV_X1 U13858 ( .A(n10631), .ZN(n10634) );
  NAND2_X1 U13859 ( .A1(n10636), .A2(n10632), .ZN(n10633) );
  INV_X1 U13860 ( .A(n10644), .ZN(n10666) );
  AOI22_X1 U13861 ( .A1(n11098), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10645) );
  NAND2_X1 U13862 ( .A1(n10646), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U13863 ( .A1(n10658), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10649) );
  AOI21_X1 U13864 ( .B1(n20912), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13865 ( .A1(n11098), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10653) );
  NAND2_X1 U13866 ( .A1(n10655), .A2(n10654), .ZN(n10656) );
  OAI22_X1 U13867 ( .A1(n11173), .A2(n16255), .B1(n17290), .B2(n17655), .ZN(
        n10660) );
  AOI21_X1 U13868 ( .B1(n11175), .B2(P2_REIP_REG_3__SCAN_IN), .A(n10660), .ZN(
        n10661) );
  XNOR2_X2 U13869 ( .A(n10667), .B(n10666), .ZN(n10685) );
  NAND2_X1 U13870 ( .A1(n13719), .A2(n10668), .ZN(n10670) );
  INV_X1 U13871 ( .A(n10668), .ZN(n10669) );
  NOR2_X1 U13872 ( .A1(n10685), .A2(n13666), .ZN(n10672) );
  NAND2_X1 U13873 ( .A1(n13719), .A2(n10672), .ZN(n10678) );
  INV_X1 U13874 ( .A(n10670), .ZN(n10671) );
  AOI22_X1 U13875 ( .A1(n10817), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n20629), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10681) );
  INV_X1 U13876 ( .A(n10672), .ZN(n10673) );
  INV_X1 U13877 ( .A(n10677), .ZN(n10674) );
  INV_X1 U13878 ( .A(n10675), .ZN(n10676) );
  INV_X1 U13879 ( .A(n10678), .ZN(n10679) );
  INV_X1 U13880 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13456) );
  INV_X1 U13881 ( .A(n13223), .ZN(n17649) );
  INV_X1 U13882 ( .A(n13244), .ZN(n20243) );
  NAND2_X1 U13883 ( .A1(n17649), .A2(n10687), .ZN(n20378) );
  NAND2_X1 U13884 ( .A1(n10686), .A2(n14039), .ZN(n20503) );
  INV_X1 U13885 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13303) );
  NAND2_X1 U13886 ( .A1(n10687), .A2(n14039), .ZN(n17230) );
  INV_X1 U13887 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U13888 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20436), .B1(
        n20560), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10692) );
  NAND2_X2 U13889 ( .A1(n9624), .A2(n14056), .ZN(n13322) );
  INV_X1 U13890 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10693) );
  OAI22_X1 U13891 ( .A1(n13322), .A2(n10693), .B1(n14041), .B2(n13303), .ZN(
        n10697) );
  INV_X1 U13892 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13893 ( .A1(n13231), .A2(n13324), .B1(n13320), .B2(n10695), .ZN(
        n10696) );
  NOR2_X1 U13894 ( .A1(n10697), .A2(n10696), .ZN(n10717) );
  AND2_X2 U13895 ( .A1(n9617), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10736) );
  NAND2_X1 U13896 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U13897 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10703) );
  NAND2_X1 U13898 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10702) );
  AND2_X2 U13899 ( .A1(n13367), .A2(n14044), .ZN(n13386) );
  AOI22_X1 U13900 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10701) );
  INV_X1 U13901 ( .A(n10706), .ZN(n10707) );
  AOI22_X1 U13902 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10715) );
  AND2_X2 U13903 ( .A1(n10709), .A2(n13367), .ZN(n13400) );
  AND2_X1 U13904 ( .A1(n10926), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17137) );
  AND2_X2 U13905 ( .A1(n17137), .A2(n13367), .ZN(n13399) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U13907 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U13908 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13909 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10710) );
  NAND4_X1 U13910 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n11333) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17198) );
  INV_X1 U13912 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10719) );
  INV_X1 U13913 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10721) );
  INV_X1 U13914 ( .A(n20629), .ZN(n10720) );
  INV_X1 U13915 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13420) );
  INV_X1 U13916 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10724) );
  INV_X1 U13917 ( .A(n20436), .ZN(n10723) );
  INV_X1 U13918 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10722) );
  OAI22_X1 U13919 ( .A1(n10724), .A2(n20319), .B1(n10723), .B2(n10722), .ZN(
        n10726) );
  INV_X1 U13920 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11374) );
  INV_X1 U13921 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10725) );
  INV_X1 U13922 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10727) );
  INV_X1 U13923 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13418) );
  OAI22_X1 U13924 ( .A1(n10727), .A2(n20503), .B1(n17230), .B2(n13418), .ZN(
        n10730) );
  INV_X1 U13925 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U13926 ( .A1(n10817), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10728) );
  OAI211_X1 U13927 ( .C1(n20378), .C2(n13410), .A(n10728), .B(n11297), .ZN(
        n10729) );
  NOR2_X1 U13928 ( .A1(n10730), .A2(n10729), .ZN(n10731) );
  NAND2_X1 U13929 ( .A1(n13389), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13930 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U13931 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10733) );
  NAND2_X1 U13932 ( .A1(n13390), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10732) );
  NAND4_X1 U13933 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n10742) );
  NAND2_X1 U13934 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13935 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10739) );
  AOI22_X1 U13936 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10738) );
  NAND2_X1 U13937 ( .A1(n10803), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10737) );
  NAND4_X1 U13938 ( .A1(n10740), .A2(n10739), .A3(n10738), .A4(n10737), .ZN(
        n10741) );
  NOR2_X1 U13939 ( .A1(n10742), .A2(n10741), .ZN(n10753) );
  AOI22_X1 U13940 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13941 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10746) );
  NAND2_X1 U13942 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U13943 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10744) );
  NAND4_X1 U13944 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10751) );
  INV_X1 U13945 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10749) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10748) );
  OAI22_X1 U13947 ( .A1(n13322), .A2(n10749), .B1(n13320), .B2(n10748), .ZN(
        n10750) );
  NOR2_X1 U13948 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  NOR2_X1 U13949 ( .A1(n11303), .A2(n11309), .ZN(n10790) );
  NAND2_X1 U13950 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10757) );
  NAND2_X1 U13951 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U13952 ( .A1(n13390), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13953 ( .A1(n13391), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10754) );
  NAND4_X1 U13954 ( .A1(n10757), .A2(n10756), .A3(n10755), .A4(n10754), .ZN(
        n10764) );
  NAND2_X1 U13955 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10762) );
  NAND2_X1 U13956 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10761) );
  AOI22_X1 U13957 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13400), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13958 ( .A1(n13389), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10759) );
  NAND4_X1 U13959 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  NOR2_X1 U13960 ( .A1(n10764), .A2(n10763), .ZN(n10771) );
  AOI22_X1 U13961 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13962 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10765), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13399), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13964 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10766) );
  INV_X1 U13965 ( .A(n10952), .ZN(n10772) );
  NAND2_X1 U13966 ( .A1(n10790), .A2(n10772), .ZN(n10794) );
  AOI22_X1 U13967 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10803), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U13968 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10777) );
  NAND2_X1 U13969 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10776) );
  NAND2_X1 U13970 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10775) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13400), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10774) );
  NAND4_X1 U13972 ( .A1(n10777), .A2(n10776), .A3(n10775), .A4(n10774), .ZN(
        n10783) );
  INV_X1 U13973 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10778) );
  INV_X1 U13974 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11396) );
  OAI22_X1 U13975 ( .A1(n13322), .A2(n10778), .B1(n13320), .B2(n11396), .ZN(
        n10781) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10779) );
  OAI22_X1 U13977 ( .A1(n13233), .A2(n13324), .B1(n14041), .B2(n10779), .ZN(
        n10780) );
  OR2_X1 U13978 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  NOR2_X1 U13979 ( .A1(n10783), .A2(n10782), .ZN(n10787) );
  AOI22_X1 U13980 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U13981 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10785) );
  AOI22_X1 U13982 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13399), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13983 ( .A1(n10794), .A2(n11320), .ZN(n10789) );
  INV_X1 U13984 ( .A(n10790), .ZN(n13631) );
  NAND2_X1 U13985 ( .A1(n13631), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13630) );
  XNOR2_X1 U13986 ( .A(n11303), .B(n10952), .ZN(n10791) );
  NOR2_X1 U13987 ( .A1(n13630), .A2(n10791), .ZN(n10793) );
  INV_X1 U13988 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20202) );
  AOI21_X1 U13989 ( .B1(n13630), .B2(n10791), .A(n10793), .ZN(n10792) );
  INV_X1 U13990 ( .A(n10792), .ZN(n20203) );
  NOR2_X1 U13991 ( .A1(n20202), .A2(n20203), .ZN(n20201) );
  NOR2_X1 U13992 ( .A1(n10793), .A2(n20201), .ZN(n10795) );
  XNOR2_X1 U13993 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10795), .ZN(
        n20191) );
  XNOR2_X1 U13994 ( .A(n10794), .B(n11320), .ZN(n20190) );
  NAND2_X1 U13995 ( .A1(n20191), .A2(n20190), .ZN(n20189) );
  INV_X1 U13996 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20234) );
  NAND2_X1 U13997 ( .A1(n20189), .A2(n10482), .ZN(n10796) );
  INV_X1 U13998 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17099) );
  XNOR2_X1 U13999 ( .A(n10796), .B(n17099), .ZN(n17104) );
  NAND2_X1 U14000 ( .A1(n10796), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10797) );
  AOI22_X1 U14001 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13399), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U14002 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10800) );
  NAND2_X1 U14003 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10799) );
  NAND2_X1 U14004 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10798) );
  NAND4_X1 U14005 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10806) );
  INV_X1 U14006 ( .A(n10802), .ZN(n11437) );
  INV_X1 U14007 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13323) );
  INV_X1 U14008 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10804) );
  NOR2_X1 U14009 ( .A1(n10806), .A2(n10805), .ZN(n10814) );
  NAND2_X1 U14010 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10810) );
  NAND2_X1 U14011 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10809) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13400), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U14013 ( .A1(n13390), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10807) );
  AOI22_X1 U14014 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13392), .B1(
        n11395), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13391), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10811) );
  INV_X1 U14016 ( .A(n10924), .ZN(n11338) );
  INV_X1 U14017 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U14018 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10816), .B1(
        n17176), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U14019 ( .A1(n10817), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n20629), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U14020 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10818), .B1(
        n10854), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U14021 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20436), .B1(
        n20560), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U14022 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20316), .B1(
        n20684), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10827) );
  INV_X1 U14023 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13507) );
  INV_X1 U14024 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10841) );
  OAI22_X1 U14025 ( .A1(n13507), .A2(n20378), .B1(n20503), .B2(n10841), .ZN(
        n10825) );
  INV_X1 U14026 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11456) );
  INV_X1 U14027 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13515) );
  OAI22_X1 U14028 ( .A1(n11456), .A2(n20257), .B1(n17230), .B2(n13515), .ZN(
        n10824) );
  NOR2_X1 U14029 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AOI22_X1 U14030 ( .A1(n13399), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U14031 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10831) );
  NAND2_X1 U14032 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10830) );
  NAND2_X1 U14033 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10829) );
  NAND4_X1 U14034 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10835) );
  INV_X1 U14035 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10833) );
  OAI22_X1 U14036 ( .A1(n13322), .A2(n10833), .B1(n13324), .B2(n11456), .ZN(
        n10834) );
  NOR2_X1 U14037 ( .A1(n10835), .A2(n10834), .ZN(n10845) );
  NAND2_X1 U14038 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10839) );
  NAND2_X1 U14039 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10838) );
  AOI22_X1 U14040 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U14041 ( .A1(n13398), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10836) );
  AOI22_X1 U14042 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11395), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10844) );
  INV_X1 U14043 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10840) );
  OAI22_X1 U14044 ( .A1(n14041), .A2(n10841), .B1(n13320), .B2(n10840), .ZN(
        n10842) );
  INV_X1 U14045 ( .A(n10842), .ZN(n10843) );
  NAND4_X1 U14046 ( .A1(n10845), .A2(n9684), .A3(n10844), .A4(n10843), .ZN(
        n11343) );
  INV_X1 U14047 ( .A(n11343), .ZN(n10846) );
  NAND2_X1 U14048 ( .A1(n10846), .A2(n16324), .ZN(n10847) );
  INV_X1 U14049 ( .A(n10849), .ZN(n10850) );
  INV_X1 U14050 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17072) );
  NAND2_X1 U14051 ( .A1(n10853), .A2(n17072), .ZN(n17062) );
  OR2_X2 U14052 ( .A1(n10853), .A2(n17072), .ZN(n17064) );
  AOI22_X1 U14053 ( .A1(n17176), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10818), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U14054 ( .A1(n10817), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n20629), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U14055 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10854), .B1(
        n20726), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U14056 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20436), .B1(
        n20684), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U14057 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20316), .B1(
        n20560), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10862) );
  INV_X1 U14058 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16413) );
  INV_X1 U14059 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10866) );
  OAI22_X1 U14060 ( .A1(n16413), .A2(n20257), .B1(n20503), .B2(n10866), .ZN(
        n10860) );
  INV_X1 U14061 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13525) );
  INV_X1 U14062 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13533) );
  OAI22_X1 U14063 ( .A1(n13525), .A2(n20378), .B1(n17230), .B2(n13533), .ZN(
        n10859) );
  NOR2_X1 U14064 ( .A1(n10860), .A2(n10859), .ZN(n10861) );
  INV_X1 U14065 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10865) );
  INV_X1 U14066 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10864) );
  OAI22_X1 U14067 ( .A1(n13322), .A2(n10865), .B1(n13320), .B2(n10864), .ZN(
        n10868) );
  OAI22_X1 U14068 ( .A1(n16413), .A2(n13324), .B1(n14041), .B2(n10866), .ZN(
        n10867) );
  NOR2_X1 U14069 ( .A1(n10868), .A2(n10867), .ZN(n10872) );
  AOI22_X1 U14070 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n11395), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U14071 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U14072 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10869) );
  NAND4_X1 U14073 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10878) );
  AOI22_X1 U14074 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U14075 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U14076 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U14077 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10873) );
  NAND4_X1 U14078 ( .A1(n10876), .A2(n10875), .A3(n10874), .A4(n10873), .ZN(
        n10877) );
  NAND2_X1 U14079 ( .A1(n10962), .A2(n16324), .ZN(n10879) );
  INV_X1 U14080 ( .A(n17063), .ZN(n10880) );
  NAND2_X1 U14081 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10887) );
  NAND2_X1 U14082 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10886) );
  NAND2_X1 U14083 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10885) );
  AOI22_X1 U14084 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10884) );
  NAND4_X1 U14085 ( .A1(n10887), .A2(n10886), .A3(n10885), .A4(n10884), .ZN(
        n10894) );
  INV_X1 U14086 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10889) );
  INV_X1 U14087 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10888) );
  OAI22_X1 U14088 ( .A1(n13322), .A2(n10889), .B1(n13320), .B2(n10888), .ZN(
        n10892) );
  INV_X1 U14089 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11492) );
  INV_X1 U14090 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10890) );
  OAI22_X1 U14091 ( .A1(n11492), .A2(n13324), .B1(n14041), .B2(n10890), .ZN(
        n10891) );
  OR2_X1 U14092 ( .A1(n10892), .A2(n10891), .ZN(n10893) );
  NOR2_X1 U14093 ( .A1(n10894), .A2(n10893), .ZN(n10904) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U14095 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10897) );
  NAND2_X1 U14096 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U14097 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10895) );
  NAND4_X1 U14098 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10902) );
  NAND2_X1 U14099 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10900) );
  NAND2_X1 U14100 ( .A1(n13398), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10899) );
  NAND2_X1 U14101 ( .A1(n10900), .A2(n10899), .ZN(n10901) );
  NOR2_X1 U14102 ( .A1(n10902), .A2(n10901), .ZN(n10903) );
  AND2_X2 U14103 ( .A1(n10904), .A2(n10903), .ZN(n11555) );
  OAI21_X1 U14104 ( .B1(n10905), .B2(n11555), .A(n17024), .ZN(n10906) );
  NAND2_X1 U14105 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U14106 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10909) );
  NOR2_X1 U14107 ( .A1(n12450), .A2(n10909), .ZN(n12468) );
  AND3_X1 U14108 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10910) );
  NAND2_X1 U14109 ( .A1(n12468), .A2(n10910), .ZN(n16584) );
  NAND3_X1 U14110 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10911) );
  NOR2_X1 U14111 ( .A1(n16584), .A2(n10911), .ZN(n10912) );
  INV_X1 U14112 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16830) );
  NAND2_X1 U14113 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U14114 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10913) );
  NOR2_X1 U14115 ( .A1(n16815), .A2(n10913), .ZN(n10914) );
  XNOR2_X1 U14116 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U14117 ( .A1(n10944), .A2(n10925), .ZN(n10916) );
  NAND2_X1 U14118 ( .A1(n17256), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10915) );
  NAND2_X1 U14119 ( .A1(n10916), .A2(n10915), .ZN(n10930) );
  NAND2_X1 U14120 ( .A1(n10930), .A2(n10928), .ZN(n10918) );
  NAND2_X1 U14121 ( .A1(n20894), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10917) );
  MUX2_X1 U14122 ( .A(n11333), .B(n11204), .S(n11192), .Z(n10958) );
  INV_X1 U14123 ( .A(n10919), .ZN(n10920) );
  NAND2_X1 U14124 ( .A1(n10921), .A2(n10920), .ZN(n10923) );
  NAND2_X1 U14125 ( .A1(n20885), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10922) );
  NAND2_X1 U14126 ( .A1(n10923), .A2(n10922), .ZN(n10939) );
  NAND2_X1 U14127 ( .A1(n10937), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10940) );
  MUX2_X1 U14128 ( .A(n10924), .B(n11208), .S(n11192), .Z(n10959) );
  NAND2_X1 U14129 ( .A1(n10958), .A2(n10959), .ZN(n11190) );
  INV_X1 U14130 ( .A(n11190), .ZN(n10934) );
  INV_X1 U14131 ( .A(n10925), .ZN(n10943) );
  NAND2_X1 U14132 ( .A1(n10926), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10927) );
  NAND2_X1 U14133 ( .A1(n10943), .A2(n10927), .ZN(n11197) );
  MUX2_X1 U14134 ( .A(n11303), .B(n11197), .S(n11192), .Z(n10980) );
  INV_X1 U14135 ( .A(n10944), .ZN(n11198) );
  INV_X1 U14136 ( .A(n10928), .ZN(n10929) );
  XNOR2_X1 U14137 ( .A(n10930), .B(n10929), .ZN(n11191) );
  INV_X1 U14138 ( .A(n11191), .ZN(n11201) );
  OAI21_X1 U14139 ( .B1(n10980), .B2(n11198), .A(n10955), .ZN(n10933) );
  NAND2_X1 U14140 ( .A1(n10934), .A2(n10933), .ZN(n17265) );
  AND2_X1 U14141 ( .A1(n16324), .A2(n17183), .ZN(n12774) );
  INV_X1 U14142 ( .A(n12774), .ZN(n10936) );
  NOR2_X1 U14143 ( .A1(n10937), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10938) );
  NOR2_X1 U14144 ( .A1(n17263), .A2(n11211), .ZN(n10942) );
  NAND2_X1 U14145 ( .A1(n17265), .A2(n10942), .ZN(n17276) );
  INV_X1 U14146 ( .A(n11211), .ZN(n17264) );
  XNOR2_X1 U14147 ( .A(n10944), .B(n10943), .ZN(n11195) );
  NAND4_X1 U14148 ( .A1(n11208), .A2(n11191), .A3(n11204), .A4(n11195), .ZN(
        n10945) );
  INV_X1 U14149 ( .A(n11197), .ZN(n11196) );
  NAND4_X1 U14150 ( .A1(n11208), .A2(n11191), .A3(n11204), .A4(n11196), .ZN(
        n10946) );
  AND2_X1 U14151 ( .A1(n13611), .A2(n10946), .ZN(n10948) );
  INV_X1 U14152 ( .A(n10947), .ZN(n14047) );
  NAND2_X1 U14153 ( .A1(n14047), .A2(n10937), .ZN(n13647) );
  INV_X1 U14154 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13618) );
  OAI21_X1 U14155 ( .B1(n11395), .B2(n13647), .A(n13618), .ZN(n17111) );
  MUX2_X1 U14156 ( .A(n10948), .B(n17111), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20898) );
  NOR2_X1 U14157 ( .A1(n10935), .A2(n11192), .ZN(n20902) );
  NAND2_X1 U14158 ( .A1(n20898), .A2(n20902), .ZN(n10949) );
  NAND2_X1 U14159 ( .A1(n17276), .A2(n10949), .ZN(n10950) );
  NOR2_X1 U14160 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10953) );
  AND2_X1 U14161 ( .A1(n20273), .A2(n10953), .ZN(n10954) );
  NOR2_X2 U14162 ( .A1(n10981), .A2(n10979), .ZN(n10974) );
  MUX2_X1 U14163 ( .A(n10958), .B(n16255), .S(n20273), .Z(n10975) );
  NAND2_X1 U14164 ( .A1(n10974), .A2(n10975), .ZN(n10973) );
  INV_X1 U14165 ( .A(n10959), .ZN(n10960) );
  INV_X1 U14166 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10961) );
  MUX2_X1 U14167 ( .A(n11343), .B(n10961), .S(n20273), .Z(n11000) );
  INV_X1 U14168 ( .A(n10964), .ZN(n11004) );
  MUX2_X1 U14169 ( .A(n10962), .B(P2_EBX_REG_6__SCAN_IN), .S(n20273), .Z(
        n10968) );
  XNOR2_X1 U14170 ( .A(n11004), .B(n10968), .ZN(n20074) );
  MUX2_X1 U14171 ( .A(n11555), .B(P2_EBX_REG_7__SCAN_IN), .S(n20273), .Z(
        n10970) );
  NOR2_X1 U14172 ( .A1(n10968), .A2(n10970), .ZN(n10963) );
  NAND2_X1 U14173 ( .A1(n10965), .A2(n10966), .ZN(n10967) );
  NAND2_X1 U14174 ( .A1(n11015), .A2(n10967), .ZN(n16179) );
  NOR2_X1 U14175 ( .A1(n16179), .A2(n11555), .ZN(n11009) );
  NAND2_X1 U14176 ( .A1(n11009), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16740) );
  INV_X1 U14177 ( .A(n10968), .ZN(n10969) );
  NAND2_X1 U14178 ( .A1(n10964), .A2(n10969), .ZN(n10972) );
  INV_X1 U14179 ( .A(n10970), .ZN(n10971) );
  XNOR2_X1 U14180 ( .A(n10972), .B(n10971), .ZN(n16193) );
  NAND2_X1 U14181 ( .A1(n16193), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16757) );
  AND2_X1 U14182 ( .A1(n16740), .A2(n16757), .ZN(n16699) );
  INV_X1 U14183 ( .A(n10974), .ZN(n10977) );
  INV_X1 U14184 ( .A(n10975), .ZN(n10976) );
  NAND2_X1 U14185 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U14186 ( .A1(n10973), .A2(n10978), .ZN(n16248) );
  XNOR2_X1 U14187 ( .A(n10979), .B(n10981), .ZN(n10987) );
  NAND2_X1 U14188 ( .A1(n10987), .A2(n20234), .ZN(n10986) );
  MUX2_X1 U14189 ( .A(n10980), .B(n10628), .S(n20273), .Z(n13627) );
  INV_X1 U14190 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17125) );
  NOR2_X1 U14191 ( .A1(n13627), .A2(n17125), .ZN(n13628) );
  INV_X1 U14192 ( .A(n10981), .ZN(n10983) );
  AND3_X1 U14193 ( .A1(n20273), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10982) );
  NOR2_X1 U14194 ( .A1(n10983), .A2(n10982), .ZN(n16276) );
  NAND2_X1 U14195 ( .A1(n13628), .A2(n16276), .ZN(n10985) );
  XOR2_X1 U14196 ( .A(n16276), .B(n13628), .Z(n20206) );
  NAND2_X1 U14197 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20206), .ZN(
        n10984) );
  NAND2_X1 U14198 ( .A1(n10985), .A2(n10984), .ZN(n20186) );
  NAND2_X1 U14199 ( .A1(n10986), .A2(n20186), .ZN(n10989) );
  INV_X1 U14200 ( .A(n10987), .ZN(n20187) );
  NAND2_X1 U14201 ( .A1(n20187), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14202 ( .A1(n10989), .A2(n10988), .ZN(n17097) );
  INV_X1 U14203 ( .A(n10990), .ZN(n11002) );
  NAND2_X1 U14204 ( .A1(n11002), .A2(n10991), .ZN(n17082) );
  NAND2_X1 U14205 ( .A1(n17082), .A2(n17071), .ZN(n10994) );
  OAI21_X1 U14206 ( .B1(n17097), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10994), .ZN(n10992) );
  INV_X1 U14207 ( .A(n10992), .ZN(n10993) );
  NAND3_X1 U14208 ( .A1(n10994), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17097), .ZN(n10997) );
  INV_X1 U14209 ( .A(n17082), .ZN(n10995) );
  NAND2_X1 U14210 ( .A1(n10995), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10996) );
  AND2_X1 U14211 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NAND2_X1 U14212 ( .A1(n10999), .A2(n10998), .ZN(n17069) );
  INV_X1 U14213 ( .A(n11000), .ZN(n11001) );
  NAND2_X1 U14214 ( .A1(n11002), .A2(n11001), .ZN(n11003) );
  NAND2_X1 U14215 ( .A1(n11004), .A2(n11003), .ZN(n17067) );
  NOR2_X1 U14216 ( .A1(n17067), .A2(n17072), .ZN(n11005) );
  NAND2_X1 U14217 ( .A1(n17067), .A2(n17072), .ZN(n11006) );
  INV_X1 U14218 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n20107) );
  NAND2_X1 U14219 ( .A1(n11028), .A2(n11095), .ZN(n11027) );
  AND3_X1 U14220 ( .A1(n9734), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n20273), .ZN(
        n11008) );
  OR2_X1 U14221 ( .A1(n11027), .A2(n11008), .ZN(n16139) );
  INV_X1 U14222 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11274) );
  OAI21_X1 U14223 ( .B1(n16139), .B2(n11555), .A(n11274), .ZN(n16703) );
  INV_X1 U14224 ( .A(n11009), .ZN(n11010) );
  NAND2_X1 U14225 ( .A1(n11010), .A2(n17024), .ZN(n16739) );
  INV_X1 U14226 ( .A(n16193), .ZN(n11011) );
  INV_X1 U14227 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17040) );
  NAND2_X1 U14228 ( .A1(n11011), .A2(n17040), .ZN(n16756) );
  AND2_X1 U14229 ( .A1(n16739), .A2(n16756), .ZN(n16697) );
  NAND2_X1 U14230 ( .A1(n20273), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11012) );
  MUX2_X1 U14231 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11012), .S(n9654), .Z(
        n11013) );
  NAND2_X1 U14232 ( .A1(n11013), .A2(n11095), .ZN(n16148) );
  OR2_X1 U14233 ( .A1(n16148), .A2(n11555), .ZN(n11014) );
  INV_X1 U14234 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16720) );
  NAND2_X1 U14235 ( .A1(n11014), .A2(n16720), .ZN(n16715) );
  NAND2_X1 U14236 ( .A1(n20273), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11016) );
  MUX2_X1 U14237 ( .A(n20273), .B(n11016), .S(n11015), .Z(n11017) );
  NAND2_X1 U14238 ( .A1(n16173), .A2(n11559), .ZN(n11018) );
  INV_X1 U14239 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U14240 ( .A1(n11018), .A2(n11023), .ZN(n16730) );
  AND4_X1 U14241 ( .A1(n16703), .A2(n16697), .A3(n16715), .A4(n16730), .ZN(
        n11019) );
  INV_X1 U14242 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16692) );
  INV_X1 U14243 ( .A(n16139), .ZN(n11021) );
  NOR2_X1 U14244 ( .A1(n11555), .A2(n11274), .ZN(n11020) );
  NAND2_X1 U14245 ( .A1(n11021), .A2(n11020), .ZN(n16702) );
  OR2_X1 U14246 ( .A1(n11555), .A2(n16720), .ZN(n11022) );
  OR2_X1 U14247 ( .A1(n16148), .A2(n11022), .ZN(n16714) );
  NOR2_X1 U14248 ( .A1(n11555), .A2(n11023), .ZN(n11024) );
  NAND2_X1 U14249 ( .A1(n16173), .A2(n11024), .ZN(n16729) );
  AND2_X1 U14250 ( .A1(n16714), .A2(n16729), .ZN(n16700) );
  AND2_X1 U14251 ( .A1(n16702), .A2(n16700), .ZN(n11025) );
  NAND2_X1 U14252 ( .A1(n20273), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U14253 ( .A1(n11027), .A2(n11026), .ZN(n11051) );
  NAND3_X1 U14254 ( .A1(n11028), .A2(n20273), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n11029) );
  NAND2_X1 U14255 ( .A1(n11051), .A2(n11029), .ZN(n16122) );
  INV_X1 U14256 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16978) );
  OR3_X1 U14257 ( .A1(n16122), .A2(n11555), .A3(n16978), .ZN(n16681) );
  INV_X1 U14258 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11031) );
  INV_X1 U14259 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11030) );
  NAND2_X1 U14260 ( .A1(n11031), .A2(n11030), .ZN(n11032) );
  INV_X1 U14261 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16360) );
  INV_X1 U14262 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16356) );
  NAND2_X1 U14263 ( .A1(n11033), .A2(n16356), .ZN(n11079) );
  NAND2_X1 U14264 ( .A1(n11079), .A2(n11095), .ZN(n11077) );
  INV_X1 U14265 ( .A(n11033), .ZN(n11037) );
  AND3_X1 U14266 ( .A1(n11037), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n20273), .ZN(
        n11034) );
  OR2_X1 U14267 ( .A1(n11077), .A2(n11034), .ZN(n15993) );
  INV_X1 U14268 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16603) );
  OAI21_X1 U14269 ( .B1(n15993), .B2(n11555), .A(n16603), .ZN(n16596) );
  INV_X1 U14270 ( .A(n11035), .ZN(n11042) );
  NAND2_X1 U14271 ( .A1(n11042), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11036) );
  MUX2_X1 U14272 ( .A(n11042), .B(n11036), .S(n20273), .Z(n11038) );
  NAND2_X1 U14273 ( .A1(n15997), .A2(n11559), .ZN(n11039) );
  INV_X1 U14274 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12469) );
  NAND2_X1 U14275 ( .A1(n11039), .A2(n12469), .ZN(n16597) );
  NAND2_X1 U14276 ( .A1(n9715), .A2(n11040), .ZN(n11041) );
  NAND2_X1 U14277 ( .A1(n11042), .A2(n11041), .ZN(n16016) );
  OR2_X1 U14278 ( .A1(n16016), .A2(n11555), .ZN(n11043) );
  INV_X1 U14279 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16615) );
  NAND2_X1 U14280 ( .A1(n11043), .A2(n16615), .ZN(n16613) );
  INV_X1 U14281 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n16379) );
  NAND2_X1 U14282 ( .A1(n10380), .A2(n16379), .ZN(n11047) );
  INV_X1 U14283 ( .A(n11095), .ZN(n11044) );
  AOI21_X1 U14284 ( .B1(n11054), .B2(n11045), .A(n11044), .ZN(n11046) );
  NAND2_X1 U14285 ( .A1(n16072), .A2(n11559), .ZN(n11048) );
  XNOR2_X1 U14286 ( .A(n11048), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16642) );
  NAND2_X1 U14287 ( .A1(n9709), .A2(n9758), .ZN(n11049) );
  NAND2_X1 U14288 ( .A1(n11060), .A2(n11049), .ZN(n16053) );
  OR2_X1 U14289 ( .A1(n16053), .A2(n11555), .ZN(n11050) );
  NAND2_X1 U14290 ( .A1(n11050), .A2(n10094), .ZN(n16632) );
  XNOR2_X1 U14291 ( .A(n11051), .B(n9761), .ZN(n16102) );
  NAND2_X1 U14292 ( .A1(n16102), .A2(n11559), .ZN(n11071) );
  INV_X1 U14293 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U14294 ( .A1(n11071), .A2(n16961), .ZN(n16670) );
  OR2_X1 U14295 ( .A1(n16122), .A2(n11555), .ZN(n11052) );
  NAND2_X1 U14296 ( .A1(n11052), .A2(n16978), .ZN(n16682) );
  AND2_X1 U14297 ( .A1(n16670), .A2(n16682), .ZN(n12451) );
  OR2_X1 U14298 ( .A1(n11056), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11058) );
  AND2_X1 U14299 ( .A1(n20273), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U14300 ( .A1(n11058), .A2(n11053), .ZN(n11055) );
  NAND2_X1 U14301 ( .A1(n11055), .A2(n11054), .ZN(n16084) );
  INV_X1 U14302 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16936) );
  OAI21_X1 U14303 ( .B1(n16084), .B2(n11555), .A(n16936), .ZN(n16651) );
  NAND2_X1 U14304 ( .A1(n20273), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11057) );
  MUX2_X1 U14305 ( .A(n20273), .B(n11057), .S(n11056), .Z(n11059) );
  NAND2_X1 U14306 ( .A1(n11059), .A2(n11058), .ZN(n16094) );
  INV_X1 U14307 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16955) );
  NAND2_X1 U14308 ( .A1(n11072), .A2(n16955), .ZN(n16661) );
  AND4_X1 U14309 ( .A1(n16632), .A2(n12451), .A3(n16651), .A4(n16661), .ZN(
        n11062) );
  XNOR2_X1 U14310 ( .A(n11060), .B(n9764), .ZN(n16036) );
  NAND2_X1 U14311 ( .A1(n16036), .A2(n11559), .ZN(n11061) );
  INV_X1 U14312 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16626) );
  NAND2_X1 U14313 ( .A1(n11061), .A2(n16626), .ZN(n16621) );
  AND4_X1 U14314 ( .A1(n16613), .A2(n16642), .A3(n11062), .A4(n16621), .ZN(
        n11063) );
  INV_X1 U14315 ( .A(n15993), .ZN(n11066) );
  NOR2_X1 U14316 ( .A1(n11555), .A2(n16603), .ZN(n11065) );
  NAND2_X1 U14317 ( .A1(n11066), .A2(n11065), .ZN(n16595) );
  INV_X1 U14318 ( .A(n16036), .ZN(n11067) );
  AND2_X1 U14319 ( .A1(n16612), .A2(n16620), .ZN(n12453) );
  OR3_X1 U14320 ( .A1(n16053), .A2(n11555), .A3(n10094), .ZN(n16631) );
  NOR2_X1 U14321 ( .A1(n11555), .A2(n10406), .ZN(n11068) );
  NAND2_X1 U14322 ( .A1(n16072), .A2(n11068), .ZN(n12452) );
  INV_X1 U14323 ( .A(n16084), .ZN(n11070) );
  NOR2_X1 U14324 ( .A1(n11555), .A2(n16936), .ZN(n11069) );
  NAND2_X1 U14325 ( .A1(n11070), .A2(n11069), .ZN(n16650) );
  NAND4_X1 U14326 ( .A1(n16631), .A2(n12452), .A3(n16650), .A4(n16671), .ZN(
        n11073) );
  NOR2_X1 U14327 ( .A1(n11072), .A2(n16955), .ZN(n16660) );
  NOR2_X1 U14328 ( .A1(n11073), .A2(n16660), .ZN(n11075) );
  NOR2_X1 U14329 ( .A1(n11555), .A2(n12469), .ZN(n11074) );
  NAND2_X1 U14330 ( .A1(n15997), .A2(n11074), .ZN(n16598) );
  AND4_X1 U14331 ( .A1(n16595), .A2(n12453), .A3(n11075), .A4(n16598), .ZN(
        n11076) );
  NAND2_X1 U14332 ( .A1(n20273), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14333 ( .A1(n11079), .A2(n10370), .ZN(n11080) );
  NAND2_X1 U14334 ( .A1(n11083), .A2(n11080), .ZN(n15979) );
  OR2_X1 U14335 ( .A1(n15979), .A2(n11555), .ZN(n11081) );
  INV_X1 U14336 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11278) );
  NAND2_X1 U14337 ( .A1(n11081), .A2(n11278), .ZN(n16586) );
  OR3_X1 U14338 ( .A1(n15979), .A2(n11555), .A3(n11278), .ZN(n16585) );
  AND2_X1 U14339 ( .A1(n20273), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11082) );
  NAND2_X1 U14340 ( .A1(n11083), .A2(n11082), .ZN(n11084) );
  NAND2_X1 U14341 ( .A1(n9682), .A2(n11084), .ZN(n15958) );
  OR2_X1 U14342 ( .A1(n15958), .A2(n11555), .ZN(n11085) );
  XNOR2_X1 U14343 ( .A(n11085), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16573) );
  INV_X1 U14344 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U14345 ( .A1(n11095), .A2(n11559), .ZN(n16564) );
  INV_X1 U14346 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16843) );
  NAND2_X1 U14347 ( .A1(n16564), .A2(n16843), .ZN(n11548) );
  NAND2_X1 U14348 ( .A1(n11551), .A2(n11548), .ZN(n16556) );
  NAND2_X1 U14349 ( .A1(n20273), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11089) );
  MUX2_X1 U14350 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n11089), .S(n11094), .Z(
        n11090) );
  NAND2_X1 U14351 ( .A1(n15917), .A2(n11559), .ZN(n11091) );
  NAND2_X1 U14352 ( .A1(n11091), .A2(n16830), .ZN(n16554) );
  INV_X1 U14353 ( .A(n16554), .ZN(n11093) );
  NOR2_X1 U14354 ( .A1(n11555), .A2(n16830), .ZN(n11092) );
  NAND2_X1 U14355 ( .A1(n15917), .A2(n11092), .ZN(n16553) );
  OAI21_X1 U14356 ( .B1(n16556), .B2(n11093), .A(n16553), .ZN(n11096) );
  INV_X1 U14357 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16330) );
  OR2_X1 U14358 ( .A1(n11543), .A2(n11555), .ZN(n11552) );
  XNOR2_X1 U14359 ( .A(n11096), .B(n11549), .ZN(n16826) );
  INV_X1 U14360 ( .A(n13617), .ZN(n11097) );
  INV_X1 U14361 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U14362 ( .A1(n11186), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11099) );
  AOI21_X1 U14363 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11100), .ZN(n11160) );
  INV_X1 U14364 ( .A(n11101), .ZN(n11102) );
  INV_X1 U14365 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14366 ( .A1(n11186), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11103) );
  AOI21_X1 U14367 ( .B1(n11185), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11105), .ZN(n16226) );
  INV_X1 U14368 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14369 ( .A1(n11098), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11106) );
  AOI21_X1 U14370 ( .B1(n9585), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11107), .ZN(n14098) );
  NAND2_X1 U14371 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11109) );
  INV_X1 U14372 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U14373 ( .A1(n11186), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11108) );
  NAND2_X1 U14374 ( .A1(n11109), .A2(n9689), .ZN(n14204) );
  AND2_X2 U14375 ( .A1(n14096), .A2(n14204), .ZN(n14203) );
  NAND2_X1 U14376 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11112) );
  INV_X1 U14377 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n16419) );
  OAI22_X1 U14378 ( .A1(n11173), .A2(n16419), .B1(n17290), .B2(n16760), .ZN(
        n11110) );
  AOI21_X1 U14379 ( .B1(n11175), .B2(P2_REIP_REG_7__SCAN_IN), .A(n11110), .ZN(
        n11111) );
  NAND2_X1 U14380 ( .A1(n11112), .A2(n11111), .ZN(n16190) );
  INV_X1 U14381 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20819) );
  AOI22_X1 U14382 ( .A1(n11098), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11113) );
  AOI21_X1 U14383 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11114), .ZN(n16177) );
  INV_X1 U14384 ( .A(n16177), .ZN(n11115) );
  INV_X1 U14385 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U14386 ( .A1(n11098), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11116) );
  AOI21_X1 U14387 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11117), .ZN(n16161) );
  INV_X1 U14388 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U14389 ( .A1(n11186), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11118) );
  AOI21_X1 U14390 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11119), .ZN(n16145) );
  NAND2_X1 U14391 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11122) );
  OAI22_X1 U14392 ( .A1(n11173), .A2(n16404), .B1(n17290), .B2(n16707), .ZN(
        n11120) );
  AOI21_X1 U14393 ( .B1(n11175), .B2(P2_REIP_REG_11__SCAN_IN), .A(n11120), 
        .ZN(n11121) );
  NAND2_X1 U14394 ( .A1(n11122), .A2(n11121), .ZN(n16133) );
  NAND2_X1 U14395 ( .A1(n16147), .A2(n16133), .ZN(n16113) );
  INV_X1 U14396 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16685) );
  AOI22_X1 U14397 ( .A1(n11186), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11123) );
  AOI21_X1 U14398 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11124), .ZN(n16115) );
  INV_X1 U14399 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16675) );
  AOI22_X1 U14400 ( .A1(n11098), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11126) );
  AOI21_X1 U14401 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11127), .ZN(n16101) );
  NAND2_X1 U14402 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11129) );
  INV_X1 U14403 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U14404 ( .A1(n11098), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11128) );
  NAND2_X1 U14405 ( .A1(n11129), .A2(n9690), .ZN(n16088) );
  NAND2_X1 U14406 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11131) );
  INV_X1 U14407 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U14408 ( .A1(n11186), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11130) );
  NAND2_X1 U14409 ( .A1(n11131), .A2(n9691), .ZN(n16076) );
  NAND2_X1 U14410 ( .A1(n16075), .A2(n16076), .ZN(n16060) );
  INV_X1 U14411 ( .A(n16060), .ZN(n11135) );
  INV_X1 U14412 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n16643) );
  AOI22_X1 U14413 ( .A1(n11098), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11132) );
  AOI21_X1 U14414 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11133), .ZN(n16061) );
  INV_X1 U14415 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U14416 ( .A1(n11098), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11136) );
  AOI21_X1 U14417 ( .B1(n9585), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11137), .ZN(n16042) );
  INV_X1 U14418 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U14419 ( .A1(n11186), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11138) );
  AOI21_X1 U14420 ( .B1(n9585), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11139), .ZN(n16029) );
  NAND2_X1 U14421 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11141) );
  INV_X1 U14422 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U14423 ( .A1(n11098), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11140) );
  NAND2_X1 U14424 ( .A1(n11141), .A2(n9692), .ZN(n16011) );
  NAND2_X1 U14425 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11144) );
  INV_X1 U14426 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12482) );
  OAI22_X1 U14427 ( .A1(n11173), .A2(n16360), .B1(n17290), .B2(n12482), .ZN(
        n11142) );
  AOI21_X1 U14428 ( .B1(n11175), .B2(P2_REIP_REG_20__SCAN_IN), .A(n11142), 
        .ZN(n11143) );
  NAND2_X1 U14429 ( .A1(n11144), .A2(n11143), .ZN(n12460) );
  AND2_X2 U14430 ( .A1(n12458), .A2(n12460), .ZN(n12457) );
  NAND2_X1 U14431 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11147) );
  INV_X1 U14432 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16605) );
  OAI22_X1 U14433 ( .A1(n11173), .A2(n16356), .B1(n17290), .B2(n16605), .ZN(
        n11145) );
  AOI21_X1 U14434 ( .B1(n11175), .B2(P2_REIP_REG_21__SCAN_IN), .A(n11145), 
        .ZN(n11146) );
  NAND2_X1 U14435 ( .A1(n11147), .A2(n11146), .ZN(n15985) );
  INV_X1 U14436 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16589) );
  AOI22_X1 U14437 ( .A1(n11186), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11148) );
  AOI21_X1 U14438 ( .B1(n9585), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11149), .ZN(n15967) );
  INV_X1 U14439 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20842) );
  AOI22_X1 U14440 ( .A1(n11186), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11150) );
  AOI21_X1 U14441 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11151), .ZN(n15949) );
  INV_X1 U14442 ( .A(n15949), .ZN(n11152) );
  AND2_X2 U14443 ( .A1(n15948), .A2(n11152), .ZN(n15932) );
  NAND2_X1 U14444 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11154) );
  INV_X1 U14445 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20844) );
  AOI22_X1 U14446 ( .A1(n11098), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11153) );
  NAND2_X1 U14447 ( .A1(n11154), .A2(n9755), .ZN(n15933) );
  NAND2_X1 U14448 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11158) );
  INV_X1 U14449 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11155) );
  OAI22_X1 U14450 ( .A1(n11173), .A2(n11155), .B1(n17290), .B2(n16557), .ZN(
        n11156) );
  AOI21_X1 U14451 ( .B1(n11175), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11156), 
        .ZN(n11157) );
  NAND2_X1 U14452 ( .A1(n11158), .A2(n11157), .ZN(n15916) );
  AOI21_X1 U14453 ( .B1(n11160), .B2(n11159), .A(n11171), .ZN(n16329) );
  OR2_X1 U14454 ( .A1(n20906), .A2(n17288), .ZN(n17109) );
  NAND2_X1 U14455 ( .A1(n17109), .A2(n20912), .ZN(n11161) );
  AND2_X1 U14456 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17120) );
  INV_X1 U14457 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U14458 ( .A1(n20050), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12834) );
  NAND2_X1 U14459 ( .A1(n17114), .A2(n12834), .ZN(n13633) );
  NAND2_X1 U14460 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12800), .ZN(
        n12799) );
  NAND2_X1 U14461 ( .A1(n12824), .A2(n11164), .ZN(n11162) );
  AND2_X1 U14462 ( .A1(n12825), .A2(n11162), .ZN(n15904) );
  NAND2_X1 U14463 ( .A1(n20209), .A2(n15904), .ZN(n11163) );
  NAND2_X1 U14464 ( .A1(n17288), .A2(n20559), .ZN(n13621) );
  NOR2_X2 U14465 ( .A1(n13621), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20179) );
  NAND2_X1 U14466 ( .A1(n20179), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16817) );
  OAI211_X1 U14467 ( .C1(n17654), .C2(n11164), .A(n11163), .B(n16817), .ZN(
        n11165) );
  INV_X1 U14468 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U14469 ( .A1(n11186), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11169) );
  AOI21_X1 U14470 ( .B1(n9626), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11170), .ZN(n15885) );
  NAND2_X1 U14471 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11177) );
  INV_X1 U14472 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15869) );
  INV_X1 U14473 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U14474 ( .A1(n11173), .A2(n15869), .B1(n17290), .B2(n11172), .ZN(
        n11174) );
  AOI21_X1 U14475 ( .B1(n11175), .B2(P2_REIP_REG_28__SCAN_IN), .A(n11174), 
        .ZN(n11176) );
  NAND2_X1 U14476 ( .A1(n11177), .A2(n11176), .ZN(n13204) );
  INV_X1 U14477 ( .A(n13204), .ZN(n11178) );
  NAND2_X1 U14478 ( .A1(n9585), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11180) );
  INV_X1 U14479 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U14480 ( .A1(n11098), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11179) );
  NAND2_X1 U14481 ( .A1(n11180), .A2(n9756), .ZN(n15850) );
  NAND2_X1 U14482 ( .A1(n13202), .A2(n15850), .ZN(n15852) );
  INV_X1 U14483 ( .A(n15852), .ZN(n11184) );
  INV_X1 U14484 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U14485 ( .A1(n11098), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11181) );
  AOI21_X1 U14486 ( .B1(n9585), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11182), .ZN(n11235) );
  INV_X1 U14487 ( .A(n11235), .ZN(n11183) );
  NAND2_X1 U14488 ( .A1(n11184), .A2(n11183), .ZN(n11237) );
  INV_X1 U14489 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20858) );
  NAND2_X1 U14490 ( .A1(n9626), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11188) );
  AOI22_X1 U14491 ( .A1(n11186), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11187) );
  XNOR2_X2 U14492 ( .A(n11237), .B(n11189), .ZN(n16530) );
  NAND2_X1 U14493 ( .A1(n11190), .A2(n11192), .ZN(n11207) );
  NAND2_X1 U14494 ( .A1(n20913), .A2(n11309), .ZN(n11193) );
  MUX2_X1 U14495 ( .A(n11193), .B(n11192), .S(n11191), .Z(n11203) );
  OAI211_X1 U14496 ( .C1(n11297), .C2(n11196), .A(n11244), .B(n11195), .ZN(
        n11200) );
  OAI21_X1 U14497 ( .B1(n11198), .B2(n11197), .A(n12775), .ZN(n11199) );
  OAI211_X1 U14498 ( .C1(n11194), .C2(n11201), .A(n11200), .B(n11199), .ZN(
        n11202) );
  NAND2_X1 U14499 ( .A1(n11203), .A2(n11202), .ZN(n11205) );
  NAND2_X1 U14500 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  INV_X1 U14501 ( .A(n11208), .ZN(n11209) );
  AOI21_X1 U14502 ( .B1(n12775), .B2(n11209), .A(n11211), .ZN(n11210) );
  NAND2_X1 U14503 ( .A1(n13680), .A2(n11211), .ZN(n11212) );
  AND2_X1 U14504 ( .A1(n11214), .A2(n11213), .ZN(n17268) );
  NAND2_X1 U14505 ( .A1(n17266), .A2(n17268), .ZN(n13637) );
  NAND2_X1 U14506 ( .A1(n11241), .A2(n10625), .ZN(n11215) );
  NAND2_X1 U14507 ( .A1(n11215), .A2(n11297), .ZN(n17129) );
  NAND2_X1 U14508 ( .A1(n11216), .A2(n10625), .ZN(n11217) );
  NAND2_X1 U14509 ( .A1(n11217), .A2(n12774), .ZN(n11248) );
  NAND2_X1 U14510 ( .A1(n17129), .A2(n11248), .ZN(n11219) );
  NAND2_X1 U14511 ( .A1(n11219), .A2(n11218), .ZN(n11231) );
  INV_X1 U14512 ( .A(n11221), .ZN(n20915) );
  AOI22_X1 U14513 ( .A1(n20915), .A2(n17205), .B1(n17183), .B2(n17239), .ZN(
        n11228) );
  NAND2_X1 U14514 ( .A1(n11222), .A2(n11223), .ZN(n11224) );
  NAND2_X1 U14515 ( .A1(n11224), .A2(n11221), .ZN(n11225) );
  NAND2_X1 U14516 ( .A1(n11225), .A2(n10622), .ZN(n11227) );
  NAND2_X1 U14517 ( .A1(n11226), .A2(n10599), .ZN(n13580) );
  AND4_X1 U14518 ( .A1(n11229), .A2(n11228), .A3(n11227), .A4(n13580), .ZN(
        n11230) );
  NAND2_X1 U14519 ( .A1(n17127), .A2(n10599), .ZN(n14040) );
  NAND2_X1 U14520 ( .A1(n13637), .A2(n14040), .ZN(n11232) );
  AND2_X1 U14521 ( .A1(n16418), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11233) );
  AOI21_X1 U14522 ( .B1(n16530), .B2(n20112), .A(n11233), .ZN(n11234) );
  NAND2_X1 U14523 ( .A1(n15852), .A2(n11235), .ZN(n11236) );
  NAND2_X1 U14524 ( .A1(n11238), .A2(n11244), .ZN(n11239) );
  NAND2_X1 U14525 ( .A1(n11239), .A2(n17205), .ZN(n11240) );
  INV_X1 U14526 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20799) );
  NAND2_X1 U14527 ( .A1(n20799), .A2(n20806), .ZN(n20049) );
  OAI211_X1 U14528 ( .C1(n20799), .C2(n20806), .A(n20789), .B(n20049), .ZN(
        n20794) );
  INV_X1 U14529 ( .A(n20917), .ZN(n20910) );
  NOR2_X1 U14530 ( .A1(n20794), .A2(n20910), .ZN(n13640) );
  NAND2_X1 U14531 ( .A1(n11241), .A2(n10596), .ZN(n11250) );
  NAND2_X1 U14532 ( .A1(n16324), .A2(n17205), .ZN(n11264) );
  NAND2_X1 U14533 ( .A1(n11264), .A2(n11244), .ZN(n11245) );
  NAND2_X1 U14534 ( .A1(n11245), .A2(n10613), .ZN(n11246) );
  NAND2_X1 U14535 ( .A1(n11246), .A2(n10596), .ZN(n11247) );
  NAND2_X1 U14536 ( .A1(n11248), .A2(n11247), .ZN(n11249) );
  AOI21_X1 U14537 ( .B1(n11250), .B2(n11243), .A(n11249), .ZN(n11266) );
  NAND3_X1 U14538 ( .A1(n11258), .A2(n13611), .A3(n13640), .ZN(n11252) );
  AND2_X1 U14539 ( .A1(n11266), .A2(n11252), .ZN(n13636) );
  NOR2_X1 U14540 ( .A1(n10935), .A2(n16324), .ZN(n11253) );
  NAND2_X1 U14541 ( .A1(n20898), .A2(n11253), .ZN(n11256) );
  MUX2_X1 U14542 ( .A(n11258), .B(n17239), .S(n16324), .Z(n11254) );
  NAND3_X1 U14543 ( .A1(n11254), .A2(n13611), .A3(n20917), .ZN(n11255) );
  NAND2_X1 U14544 ( .A1(n11258), .A2(n17183), .ZN(n12838) );
  NAND2_X1 U14545 ( .A1(n11259), .A2(n12838), .ZN(n17161) );
  NAND2_X1 U14546 ( .A1(n17161), .A2(n16324), .ZN(n11261) );
  NAND2_X1 U14547 ( .A1(n11261), .A2(n11260), .ZN(n11262) );
  NAND2_X1 U14548 ( .A1(n17127), .A2(n11223), .ZN(n11263) );
  NOR2_X1 U14549 ( .A1(n16909), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20231) );
  INV_X1 U14550 ( .A(n11264), .ZN(n11265) );
  NAND2_X1 U14551 ( .A1(n11266), .A2(n11265), .ZN(n14043) );
  INV_X1 U14552 ( .A(n14043), .ZN(n17267) );
  NOR2_X1 U14553 ( .A1(n20202), .A2(n17125), .ZN(n20250) );
  NOR2_X1 U14554 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20250), .ZN(
        n11281) );
  INV_X1 U14555 ( .A(n11281), .ZN(n11267) );
  NOR2_X1 U14556 ( .A1(n20217), .A2(n11267), .ZN(n20230) );
  NOR2_X1 U14557 ( .A1(n20231), .A2(n20230), .ZN(n11270) );
  OR2_X1 U14558 ( .A1(n16909), .A2(n20250), .ZN(n11269) );
  INV_X2 U14559 ( .A(n20179), .ZN(n20207) );
  NAND2_X1 U14560 ( .A1(n11268), .A2(n20207), .ZN(n17657) );
  AND2_X1 U14561 ( .A1(n11269), .A2(n17657), .ZN(n20235) );
  NAND2_X1 U14562 ( .A1(n20236), .A2(n17099), .ZN(n11271) );
  NOR2_X1 U14563 ( .A1(n17072), .A2(n17071), .ZN(n17070) );
  NAND2_X1 U14564 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17070), .ZN(
        n11284) );
  AND2_X1 U14565 ( .A1(n20236), .A2(n11284), .ZN(n11272) );
  NOR2_X1 U14566 ( .A1(n17024), .A2(n17040), .ZN(n17013) );
  INV_X1 U14567 ( .A(n17013), .ZN(n17026) );
  NAND2_X1 U14568 ( .A1(n20236), .A2(n17026), .ZN(n11273) );
  NOR2_X1 U14569 ( .A1(n11274), .A2(n16720), .ZN(n11286) );
  NAND2_X1 U14570 ( .A1(n17015), .A2(n11286), .ZN(n11275) );
  INV_X1 U14571 ( .A(n20236), .ZN(n16914) );
  NAND2_X1 U14572 ( .A1(n17098), .A2(n16914), .ZN(n16999) );
  NAND2_X1 U14573 ( .A1(n11275), .A2(n16999), .ZN(n16979) );
  NAND2_X1 U14574 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16947) );
  OAI21_X1 U14575 ( .B1(n16955), .B2(n16947), .A(n16999), .ZN(n11276) );
  AND2_X1 U14576 ( .A1(n16999), .A2(n16584), .ZN(n11277) );
  NOR2_X1 U14577 ( .A1(n11279), .A2(n11278), .ZN(n11292) );
  INV_X1 U14578 ( .A(n11292), .ZN(n16854) );
  AND2_X1 U14579 ( .A1(n20236), .A2(n16854), .ZN(n11280) );
  INV_X1 U14580 ( .A(n16584), .ZN(n11288) );
  NAND2_X1 U14581 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20250), .ZN(
        n20218) );
  NAND2_X1 U14582 ( .A1(n11283), .A2(n11282), .ZN(n17100) );
  NAND2_X1 U14583 ( .A1(n17100), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17086) );
  NOR2_X2 U14584 ( .A1(n17086), .A2(n11284), .ZN(n17041) );
  AND2_X1 U14585 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17013), .ZN(
        n11285) );
  NAND2_X1 U14586 ( .A1(n17041), .A2(n11285), .ZN(n17001) );
  INV_X1 U14587 ( .A(n11286), .ZN(n16985) );
  NOR2_X2 U14588 ( .A1(n17001), .A2(n16985), .ZN(n16975) );
  NAND2_X1 U14589 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16975), .ZN(
        n16962) );
  INV_X1 U14590 ( .A(n16962), .ZN(n11287) );
  AND2_X2 U14591 ( .A1(n16951), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16937) );
  AND2_X2 U14592 ( .A1(n11288), .A2(n16937), .ZN(n16865) );
  NOR2_X1 U14593 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16854), .ZN(
        n11289) );
  NAND2_X1 U14594 ( .A1(n16865), .A2(n11289), .ZN(n16842) );
  NAND2_X1 U14595 ( .A1(n20236), .A2(n16815), .ZN(n11290) );
  INV_X1 U14596 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16775) );
  NAND2_X1 U14597 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11546) );
  OAI21_X1 U14598 ( .B1(n16775), .B2(n11546), .A(n20236), .ZN(n11291) );
  AND2_X1 U14599 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11292), .ZN(
        n11293) );
  NAND2_X1 U14600 ( .A1(n16865), .A2(n11293), .ZN(n16814) );
  NOR2_X1 U14601 ( .A1(n16789), .A2(n11546), .ZN(n16776) );
  INV_X1 U14602 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12494) );
  NAND3_X1 U14603 ( .A1(n16776), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12494), .ZN(n11294) );
  OR2_X1 U14604 ( .A1(n20207), .A2(n12844), .ZN(n12439) );
  NAND2_X1 U14605 ( .A1(n11294), .A2(n12439), .ZN(n11295) );
  AOI21_X1 U14606 ( .B1(n12493), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11295), .ZN(n11296) );
  OAI21_X1 U14607 ( .B1(n13602), .B2(n20242), .A(n11296), .ZN(n11542) );
  AND2_X4 U14608 ( .A1(n13594), .A2(n11304), .ZN(n12490) );
  NAND2_X1 U14609 ( .A1(n12490), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11302) );
  INV_X1 U14610 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11299) );
  OAI211_X1 U14611 ( .C1(n10625), .C2(n11299), .A(n11298), .B(n11308), .ZN(
        n11300) );
  INV_X1 U14612 ( .A(n11300), .ZN(n11301) );
  NAND2_X1 U14613 ( .A1(n11302), .A2(n11301), .ZN(n14167) );
  INV_X1 U14614 ( .A(n11303), .ZN(n11306) );
  NAND2_X1 U14615 ( .A1(n11304), .A2(n9914), .ZN(n11488) );
  MUX2_X1 U14616 ( .A(n10625), .B(n20679), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11310) );
  NAND2_X1 U14617 ( .A1(n11309), .A2(n11308), .ZN(n11312) );
  NAND3_X1 U14618 ( .A1(n11311), .A2(n11310), .A3(n11321), .ZN(n14166) );
  NAND2_X1 U14619 ( .A1(n14167), .A2(n14166), .ZN(n11316) );
  AOI22_X1 U14620 ( .A1(n11323), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11313) );
  XNOR2_X1 U14621 ( .A(n11316), .B(n11317), .ZN(n14178) );
  AOI22_X1 U14622 ( .A1(n11314), .A2(n16324), .B1(n11307), .B2(n10625), .ZN(
        n11315) );
  MUX2_X1 U14623 ( .A(n17256), .B(n11315), .S(n11308), .Z(n14177) );
  NAND2_X1 U14624 ( .A1(n14178), .A2(n14177), .ZN(n14176) );
  INV_X1 U14625 ( .A(n11317), .ZN(n11318) );
  NAND2_X1 U14626 ( .A1(n11316), .A2(n11318), .ZN(n11319) );
  NAND2_X1 U14627 ( .A1(n14176), .A2(n11319), .ZN(n11329) );
  OR2_X1 U14628 ( .A1(n11488), .A2(n11320), .ZN(n11322) );
  OAI211_X1 U14629 ( .C1(n11308), .C2(n20894), .A(n11322), .B(n11321), .ZN(
        n11327) );
  XNOR2_X1 U14630 ( .A(n11329), .B(n11327), .ZN(n14173) );
  NAND2_X1 U14631 ( .A1(n12490), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14632 ( .A1(n12489), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11325) );
  AND2_X1 U14633 ( .A1(n11326), .A2(n11325), .ZN(n14172) );
  NAND2_X2 U14634 ( .A1(n14173), .A2(n14172), .ZN(n14175) );
  INV_X1 U14635 ( .A(n11327), .ZN(n11328) );
  NAND2_X1 U14636 ( .A1(n11329), .A2(n11328), .ZN(n11330) );
  AOI22_X1 U14637 ( .A1(n11324), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11332) );
  NAND2_X1 U14638 ( .A1(n12489), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11331) );
  AND2_X1 U14639 ( .A1(n11332), .A2(n11331), .ZN(n11336) );
  NAND2_X1 U14640 ( .A1(n12490), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U14641 ( .A1(n11305), .A2(n11333), .ZN(n11334) );
  INV_X1 U14642 ( .A(n16245), .ZN(n11337) );
  NAND2_X1 U14643 ( .A1(n12490), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14644 ( .A1(n12489), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11340) );
  OR2_X1 U14645 ( .A1(n11488), .A2(n11338), .ZN(n11339) );
  AOI22_X1 U14646 ( .A1(n12489), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11345) );
  NAND2_X1 U14647 ( .A1(n11305), .A2(n11343), .ZN(n11344) );
  OAI211_X1 U14648 ( .C1(n11342), .C2(n11346), .A(n11345), .B(n11344), .ZN(
        n16203) );
  NAND2_X1 U14649 ( .A1(n16204), .A2(n16203), .ZN(n16206) );
  NAND2_X1 U14650 ( .A1(n11305), .A2(n11347), .ZN(n11348) );
  AOI22_X1 U14651 ( .A1(n12489), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11349) );
  OAI21_X1 U14652 ( .B1(n11342), .B2(n20815), .A(n11349), .ZN(n14345) );
  AOI21_X1 U14653 ( .B1(n14344), .B2(n14345), .A(n9769), .ZN(n11350) );
  INV_X1 U14654 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20817) );
  AOI22_X1 U14655 ( .A1(n12489), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11351) );
  OAI21_X1 U14656 ( .B1(n11342), .B2(n20817), .A(n11351), .ZN(n14347) );
  NAND2_X1 U14657 ( .A1(n12490), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14658 ( .A1(n12489), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11371) );
  INV_X1 U14659 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11353) );
  INV_X1 U14660 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11352) );
  OAI22_X1 U14661 ( .A1(n13322), .A2(n11353), .B1(n13320), .B2(n11352), .ZN(
        n11356) );
  INV_X1 U14662 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11354) );
  INV_X1 U14663 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17191) );
  OAI22_X1 U14664 ( .A1(n14041), .A2(n11354), .B1(n13324), .B2(n17191), .ZN(
        n11355) );
  NOR2_X1 U14665 ( .A1(n11356), .A2(n11355), .ZN(n11368) );
  NAND2_X1 U14666 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11360) );
  NAND2_X1 U14667 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11359) );
  NAND2_X1 U14668 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11358) );
  AOI22_X1 U14669 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11357) );
  AND4_X1 U14670 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n11367) );
  AOI22_X1 U14671 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14672 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14673 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14674 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14675 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11361) );
  AND4_X1 U14676 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  NAND4_X1 U14677 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n16409) );
  INV_X1 U14678 ( .A(n16409), .ZN(n11369) );
  OR2_X1 U14679 ( .A1(n11488), .A2(n11369), .ZN(n11370) );
  NAND2_X1 U14680 ( .A1(n12490), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14681 ( .A1(n12489), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11324), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11391) );
  INV_X1 U14682 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11375) );
  OAI22_X1 U14683 ( .A1(n13322), .A2(n11375), .B1(n13320), .B2(n11374), .ZN(
        n11377) );
  OAI22_X1 U14684 ( .A1(n17198), .A2(n13324), .B1(n14041), .B2(n13420), .ZN(
        n11376) );
  NOR2_X1 U14685 ( .A1(n11377), .A2(n11376), .ZN(n11389) );
  NAND2_X1 U14686 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14687 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11380) );
  NAND2_X1 U14688 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11379) );
  AOI22_X1 U14689 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11378) );
  AND4_X1 U14690 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11388) );
  AOI22_X1 U14691 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14693 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14694 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14695 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11382) );
  AND4_X1 U14696 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  NAND4_X1 U14697 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n13258) );
  INV_X1 U14698 ( .A(n13258), .ZN(n16405) );
  OR2_X1 U14699 ( .A1(n11488), .A2(n16405), .ZN(n11390) );
  NAND2_X1 U14700 ( .A1(n11394), .A2(n11393), .ZN(n14259) );
  INV_X1 U14701 ( .A(n14259), .ZN(n11417) );
  NAND2_X1 U14702 ( .A1(n12490), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14703 ( .A1(n12489), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11414) );
  INV_X1 U14704 ( .A(n11395), .ZN(n11439) );
  OAI22_X1 U14705 ( .A1(n11439), .A2(n11396), .B1(n13320), .B2(n13233), .ZN(
        n11400) );
  INV_X1 U14706 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11398) );
  INV_X1 U14707 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11397) );
  OAI22_X1 U14708 ( .A1(n13322), .A2(n11398), .B1(n14041), .B2(n11397), .ZN(
        n11399) );
  NOR2_X1 U14709 ( .A1(n11400), .A2(n11399), .ZN(n11412) );
  NAND2_X1 U14710 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14711 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11403) );
  AOI22_X1 U14712 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14713 ( .A1(n13398), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11401) );
  AND4_X1 U14714 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n11411) );
  AOI22_X1 U14715 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11408) );
  NAND2_X1 U14716 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11407) );
  NAND2_X1 U14717 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11406) );
  NAND2_X1 U14718 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11405) );
  AND4_X1 U14719 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(
        n11410) );
  AOI22_X1 U14720 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13390), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14721 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n16392) );
  INV_X1 U14722 ( .A(n16392), .ZN(n20103) );
  OR2_X1 U14723 ( .A1(n11488), .A2(n20103), .ZN(n11413) );
  NAND2_X1 U14724 ( .A1(n11417), .A2(n11416), .ZN(n14258) );
  NAND2_X1 U14725 ( .A1(n12490), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14726 ( .A1(n12489), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11434) );
  INV_X1 U14727 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11418) );
  OAI22_X1 U14728 ( .A1(n13322), .A2(n11418), .B1(n13320), .B2(n13231), .ZN(
        n11420) );
  INV_X1 U14729 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13458) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13465) );
  OAI22_X1 U14731 ( .A1(n13458), .A2(n13324), .B1(n14041), .B2(n13465), .ZN(
        n11419) );
  NOR2_X1 U14732 ( .A1(n11420), .A2(n11419), .ZN(n11432) );
  NAND2_X1 U14733 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11424) );
  NAND2_X1 U14734 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11423) );
  NAND2_X1 U14735 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11422) );
  AOI22_X1 U14736 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11421) );
  AND4_X1 U14737 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11431) );
  AOI22_X1 U14738 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14740 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11427) );
  NAND2_X1 U14741 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11426) );
  NAND2_X1 U14742 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11425) );
  AND4_X1 U14743 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11429) );
  NAND4_X1 U14744 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n16401) );
  INV_X1 U14745 ( .A(n16401), .ZN(n16393) );
  OR2_X1 U14746 ( .A1(n11488), .A2(n16393), .ZN(n11433) );
  AOI22_X1 U14747 ( .A1(n12489), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11455) );
  INV_X1 U14748 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11436) );
  INV_X1 U14749 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13493) );
  OAI22_X1 U14750 ( .A1(n11437), .A2(n11436), .B1(n14041), .B2(n13493), .ZN(
        n11441) );
  INV_X1 U14751 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11438) );
  INV_X1 U14752 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14093) );
  OAI22_X1 U14753 ( .A1(n11439), .A2(n11438), .B1(n13320), .B2(n14093), .ZN(
        n11440) );
  NOR2_X1 U14754 ( .A1(n11441), .A2(n11440), .ZN(n11453) );
  NAND2_X1 U14755 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11445) );
  NAND2_X1 U14756 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11444) );
  AOI22_X1 U14757 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11443) );
  NAND2_X1 U14758 ( .A1(n13390), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11442) );
  AND4_X1 U14759 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11452) );
  AOI22_X1 U14760 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U14761 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11448) );
  NAND2_X1 U14762 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11447) );
  NAND2_X1 U14763 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11446) );
  AND4_X1 U14764 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11451) );
  AOI22_X1 U14765 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11450) );
  NAND4_X1 U14766 ( .A1(n11453), .A2(n11452), .A3(n11451), .A4(n11450), .ZN(
        n13257) );
  INV_X1 U14767 ( .A(n13257), .ZN(n20093) );
  OR2_X1 U14768 ( .A1(n11488), .A2(n20093), .ZN(n11454) );
  OAI211_X1 U14769 ( .C1(n11342), .C2(n16685), .A(n11455), .B(n11454), .ZN(
        n14264) );
  NAND2_X1 U14770 ( .A1(n12490), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14771 ( .A1(n12489), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11473) );
  INV_X1 U14772 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11457) );
  OAI22_X1 U14773 ( .A1(n13322), .A2(n11457), .B1(n13320), .B2(n11456), .ZN(
        n11459) );
  INV_X1 U14774 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13517) );
  INV_X1 U14775 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13509) );
  OAI22_X1 U14776 ( .A1(n14041), .A2(n13517), .B1(n13324), .B2(n13509), .ZN(
        n11458) );
  NOR2_X1 U14777 ( .A1(n11459), .A2(n11458), .ZN(n11471) );
  NAND2_X1 U14778 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U14779 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14780 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11461) );
  AOI22_X1 U14781 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11460) );
  AND4_X1 U14782 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11470) );
  AOI22_X1 U14783 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14784 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U14785 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14786 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U14787 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11464) );
  AND4_X1 U14788 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11468) );
  NAND4_X1 U14789 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n16394) );
  NAND2_X1 U14790 ( .A1(n11305), .A2(n16394), .ZN(n11472) );
  NAND2_X1 U14791 ( .A1(n12490), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14792 ( .A1(n12489), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11490) );
  NAND2_X1 U14793 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11477) );
  AOI22_X1 U14794 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11476) );
  AND2_X1 U14795 ( .A1(n11477), .A2(n11476), .ZN(n11481) );
  AOI22_X1 U14796 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13390), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14797 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14798 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14799 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11487) );
  AOI22_X1 U14800 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14801 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14802 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U14803 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11482) );
  NAND4_X1 U14804 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11486) );
  OR2_X1 U14805 ( .A1(n11488), .A2(n16387), .ZN(n11489) );
  AOI22_X1 U14806 ( .A1(n12489), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11510) );
  INV_X1 U14807 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11493) );
  OAI22_X1 U14808 ( .A1(n13322), .A2(n11493), .B1(n13320), .B2(n11492), .ZN(
        n11496) );
  INV_X1 U14809 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13563) );
  INV_X1 U14810 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11494) );
  OAI22_X1 U14811 ( .A1(n13563), .A2(n13324), .B1(n14041), .B2(n11494), .ZN(
        n11495) );
  NOR2_X1 U14812 ( .A1(n11496), .A2(n11495), .ZN(n11508) );
  NAND2_X1 U14813 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14814 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14815 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11498) );
  AOI22_X1 U14816 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10758), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11497) );
  AND4_X1 U14817 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11507) );
  AOI22_X1 U14818 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14819 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14820 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14821 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14822 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11501) );
  AND4_X1 U14823 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  NAND4_X1 U14824 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n16383) );
  NAND2_X1 U14825 ( .A1(n11305), .A2(n16383), .ZN(n11509) );
  OAI211_X1 U14826 ( .C1(n11342), .C2(n20829), .A(n11510), .B(n11509), .ZN(
        n14476) );
  AOI22_X1 U14827 ( .A1(n12489), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11511) );
  OAI21_X1 U14828 ( .B1(n11342), .B2(n16643), .A(n11511), .ZN(n16059) );
  INV_X1 U14829 ( .A(n16045), .ZN(n11515) );
  NAND2_X1 U14830 ( .A1(n12490), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14831 ( .A1(n12489), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U14832 ( .A1(n12490), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14833 ( .A1(n12489), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11516) );
  INV_X1 U14834 ( .A(n16039), .ZN(n11518) );
  NAND2_X1 U14835 ( .A1(n12490), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14836 ( .A1(n12489), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11519) );
  INV_X1 U14837 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n16000) );
  AOI22_X1 U14838 ( .A1(n12489), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11521) );
  OAI21_X1 U14839 ( .B1(n11342), .B2(n16000), .A(n11521), .ZN(n12464) );
  NAND2_X1 U14840 ( .A1(n12463), .A2(n12464), .ZN(n12462) );
  NAND2_X1 U14841 ( .A1(n12490), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14842 ( .A1(n12489), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14843 ( .A1(n12490), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14844 ( .A1(n12489), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14845 ( .A1(n12489), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11526) );
  OAI21_X1 U14846 ( .B1(n11342), .B2(n20842), .A(n11526), .ZN(n15946) );
  AOI22_X1 U14847 ( .A1(n12489), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11527) );
  OAI21_X1 U14848 ( .B1(n11342), .B2(n20844), .A(n11527), .ZN(n15931) );
  NAND2_X1 U14849 ( .A1(n15930), .A2(n15931), .ZN(n15912) );
  NAND2_X1 U14850 ( .A1(n12490), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14851 ( .A1(n12489), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11528) );
  NOR2_X2 U14852 ( .A1(n15912), .A2(n15914), .ZN(n15897) );
  NAND2_X1 U14853 ( .A1(n12490), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14854 ( .A1(n12489), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11530) );
  AND2_X1 U14855 ( .A1(n11531), .A2(n11530), .ZN(n15898) );
  INV_X1 U14856 ( .A(n15898), .ZN(n11532) );
  AOI22_X1 U14857 ( .A1(n12489), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11533) );
  OAI21_X1 U14858 ( .B1(n11342), .B2(n20851), .A(n11533), .ZN(n15883) );
  NAND2_X1 U14859 ( .A1(n12490), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14860 ( .A1(n11323), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11534) );
  AOI222_X1 U14861 ( .A1(n12490), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n12489), 
        .B2(P2_EAX_REG_29__SCAN_IN), .C1(n11324), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U14862 ( .A1(n11323), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11324), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11537) );
  OAI21_X1 U14863 ( .B1(n11342), .B2(n12844), .A(n11537), .ZN(n11538) );
  INV_X1 U14864 ( .A(n17268), .ZN(n14042) );
  NAND2_X1 U14865 ( .A1(n12838), .A2(n11243), .ZN(n17271) );
  NAND2_X1 U14866 ( .A1(n17271), .A2(n11309), .ZN(n11539) );
  NAND2_X1 U14867 ( .A1(n14042), .A2(n11539), .ZN(n11540) );
  NOR2_X1 U14868 ( .A1(n13583), .A2(n20227), .ZN(n11541) );
  NAND2_X1 U14869 ( .A1(n20273), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13188) );
  AND2_X1 U14870 ( .A1(n20273), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11544) );
  NAND2_X1 U14871 ( .A1(n13191), .A2(n11544), .ZN(n11545) );
  NOR2_X2 U14872 ( .A1(n15877), .A2(n11555), .ZN(n13192) );
  INV_X1 U14873 ( .A(n11546), .ZN(n11547) );
  NOR2_X1 U14874 ( .A1(n13192), .A2(n11547), .ZN(n12496) );
  INV_X1 U14875 ( .A(n12496), .ZN(n11554) );
  INV_X1 U14876 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16818) );
  OR2_X1 U14877 ( .A1(n11552), .A2(n16818), .ZN(n11553) );
  NAND2_X1 U14878 ( .A1(n20273), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11556) );
  XOR2_X1 U14879 ( .A(n11556), .B(n11557), .Z(n15860) );
  AOI21_X1 U14880 ( .B1(n15860), .B2(n11559), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16533) );
  NAND3_X1 U14881 ( .A1(n15860), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11559), .ZN(n16534) );
  NAND2_X1 U14882 ( .A1(n20273), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11558) );
  AOI21_X1 U14883 ( .B1(n12850), .B2(n11559), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12497) );
  INV_X1 U14884 ( .A(n12497), .ZN(n11560) );
  NAND3_X1 U14885 ( .A1(n12850), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11559), .ZN(n12499) );
  NAND2_X1 U14886 ( .A1(n11560), .A2(n12499), .ZN(n11561) );
  INV_X1 U14887 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16805) );
  INV_X1 U14888 ( .A(n17263), .ZN(n11562) );
  NAND3_X1 U14889 ( .A1(n11566), .A2(n11565), .A3(n11564), .ZN(P2_U3016) );
  AND2_X4 U14890 ( .A1(n11573), .A2(n14224), .ZN(n12324) );
  AOI22_X1 U14891 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12324), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11571) );
  AND2_X2 U14892 ( .A1(n14224), .A2(n14214), .ZN(n12332) );
  NOR2_X2 U14893 ( .A1(n11567), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11572) );
  AND2_X4 U14894 ( .A1(n11572), .A2(n14214), .ZN(n14223) );
  AOI22_X1 U14895 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11570) );
  NOR2_X4 U14896 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14215) );
  AND2_X2 U14897 ( .A1(n11573), .A2(n14215), .ZN(n11728) );
  AOI22_X1 U14898 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11728), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11569) );
  AND2_X4 U14899 ( .A1(n11574), .A2(n14215), .ZN(n12321) );
  AND2_X4 U14900 ( .A1(n14215), .A2(n14214), .ZN(n12323) );
  AOI22_X1 U14901 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11568) );
  AND2_X2 U14902 ( .A1(n11572), .A2(n14245), .ZN(n12257) );
  AND2_X2 U14903 ( .A1(n11573), .A2(n14216), .ZN(n11734) );
  AOI22_X1 U14904 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11579) );
  AND2_X2 U14905 ( .A1(n14245), .A2(n14215), .ZN(n11746) );
  AOI22_X1 U14906 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11578) );
  AND2_X2 U14907 ( .A1(n14221), .A2(n11575), .ZN(n12018) );
  AOI22_X1 U14908 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11577) );
  AND2_X4 U14909 ( .A1(n14216), .A2(n14245), .ZN(n12335) );
  AOI22_X1 U14910 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14911 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14912 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14913 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14914 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14915 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AOI22_X1 U14916 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14917 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14918 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14919 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14920 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  AOI22_X1 U14921 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14922 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14923 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14924 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11591) );
  NAND4_X1 U14925 ( .A1(n11594), .A2(n11593), .A3(n11592), .A4(n11591), .ZN(
        n11600) );
  AOI22_X1 U14926 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14927 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14928 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14929 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11595) );
  NAND4_X1 U14930 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11599) );
  AOI22_X1 U14931 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14932 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14933 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14934 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14935 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14936 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14937 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14938 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14939 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14940 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14941 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14942 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11610) );
  NAND4_X1 U14943 ( .A1(n11613), .A2(n11612), .A3(n11611), .A4(n11610), .ZN(
        n11619) );
  AOI22_X1 U14944 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14945 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14946 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14947 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U14948 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11618) );
  NAND2_X1 U14949 ( .A1(n11657), .A2(n12432), .ZN(n11620) );
  AOI22_X1 U14950 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14951 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14952 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14953 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14954 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14955 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14956 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14957 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11626) );
  AND2_X1 U14958 ( .A1(n11660), .A2(n14568), .ZN(n11630) );
  INV_X1 U14959 ( .A(n14299), .ZN(n11664) );
  AOI22_X1 U14960 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14961 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11734), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14962 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14963 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11633) );
  NAND4_X1 U14964 ( .A1(n11636), .A2(n11635), .A3(n11634), .A4(n11633), .ZN(
        n11642) );
  AOI22_X1 U14965 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14966 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14967 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14968 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11637) );
  NAND4_X1 U14969 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11641) );
  INV_X1 U14970 ( .A(n11810), .ZN(n11721) );
  AOI22_X1 U14971 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11745), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14972 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11746), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14973 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14974 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14975 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11652) );
  AOI22_X1 U14976 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14977 ( .A1(n11734), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14978 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11728), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14979 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12117), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14980 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11651) );
  OR2_X4 U14981 ( .A1(n11652), .A2(n11651), .ZN(n14542) );
  XNOR2_X1 U14982 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12599) );
  INV_X1 U14983 ( .A(n12599), .ZN(n11653) );
  OAI21_X1 U14984 ( .B1(n14542), .B2(n11653), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11654) );
  NOR2_X1 U14985 ( .A1(n11674), .A2(n11654), .ZN(n11655) );
  NOR2_X1 U14986 ( .A1(n11656), .A2(n11655), .ZN(n11670) );
  NAND2_X1 U14987 ( .A1(n12613), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11669) );
  NAND2_X1 U14988 ( .A1(n11659), .A2(n14325), .ZN(n11661) );
  NAND2_X1 U14989 ( .A1(n11661), .A2(n14317), .ZN(n11686) );
  NAND2_X1 U14990 ( .A1(n12615), .A2(n15500), .ZN(n11666) );
  NAND2_X1 U14991 ( .A1(n14309), .A2(n14304), .ZN(n12731) );
  NAND2_X1 U14992 ( .A1(n11667), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11668) );
  NAND3_X1 U14993 ( .A1(n11670), .A2(n11669), .A3(n11668), .ZN(n11698) );
  NAND2_X1 U14994 ( .A1(n11698), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11673) );
  NAND2_X1 U14995 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11701) );
  OAI21_X1 U14996 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11701), .ZN(n15722) );
  NAND2_X1 U14997 ( .A1(n17527), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11695) );
  INV_X1 U14998 ( .A(n11671), .ZN(n11672) );
  NAND2_X1 U14999 ( .A1(n11673), .A2(n11672), .ZN(n11677) );
  INV_X1 U15000 ( .A(n14222), .ZN(n11684) );
  INV_X1 U15001 ( .A(n12432), .ZN(n12605) );
  NAND2_X1 U15002 ( .A1(n13842), .A2(n12605), .ZN(n12727) );
  OR2_X1 U15003 ( .A1(n11674), .A2(n14546), .ZN(n11675) );
  OAI21_X2 U15004 ( .B1(n11676), .B2(n12624), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11697) );
  XNOR2_X2 U15005 ( .A(n11677), .B(n11697), .ZN(n14291) );
  NAND2_X1 U15006 ( .A1(n11698), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11679) );
  MUX2_X1 U15007 ( .A(n17525), .B(n12996), .S(n21307), .Z(n11678) );
  INV_X1 U15008 ( .A(n11680), .ZN(n11681) );
  OAI21_X1 U15009 ( .B1(n9625), .B2(n11682), .A(n11681), .ZN(n11693) );
  INV_X1 U15010 ( .A(n11683), .ZN(n11690) );
  NAND2_X1 U15011 ( .A1(n11684), .A2(n9602), .ZN(n12741) );
  NAND2_X1 U15012 ( .A1(n11686), .A2(n14436), .ZN(n11688) );
  NAND2_X1 U15013 ( .A1(n15504), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20930) );
  INV_X1 U15014 ( .A(n20930), .ZN(n11687) );
  NAND3_X1 U15015 ( .A1(n12741), .A2(n11688), .A3(n11687), .ZN(n11689) );
  NOR2_X1 U15016 ( .A1(n11690), .A2(n11689), .ZN(n11692) );
  NAND3_X1 U15017 ( .A1(n12615), .A2(n14542), .A3(n15500), .ZN(n11691) );
  NAND3_X1 U15018 ( .A1(n11693), .A2(n11692), .A3(n11691), .ZN(n11742) );
  NAND2_X2 U15019 ( .A1(n14291), .A2(n11725), .ZN(n11724) );
  AND2_X1 U15020 ( .A1(n11695), .A2(n11694), .ZN(n11696) );
  NAND2_X1 U15021 ( .A1(n11724), .A2(n11707), .ZN(n11705) );
  NAND2_X1 U15022 ( .A1(n11699), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11704) );
  INV_X1 U15023 ( .A(n12996), .ZN(n11806) );
  INV_X1 U15024 ( .A(n11701), .ZN(n11700) );
  NAND2_X1 U15025 ( .A1(n11700), .A2(n21203), .ZN(n14355) );
  NAND2_X1 U15026 ( .A1(n11701), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11702) );
  NAND2_X1 U15027 ( .A1(n14355), .A2(n11702), .ZN(n15538) );
  NAND2_X1 U15028 ( .A1(n11806), .A2(n15538), .ZN(n11703) );
  INV_X1 U15029 ( .A(n11706), .ZN(n11708) );
  NAND3_X1 U15030 ( .A1(n11724), .A2(n11708), .A3(n11707), .ZN(n11709) );
  INV_X1 U15031 ( .A(n14223), .ZN(n11733) );
  AOI22_X1 U15032 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U15033 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U15034 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U15035 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11710) );
  NAND4_X1 U15036 ( .A1(n11713), .A2(n11712), .A3(n11711), .A4(n11710), .ZN(
        n11719) );
  AOI22_X1 U15037 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U15038 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U15039 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U15040 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11714) );
  NAND4_X1 U15041 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11718) );
  AOI22_X1 U15042 ( .A1(n11721), .A2(n11720), .B1(n12397), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11722) );
  INV_X1 U15043 ( .A(n14291), .ZN(n11727) );
  AOI22_X1 U15044 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U15045 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U15046 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U15047 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U15048 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11740) );
  AOI22_X1 U15049 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U15050 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U15051 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U15052 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11735) );
  NAND4_X1 U15053 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11739) );
  NAND2_X1 U15054 ( .A1(n11767), .A2(n12525), .ZN(n11741) );
  INV_X1 U15055 ( .A(n11742), .ZN(n11743) );
  AOI22_X1 U15056 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U15057 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U15058 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U15059 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U15060 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11756) );
  AOI22_X1 U15061 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U15062 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U15063 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U15064 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U15065 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11755) );
  AOI22_X1 U15066 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12331), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15067 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11835), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U15068 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12322), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U15069 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11757) );
  NAND4_X1 U15070 ( .A1(n11760), .A2(n11759), .A3(n11758), .A4(n11757), .ZN(
        n11766) );
  AOI22_X1 U15071 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U15072 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12256), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U15073 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U15074 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U15075 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11765) );
  XNOR2_X1 U15076 ( .A(n12506), .B(n12531), .ZN(n11768) );
  NAND2_X1 U15077 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  INV_X1 U15078 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11771) );
  NOR2_X1 U15079 ( .A1(n12387), .A2(n11771), .ZN(n11774) );
  INV_X1 U15080 ( .A(n12525), .ZN(n11772) );
  OAI21_X1 U15081 ( .B1(n11772), .B2(n11810), .A(n11809), .ZN(n11773) );
  INV_X2 U15082 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U15083 ( .A1(n12605), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11851) );
  INV_X2 U15084 ( .A(n12295), .ZN(n14538) );
  XNOR2_X1 U15085 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21015) );
  AOI21_X1 U15086 ( .B1(n14538), .B2(n21015), .A(n12351), .ZN(n11777) );
  NAND2_X1 U15087 ( .A1(n12352), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11776) );
  OAI211_X1 U15088 ( .C1(n11851), .C2(n14233), .A(n11777), .B(n11776), .ZN(
        n11778) );
  INV_X1 U15089 ( .A(n11778), .ZN(n11779) );
  NAND2_X1 U15090 ( .A1(n12351), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11801) );
  AOI22_X1 U15091 ( .A1(n12352), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11775), .ZN(n11783) );
  INV_X1 U15092 ( .A(n11851), .ZN(n11792) );
  NAND2_X1 U15093 ( .A1(n11792), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11782) );
  AND2_X1 U15094 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  INV_X1 U15095 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15544) );
  NAND2_X1 U15096 ( .A1(n14541), .A2(n12531), .ZN(n11785) );
  OAI211_X1 U15097 ( .C1(n12387), .C2(n15544), .A(n11786), .B(n11785), .ZN(
        n11787) );
  NAND2_X1 U15098 ( .A1(n15559), .A2(n9602), .ZN(n11789) );
  NAND2_X1 U15099 ( .A1(n11789), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U15100 ( .A1(n14290), .A2(n12027), .ZN(n11794) );
  AOI22_X1 U15101 ( .A1(n11792), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n11791), .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U15102 ( .A1(n11794), .A2(n11793), .ZN(n13818) );
  AND2_X1 U15103 ( .A1(n11775), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U15104 ( .A1(n13819), .A2(n11796), .ZN(n13817) );
  INV_X1 U15105 ( .A(n11796), .ZN(n11797) );
  NAND2_X1 U15106 ( .A1(n11797), .A2(n12295), .ZN(n11798) );
  INV_X1 U15107 ( .A(n11802), .ZN(n11803) );
  NAND2_X1 U15108 ( .A1(n11699), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11808) );
  NAND3_X1 U15109 ( .A1(n17510), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15641) );
  INV_X1 U15110 ( .A(n15641), .ZN(n11804) );
  NAND2_X1 U15111 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11804), .ZN(
        n14394) );
  NAND2_X1 U15112 ( .A1(n17510), .A2(n14394), .ZN(n11805) );
  NOR3_X1 U15113 ( .A1(n17510), .A2(n21203), .A3(n14356), .ZN(n14289) );
  NAND2_X1 U15114 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14289), .ZN(
        n14293) );
  AOI22_X1 U15115 ( .A1(n11806), .A2(n15681), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17527), .ZN(n11807) );
  AOI22_X1 U15116 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15117 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U15118 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15119 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U15120 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11820) );
  AOI22_X1 U15121 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U15122 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U15123 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U15124 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11815) );
  NAND4_X1 U15125 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11819) );
  AOI22_X1 U15126 ( .A1(n12405), .A2(n12518), .B1(n12397), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11821) );
  NAND2_X1 U15127 ( .A1(n15526), .A2(n12027), .ZN(n11832) );
  NAND2_X1 U15128 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11825) );
  INV_X1 U15129 ( .A(n11825), .ZN(n11824) );
  INV_X1 U15130 ( .A(n11852), .ZN(n11827) );
  INV_X1 U15131 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U15132 ( .A1(n14889), .A2(n11825), .ZN(n11826) );
  NAND2_X1 U15133 ( .A1(n11827), .A2(n11826), .ZN(n14890) );
  AOI22_X1 U15134 ( .A1(n14890), .A2(n14538), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11829) );
  NAND2_X1 U15135 ( .A1(n12352), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11828) );
  OAI211_X1 U15136 ( .C1(n11851), .C2(n11823), .A(n11829), .B(n11828), .ZN(
        n11830) );
  INV_X1 U15137 ( .A(n11830), .ZN(n11831) );
  AOI22_X1 U15138 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15139 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U15140 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15141 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11836) );
  NAND4_X1 U15142 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11845) );
  AOI22_X1 U15143 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U15144 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U15145 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U15146 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11840) );
  NAND4_X1 U15147 ( .A1(n11843), .A2(n11842), .A3(n11841), .A4(n11840), .ZN(
        n11844) );
  NAND2_X1 U15148 ( .A1(n12405), .A2(n12520), .ZN(n11847) );
  NAND2_X1 U15149 ( .A1(n12397), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U15150 ( .A1(n11847), .A2(n11846), .ZN(n11858) );
  XNOR2_X1 U15151 ( .A(n11857), .B(n11858), .ZN(n12517) );
  INV_X1 U15152 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11850) );
  NAND2_X1 U15153 ( .A1(n11775), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11849) );
  NAND2_X1 U15154 ( .A1(n12352), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11848) );
  OAI211_X1 U15155 ( .C1(n11851), .C2(n11850), .A(n11849), .B(n11848), .ZN(
        n11853) );
  OAI21_X1 U15156 ( .B1(n11852), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11871), .ZN(n21105) );
  MUX2_X1 U15157 ( .A(n11853), .B(n21105), .S(n14538), .Z(n11854) );
  AOI21_X1 U15158 ( .B1(n12517), .B2(n12027), .A(n11854), .ZN(n14387) );
  AOI22_X1 U15159 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U15160 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11861) );
  INV_X1 U15161 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U15162 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U15163 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U15164 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11868) );
  AOI22_X1 U15165 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U15166 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15167 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U15168 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11863) );
  NAND4_X1 U15169 ( .A1(n11866), .A2(n11865), .A3(n11864), .A4(n11863), .ZN(
        n11867) );
  NAND2_X1 U15170 ( .A1(n12405), .A2(n12565), .ZN(n11870) );
  NAND2_X1 U15171 ( .A1(n12397), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U15172 ( .A1(n11870), .A2(n11869), .ZN(n11877) );
  INV_X1 U15173 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11875) );
  AND2_X1 U15174 ( .A1(n11871), .A2(n14877), .ZN(n11872) );
  OR2_X1 U15175 ( .A1(n11872), .A2(n11891), .ZN(n17590) );
  INV_X1 U15176 ( .A(n12351), .ZN(n11904) );
  NOR2_X1 U15177 ( .A1(n11904), .A2(n14877), .ZN(n11873) );
  AOI21_X1 U15178 ( .B1(n17590), .B2(n14538), .A(n11873), .ZN(n11874) );
  OAI21_X1 U15179 ( .B1(n12346), .B2(n11875), .A(n11874), .ZN(n11876) );
  AOI21_X1 U15180 ( .B1(n12508), .B2(n12027), .A(n11876), .ZN(n14485) );
  INV_X1 U15181 ( .A(n11877), .ZN(n11878) );
  AOI22_X1 U15182 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15183 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U15184 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15185 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U15186 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11888) );
  AOI22_X1 U15187 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U15188 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U15189 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15190 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U15191 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  NAND2_X1 U15192 ( .A1(n12405), .A2(n12564), .ZN(n11890) );
  NAND2_X1 U15193 ( .A1(n12397), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U15194 ( .A1(n9712), .A2(n11895), .ZN(n12553) );
  INV_X1 U15195 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21057) );
  OR2_X1 U15196 ( .A1(n11891), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11892) );
  NAND2_X1 U15197 ( .A1(n11900), .A2(n11892), .ZN(n20982) );
  AOI22_X1 U15198 ( .A1(n20982), .A2(n14538), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11893) );
  OAI21_X1 U15199 ( .B1(n12346), .B2(n21057), .A(n11893), .ZN(n11894) );
  INV_X1 U15200 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U15201 ( .A1(n12405), .A2(n12572), .ZN(n11897) );
  OAI21_X1 U15202 ( .B1(n11898), .B2(n12387), .A(n11897), .ZN(n11899) );
  XNOR2_X1 U15203 ( .A(n12554), .B(n11899), .ZN(n12563) );
  NAND2_X1 U15204 ( .A1(n12563), .A2(n12027), .ZN(n11907) );
  NAND2_X1 U15205 ( .A1(n11900), .A2(n20981), .ZN(n11902) );
  INV_X1 U15206 ( .A(n11931), .ZN(n11901) );
  NAND2_X1 U15207 ( .A1(n11902), .A2(n11901), .ZN(n20967) );
  NAND2_X1 U15208 ( .A1(n20967), .A2(n14538), .ZN(n11903) );
  OAI21_X1 U15209 ( .B1(n20981), .B2(n11904), .A(n11903), .ZN(n11905) );
  AOI21_X1 U15210 ( .B1(n12352), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11905), .ZN(
        n11906) );
  AOI22_X1 U15211 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15212 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12256), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15213 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11835), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15214 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U15215 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U15216 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n12333), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15217 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12322), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15218 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15219 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U15220 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  OAI21_X1 U15221 ( .B1(n11917), .B2(n11916), .A(n12027), .ZN(n11920) );
  XNOR2_X1 U15222 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11931), .ZN(
        n15259) );
  AOI22_X1 U15223 ( .A1(n14538), .A2(n15259), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U15224 ( .A1(n12352), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15225 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15226 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15227 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15228 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U15229 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11930) );
  AOI22_X1 U15230 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15231 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15232 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15233 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11925) );
  NAND4_X1 U15234 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11929) );
  OAI21_X1 U15235 ( .B1(n11930), .B2(n11929), .A(n12027), .ZN(n11935) );
  INV_X1 U15236 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15248) );
  XOR2_X1 U15237 ( .A(n15248), .B(n11946), .Z(n20951) );
  INV_X1 U15238 ( .A(n20951), .ZN(n11932) );
  AOI22_X1 U15239 ( .A1(n12351), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14538), .B2(n11932), .ZN(n11934) );
  NAND2_X1 U15240 ( .A1(n12352), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15241 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15242 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15243 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15244 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11936) );
  NAND4_X1 U15245 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11945) );
  AOI22_X1 U15246 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15247 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15248 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15249 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11940) );
  NAND4_X1 U15250 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11944) );
  NOR2_X1 U15251 ( .A1(n11945), .A2(n11944), .ZN(n11951) );
  INV_X1 U15252 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11948) );
  XNOR2_X1 U15253 ( .A(n11948), .B(n11952), .ZN(n15241) );
  AOI22_X1 U15254 ( .A1(n15241), .A2(n14538), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U15255 ( .A1(n12352), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11949) );
  OAI211_X1 U15256 ( .C1(n9890), .C2(n11951), .A(n11950), .B(n11949), .ZN(
        n14849) );
  NAND2_X1 U15257 ( .A1(n12352), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11959) );
  INV_X1 U15258 ( .A(n11954), .ZN(n11956) );
  INV_X1 U15259 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U15260 ( .A1(n11956), .A2(n11955), .ZN(n11957) );
  NAND2_X1 U15261 ( .A1(n12030), .A2(n11957), .ZN(n17562) );
  AOI22_X1 U15262 ( .A1(n17562), .A2(n14538), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U15263 ( .A1(n11959), .A2(n11958), .ZN(n14786) );
  AOI22_X1 U15264 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15265 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15266 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15267 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U15268 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11969) );
  AOI22_X1 U15269 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15270 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15271 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15272 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U15273 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11968) );
  OR2_X1 U15274 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AND2_X1 U15275 ( .A1(n12027), .A2(n11970), .ZN(n14809) );
  AOI22_X1 U15276 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15277 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15278 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15279 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U15280 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11980) );
  AOI22_X1 U15281 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15282 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15283 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15284 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15285 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  OAI21_X1 U15286 ( .B1(n11980), .B2(n11979), .A(n12027), .ZN(n11986) );
  NAND2_X1 U15287 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U15288 ( .A1(n12053), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11982) );
  INV_X1 U15289 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14796) );
  XNOR2_X1 U15290 ( .A(n11982), .B(n14796), .ZN(n15189) );
  NAND2_X1 U15291 ( .A1(n15189), .A2(n14538), .ZN(n11985) );
  NAND2_X1 U15292 ( .A1(n12352), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U15293 ( .A1(n12351), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11983) );
  NAND4_X1 U15294 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n14792) );
  INV_X1 U15295 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21043) );
  INV_X1 U15296 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14836) );
  XNOR2_X1 U15297 ( .A(n12030), .B(n14836), .ZN(n15219) );
  AOI22_X1 U15298 ( .A1(n15219), .A2(n14538), .B1(n12351), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15299 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15300 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15301 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15302 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U15303 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11996) );
  AOI22_X1 U15304 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15305 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15306 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15307 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U15308 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  OR2_X1 U15309 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  NAND2_X1 U15310 ( .A1(n12027), .A2(n11997), .ZN(n11998) );
  OAI211_X1 U15311 ( .C1(n12346), .C2(n21043), .A(n11999), .B(n11998), .ZN(
        n14810) );
  OAI211_X1 U15312 ( .C1(n14786), .C2(n14809), .A(n14792), .B(n14810), .ZN(
        n12000) );
  INV_X1 U15313 ( .A(n12000), .ZN(n12037) );
  AOI22_X1 U15314 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15315 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15316 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15317 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12001) );
  NAND4_X1 U15318 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12010) );
  AOI22_X1 U15319 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15320 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15321 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15322 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U15323 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12009) );
  OAI21_X1 U15324 ( .B1(n12010), .B2(n12009), .A(n12027), .ZN(n12016) );
  INV_X1 U15325 ( .A(n12053), .ZN(n12012) );
  INV_X1 U15326 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12011) );
  XNOR2_X1 U15327 ( .A(n12012), .B(n12011), .ZN(n17547) );
  NAND2_X1 U15328 ( .A1(n17547), .A2(n14538), .ZN(n12015) );
  NAND2_X1 U15329 ( .A1(n12352), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U15330 ( .A1(n12351), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12013) );
  NAND4_X1 U15331 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n14791) );
  AOI22_X1 U15332 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15333 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15334 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12018), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15335 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15336 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12029) );
  AOI22_X1 U15337 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15338 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15339 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15340 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12023) );
  NAND4_X1 U15341 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12028) );
  OAI21_X1 U15342 ( .B1(n12029), .B2(n12028), .A(n12027), .ZN(n12036) );
  NAND2_X1 U15343 ( .A1(n12351), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U15344 ( .A1(n12352), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12034) );
  INV_X1 U15345 ( .A(n12030), .ZN(n12031) );
  NAND2_X1 U15346 ( .A1(n12031), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12032) );
  INV_X1 U15347 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14817) );
  XNOR2_X1 U15348 ( .A(n12032), .B(n14817), .ZN(n15212) );
  NAND2_X1 U15349 ( .A1(n15212), .A2(n14538), .ZN(n12033) );
  NAND4_X1 U15350 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n14811) );
  AOI22_X1 U15351 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n9607), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15352 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12322), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15353 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15354 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12333), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15355 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12048) );
  AOI22_X1 U15356 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15357 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15358 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15359 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15360 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12047) );
  NOR2_X1 U15361 ( .A1(n12048), .A2(n12047), .ZN(n12051) );
  AOI21_X1 U15362 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15177), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12049) );
  AOI21_X1 U15363 ( .B1(n12352), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12049), .ZN(
        n12050) );
  OAI21_X1 U15364 ( .B1(n12310), .B2(n12051), .A(n12050), .ZN(n12055) );
  XNOR2_X1 U15365 ( .A(n12067), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15179) );
  NAND2_X1 U15366 ( .A1(n15179), .A2(n14538), .ZN(n12054) );
  NAND2_X1 U15367 ( .A1(n12055), .A2(n12054), .ZN(n14772) );
  INV_X1 U15368 ( .A(n14772), .ZN(n12056) );
  AOI22_X1 U15369 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15370 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15371 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15372 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12057) );
  NAND4_X1 U15373 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n12057), .ZN(
        n12066) );
  AOI22_X1 U15374 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15375 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15376 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15377 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12061) );
  NAND4_X1 U15378 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12065) );
  NOR2_X1 U15379 ( .A1(n12066), .A2(n12065), .ZN(n12070) );
  AOI22_X1 U15380 ( .A1(n12352), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12351), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12069) );
  INV_X1 U15381 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14761) );
  XNOR2_X1 U15382 ( .A(n12084), .B(n14761), .ZN(n15164) );
  NAND2_X1 U15383 ( .A1(n15164), .A2(n14538), .ZN(n12068) );
  OAI211_X1 U15384 ( .C1(n12310), .C2(n12070), .A(n12069), .B(n12068), .ZN(
        n14755) );
  NAND2_X1 U15385 ( .A1(n12310), .A2(n12295), .ZN(n12270) );
  AOI22_X1 U15386 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15387 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15388 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15389 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12072) );
  AOI21_X1 U15390 ( .B1(n12325), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n14538), .ZN(n12071) );
  AND2_X1 U15391 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  NAND4_X1 U15392 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12082) );
  AOI22_X1 U15393 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15394 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15395 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15396 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15397 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12081) );
  OR2_X1 U15398 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  NAND2_X1 U15399 ( .A1(n12270), .A2(n12083), .ZN(n12088) );
  AOI22_X1 U15400 ( .A1(n12352), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11775), .ZN(n12087) );
  XNOR2_X1 U15401 ( .A(n12103), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14742) );
  AND2_X1 U15402 ( .A1(n14742), .A2(n14538), .ZN(n12086) );
  AOI21_X1 U15403 ( .B1(n12088), .B2(n12087), .A(n12086), .ZN(n14741) );
  AOI22_X1 U15404 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12334), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15405 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15406 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15407 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U15408 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12098) );
  AOI22_X1 U15409 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15410 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15411 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15412 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12093) );
  NAND4_X1 U15413 ( .A1(n12096), .A2(n12095), .A3(n12094), .A4(n12093), .ZN(
        n12097) );
  NOR2_X1 U15414 ( .A1(n12098), .A2(n12097), .ZN(n12102) );
  OAI21_X1 U15415 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21204), .A(
        n11775), .ZN(n12099) );
  INV_X1 U15416 ( .A(n12099), .ZN(n12100) );
  AOI21_X1 U15417 ( .B1(n12352), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12100), .ZN(
        n12101) );
  OAI21_X1 U15418 ( .B1(n12310), .B2(n12102), .A(n12101), .ZN(n12110) );
  INV_X1 U15419 ( .A(n12103), .ZN(n12104) );
  INV_X1 U15420 ( .A(n12105), .ZN(n12107) );
  INV_X1 U15421 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12106) );
  NAND2_X1 U15422 ( .A1(n12107), .A2(n12106), .ZN(n12108) );
  NAND2_X1 U15423 ( .A1(n12129), .A2(n12108), .ZN(n15142) );
  NAND2_X1 U15424 ( .A1(n12110), .A2(n12109), .ZN(n14728) );
  AOI22_X1 U15425 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15426 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15427 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15428 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U15429 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n12123) );
  AOI22_X1 U15430 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15431 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12120) );
  NAND2_X1 U15432 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12116) );
  AOI21_X1 U15433 ( .B1(n12325), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n14538), .ZN(n12115) );
  AND2_X1 U15434 ( .A1(n12116), .A2(n12115), .ZN(n12119) );
  AOI22_X1 U15435 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12118) );
  NAND4_X1 U15436 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12122) );
  OAI21_X1 U15437 ( .B1(n12123), .B2(n12122), .A(n12270), .ZN(n12125) );
  AOI22_X1 U15438 ( .A1(n12352), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11775), .ZN(n12124) );
  NAND2_X1 U15439 ( .A1(n12125), .A2(n12124), .ZN(n12127) );
  XNOR2_X1 U15440 ( .A(n12129), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15134) );
  NAND2_X1 U15441 ( .A1(n15134), .A2(n14538), .ZN(n12126) );
  NAND2_X1 U15442 ( .A1(n12127), .A2(n12126), .ZN(n14713) );
  INV_X1 U15443 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12130) );
  NAND2_X1 U15444 ( .A1(n12131), .A2(n12130), .ZN(n12132) );
  NAND2_X1 U15445 ( .A1(n12254), .A2(n12132), .ZN(n15124) );
  AOI22_X1 U15446 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15447 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15448 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15449 ( .A1(n12176), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12133) );
  NAND4_X1 U15450 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12142) );
  AOI22_X1 U15451 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15452 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15453 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15454 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12137) );
  NAND4_X1 U15455 ( .A1(n12140), .A2(n12139), .A3(n12138), .A4(n12137), .ZN(
        n12141) );
  NOR2_X1 U15456 ( .A1(n12142), .A2(n12141), .ZN(n12144) );
  AOI22_X1 U15457 ( .A1(n12352), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11775), .ZN(n12143) );
  OAI21_X1 U15458 ( .B1(n12310), .B2(n12144), .A(n12143), .ZN(n12145) );
  MUX2_X1 U15459 ( .A(n15124), .B(n12145), .S(n12295), .Z(n14700) );
  AOI22_X1 U15460 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15461 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15462 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15463 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12146) );
  NAND4_X1 U15464 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12155) );
  AOI22_X1 U15465 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15466 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15467 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15468 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15469 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12154) );
  NOR2_X1 U15470 ( .A1(n12155), .A2(n12154), .ZN(n12278) );
  AOI22_X1 U15471 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15472 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15473 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15474 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15475 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12165) );
  AOI22_X1 U15476 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15477 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15478 ( .A1(n12284), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15479 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15480 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12164) );
  NOR2_X1 U15481 ( .A1(n12165), .A2(n12164), .ZN(n12243) );
  AOI22_X1 U15482 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15483 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15484 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15485 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15486 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12175) );
  AOI22_X1 U15487 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15488 ( .A1(n12330), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15489 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15490 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U15491 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12174) );
  NOR2_X1 U15492 ( .A1(n12175), .A2(n12174), .ZN(n12231) );
  AOI22_X1 U15493 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n12017), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15494 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15495 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12176), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15496 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15497 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12186) );
  AOI22_X1 U15498 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12334), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15499 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12322), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15500 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12279), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15501 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12181) );
  NAND4_X1 U15502 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12185) );
  NOR2_X1 U15503 ( .A1(n12186), .A2(n12185), .ZN(n12232) );
  NOR2_X1 U15504 ( .A1(n12231), .A2(n12232), .ZN(n12225) );
  AOI22_X1 U15505 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15506 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15507 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15508 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15509 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12196) );
  AOI22_X1 U15510 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15511 ( .A1(n9623), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15512 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15513 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12191) );
  NAND4_X1 U15514 ( .A1(n12194), .A2(n12193), .A3(n12192), .A4(n12191), .ZN(
        n12195) );
  OR2_X1 U15515 ( .A1(n12196), .A2(n12195), .ZN(n12223) );
  NAND2_X1 U15516 ( .A1(n12225), .A2(n12223), .ZN(n12242) );
  NOR2_X1 U15517 ( .A1(n12243), .A2(n12242), .ZN(n12218) );
  AOI22_X1 U15518 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15519 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15520 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12263), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15521 ( .A1(n12335), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15522 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12207) );
  AOI22_X1 U15523 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15524 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15525 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15526 ( .A1(n12201), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15527 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12206) );
  OR2_X1 U15528 ( .A1(n12207), .A2(n12206), .ZN(n12217) );
  NAND2_X1 U15529 ( .A1(n12218), .A2(n12217), .ZN(n12277) );
  XNOR2_X1 U15530 ( .A(n12278), .B(n12277), .ZN(n12209) );
  AOI22_X1 U15531 ( .A1(n12352), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11775), .ZN(n12208) );
  OAI21_X1 U15532 ( .B1(n12209), .B2(n12310), .A(n12208), .ZN(n12216) );
  INV_X1 U15533 ( .A(n12213), .ZN(n12214) );
  INV_X1 U15534 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U15535 ( .A1(n12214), .A2(n14625), .ZN(n12215) );
  NAND2_X1 U15536 ( .A1(n12312), .A2(n12215), .ZN(n15073) );
  MUX2_X1 U15537 ( .A(n12216), .B(n15073), .S(n14538), .Z(n14623) );
  XNOR2_X1 U15538 ( .A(n12218), .B(n12217), .ZN(n12220) );
  AOI22_X1 U15539 ( .A1(n12352), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n11775), .ZN(n12219) );
  OAI21_X1 U15540 ( .B1(n12220), .B2(n12310), .A(n12219), .ZN(n12222) );
  INV_X1 U15541 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12221) );
  XNOR2_X1 U15542 ( .A(n12250), .B(n12221), .ZN(n15082) );
  MUX2_X1 U15543 ( .A(n12222), .B(n15082), .S(n14538), .Z(n14637) );
  INV_X1 U15544 ( .A(n14637), .ZN(n12253) );
  INV_X1 U15545 ( .A(n12223), .ZN(n12224) );
  XNOR2_X1 U15546 ( .A(n12225), .B(n12224), .ZN(n12229) );
  INV_X1 U15547 ( .A(n12310), .ZN(n12348) );
  INV_X1 U15548 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12227) );
  INV_X1 U15549 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12226) );
  OAI22_X1 U15550 ( .A1(n12346), .A2(n12227), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12226), .ZN(n12228) );
  AOI21_X1 U15551 ( .B1(n12229), .B2(n12348), .A(n12228), .ZN(n12230) );
  XNOR2_X1 U15552 ( .A(n12240), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15088) );
  MUX2_X1 U15553 ( .A(n12230), .B(n15088), .S(n14538), .Z(n14666) );
  XNOR2_X1 U15554 ( .A(n12232), .B(n12231), .ZN(n12234) );
  AOI22_X1 U15555 ( .A1(n12352), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n11775), .ZN(n12233) );
  OAI21_X1 U15556 ( .B1(n12234), .B2(n12310), .A(n12233), .ZN(n12235) );
  INV_X1 U15557 ( .A(n12235), .ZN(n12241) );
  INV_X1 U15558 ( .A(n12236), .ZN(n12238) );
  INV_X1 U15559 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15560 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  AND2_X1 U15561 ( .A1(n12240), .A2(n12239), .ZN(n15096) );
  MUX2_X1 U15562 ( .A(n12241), .B(n15096), .S(n14538), .Z(n12854) );
  XNOR2_X1 U15563 ( .A(n12243), .B(n12242), .ZN(n12245) );
  AOI22_X1 U15564 ( .A1(n12352), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11775), .ZN(n12244) );
  OAI21_X1 U15565 ( .B1(n12245), .B2(n12310), .A(n12244), .ZN(n12251) );
  INV_X1 U15566 ( .A(n12246), .ZN(n12248) );
  INV_X1 U15567 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12247) );
  NAND2_X1 U15568 ( .A1(n12248), .A2(n12247), .ZN(n12249) );
  NAND2_X1 U15569 ( .A1(n12250), .A2(n12249), .ZN(n14656) );
  MUX2_X1 U15570 ( .A(n12251), .B(n14656), .S(n14538), .Z(n12985) );
  INV_X1 U15571 ( .A(n12985), .ZN(n12252) );
  NOR2_X1 U15572 ( .A1(n12253), .A2(n12986), .ZN(n14621) );
  AND2_X1 U15573 ( .A1(n14623), .A2(n14621), .ZN(n12275) );
  XNOR2_X1 U15574 ( .A(n12254), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15106) );
  AOI22_X1 U15575 ( .A1(n12352), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11775), .ZN(n12274) );
  AOI22_X1 U15576 ( .A1(n9607), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15577 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15578 ( .A1(n12257), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12279), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15579 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15580 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12272) );
  AOI22_X1 U15581 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15582 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15583 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U15584 ( .A1(n12263), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12265) );
  AOI21_X1 U15585 ( .B1(n12325), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n14538), .ZN(n12264) );
  AND2_X1 U15586 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  NAND4_X1 U15587 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12271) );
  OAI21_X1 U15588 ( .B1(n12272), .B2(n12271), .A(n12270), .ZN(n12273) );
  INV_X1 U15589 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14614) );
  XNOR2_X1 U15590 ( .A(n12312), .B(n14614), .ZN(n15064) );
  NOR2_X1 U15591 ( .A1(n12278), .A2(n12277), .ZN(n12308) );
  AOI22_X1 U15592 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15593 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15594 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15595 ( .A1(n12279), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12280) );
  NAND4_X1 U15596 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12290) );
  AOI22_X1 U15597 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12288) );
  INV_X1 U15598 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U15599 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15600 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15601 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15602 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12289) );
  OR2_X1 U15603 ( .A1(n12290), .A2(n12289), .ZN(n12307) );
  XNOR2_X1 U15604 ( .A(n12308), .B(n12307), .ZN(n12293) );
  NAND2_X1 U15605 ( .A1(n12352), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12292) );
  OAI21_X1 U15606 ( .B1(n21204), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n11775), .ZN(n12291) );
  OAI211_X1 U15607 ( .C1(n12293), .C2(n12310), .A(n12292), .B(n12291), .ZN(
        n12294) );
  OAI21_X1 U15608 ( .B1(n15064), .B2(n12295), .A(n12294), .ZN(n14613) );
  AOI22_X1 U15609 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15610 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15611 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15612 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15613 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12306) );
  AOI22_X1 U15614 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9607), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15615 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11835), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15616 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15617 ( .A1(n12333), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U15618 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12305) );
  NOR2_X1 U15619 ( .A1(n12306), .A2(n12305), .ZN(n12320) );
  NAND2_X1 U15620 ( .A1(n12308), .A2(n12307), .ZN(n12319) );
  XNOR2_X1 U15621 ( .A(n12320), .B(n12319), .ZN(n12311) );
  AOI22_X1 U15622 ( .A1(n12352), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11775), .ZN(n12309) );
  OAI21_X1 U15623 ( .B1(n12311), .B2(n12310), .A(n12309), .ZN(n12318) );
  INV_X1 U15624 ( .A(n12312), .ZN(n12313) );
  INV_X1 U15625 ( .A(n12314), .ZN(n12316) );
  INV_X1 U15626 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15627 ( .A1(n12316), .A2(n12315), .ZN(n12317) );
  NAND2_X1 U15628 ( .A1(n14533), .A2(n12317), .ZN(n15049) );
  MUX2_X1 U15629 ( .A(n12318), .B(n15049), .S(n14538), .Z(n14595) );
  XNOR2_X1 U15630 ( .A(n14533), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14562) );
  NOR2_X1 U15631 ( .A1(n12320), .A2(n12319), .ZN(n12343) );
  AOI22_X1 U15632 ( .A1(n12322), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12321), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15633 ( .A1(n12324), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12323), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15634 ( .A1(n11625), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15635 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12284), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15636 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12341) );
  AOI22_X1 U15637 ( .A1(n12262), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15638 ( .A1(n12332), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12331), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15639 ( .A1(n12334), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12333), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15640 ( .A1(n11835), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12335), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15641 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12340) );
  NOR2_X1 U15642 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  XNOR2_X1 U15643 ( .A(n12343), .B(n12342), .ZN(n12349) );
  INV_X1 U15644 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12345) );
  OAI21_X1 U15645 ( .B1(n21204), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n11775), .ZN(n12344) );
  OAI21_X1 U15646 ( .B1(n12346), .B2(n12345), .A(n12344), .ZN(n12347) );
  AOI21_X1 U15647 ( .B1(n12349), .B2(n12348), .A(n12347), .ZN(n12350) );
  AOI21_X1 U15648 ( .B1(n14562), .B2(n14538), .A(n12350), .ZN(n13214) );
  NAND2_X1 U15649 ( .A1(n14597), .A2(n13214), .ZN(n12355) );
  AOI22_X1 U15650 ( .A1(n12352), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12351), .ZN(n12353) );
  INV_X1 U15651 ( .A(n12353), .ZN(n12354) );
  INV_X1 U15652 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12356) );
  AND2_X1 U15653 ( .A1(n12356), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12357) );
  NOR2_X1 U15654 ( .A1(n12370), .A2(n12357), .ZN(n12359) );
  NAND2_X1 U15655 ( .A1(n11659), .A2(n14304), .ZN(n12358) );
  NAND2_X1 U15656 ( .A1(n12358), .A2(n14546), .ZN(n12377) );
  XNOR2_X1 U15657 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12369) );
  XNOR2_X1 U15658 ( .A(n12369), .B(n12370), .ZN(n12412) );
  INV_X1 U15659 ( .A(n12412), .ZN(n12364) );
  NAND2_X1 U15660 ( .A1(n12405), .A2(n14542), .ZN(n12361) );
  NAND2_X1 U15661 ( .A1(n11659), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12362) );
  OAI211_X1 U15662 ( .C1(n12364), .C2(n12387), .A(n12361), .B(n12362), .ZN(
        n12365) );
  NAND2_X1 U15663 ( .A1(n12362), .A2(n14542), .ZN(n12363) );
  OAI22_X1 U15664 ( .A1(n12366), .A2(n12365), .B1(n12396), .B2(n12364), .ZN(
        n12368) );
  NAND2_X1 U15665 ( .A1(n12366), .A2(n12365), .ZN(n12367) );
  NAND2_X1 U15666 ( .A1(n12368), .A2(n12367), .ZN(n12376) );
  NAND2_X1 U15667 ( .A1(n12370), .A2(n12369), .ZN(n12372) );
  NAND2_X1 U15668 ( .A1(n14356), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12371) );
  NAND2_X1 U15669 ( .A1(n12372), .A2(n12371), .ZN(n12381) );
  XNOR2_X1 U15670 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12373) );
  XNOR2_X1 U15671 ( .A(n12381), .B(n12373), .ZN(n12414) );
  INV_X1 U15672 ( .A(n12414), .ZN(n12378) );
  NAND2_X1 U15673 ( .A1(n12405), .A2(n12378), .ZN(n12374) );
  OAI211_X1 U15674 ( .C1(n12378), .C2(n12387), .A(n12374), .B(n12377), .ZN(
        n12375) );
  NAND2_X1 U15675 ( .A1(n12376), .A2(n12375), .ZN(n12389) );
  INV_X1 U15676 ( .A(n12377), .ZN(n12379) );
  NAND3_X1 U15677 ( .A1(n12379), .A2(n12378), .A3(n12405), .ZN(n12388) );
  NOR2_X1 U15678 ( .A1(n14233), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12380) );
  NAND2_X1 U15679 ( .A1(n14233), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12382) );
  AND2_X1 U15680 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  OR2_X1 U15681 ( .A1(n12386), .A2(n12391), .ZN(n12413) );
  AOI22_X1 U15682 ( .A1(n12389), .A2(n12388), .B1(n12387), .B2(n12413), .ZN(
        n12395) );
  INV_X1 U15683 ( .A(n12413), .ZN(n12390) );
  NOR2_X1 U15684 ( .A1(n12402), .A2(n12390), .ZN(n12394) );
  NAND2_X1 U15685 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12401), .ZN(
        n12392) );
  INV_X1 U15686 ( .A(n12415), .ZN(n12393) );
  OAI22_X1 U15687 ( .A1(n12395), .A2(n12394), .B1(n12397), .B2(n12393), .ZN(
        n12400) );
  NAND2_X1 U15688 ( .A1(n21369), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12399) );
  NAND3_X1 U15689 ( .A1(n12415), .A2(n12397), .A3(n12396), .ZN(n12398) );
  AOI222_X1 U15690 ( .A1(n12401), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12401), .B2(n11850), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n11850), .ZN(n12416) );
  INV_X1 U15691 ( .A(n12402), .ZN(n12403) );
  NAND2_X1 U15692 ( .A1(n12416), .A2(n12403), .ZN(n12404) );
  NAND2_X1 U15693 ( .A1(n12416), .A2(n12405), .ZN(n12406) );
  NAND2_X1 U15694 ( .A1(n13842), .A2(n12855), .ZN(n12407) );
  NAND2_X1 U15695 ( .A1(n12408), .A2(n12407), .ZN(n12419) );
  NAND3_X1 U15696 ( .A1(n12737), .A2(n12526), .A3(n12411), .ZN(n12995) );
  INV_X1 U15697 ( .A(n9625), .ZN(n14872) );
  NOR4_X1 U15698 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12417) );
  NOR2_X1 U15699 ( .A1(n12417), .A2(n12416), .ZN(n13657) );
  NAND2_X1 U15700 ( .A1(n13657), .A2(n21389), .ZN(n12600) );
  OAI22_X1 U15701 ( .A1(n17532), .A2(n14218), .B1(n12600), .B2(n13849), .ZN(
        n13836) );
  AND2_X1 U15702 ( .A1(n15029), .A2(n14569), .ZN(n12421) );
  NAND2_X1 U15703 ( .A1(n15042), .A2(n12421), .ZN(n12438) );
  NOR4_X1 U15704 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12425) );
  NOR4_X1 U15705 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12424) );
  NOR4_X1 U15706 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12423) );
  NOR4_X1 U15707 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12422) );
  AND4_X1 U15708 ( .A1(n12425), .A2(n12424), .A3(n12423), .A4(n12422), .ZN(
        n12430) );
  NOR4_X1 U15709 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12428) );
  NOR4_X1 U15710 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12427) );
  NOR4_X1 U15711 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12426) );
  AND4_X1 U15712 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n21400), .ZN(
        n12429) );
  NAND2_X1 U15713 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  NOR3_X1 U15714 ( .A1(n15022), .A2(n14974), .A3(n12432), .ZN(n12433) );
  AOI22_X1 U15715 ( .A1(n15006), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15022), .ZN(n12434) );
  INV_X1 U15716 ( .A(n12434), .ZN(n12436) );
  NAND3_X1 U15717 ( .A1(n15029), .A2(n12605), .A3(n14974), .ZN(n14567) );
  INV_X1 U15718 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20286) );
  NOR2_X1 U15719 ( .A1(n14567), .A2(n20286), .ZN(n12435) );
  NOR2_X1 U15720 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  NAND2_X1 U15721 ( .A1(n12438), .A2(n12437), .ZN(P1_U2873) );
  INV_X1 U15722 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12953) );
  XOR2_X1 U15723 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12832), .Z(
        n15840) );
  INV_X1 U15724 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12440) );
  OAI21_X1 U15725 ( .B1(n17654), .B2(n12440), .A(n12439), .ZN(n12441) );
  AOI21_X1 U15726 ( .B1(n20209), .B2(n15840), .A(n12441), .ZN(n12442) );
  OAI21_X1 U15727 ( .B1(n13602), .B2(n20194), .A(n12442), .ZN(n12443) );
  OR2_X1 U15728 ( .A1(n12445), .A2(n16773), .ZN(n12446) );
  NAND3_X1 U15729 ( .A1(n12448), .A2(n12447), .A3(n12446), .ZN(P2_U2984) );
  OAI21_X1 U15730 ( .B1(n16614), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16604), .ZN(n12477) );
  INV_X1 U15731 ( .A(n12453), .ZN(n12455) );
  NAND2_X1 U15732 ( .A1(n16597), .A2(n16598), .ZN(n12456) );
  XNOR2_X1 U15733 ( .A(n16599), .B(n12456), .ZN(n12486) );
  NOR2_X1 U15734 ( .A1(n12459), .A2(n12460), .ZN(n12461) );
  OR2_X1 U15735 ( .A1(n12457), .A2(n12461), .ZN(n16361) );
  NOR2_X1 U15736 ( .A1(n16361), .A2(n20242), .ZN(n12473) );
  OR2_X1 U15737 ( .A1(n12463), .A2(n12464), .ZN(n12465) );
  NAND2_X1 U15738 ( .A1(n12462), .A2(n12465), .ZN(n16493) );
  INV_X1 U15739 ( .A(n12468), .ZN(n12466) );
  AND2_X1 U15740 ( .A1(n16999), .A2(n12466), .ZN(n12467) );
  OR2_X1 U15741 ( .A1(n16942), .A2(n12467), .ZN(n16903) );
  AND3_X1 U15742 ( .A1(n16937), .A2(n12468), .A3(n16615), .ZN(n16890) );
  OAI21_X1 U15743 ( .B1(n16903), .B2(n16890), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12471) );
  OR2_X1 U15744 ( .A1(n20207), .A2(n16000), .ZN(n12480) );
  AND3_X1 U15745 ( .A1(n16937), .A2(n12468), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16877) );
  NAND2_X1 U15746 ( .A1(n16877), .A2(n12469), .ZN(n12470) );
  NAND2_X1 U15747 ( .A1(n10458), .A2(n10460), .ZN(n12472) );
  OAI21_X1 U15748 ( .B1(n12486), .B2(n20241), .A(n12474), .ZN(n12475) );
  NAND2_X1 U15749 ( .A1(n10461), .A2(n12476), .ZN(P2_U3026) );
  INV_X1 U15750 ( .A(n16361), .ZN(n12484) );
  OAI21_X1 U15751 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12813), .A(
        n12478), .ZN(n15999) );
  INV_X1 U15752 ( .A(n15999), .ZN(n12479) );
  NAND2_X1 U15753 ( .A1(n20209), .A2(n12479), .ZN(n12481) );
  OAI211_X1 U15754 ( .C1(n17654), .C2(n12482), .A(n12481), .B(n12480), .ZN(
        n12483) );
  OAI21_X1 U15755 ( .B1(n12486), .B2(n20211), .A(n12485), .ZN(n12487) );
  NAND2_X1 U15756 ( .A1(n10485), .A2(n12488), .ZN(P2_U2994) );
  AOI222_X1 U15757 ( .A1(n12490), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12489), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11324), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12491) );
  INV_X1 U15758 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U15759 ( .A1(n20179), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n16527) );
  INV_X1 U15760 ( .A(n20219), .ZN(n12495) );
  NOR2_X1 U15761 ( .A1(n12497), .A2(n12496), .ZN(n12498) );
  OAI211_X1 U15762 ( .C1(n13196), .C2(n10221), .A(n12498), .B(n10218), .ZN(
        n12500) );
  INV_X1 U15763 ( .A(n12501), .ZN(n12502) );
  INV_X1 U15764 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12845) );
  NAND2_X1 U15765 ( .A1(n12502), .A2(n12845), .ZN(n12503) );
  MUX2_X1 U15766 ( .A(n11543), .B(n12503), .S(n20273), .Z(n15845) );
  XNOR2_X1 U15767 ( .A(n12504), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12505) );
  INV_X1 U15768 ( .A(n12562), .ZN(n13807) );
  INV_X1 U15769 ( .A(n15045), .ZN(n12596) );
  NAND2_X1 U15770 ( .A1(n12525), .A2(n12531), .ZN(n12541) );
  NAND2_X1 U15771 ( .A1(n12541), .A2(n12540), .ZN(n12519) );
  AND2_X1 U15772 ( .A1(n12518), .A2(n12520), .ZN(n12509) );
  NAND2_X1 U15773 ( .A1(n12519), .A2(n12509), .ZN(n12567) );
  XNOR2_X1 U15774 ( .A(n12567), .B(n12565), .ZN(n12510) );
  NAND2_X1 U15775 ( .A1(n12510), .A2(n14436), .ZN(n12511) );
  INV_X1 U15776 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17627) );
  NAND2_X1 U15777 ( .A1(n12512), .A2(n12562), .ZN(n12516) );
  INV_X1 U15778 ( .A(n12518), .ZN(n12513) );
  XNOR2_X1 U15779 ( .A(n12519), .B(n12513), .ZN(n12514) );
  NAND2_X1 U15780 ( .A1(n12514), .A2(n14436), .ZN(n12515) );
  NAND2_X1 U15781 ( .A1(n12517), .A2(n12562), .ZN(n12524) );
  NAND2_X1 U15782 ( .A1(n12519), .A2(n12518), .ZN(n12521) );
  XNOR2_X1 U15783 ( .A(n12521), .B(n12520), .ZN(n12522) );
  NAND2_X1 U15784 ( .A1(n12522), .A2(n14436), .ZN(n12523) );
  XNOR2_X1 U15785 ( .A(n12525), .B(n12531), .ZN(n12527) );
  INV_X1 U15786 ( .A(n14436), .ZN(n21470) );
  OAI211_X1 U15787 ( .C1(n12527), .C2(n21470), .A(n12526), .B(n14568), .ZN(
        n12528) );
  INV_X1 U15788 ( .A(n12528), .ZN(n12529) );
  NAND2_X1 U15789 ( .A1(n14541), .A2(n14299), .ZN(n12542) );
  OR2_X1 U15790 ( .A1(n21470), .A2(n12531), .ZN(n13805) );
  NAND3_X1 U15791 ( .A1(n12532), .A2(n12542), .A3(n13805), .ZN(n12535) );
  AND2_X1 U15792 ( .A1(n12542), .A2(n13807), .ZN(n12533) );
  INV_X1 U15793 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12748) );
  AOI21_X1 U15794 ( .B1(n12533), .B2(n13805), .A(n12748), .ZN(n12534) );
  XNOR2_X1 U15795 ( .A(n12537), .B(n13808), .ZN(n14110) );
  NAND2_X1 U15796 ( .A1(n14110), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14109) );
  INV_X1 U15797 ( .A(n13808), .ZN(n12536) );
  NAND2_X1 U15798 ( .A1(n12537), .A2(n12536), .ZN(n12538) );
  INV_X1 U15799 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21123) );
  NAND2_X1 U15800 ( .A1(n12539), .A2(n12562), .ZN(n12545) );
  XNOR2_X1 U15801 ( .A(n12541), .B(n12540), .ZN(n12543) );
  INV_X1 U15802 ( .A(n12542), .ZN(n13804) );
  AOI21_X1 U15803 ( .B1(n12543), .B2(n14436), .A(n13804), .ZN(n12544) );
  NAND2_X1 U15804 ( .A1(n12545), .A2(n12544), .ZN(n14194) );
  NAND2_X1 U15805 ( .A1(n14195), .A2(n14194), .ZN(n14193) );
  NAND2_X1 U15806 ( .A1(n12546), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12547) );
  NAND3_X1 U15807 ( .A1(n12548), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U15808 ( .A1(n12551), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U15809 ( .A1(n17583), .A2(n12552), .ZN(n17577) );
  NAND3_X1 U15810 ( .A1(n12554), .A2(n12562), .A3(n12553), .ZN(n12559) );
  INV_X1 U15811 ( .A(n12567), .ZN(n12555) );
  NAND2_X1 U15812 ( .A1(n12555), .A2(n12565), .ZN(n12556) );
  XNOR2_X1 U15813 ( .A(n12556), .B(n12564), .ZN(n12557) );
  NAND2_X1 U15814 ( .A1(n12557), .A2(n14436), .ZN(n12558) );
  OR2_X1 U15815 ( .A1(n17578), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12560) );
  NAND2_X1 U15816 ( .A1(n17578), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U15817 ( .A1(n12563), .A2(n12562), .ZN(n12570) );
  NAND2_X1 U15818 ( .A1(n12565), .A2(n12564), .ZN(n12566) );
  OR2_X1 U15819 ( .A1(n12567), .A2(n12566), .ZN(n12574) );
  XNOR2_X1 U15820 ( .A(n12574), .B(n12572), .ZN(n12568) );
  NAND2_X1 U15821 ( .A1(n12568), .A2(n14436), .ZN(n12569) );
  NAND2_X1 U15822 ( .A1(n12570), .A2(n12569), .ZN(n12571) );
  NAND2_X1 U15823 ( .A1(n12571), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17570) );
  NAND2_X1 U15824 ( .A1(n14436), .A2(n12572), .ZN(n12573) );
  NOR2_X1 U15825 ( .A1(n12574), .A2(n12573), .ZN(n15224) );
  NAND2_X1 U15826 ( .A1(n15224), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12576) );
  NOR2_X1 U15827 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12575) );
  AOI21_X1 U15828 ( .B1(n15245), .B2(n12576), .A(n12575), .ZN(n12581) );
  INV_X1 U15829 ( .A(n15224), .ZN(n12577) );
  INV_X1 U15830 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15255) );
  NAND2_X1 U15831 ( .A1(n12577), .A2(n15255), .ZN(n12578) );
  NAND2_X1 U15832 ( .A1(n12578), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12579) );
  NAND2_X1 U15833 ( .A1(n15245), .A2(n12579), .ZN(n12580) );
  INV_X1 U15834 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15159) );
  INV_X1 U15835 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15408) );
  INV_X1 U15836 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15395) );
  INV_X1 U15837 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15449) );
  INV_X1 U15838 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15435) );
  NAND3_X1 U15839 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12584) );
  INV_X1 U15840 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15427) );
  OR2_X1 U15841 ( .A1(n15245), .A2(n15427), .ZN(n12587) );
  NAND2_X1 U15842 ( .A1(n12586), .A2(n12587), .ZN(n12592) );
  NOR2_X1 U15843 ( .A1(n15227), .A2(n15408), .ZN(n15169) );
  INV_X1 U15844 ( .A(n15158), .ZN(n12590) );
  NAND2_X1 U15845 ( .A1(n15173), .A2(n15171), .ZN(n12589) );
  INV_X1 U15846 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15459) );
  INV_X1 U15847 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15478) );
  NAND2_X1 U15848 ( .A1(n15459), .A2(n15478), .ZN(n15202) );
  NOR2_X1 U15849 ( .A1(n15202), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12591) );
  NOR2_X1 U15850 ( .A1(n15227), .A2(n12591), .ZN(n15155) );
  AND2_X1 U15851 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12762) );
  INV_X1 U15852 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15120) );
  INV_X1 U15853 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15366) );
  INV_X1 U15854 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15361) );
  INV_X1 U15855 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15113) );
  INV_X1 U15856 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15323) );
  INV_X1 U15857 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15315) );
  INV_X1 U15858 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15086) );
  NAND3_X1 U15859 ( .A1(n15323), .A2(n15315), .A3(n15086), .ZN(n12594) );
  NOR2_X1 U15860 ( .A1(n12594), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15055) );
  INV_X1 U15861 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15060) );
  NAND2_X1 U15862 ( .A1(n15055), .A2(n15060), .ZN(n12593) );
  NOR2_X1 U15863 ( .A1(n15053), .A2(n12593), .ZN(n15034) );
  AND3_X1 U15864 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U15865 ( .A1(n12595), .A2(n15245), .ZN(n15084) );
  AND2_X1 U15866 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U15867 ( .A1(n15227), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15044) );
  INV_X1 U15868 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12597) );
  NOR2_X1 U15869 ( .A1(n12599), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n17543) );
  INV_X1 U15870 ( .A(n17543), .ZN(n14545) );
  NAND2_X1 U15871 ( .A1(n14542), .A2(n14545), .ZN(n12602) );
  INV_X1 U15872 ( .A(n12600), .ZN(n12601) );
  NAND2_X1 U15873 ( .A1(n12602), .A2(n12601), .ZN(n12611) );
  NAND2_X1 U15874 ( .A1(n12603), .A2(n21389), .ZN(n12604) );
  NAND2_X1 U15875 ( .A1(n12604), .A2(n14304), .ZN(n12607) );
  NAND2_X1 U15876 ( .A1(n14436), .A2(n14545), .ZN(n12606) );
  AOI21_X1 U15877 ( .B1(n12607), .B2(n12606), .A(n12605), .ZN(n12608) );
  MUX2_X1 U15878 ( .A(n12611), .B(n12610), .S(n12609), .Z(n12620) );
  NAND2_X1 U15879 ( .A1(n12612), .A2(n14542), .ZN(n12744) );
  INV_X1 U15880 ( .A(n12744), .ZN(n12618) );
  NAND3_X1 U15881 ( .A1(n12615), .A2(n14304), .A3(n12744), .ZN(n12736) );
  INV_X1 U15882 ( .A(n12736), .ZN(n12616) );
  NOR2_X1 U15883 ( .A1(n12995), .A2(n12616), .ZN(n12617) );
  NOR2_X1 U15884 ( .A1(n12614), .A2(n12617), .ZN(n13834) );
  AOI21_X1 U15885 ( .B1(n17532), .B2(n12618), .A(n13834), .ZN(n12619) );
  NOR2_X1 U15886 ( .A1(n12621), .A2(n9625), .ZN(n12622) );
  OR2_X1 U15887 ( .A1(n12995), .A2(n12622), .ZN(n13653) );
  NOR2_X1 U15888 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  NAND2_X1 U15889 ( .A1(n12714), .A2(n14899), .ZN(n12629) );
  NAND2_X1 U15890 ( .A1(n12626), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12627) );
  OAI211_X1 U15891 ( .C1(n14579), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12637), .B(
        n12627), .ZN(n12628) );
  NAND2_X1 U15892 ( .A1(n12629), .A2(n12628), .ZN(n12633) );
  INV_X1 U15893 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12630) );
  OR2_X1 U15894 ( .A1(n12637), .A2(n12630), .ZN(n12632) );
  NAND2_X1 U15895 ( .A1(n10323), .A2(n12630), .ZN(n12631) );
  NAND2_X1 U15896 ( .A1(n12632), .A2(n12631), .ZN(n13811) );
  XNOR2_X1 U15897 ( .A(n12633), .B(n13811), .ZN(n14907) );
  NAND2_X1 U15898 ( .A1(n14907), .A2(n13829), .ZN(n12635) );
  INV_X1 U15899 ( .A(n12633), .ZN(n12634) );
  NAND2_X1 U15900 ( .A1(n12635), .A2(n12634), .ZN(n14209) );
  MUX2_X1 U15901 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n12636) );
  OAI21_X1 U15902 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14580), .A(
        n12636), .ZN(n14208) );
  INV_X1 U15903 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21007) );
  NAND2_X1 U15904 ( .A1(n12714), .A2(n21007), .ZN(n12640) );
  NAND2_X1 U15905 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12638) );
  OAI211_X1 U15906 ( .C1(n14579), .C2(P1_EBX_REG_4__SCAN_IN), .A(n12682), .B(
        n12638), .ZN(n12639) );
  AND2_X1 U15907 ( .A1(n12640), .A2(n12639), .ZN(n14430) );
  INV_X1 U15908 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14257) );
  NAND2_X1 U15909 ( .A1(n9610), .A2(n14257), .ZN(n12645) );
  INV_X2 U15910 ( .A(n10323), .ZN(n14576) );
  NAND2_X1 U15911 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U15912 ( .A1(n12682), .A2(n12642), .ZN(n12643) );
  OAI21_X1 U15913 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n14579), .A(n12643), .ZN(
        n12644) );
  NAND2_X1 U15914 ( .A1(n12645), .A2(n12644), .ZN(n14431) );
  NAND2_X1 U15915 ( .A1(n14430), .A2(n14431), .ZN(n12646) );
  NAND2_X1 U15916 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12647) );
  NAND2_X1 U15917 ( .A1(n12682), .A2(n12647), .ZN(n12648) );
  OAI21_X1 U15918 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14579), .A(n12648), .ZN(
        n12649) );
  OAI21_X1 U15919 ( .B1(n12720), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12649), .ZN(
        n14486) );
  AND2_X2 U15920 ( .A1(n14487), .A2(n14486), .ZN(n17612) );
  INV_X1 U15921 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21034) );
  NAND2_X1 U15922 ( .A1(n12714), .A2(n21034), .ZN(n12652) );
  NAND2_X1 U15923 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12650) );
  OAI211_X1 U15924 ( .C1(n14579), .C2(P1_EBX_REG_6__SCAN_IN), .A(n12682), .B(
        n12650), .ZN(n12651) );
  AND2_X1 U15925 ( .A1(n12652), .A2(n12651), .ZN(n17611) );
  INV_X1 U15926 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12653) );
  NAND2_X1 U15927 ( .A1(n12714), .A2(n12653), .ZN(n12656) );
  NAND2_X1 U15928 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12654) );
  OAI211_X1 U15929 ( .C1(n14579), .C2(P1_EBX_REG_8__SCAN_IN), .A(n12682), .B(
        n12654), .ZN(n12655) );
  AND2_X1 U15930 ( .A1(n12656), .A2(n12655), .ZN(n14861) );
  INV_X1 U15931 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20964) );
  NAND2_X1 U15932 ( .A1(n9610), .A2(n20964), .ZN(n12660) );
  NAND2_X1 U15933 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12657) );
  NAND2_X1 U15934 ( .A1(n12682), .A2(n12657), .ZN(n12658) );
  OAI21_X1 U15935 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n14579), .A(n12658), .ZN(
        n12659) );
  NAND2_X1 U15936 ( .A1(n12660), .A2(n12659), .ZN(n14862) );
  INV_X1 U15937 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20954) );
  NAND2_X1 U15938 ( .A1(n9610), .A2(n20954), .ZN(n12664) );
  NAND2_X1 U15939 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12661) );
  NAND2_X1 U15940 ( .A1(n12682), .A2(n12661), .ZN(n12662) );
  OAI21_X1 U15941 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14579), .A(n12662), .ZN(
        n12663) );
  MUX2_X1 U15942 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12665) );
  INV_X1 U15943 ( .A(n12665), .ZN(n12667) );
  NOR2_X1 U15944 ( .A1(n14580), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12666) );
  NOR2_X1 U15945 ( .A1(n12667), .A2(n12666), .ZN(n14851) );
  NAND2_X1 U15946 ( .A1(n14957), .A2(n14851), .ZN(n14948) );
  INV_X1 U15947 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14953) );
  NAND2_X1 U15948 ( .A1(n9610), .A2(n14953), .ZN(n12671) );
  NAND2_X1 U15949 ( .A1(n12682), .A2(n15459), .ZN(n12669) );
  NAND2_X1 U15950 ( .A1(n13829), .A2(n14953), .ZN(n12668) );
  NAND3_X1 U15951 ( .A1(n12669), .A2(n14576), .A3(n12668), .ZN(n12670) );
  NAND2_X1 U15952 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12673) );
  OAI211_X1 U15953 ( .C1(n14579), .C2(P1_EBX_REG_12__SCAN_IN), .A(n12682), .B(
        n12673), .ZN(n12674) );
  OAI21_X1 U15954 ( .B1(n12711), .B2(P1_EBX_REG_12__SCAN_IN), .A(n12674), .ZN(
        n14837) );
  INV_X1 U15955 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14814) );
  NAND2_X1 U15956 ( .A1(n9610), .A2(n14814), .ZN(n12678) );
  NAND2_X1 U15957 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12675) );
  NAND2_X1 U15958 ( .A1(n12682), .A2(n12675), .ZN(n12676) );
  OAI21_X1 U15959 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(n14579), .A(n12676), .ZN(
        n12677) );
  MUX2_X1 U15960 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12679) );
  INV_X1 U15961 ( .A(n12679), .ZN(n12681) );
  NOR2_X1 U15962 ( .A1(n14580), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12680) );
  NOR2_X1 U15963 ( .A1(n12681), .A2(n12680), .ZN(n14939) );
  NAND2_X1 U15964 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  INV_X1 U15965 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14934) );
  NAND2_X1 U15966 ( .A1(n9610), .A2(n14934), .ZN(n12685) );
  NAND2_X1 U15967 ( .A1(n12682), .A2(n15408), .ZN(n12683) );
  OAI211_X1 U15968 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n14579), .A(n12683), .B(
        n14576), .ZN(n12684) );
  NOR2_X2 U15969 ( .A1(n14941), .A2(n14800), .ZN(n14773) );
  MUX2_X1 U15970 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12686) );
  OAI21_X1 U15971 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14580), .A(
        n12686), .ZN(n14774) );
  INV_X1 U15972 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U15973 ( .A1(n9610), .A2(n12688), .ZN(n12691) );
  NAND2_X1 U15974 ( .A1(n12682), .A2(n15395), .ZN(n12689) );
  OAI211_X1 U15975 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n14579), .A(n12689), .B(
        n14576), .ZN(n12690) );
  MUX2_X1 U15976 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12692) );
  OAI21_X1 U15977 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14580), .A(
        n12692), .ZN(n14752) );
  NOR2_X1 U15978 ( .A1(n14767), .A2(n14752), .ZN(n12693) );
  NAND2_X1 U15979 ( .A1(n12682), .A2(n15361), .ZN(n12694) );
  OAI211_X1 U15980 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n14579), .A(n12694), .B(
        n14576), .ZN(n12695) );
  OAI21_X1 U15981 ( .B1(n12720), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12695), .ZN(
        n14726) );
  NAND2_X1 U15982 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12696) );
  OAI211_X1 U15983 ( .C1(n14579), .C2(P1_EBX_REG_20__SCAN_IN), .A(n12682), .B(
        n12696), .ZN(n12697) );
  OAI21_X1 U15984 ( .B1(n12711), .B2(P1_EBX_REG_20__SCAN_IN), .A(n12697), .ZN(
        n14714) );
  INV_X1 U15985 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U15986 ( .A1(n9610), .A2(n14706), .ZN(n12700) );
  NAND2_X1 U15987 ( .A1(n12682), .A2(n15120), .ZN(n12698) );
  OAI211_X1 U15988 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n14579), .A(n12698), .B(
        n14576), .ZN(n12699) );
  NOR2_X2 U15989 ( .A1(n14716), .A2(n14709), .ZN(n14696) );
  MUX2_X1 U15990 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12701) );
  OAI21_X1 U15991 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14580), .A(
        n12701), .ZN(n12702) );
  INV_X1 U15992 ( .A(n12702), .ZN(n14695) );
  NAND2_X1 U15993 ( .A1(n12682), .A2(n15323), .ZN(n12703) );
  OAI211_X1 U15994 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n14579), .A(n12703), .B(
        n14576), .ZN(n12704) );
  OAI21_X1 U15995 ( .B1(n12720), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12704), .ZN(
        n12861) );
  MUX2_X1 U15996 ( .A(n12711), .B(n14576), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12705) );
  OAI21_X1 U15997 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14580), .A(
        n12705), .ZN(n14676) );
  INV_X1 U15998 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U15999 ( .A1(n9610), .A2(n14925), .ZN(n12708) );
  NAND2_X1 U16000 ( .A1(n12682), .A2(n15315), .ZN(n12706) );
  OAI211_X1 U16001 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14579), .A(n12706), .B(
        n14576), .ZN(n12707) );
  NAND2_X1 U16002 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12709) );
  OAI211_X1 U16003 ( .C1(n14579), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12682), .B(
        n12709), .ZN(n12710) );
  OAI21_X1 U16004 ( .B1(n12711), .B2(P1_EBX_REG_26__SCAN_IN), .A(n12710), .ZN(
        n14638) );
  INV_X1 U16005 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U16006 ( .A1(n12682), .A2(n15297), .ZN(n12712) );
  OAI211_X1 U16007 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14579), .A(n12712), .B(
        n14576), .ZN(n12713) );
  OAI21_X1 U16008 ( .B1(n12720), .B2(P1_EBX_REG_27__SCAN_IN), .A(n12713), .ZN(
        n14629) );
  INV_X1 U16009 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U16010 ( .A1(n12714), .A2(n14921), .ZN(n12717) );
  NAND2_X1 U16011 ( .A1(n14576), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12715) );
  OAI211_X1 U16012 ( .C1(n14579), .C2(P1_EBX_REG_28__SCAN_IN), .A(n12682), .B(
        n12715), .ZN(n12716) );
  AND2_X1 U16013 ( .A1(n12717), .A2(n12716), .ZN(n14609) );
  OR2_X1 U16014 ( .A1(n14580), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12719) );
  INV_X1 U16015 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14920) );
  NAND2_X1 U16016 ( .A1(n13829), .A2(n14920), .ZN(n12718) );
  NAND2_X1 U16017 ( .A1(n12719), .A2(n12718), .ZN(n12721) );
  OAI22_X1 U16018 ( .A1(n12721), .A2(n10323), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12720), .ZN(n14594) );
  NAND2_X1 U16019 ( .A1(n14611), .A2(n14594), .ZN(n14593) );
  NAND2_X1 U16020 ( .A1(n14593), .A2(n10323), .ZN(n12724) );
  INV_X1 U16021 ( .A(n12721), .ZN(n12722) );
  NAND2_X1 U16022 ( .A1(n14611), .A2(n12722), .ZN(n12723) );
  NAND2_X1 U16023 ( .A1(n12724), .A2(n12723), .ZN(n12725) );
  AOI22_X1 U16024 ( .A1(n14580), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14579), .ZN(n14581) );
  INV_X1 U16025 ( .A(n12749), .ZN(n12729) );
  NAND2_X1 U16026 ( .A1(n12603), .A2(n14436), .ZN(n12726) );
  OAI21_X1 U16027 ( .B1(n12727), .B2(n14294), .A(n12726), .ZN(n12728) );
  NAND2_X1 U16028 ( .A1(n12614), .A2(n14542), .ZN(n15501) );
  INV_X1 U16029 ( .A(n14885), .ZN(n12733) );
  INV_X1 U16030 ( .A(n12731), .ZN(n12732) );
  AND3_X1 U16031 ( .A1(n12736), .A2(n12735), .A3(n12734), .ZN(n12740) );
  NAND2_X1 U16032 ( .A1(n12737), .A2(n14222), .ZN(n12738) );
  NAND2_X1 U16033 ( .A1(n12738), .A2(n14542), .ZN(n12739) );
  OAI211_X1 U16034 ( .C1(n11680), .C2(n14872), .A(n12740), .B(n12739), .ZN(
        n13847) );
  OAI21_X1 U16035 ( .B1(n13843), .B2(n14304), .A(n12741), .ZN(n12742) );
  NOR2_X1 U16036 ( .A1(n13847), .A2(n12742), .ZN(n12743) );
  INV_X1 U16037 ( .A(n14220), .ZN(n12745) );
  NAND2_X1 U16038 ( .A1(n21130), .A2(n17600), .ZN(n21148) );
  INV_X1 U16039 ( .A(n12766), .ZN(n12757) );
  INV_X1 U16040 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15491) );
  INV_X1 U16041 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17619) );
  INV_X1 U16042 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12747) );
  INV_X1 U16043 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12746) );
  NOR2_X1 U16044 ( .A1(n12747), .A2(n12746), .ZN(n21112) );
  NAND2_X1 U16045 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21112), .ZN(
        n17614) );
  NOR2_X1 U16046 ( .A1(n17619), .A2(n17614), .ZN(n17593) );
  NAND3_X1 U16047 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n17593), .ZN(n12750) );
  NAND2_X1 U16048 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15467) );
  OR4_X1 U16049 ( .A1(n15478), .A2(n15491), .A3(n12750), .A4(n15467), .ZN(
        n15448) );
  NOR3_X1 U16050 ( .A1(n15449), .A2(n15459), .A3(n15448), .ZN(n15442) );
  NOR4_X1 U16051 ( .A1(n15427), .A2(n15408), .A3(n15159), .A4(n15395), .ZN(
        n15387) );
  INV_X1 U16052 ( .A(n15387), .ZN(n15388) );
  NOR2_X1 U16053 ( .A1(n15113), .A2(n15388), .ZN(n12760) );
  AND2_X1 U16054 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12760), .ZN(
        n15343) );
  AND2_X1 U16055 ( .A1(n15442), .A2(n15343), .ZN(n15344) );
  OR2_X2 U16056 ( .A1(n12996), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15176) );
  AOI21_X1 U16057 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17597) );
  NOR2_X1 U16058 ( .A1(n12750), .A2(n17597), .ZN(n15484) );
  NAND2_X1 U16059 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15193) );
  NOR2_X1 U16060 ( .A1(n15193), .A2(n15491), .ZN(n12751) );
  AND2_X1 U16061 ( .A1(n15484), .A2(n12751), .ZN(n15450) );
  AND2_X1 U16062 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12752) );
  AND2_X1 U16063 ( .A1(n15450), .A2(n12752), .ZN(n15424) );
  NAND2_X1 U16064 ( .A1(n15424), .A2(n12760), .ZN(n12753) );
  NAND2_X1 U16065 ( .A1(n21127), .A2(n12753), .ZN(n12754) );
  OAI211_X1 U16066 ( .C1(n21130), .C2(n15344), .A(n21129), .B(n12754), .ZN(
        n15376) );
  INV_X1 U16067 ( .A(n12762), .ZN(n15353) );
  OR2_X1 U16068 ( .A1(n21148), .A2(n9895), .ZN(n15471) );
  NAND2_X1 U16069 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U16070 ( .A1(n21148), .A2(n12759), .ZN(n12755) );
  NOR2_X1 U16071 ( .A1(n15334), .A2(n21148), .ZN(n12756) );
  INV_X1 U16072 ( .A(n12756), .ZN(n15266) );
  OAI21_X1 U16073 ( .B1(n15303), .B2(n17601), .A(n15321), .ZN(n15312) );
  INV_X1 U16074 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12764) );
  NOR2_X1 U16075 ( .A1(n15312), .A2(n12764), .ZN(n15305) );
  NOR2_X1 U16076 ( .A1(n15305), .A2(n12756), .ZN(n15293) );
  AOI21_X1 U16077 ( .B1(n12757), .B2(n15266), .A(n15293), .ZN(n15278) );
  OAI211_X1 U16078 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n17601), .A(
        n15278), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15267) );
  INV_X1 U16079 ( .A(n15267), .ZN(n12768) );
  NAND2_X1 U16080 ( .A1(n12748), .A2(n15434), .ZN(n21147) );
  NAND2_X1 U16081 ( .A1(n15468), .A2(n21147), .ZN(n21134) );
  NAND2_X1 U16082 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15442), .ZN(
        n15383) );
  OR2_X1 U16083 ( .A1(n21134), .A2(n15383), .ZN(n15322) );
  NAND2_X1 U16084 ( .A1(n21127), .A2(n15424), .ZN(n12758) );
  NAND2_X1 U16085 ( .A1(n15322), .A2(n12758), .ZN(n15410) );
  INV_X1 U16086 ( .A(n12759), .ZN(n12761) );
  AND3_X1 U16087 ( .A1(n12762), .A2(n12761), .A3(n12760), .ZN(n12763) );
  NAND2_X1 U16088 ( .A1(n15410), .A2(n12763), .ZN(n15331) );
  INV_X1 U16089 ( .A(n15303), .ZN(n12765) );
  NOR3_X1 U16090 ( .A1(n15331), .A2(n12765), .A3(n12764), .ZN(n15295) );
  NAND2_X1 U16091 ( .A1(n15295), .A2(n12766), .ZN(n15270) );
  INV_X1 U16092 ( .A(n15270), .ZN(n15275) );
  AOI21_X1 U16093 ( .B1(n15275), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U16094 ( .A1(n21133), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13215) );
  OAI21_X1 U16095 ( .B1(n12768), .B2(n12767), .A(n13215), .ZN(n12769) );
  AOI21_X1 U16096 ( .B1(n14573), .B2(n21142), .A(n12769), .ZN(n12770) );
  OAI21_X1 U16097 ( .B1(n13222), .B2(n15482), .A(n12770), .ZN(P1_U3001) );
  NAND2_X1 U16098 ( .A1(n20917), .A2(n20050), .ZN(n12839) );
  INV_X1 U16099 ( .A(n12839), .ZN(n12771) );
  NAND2_X1 U16100 ( .A1(n12775), .A2(n12771), .ZN(n12772) );
  NOR2_X2 U16101 ( .A1(n20908), .A2(n12772), .ZN(n16301) );
  INV_X1 U16102 ( .A(n20908), .ZN(n13620) );
  NAND2_X1 U16103 ( .A1(n13640), .A2(n20050), .ZN(n15838) );
  INV_X1 U16104 ( .A(n15838), .ZN(n12773) );
  AND2_X1 U16105 ( .A1(n12774), .A2(n12773), .ZN(n17287) );
  NAND3_X1 U16106 ( .A1(n12775), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12839), 
        .ZN(n12776) );
  NAND2_X1 U16107 ( .A1(n12832), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12778) );
  INV_X1 U16108 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12777) );
  AND2_X1 U16109 ( .A1(n12816), .A2(n16576), .ZN(n12780) );
  AND2_X1 U16110 ( .A1(n12784), .A2(n12781), .ZN(n12782) );
  OR2_X1 U16111 ( .A1(n12782), .A2(n9633), .ZN(n16625) );
  NAND2_X1 U16112 ( .A1(n12811), .A2(n16635), .ZN(n12783) );
  AND2_X1 U16113 ( .A1(n12784), .A2(n12783), .ZN(n16638) );
  INV_X1 U16114 ( .A(n12807), .ZN(n12786) );
  NAND2_X1 U16115 ( .A1(n12806), .A2(n16093), .ZN(n12785) );
  NAND2_X1 U16116 ( .A1(n12786), .A2(n12785), .ZN(n16664) );
  OR2_X1 U16117 ( .A1(n12789), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12787) );
  NAND2_X1 U16118 ( .A1(n12804), .A2(n12787), .ZN(n16687) );
  AND2_X1 U16119 ( .A1(n12792), .A2(n16707), .ZN(n12788) );
  NOR2_X1 U16120 ( .A1(n12789), .A2(n12788), .ZN(n16709) );
  NAND2_X1 U16121 ( .A1(n12794), .A2(n12790), .ZN(n12791) );
  NAND2_X1 U16122 ( .A1(n12792), .A2(n12791), .ZN(n16724) );
  NAND2_X1 U16123 ( .A1(n12796), .A2(n16733), .ZN(n12793) );
  AND2_X1 U16124 ( .A1(n12794), .A2(n12793), .ZN(n16735) );
  OR2_X1 U16125 ( .A1(n12797), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12795) );
  NAND2_X1 U16126 ( .A1(n12796), .A2(n12795), .ZN(n16745) );
  AOI21_X1 U16127 ( .B1(n16760), .B2(n12801), .A(n12797), .ZN(n16762) );
  AOI21_X1 U16128 ( .B1(n17644), .B2(n12799), .A(n12802), .ZN(n17638) );
  AOI21_X1 U16129 ( .B1(n17655), .B2(n12798), .A(n12800), .ZN(n17645) );
  OAI21_X1 U16130 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12798), .ZN(n20200) );
  MUX2_X1 U16131 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16289) );
  INV_X1 U16132 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20208) );
  MUX2_X1 U16133 ( .A(n20208), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n16269) );
  NOR2_X1 U16134 ( .A1(n16289), .A2(n16269), .ZN(n16271) );
  NAND2_X1 U16135 ( .A1(n20200), .A2(n16271), .ZN(n16251) );
  NOR2_X1 U16136 ( .A1(n17645), .A2(n16251), .ZN(n16232) );
  OAI21_X1 U16137 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12800), .A(
        n12799), .ZN(n20185) );
  NAND2_X1 U16138 ( .A1(n16232), .A2(n20185), .ZN(n16208) );
  OAI21_X1 U16139 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12802), .A(
        n12801), .ZN(n20081) );
  NOR2_X1 U16140 ( .A1(n16735), .A2(n16167), .ZN(n16152) );
  NAND2_X1 U16141 ( .A1(n16724), .A2(n16152), .ZN(n16136) );
  NAND2_X1 U16142 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  NAND2_X1 U16143 ( .A1(n12806), .A2(n12805), .ZN(n16678) );
  NOR2_X1 U16144 ( .A1(n12807), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12808) );
  OR2_X1 U16145 ( .A1(n12809), .A2(n12808), .ZN(n16654) );
  AND2_X1 U16146 ( .A1(n16077), .A2(n16654), .ZN(n16065) );
  OR2_X1 U16147 ( .A1(n12809), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12810) );
  NAND2_X1 U16148 ( .A1(n12811), .A2(n12810), .ZN(n16645) );
  NOR2_X1 U16149 ( .A1(n9633), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12812) );
  OR2_X1 U16150 ( .A1(n12813), .A2(n12812), .ZN(n16617) );
  AND2_X1 U16151 ( .A1(n16017), .A2(n16617), .ZN(n16005) );
  INV_X1 U16152 ( .A(n12820), .ZN(n12815) );
  INV_X1 U16153 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U16154 ( .A1(n12815), .A2(n12814), .ZN(n12817) );
  AND2_X1 U16155 ( .A1(n12817), .A2(n12816), .ZN(n16590) );
  NOR2_X1 U16156 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12818), .ZN(
        n12819) );
  NOR2_X1 U16157 ( .A1(n12820), .A2(n12819), .ZN(n16607) );
  OR2_X1 U16158 ( .A1(n16590), .A2(n16607), .ZN(n15951) );
  OR2_X1 U16159 ( .A1(n9680), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12821) );
  NAND2_X1 U16160 ( .A1(n12822), .A2(n12821), .ZN(n15941) );
  NAND2_X1 U16161 ( .A1(n15936), .A2(n15941), .ZN(n15918) );
  NAND2_X1 U16162 ( .A1(n12822), .A2(n16557), .ZN(n12823) );
  AND2_X1 U16163 ( .A1(n12824), .A2(n12823), .ZN(n16560) );
  INV_X1 U16164 ( .A(n12828), .ZN(n12827) );
  NAND2_X1 U16165 ( .A1(n12825), .A2(n12953), .ZN(n12826) );
  NAND2_X1 U16166 ( .A1(n12827), .A2(n12826), .ZN(n16549) );
  NOR2_X1 U16167 ( .A1(n12828), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12829) );
  OR2_X1 U16168 ( .A1(n12830), .A2(n12829), .ZN(n13208) );
  INV_X1 U16169 ( .A(n13208), .ZN(n15873) );
  NOR2_X1 U16170 ( .A1(n12830), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12831) );
  OR2_X1 U16171 ( .A1(n12832), .A2(n12831), .ZN(n16538) );
  AOI21_X1 U16172 ( .B1(n15855), .B2(n16538), .A(n20080), .ZN(n15841) );
  XNOR2_X1 U16173 ( .A(n15841), .B(n15840), .ZN(n12848) );
  NAND2_X1 U16174 ( .A1(n20912), .A2(n20559), .ZN(n12833) );
  NOR2_X1 U16175 ( .A1(n11308), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20463) );
  INV_X1 U16176 ( .A(n20463), .ZN(n12835) );
  NOR2_X1 U16177 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n12835), .ZN(n12836) );
  NAND2_X1 U16178 ( .A1(n12836), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17665) );
  AND3_X1 U16179 ( .A1(n20207), .A2(n16274), .A3(n17665), .ZN(n12837) );
  NAND2_X2 U16180 ( .A1(n20908), .A2(n12837), .ZN(n16262) );
  INV_X1 U16181 ( .A(n13611), .ZN(n17272) );
  NAND2_X1 U16182 ( .A1(n13791), .A2(n15838), .ZN(n12843) );
  INV_X1 U16183 ( .A(n13668), .ZN(n12841) );
  INV_X1 U16184 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12840) );
  NAND3_X1 U16185 ( .A1(n12841), .A2(n12840), .A3(n12839), .ZN(n12842) );
  OAI22_X1 U16186 ( .A1(n20072), .A2(n12845), .B1(n12844), .B2(n16262), .ZN(
        n12846) );
  AOI21_X1 U16187 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16275), .A(
        n12846), .ZN(n12847) );
  OAI21_X1 U16188 ( .B1(n12848), .B2(n16274), .A(n12847), .ZN(n12849) );
  NAND2_X1 U16189 ( .A1(n10483), .A2(n12853), .ZN(P2_U2825) );
  NAND2_X1 U16190 ( .A1(n17532), .A2(n14220), .ZN(n12858) );
  NAND3_X1 U16191 ( .A1(n12856), .A2(n13829), .A3(n12855), .ZN(n12857) );
  NAND2_X1 U16192 ( .A1(n12858), .A2(n12857), .ZN(n12859) );
  INV_X1 U16193 ( .A(n14963), .ZN(n21031) );
  OAI21_X1 U16194 ( .B1(n12860), .B2(n12861), .A(n14675), .ZN(n12862) );
  INV_X1 U16195 ( .A(n12862), .ZN(n15335) );
  INV_X1 U16196 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n21046) );
  INV_X1 U16197 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U16198 ( .A1(n21046), .A2(keyinput10), .B1(keyinput28), .B2(n19983), 
        .ZN(n12865) );
  OAI221_X1 U16199 ( .B1(n21046), .B2(keyinput10), .C1(n19983), .C2(keyinput28), .A(n12865), .ZN(n12872) );
  INV_X1 U16200 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21375) );
  AOI22_X1 U16201 ( .A1(n21375), .A2(keyinput53), .B1(n21043), .B2(keyinput51), 
        .ZN(n12866) );
  OAI221_X1 U16202 ( .B1(n21375), .B2(keyinput53), .C1(n21043), .C2(keyinput51), .A(n12866), .ZN(n12871) );
  INV_X1 U16203 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20035) );
  INV_X1 U16204 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18466) );
  AOI22_X1 U16205 ( .A1(n20035), .A2(keyinput27), .B1(keyinput26), .B2(n18466), 
        .ZN(n12867) );
  OAI221_X1 U16206 ( .B1(n20035), .B2(keyinput27), .C1(n18466), .C2(keyinput26), .A(n12867), .ZN(n12870) );
  INV_X1 U16207 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18869) );
  AOI22_X1 U16208 ( .A1(n19918), .A2(keyinput52), .B1(keyinput18), .B2(n18869), 
        .ZN(n12868) );
  OAI221_X1 U16209 ( .B1(n19918), .B2(keyinput52), .C1(n18869), .C2(keyinput18), .A(n12868), .ZN(n12869) );
  NOR4_X1 U16210 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n12869), .ZN(
        n12946) );
  INV_X1 U16211 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12951) );
  INV_X1 U16212 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19966) );
  NOR4_X1 U16213 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .A3(n12951), .A4(n19966), .ZN(n12876)
         );
  NOR4_X1 U16214 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_13__2__SCAN_IN), .A3(P2_UWORD_REG_11__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12875) );
  INV_X1 U16215 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12971) );
  NOR4_X1 U16216 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_EBX_REG_11__SCAN_IN), .A3(P1_LWORD_REG_11__SCAN_IN), .A4(n12971), 
        .ZN(n12874) );
  NOR4_X1 U16217 ( .A1(P3_ADDRESS_REG_24__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .A3(n19918), .A4(n18869), .ZN(n12873)
         );
  NAND4_X1 U16218 ( .A1(n12876), .A2(n12875), .A3(n12874), .A4(n12873), .ZN(
        n12892) );
  INV_X1 U16219 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n12880) );
  INV_X1 U16220 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12909) );
  INV_X1 U16221 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17789) );
  NOR4_X1 U16222 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(P1_EBX_REG_28__SCAN_IN), 
        .A3(n12909), .A4(n17789), .ZN(n12879) );
  INV_X1 U16223 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16494) );
  NAND4_X1 U16224 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_8__5__SCAN_IN), .A3(P2_REIP_REG_31__SCAN_IN), .A4(
        n16494), .ZN(n12877) );
  INV_X1 U16225 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n20306) );
  NOR2_X1 U16226 ( .A1(n12877), .A2(n20306), .ZN(n12878) );
  AND4_X1 U16227 ( .A1(n13410), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12883) );
  INV_X1 U16228 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n12881) );
  INV_X1 U16229 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15975) );
  AND4_X1 U16230 ( .A1(n12881), .A2(n15975), .A3(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .A4(P2_INSTQUEUE_REG_7__3__SCAN_IN), 
        .ZN(n12882) );
  AND4_X1 U16231 ( .A1(READY21_REG_SCAN_IN), .A2(n12883), .A3(n13166), .A4(
        n12882), .ZN(n12890) );
  INV_X1 U16232 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20061) );
  INV_X1 U16233 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20291) );
  NAND4_X1 U16234 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P1_ADDRESS_REG_7__SCAN_IN), .A3(n20061), .A4(n20291), .ZN(n12885) );
  INV_X1 U16235 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n18702) );
  NAND4_X1 U16236 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(
        P3_ADS_N_REG_SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(n18702), 
        .ZN(n12884) );
  NOR2_X1 U16237 ( .A1(n12885), .A2(n12884), .ZN(n12889) );
  INV_X1 U16238 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12898) );
  NAND4_X1 U16239 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(n12898), .A4(n13515), .ZN(
        n12887) );
  INV_X1 U16240 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12924) );
  NAND4_X1 U16241 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(n12959), .A4(n12924), .ZN(
        n12886) );
  NOR2_X1 U16242 ( .A1(n12887), .A2(n12886), .ZN(n12888) );
  NOR2_X1 U16243 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20936) );
  NAND4_X1 U16244 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n20936), .ZN(
        n12891) );
  NOR2_X1 U16245 ( .A1(n12892), .A2(n12891), .ZN(n12896) );
  INV_X1 U16246 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13920) );
  INV_X1 U16247 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21376) );
  NOR4_X1 U16248 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n15060), .A3(n13920), .A4(
        n21376), .ZN(n12895) );
  INV_X1 U16249 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21052) );
  NOR4_X1 U16250 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(P1_EAX_REG_12__SCAN_IN), 
        .A3(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A4(n21052), .ZN(n12894) );
  NOR4_X1 U16251 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(P3_EBX_REG_31__SCAN_IN), .A4(
        n13533), .ZN(n12893) );
  NAND4_X1 U16252 ( .A1(n12896), .A2(n12895), .A3(n12894), .A4(n12893), .ZN(
        n12922) );
  AOI22_X1 U16253 ( .A1(n12898), .A2(keyinput14), .B1(keyinput17), .B2(n18899), 
        .ZN(n12897) );
  OAI221_X1 U16254 ( .B1(n12898), .B2(keyinput14), .C1(n18899), .C2(keyinput17), .A(n12897), .ZN(n12906) );
  INV_X1 U16255 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16256 ( .A1(n20291), .A2(keyinput57), .B1(n12900), .B2(keyinput0), 
        .ZN(n12899) );
  OAI221_X1 U16257 ( .B1(n20291), .B2(keyinput57), .C1(n12900), .C2(keyinput0), 
        .A(n12899), .ZN(n12905) );
  XNOR2_X1 U16258 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B(keyinput48), .ZN(
        n12903) );
  XNOR2_X1 U16259 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput36), .ZN(
        n12902) );
  XNOR2_X1 U16260 ( .A(keyinput15), .B(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12901) );
  NAND3_X1 U16261 ( .A1(n12903), .A2(n12902), .A3(n12901), .ZN(n12904) );
  NOR3_X1 U16262 ( .A1(n12906), .A2(n12905), .A3(n12904), .ZN(n12921) );
  INV_X1 U16263 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21373) );
  AOI22_X1 U16264 ( .A1(n12880), .A2(keyinput62), .B1(n21373), .B2(keyinput32), 
        .ZN(n12907) );
  OAI221_X1 U16265 ( .B1(n12880), .B2(keyinput62), .C1(n21373), .C2(keyinput32), .A(n12907), .ZN(n12914) );
  AOI22_X1 U16266 ( .A1(n13410), .A2(keyinput56), .B1(keyinput33), .B2(n15975), 
        .ZN(n12908) );
  OAI221_X1 U16267 ( .B1(n13410), .B2(keyinput56), .C1(n15975), .C2(keyinput33), .A(n12908), .ZN(n12913) );
  XNOR2_X1 U16268 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B(keyinput2), .ZN(
        n12911) );
  XNOR2_X1 U16269 ( .A(keyinput55), .B(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12910) );
  NAND2_X1 U16270 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  NOR3_X1 U16271 ( .A1(n12914), .A2(n12913), .A3(n12912), .ZN(n12920) );
  AOI22_X1 U16272 ( .A1(n20861), .A2(keyinput35), .B1(keyinput23), .B2(n20061), 
        .ZN(n12915) );
  OAI221_X1 U16273 ( .B1(n20861), .B2(keyinput35), .C1(n20061), .C2(keyinput23), .A(n12915), .ZN(n12918) );
  INV_X1 U16274 ( .A(READY21_REG_SCAN_IN), .ZN(n12916) );
  XNOR2_X1 U16275 ( .A(n12916), .B(keyinput44), .ZN(n12917) );
  NOR2_X1 U16276 ( .A1(n12918), .A2(n12917), .ZN(n12919) );
  AND4_X1 U16277 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12945) );
  INV_X1 U16278 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18630) );
  AOI22_X1 U16279 ( .A1(n18630), .A2(keyinput12), .B1(n12924), .B2(keyinput45), 
        .ZN(n12923) );
  OAI221_X1 U16280 ( .B1(n18630), .B2(keyinput12), .C1(n12924), .C2(keyinput45), .A(n12923), .ZN(n12933) );
  INV_X1 U16281 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U16282 ( .A1(n21052), .A2(keyinput7), .B1(keyinput4), .B2(n12926), 
        .ZN(n12925) );
  OAI221_X1 U16283 ( .B1(n21052), .B2(keyinput7), .C1(n12926), .C2(keyinput4), 
        .A(n12925), .ZN(n12932) );
  INV_X1 U16284 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U16285 ( .A1(n12928), .A2(keyinput11), .B1(keyinput29), .B2(n20995), 
        .ZN(n12927) );
  OAI221_X1 U16286 ( .B1(n12928), .B2(keyinput11), .C1(n20995), .C2(keyinput29), .A(n12927), .ZN(n12931) );
  AOI22_X1 U16287 ( .A1(n20306), .A2(keyinput34), .B1(keyinput60), .B2(n12881), 
        .ZN(n12929) );
  OAI221_X1 U16288 ( .B1(n20306), .B2(keyinput34), .C1(n12881), .C2(keyinput60), .A(n12929), .ZN(n12930) );
  NOR4_X1 U16289 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12944) );
  INV_X1 U16290 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16291 ( .A1(n17789), .A2(keyinput25), .B1(n12935), .B2(keyinput43), 
        .ZN(n12934) );
  OAI221_X1 U16292 ( .B1(n17789), .B2(keyinput25), .C1(n12935), .C2(keyinput43), .A(n12934), .ZN(n12942) );
  AOI22_X1 U16293 ( .A1(n14921), .A2(keyinput22), .B1(n13533), .B2(keyinput37), 
        .ZN(n12936) );
  OAI221_X1 U16294 ( .B1(n14921), .B2(keyinput22), .C1(n13533), .C2(keyinput37), .A(n12936), .ZN(n12941) );
  INV_X1 U16295 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19082) );
  INV_X1 U16296 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16297 ( .A1(n19082), .A2(keyinput42), .B1(keyinput30), .B2(n13179), 
        .ZN(n12937) );
  OAI221_X1 U16298 ( .B1(n19082), .B2(keyinput42), .C1(n13179), .C2(keyinput30), .A(n12937), .ZN(n12940) );
  AOI22_X1 U16299 ( .A1(n20030), .A2(keyinput13), .B1(n13303), .B2(keyinput19), 
        .ZN(n12938) );
  OAI221_X1 U16300 ( .B1(n20030), .B2(keyinput13), .C1(n13303), .C2(keyinput19), .A(n12938), .ZN(n12939) );
  NOR4_X1 U16301 ( .A1(n12942), .A2(n12941), .A3(n12940), .A4(n12939), .ZN(
        n12943) );
  NAND4_X1 U16302 ( .A1(n12946), .A2(n12945), .A3(n12944), .A4(n12943), .ZN(
        n12981) );
  INV_X1 U16303 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n18389) );
  AOI22_X1 U16304 ( .A1(n18389), .A2(keyinput20), .B1(n15060), .B2(keyinput6), 
        .ZN(n12947) );
  OAI221_X1 U16305 ( .B1(n18389), .B2(keyinput20), .C1(n15060), .C2(keyinput6), 
        .A(n12947), .ZN(n12957) );
  AOI22_X1 U16306 ( .A1(n13920), .A2(keyinput5), .B1(keyinput39), .B2(n21376), 
        .ZN(n12948) );
  OAI221_X1 U16307 ( .B1(n13920), .B2(keyinput5), .C1(n21376), .C2(keyinput39), 
        .A(n12948), .ZN(n12956) );
  INV_X1 U16308 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16309 ( .A1(n12951), .A2(keyinput46), .B1(keyinput41), .B2(n12950), 
        .ZN(n12949) );
  OAI221_X1 U16310 ( .B1(n12951), .B2(keyinput46), .C1(n12950), .C2(keyinput41), .A(n12949), .ZN(n12955) );
  AOI22_X1 U16311 ( .A1(n12953), .A2(keyinput40), .B1(keyinput1), .B2(n19966), 
        .ZN(n12952) );
  OAI221_X1 U16312 ( .B1(n12953), .B2(keyinput40), .C1(n19966), .C2(keyinput1), 
        .A(n12952), .ZN(n12954) );
  NOR4_X1 U16313 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12979) );
  INV_X1 U16314 ( .A(P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21374) );
  AOI22_X1 U16315 ( .A1(n21374), .A2(keyinput31), .B1(n12959), .B2(keyinput24), 
        .ZN(n12958) );
  OAI221_X1 U16316 ( .B1(n21374), .B2(keyinput31), .C1(n12959), .C2(keyinput24), .A(n12958), .ZN(n12966) );
  INV_X1 U16317 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17805) );
  AOI22_X1 U16318 ( .A1(n18702), .A2(keyinput38), .B1(keyinput8), .B2(n17805), 
        .ZN(n12960) );
  OAI221_X1 U16319 ( .B1(n18702), .B2(keyinput38), .C1(n17805), .C2(keyinput8), 
        .A(n12960), .ZN(n12965) );
  AOI22_X1 U16320 ( .A1(n16494), .A2(keyinput47), .B1(n20063), .B2(keyinput61), 
        .ZN(n12961) );
  OAI221_X1 U16321 ( .B1(n16494), .B2(keyinput47), .C1(n20063), .C2(keyinput61), .A(n12961), .ZN(n12964) );
  AOI22_X1 U16322 ( .A1(n10841), .A2(keyinput3), .B1(keyinput54), .B2(n20858), 
        .ZN(n12962) );
  OAI221_X1 U16323 ( .B1(n10841), .B2(keyinput3), .C1(n20858), .C2(keyinput54), 
        .A(n12962), .ZN(n12963) );
  NOR4_X1 U16324 ( .A1(n12966), .A2(n12965), .A3(n12964), .A4(n12963), .ZN(
        n12978) );
  INV_X1 U16325 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U16326 ( .A1(n20829), .A2(keyinput59), .B1(keyinput9), .B2(n13699), 
        .ZN(n12967) );
  OAI221_X1 U16327 ( .B1(n20829), .B2(keyinput59), .C1(n13699), .C2(keyinput9), 
        .A(n12967), .ZN(n12976) );
  INV_X1 U16328 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16329 ( .A1(n20039), .A2(keyinput50), .B1(keyinput58), .B2(n12969), 
        .ZN(n12968) );
  OAI221_X1 U16330 ( .B1(n20039), .B2(keyinput50), .C1(n12969), .C2(keyinput58), .A(n12968), .ZN(n12975) );
  INV_X1 U16331 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U16332 ( .A1(n17318), .A2(keyinput16), .B1(n12971), .B2(keyinput49), 
        .ZN(n12970) );
  OAI221_X1 U16333 ( .B1(n17318), .B2(keyinput16), .C1(n12971), .C2(keyinput49), .A(n12970), .ZN(n12974) );
  AOI22_X1 U16334 ( .A1(n19228), .A2(keyinput63), .B1(n16404), .B2(keyinput21), 
        .ZN(n12972) );
  OAI221_X1 U16335 ( .B1(n19228), .B2(keyinput63), .C1(n16404), .C2(keyinput21), .A(n12972), .ZN(n12973) );
  NOR4_X1 U16336 ( .A1(n12976), .A2(n12975), .A3(n12974), .A4(n12973), .ZN(
        n12977) );
  NAND3_X1 U16337 ( .A1(n12979), .A2(n12978), .A3(n12977), .ZN(n12980) );
  NOR2_X1 U16338 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  XNOR2_X1 U16339 ( .A(n12983), .B(n12982), .ZN(P1_U2849) );
  INV_X1 U16340 ( .A(n14634), .ZN(n12987) );
  INV_X1 U16341 ( .A(n14650), .ZN(n12990) );
  NAND3_X1 U16342 ( .A1(n21369), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17630) );
  INV_X1 U16343 ( .A(n17630), .ZN(n12989) );
  NAND2_X1 U16344 ( .A1(n12990), .A2(n21101), .ZN(n13004) );
  MUX2_X1 U16345 ( .A(n15323), .B(n15227), .S(n15086), .Z(n12993) );
  XNOR2_X1 U16346 ( .A(n12994), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15320) );
  NAND2_X1 U16347 ( .A1(n21311), .A2(n12996), .ZN(n21463) );
  NAND2_X1 U16348 ( .A1(n21463), .A2(n21369), .ZN(n12997) );
  NAND2_X1 U16349 ( .A1(n21369), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16350 ( .A1(n21204), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12998) );
  AND2_X1 U16351 ( .A1(n12999), .A2(n12998), .ZN(n13824) );
  INV_X1 U16352 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21429) );
  NOR2_X1 U16353 ( .A1(n15176), .A2(n21429), .ZN(n15317) );
  AOI21_X1 U16354 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15317), .ZN(n13000) );
  OAI21_X1 U16355 ( .B1(n21106), .B2(n14656), .A(n13000), .ZN(n13001) );
  INV_X1 U16356 ( .A(n13001), .ZN(n13002) );
  INV_X1 U16357 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17836) );
  INV_X1 U16358 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13024) );
  NAND2_X1 U16359 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19012) );
  INV_X1 U16360 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16361 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18943) );
  NAND2_X1 U16362 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18855) );
  NAND2_X1 U16363 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18822) );
  NAND2_X1 U16364 ( .A1(n18797), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13007) );
  NAND2_X1 U16365 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18776) );
  XNOR2_X1 U16366 ( .A(n17836), .B(n13022), .ZN(n17835) );
  INV_X1 U16367 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13019) );
  NOR2_X1 U16368 ( .A1(n13007), .A2(n10189), .ZN(n13010) );
  INV_X1 U16369 ( .A(n13010), .ZN(n13011) );
  NOR2_X1 U16370 ( .A1(n18776), .A2(n13011), .ZN(n18745) );
  INV_X1 U16371 ( .A(n18745), .ZN(n13018) );
  NOR2_X1 U16372 ( .A1(n13019), .A2(n13018), .ZN(n13017) );
  NAND2_X1 U16373 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n13017), .ZN(
        n13008) );
  INV_X1 U16374 ( .A(n13023), .ZN(n17345) );
  AOI21_X1 U16375 ( .B1(n17859), .B2(n13008), .A(n17345), .ZN(n18735) );
  OAI21_X1 U16376 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n13017), .A(
        n13008), .ZN(n18756) );
  INV_X1 U16377 ( .A(n18756), .ZN(n17862) );
  INV_X1 U16378 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18790) );
  NOR2_X1 U16379 ( .A1(n18790), .A2(n13011), .ZN(n13009) );
  OAI21_X1 U16380 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13009), .A(
        n13018), .ZN(n18778) );
  INV_X1 U16381 ( .A(n18778), .ZN(n17890) );
  AOI22_X1 U16382 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13011), .B1(
        n13010), .B2(n18790), .ZN(n18787) );
  INV_X1 U16383 ( .A(n18787), .ZN(n17903) );
  AND2_X1 U16384 ( .A1(n18797), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18802) );
  OAI21_X1 U16385 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18802), .A(
        n13011), .ZN(n18798) );
  INV_X1 U16386 ( .A(n18798), .ZN(n17913) );
  INV_X1 U16387 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17933) );
  INV_X1 U16388 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16389 ( .A1(n18878), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17989) );
  INV_X1 U16390 ( .A(n17989), .ZN(n17977) );
  NAND2_X1 U16391 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17977), .ZN(
        n17976) );
  NOR2_X1 U16392 ( .A1(n18855), .A2(n17976), .ZN(n18813) );
  INV_X1 U16393 ( .A(n18813), .ZN(n17955) );
  NOR2_X1 U16394 ( .A1(n13016), .A2(n17955), .ZN(n13015) );
  NAND2_X1 U16395 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13015), .ZN(
        n13012) );
  AOI21_X1 U16396 ( .B1(n17933), .B2(n13012), .A(n18802), .ZN(n18815) );
  OAI21_X1 U16397 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n13015), .A(
        n13012), .ZN(n18826) );
  INV_X1 U16398 ( .A(n18826), .ZN(n17936) );
  NAND2_X1 U16399 ( .A1(n13022), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13013) );
  INV_X1 U16400 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18190) );
  AND2_X1 U16401 ( .A1(n18813), .A2(n18190), .ZN(n13014) );
  AOI21_X1 U16402 ( .B1(n13016), .B2(n17955), .A(n13015), .ZN(n18846) );
  NOR2_X1 U16403 ( .A1(n17934), .A2(n9628), .ZN(n17928) );
  NOR2_X1 U16404 ( .A1(n18815), .A2(n17928), .ZN(n17927) );
  NOR2_X1 U16405 ( .A1(n17927), .A2(n9628), .ZN(n17912) );
  NOR2_X1 U16406 ( .A1(n17913), .A2(n17912), .ZN(n17911) );
  NOR2_X1 U16407 ( .A1(n17911), .A2(n9628), .ZN(n17902) );
  NOR2_X1 U16408 ( .A1(n17903), .A2(n17902), .ZN(n17901) );
  NOR2_X1 U16409 ( .A1(n17901), .A2(n9628), .ZN(n17889) );
  NOR2_X1 U16410 ( .A1(n17890), .A2(n17889), .ZN(n17888) );
  NOR2_X1 U16411 ( .A1(n17888), .A2(n9628), .ZN(n17874) );
  INV_X1 U16412 ( .A(n17874), .ZN(n13021) );
  AOI21_X1 U16413 ( .B1(n13019), .B2(n13018), .A(n13017), .ZN(n18768) );
  NOR2_X1 U16414 ( .A1(n17852), .A2(n9628), .ZN(n17843) );
  INV_X1 U16415 ( .A(n17843), .ZN(n13026) );
  AOI21_X1 U16416 ( .B1(n13024), .B2(n13023), .A(n13022), .ZN(n17844) );
  INV_X1 U16417 ( .A(n17844), .ZN(n13025) );
  INV_X1 U16418 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17812) );
  NAND2_X1 U16419 ( .A1(n13166), .A2(n17812), .ZN(n19915) );
  NOR2_X2 U16420 ( .A1(n19895), .A2(n19915), .ZN(n18097) );
  NOR2_X1 U16421 ( .A1(n9628), .A2(n19913), .ZN(n18177) );
  INV_X1 U16422 ( .A(n18177), .ZN(n18113) );
  NOR3_X1 U16423 ( .A1(n17835), .A2(n17834), .A3(n18113), .ZN(n13187) );
  INV_X1 U16424 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19991) );
  AND2_X2 U16425 ( .A1(n14143), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13042) );
  NAND2_X1 U16426 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13030) );
  NAND2_X1 U16427 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13029) );
  AND2_X2 U16428 ( .A1(n14077), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13031) );
  NAND2_X1 U16429 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13028) );
  NAND2_X1 U16430 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13027) );
  AND2_X2 U16431 ( .A1(n13042), .A2(n13031), .ZN(n13069) );
  NAND2_X1 U16432 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13035) );
  NAND2_X1 U16433 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13034) );
  NAND2_X1 U16434 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13033) );
  INV_X2 U16435 ( .A(n13057), .ZN(n17436) );
  INV_X2 U16436 ( .A(n17436), .ZN(n18426) );
  NAND2_X1 U16437 ( .A1(n18426), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13032) );
  NAND2_X1 U16438 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13041) );
  NAND2_X1 U16439 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13040) );
  NAND2_X1 U16440 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13039) );
  BUF_X2 U16441 ( .A(n13103), .Z(n18427) );
  NAND2_X1 U16442 ( .A1(n18427), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13038) );
  NAND2_X1 U16443 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13048) );
  NAND2_X1 U16444 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13047) );
  AND2_X4 U16445 ( .A1(n13044), .A2(n14132), .ZN(n18286) );
  NAND2_X1 U16446 ( .A1(n18286), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13046) );
  NAND2_X1 U16447 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13045) );
  INV_X2 U16448 ( .A(n20037), .ZN(n20018) );
  NOR2_X1 U16449 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17811) );
  INV_X1 U16450 ( .A(n17811), .ZN(n19917) );
  NAND3_X1 U16451 ( .A1(n19932), .A2(n19996), .A3(n19917), .ZN(n19922) );
  AOI22_X1 U16452 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13069), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13056) );
  BUF_X2 U16453 ( .A(n13110), .Z(n17460) );
  AOI22_X1 U16454 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16455 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16456 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13053) );
  NAND4_X1 U16457 ( .A1(n13056), .A2(n13055), .A3(n13054), .A4(n13053), .ZN(
        n13063) );
  AOI22_X1 U16458 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9590), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16459 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13860), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13060) );
  CLKBUF_X3 U16460 ( .A(n13081), .Z(n18428) );
  AOI22_X1 U16461 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16462 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13058) );
  NAND4_X1 U16463 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13058), .ZN(
        n13062) );
  AOI22_X1 U16464 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16465 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16466 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16467 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13065) );
  NAND4_X1 U16468 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13065), .ZN(
        n13075) );
  AOI22_X1 U16469 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16470 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U16471 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16472 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13070) );
  NAND4_X1 U16473 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13074) );
  AOI22_X1 U16475 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16476 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16477 ( .A1(n18410), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16478 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13077) );
  NAND4_X1 U16479 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        n13087) );
  AOI22_X1 U16480 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16481 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16482 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16483 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13082) );
  NAND4_X1 U16484 ( .A1(n13085), .A2(n13084), .A3(n13083), .A4(n13082), .ZN(
        n13086) );
  AOI22_X1 U16485 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9597), .B1(
        n9619), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16486 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9592), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16487 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13860), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16488 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13088) );
  NAND4_X1 U16489 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        n13098) );
  AOI22_X1 U16490 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n17460), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16491 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n9595), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16492 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16493 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13093) );
  NAND4_X1 U16494 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13093), .ZN(
        n13097) );
  AOI22_X1 U16495 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16496 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16497 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16498 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13099) );
  NAND4_X1 U16499 ( .A1(n13102), .A2(n13101), .A3(n13100), .A4(n13099), .ZN(
        n13109) );
  AOI22_X1 U16500 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16501 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16502 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16503 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13104) );
  NAND4_X1 U16504 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13108) );
  AOI22_X1 U16505 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13110), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U16506 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13113) );
  AOI22_X1 U16507 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U16508 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16509 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16510 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16511 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13860), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16512 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13115) );
  NOR2_X1 U16513 ( .A1(n19449), .A2(n18479), .ZN(n13969) );
  NAND2_X1 U16514 ( .A1(n14069), .A2(n13969), .ZN(n14083) );
  NAND2_X1 U16515 ( .A1(n19426), .A2(n14057), .ZN(n13958) );
  NOR2_X2 U16516 ( .A1(n19446), .A2(n19449), .ZN(n13143) );
  AOI22_X1 U16517 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16518 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16519 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16520 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13119) );
  NAND4_X1 U16521 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13128) );
  AOI22_X1 U16522 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13126) );
  AOI22_X1 U16523 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U16524 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13860), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16525 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13123) );
  NAND4_X1 U16526 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13127) );
  NAND3_X1 U16527 ( .A1(n19434), .A2(n19442), .A3(n19449), .ZN(n13141) );
  NAND2_X1 U16528 ( .A1(n18479), .A2(n19434), .ZN(n13140) );
  NOR2_X1 U16529 ( .A1(n10457), .A2(n14103), .ZN(n14088) );
  NAND2_X1 U16530 ( .A1(n19430), .A2(n18620), .ZN(n13957) );
  NOR2_X1 U16531 ( .A1(n14088), .A2(n13957), .ZN(n13968) );
  AOI21_X1 U16532 ( .B1(n13140), .B2(n13141), .A(n13968), .ZN(n13134) );
  NOR2_X1 U16533 ( .A1(n13134), .A2(n19438), .ZN(n13139) );
  AND2_X1 U16534 ( .A1(n13958), .A2(n19434), .ZN(n13967) );
  NAND2_X1 U16535 ( .A1(n13135), .A2(n19438), .ZN(n13137) );
  NAND2_X1 U16536 ( .A1(n19442), .A2(n14103), .ZN(n13136) );
  INV_X1 U16537 ( .A(n13140), .ZN(n13972) );
  NAND2_X1 U16538 ( .A1(n13972), .A2(n18476), .ZN(n13980) );
  AOI21_X1 U16539 ( .B1(n13141), .B2(n13980), .A(n18620), .ZN(n13142) );
  AOI221_X1 U16540 ( .B1(n10457), .B2(n13129), .C1(n13143), .C2(n13129), .A(
        n13142), .ZN(n13144) );
  NAND2_X1 U16541 ( .A1(n13145), .A2(n13961), .ZN(n13959) );
  INV_X1 U16542 ( .A(n13959), .ZN(n13146) );
  MUX2_X1 U16543 ( .A(n19866), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13975) );
  NAND2_X1 U16544 ( .A1(n13975), .A2(n13974), .ZN(n13163) );
  NAND2_X1 U16545 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19866), .ZN(
        n13149) );
  NAND2_X1 U16546 ( .A1(n13163), .A2(n13149), .ZN(n13161) );
  MUX2_X1 U16547 ( .A(n19882), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13159) );
  NAND2_X1 U16548 ( .A1(n13161), .A2(n13159), .ZN(n13151) );
  NAND2_X1 U16549 ( .A1(n19882), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13150) );
  NAND2_X1 U16550 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U16551 ( .A1(n13152), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13156) );
  OAI22_X1 U16552 ( .A1(n13152), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19861), .ZN(n13154) );
  AOI21_X1 U16553 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13156), .A(
        n13154), .ZN(n13153) );
  NAND2_X1 U16554 ( .A1(n13154), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13158) );
  NOR2_X1 U16555 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19861), .ZN(
        n13155) );
  NAND2_X1 U16556 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  INV_X1 U16557 ( .A(n13159), .ZN(n13160) );
  XNOR2_X1 U16558 ( .A(n13161), .B(n13160), .ZN(n13162) );
  NAND2_X1 U16559 ( .A1(n13979), .A2(n13162), .ZN(n13976) );
  OAI21_X1 U16560 ( .B1(n13974), .B2(n13975), .A(n13163), .ZN(n13164) );
  NAND2_X1 U16561 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n13169) );
  INV_X1 U16562 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19954) );
  INV_X1 U16563 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19940) );
  NAND3_X1 U16564 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n18145) );
  NOR2_X1 U16565 ( .A1(n19940), .A2(n18145), .ZN(n18120) );
  NAND2_X1 U16566 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18120), .ZN(n18065) );
  INV_X1 U16567 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19949) );
  NAND2_X1 U16568 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n18105) );
  NOR2_X1 U16569 ( .A1(n19949), .A2(n18105), .ZN(n18066) );
  NAND3_X1 U16570 ( .A1(n18066), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n18055) );
  NOR3_X1 U16571 ( .A1(n19954), .A2(n18065), .A3(n18055), .ZN(n18025) );
  NAND2_X1 U16572 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18025), .ZN(n18033) );
  NOR2_X1 U16573 ( .A1(n19958), .A2(n18033), .ZN(n18016) );
  NAND2_X1 U16574 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18016), .ZN(n17996) );
  NAND2_X1 U16575 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17909) );
  NOR2_X1 U16576 ( .A1(n19966), .A2(n17909), .ZN(n17923) );
  INV_X1 U16577 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19972) );
  INV_X1 U16578 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19970) );
  INV_X1 U16579 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19968) );
  NOR3_X1 U16580 ( .A1(n19972), .A2(n19970), .A3(n19968), .ZN(n17924) );
  INV_X1 U16581 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19976) );
  INV_X1 U16582 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19974) );
  NOR2_X1 U16583 ( .A1(n19976), .A2(n19974), .ZN(n17926) );
  NAND4_X1 U16584 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17923), .A3(n17924), 
        .A4(n17926), .ZN(n17883) );
  NOR2_X1 U16585 ( .A1(n17996), .A2(n17883), .ZN(n17898) );
  NAND2_X1 U16586 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17898), .ZN(n13170) );
  NAND2_X1 U16587 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n13167) );
  NAND2_X1 U16588 ( .A1(n20039), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19729) );
  NOR2_X1 U16589 ( .A1(n19910), .A2(n19729), .ZN(n19903) );
  NOR4_X4 U16590 ( .A1(n19402), .A2(n20042), .A3(n18097), .A4(n19903), .ZN(
        n18189) );
  AOI221_X1 U16591 ( .B1(n18167), .B2(n13170), .C1(n18167), .C2(n13167), .A(
        n18189), .ZN(n17880) );
  INV_X1 U16592 ( .A(n17880), .ZN(n13168) );
  AOI221_X1 U16593 ( .B1(n19991), .B2(n18167), .C1(n13169), .C2(n18167), .A(
        n13168), .ZN(n17849) );
  INV_X1 U16594 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19990) );
  INV_X1 U16595 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19987) );
  NAND3_X1 U16596 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n17881), .ZN(n17863) );
  NOR3_X1 U16597 ( .A1(n19990), .A2(n19987), .A3(n17863), .ZN(n17847) );
  NAND2_X1 U16598 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17847), .ZN(n13174) );
  NOR2_X1 U16599 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n13174), .ZN(n17838) );
  INV_X1 U16600 ( .A(n17838), .ZN(n13171) );
  INV_X1 U16601 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19993) );
  AOI21_X1 U16602 ( .B1(n17849), .B2(n13171), .A(n19993), .ZN(n13172) );
  INV_X1 U16603 ( .A(n13172), .ZN(n13185) );
  OAI211_X2 U16604 ( .C1(n13179), .C2(n19430), .A(n19898), .B(n13181), .ZN(
        n18186) );
  INV_X1 U16605 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19995) );
  NOR3_X1 U16606 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19995), .A3(n13174), 
        .ZN(n13175) );
  AOI21_X1 U16607 ( .B1(n18132), .B2(P3_EBX_REG_31__SCAN_IN), .A(n13175), .ZN(
        n13176) );
  INV_X1 U16608 ( .A(n13176), .ZN(n13178) );
  INV_X1 U16609 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17346) );
  NOR2_X1 U16610 ( .A1(n13178), .A2(n13177), .ZN(n13184) );
  INV_X1 U16611 ( .A(n20023), .ZN(n20028) );
  NOR2_X1 U16612 ( .A1(n13179), .A2(n19430), .ZN(n13180) );
  INV_X1 U16613 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18453) );
  NAND2_X1 U16614 ( .A1(n18168), .A2(n18453), .ZN(n18154) );
  INV_X1 U16615 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18102) );
  INV_X1 U16616 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18402) );
  NAND2_X1 U16617 ( .A1(n18084), .A2(n18402), .ZN(n18077) );
  INV_X1 U16618 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18062) );
  INV_X1 U16619 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18006) );
  NAND2_X1 U16620 ( .A1(n18014), .A2(n18006), .ZN(n18005) );
  INV_X1 U16621 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17984) );
  NAND2_X1 U16622 ( .A1(n17992), .A2(n17984), .ZN(n17983) );
  INV_X1 U16623 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n18306) );
  INV_X1 U16624 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18279) );
  INV_X1 U16625 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n18241) );
  NAND2_X1 U16626 ( .A1(n17921), .A2(n18241), .ZN(n17916) );
  INV_X1 U16627 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17892) );
  INV_X1 U16628 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17867) );
  INV_X1 U16629 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U16630 ( .A1(n17851), .A2(n14514), .ZN(n17833) );
  NOR2_X1 U16631 ( .A1(n18185), .A2(n17833), .ZN(n17839) );
  INV_X1 U16632 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U16633 ( .A1(n17839), .A2(n13182), .ZN(n13183) );
  NAND3_X1 U16634 ( .A1(n13185), .A2(n13184), .A3(n13183), .ZN(n13186) );
  NAND2_X1 U16635 ( .A1(n13189), .A2(n10365), .ZN(n13190) );
  NAND2_X1 U16636 ( .A1(n13191), .A2(n13190), .ZN(n15894) );
  INV_X1 U16637 ( .A(n13194), .ZN(n13195) );
  NOR2_X1 U16638 ( .A1(n16545), .A2(n13197), .ZN(n13200) );
  NAND2_X1 U16639 ( .A1(n13200), .A2(n13198), .ZN(n13199) );
  OAI21_X1 U16640 ( .B1(n13200), .B2(n10469), .A(n13199), .ZN(n13201) );
  NAND2_X1 U16641 ( .A1(n16788), .A2(n20196), .ZN(n13213) );
  NOR2_X1 U16642 ( .A1(n13205), .A2(n13204), .ZN(n13206) );
  INV_X1 U16643 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15868) );
  NOR2_X1 U16644 ( .A1(n20207), .A2(n15868), .ZN(n16791) );
  AOI21_X1 U16645 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16791), .ZN(n13207) );
  OAI21_X1 U16646 ( .B1(n20199), .B2(n13208), .A(n13207), .ZN(n13209) );
  AOI21_X1 U16647 ( .B1(n15879), .B2(n20213), .A(n13209), .ZN(n13211) );
  NAND2_X1 U16648 ( .A1(n13213), .A2(n13212), .ZN(P2_U2986) );
  NOR2_X1 U16649 ( .A1(n14531), .A2(n15264), .ZN(n13220) );
  INV_X1 U16650 ( .A(n21106), .ZN(n15251) );
  NAND2_X1 U16651 ( .A1(n14562), .A2(n15251), .ZN(n13218) );
  INV_X1 U16652 ( .A(n21094), .ZN(n15249) );
  INV_X1 U16653 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14532) );
  OAI21_X1 U16654 ( .B1(n15249), .B2(n14532), .A(n13215), .ZN(n13216) );
  INV_X1 U16655 ( .A(n13216), .ZN(n13217) );
  OAI21_X1 U16656 ( .B1(n13222), .B2(n20932), .A(n13221), .ZN(P1_U2969) );
  NAND2_X1 U16657 ( .A1(n13223), .A2(n13679), .ZN(n13228) );
  NAND2_X1 U16658 ( .A1(n13254), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13224) );
  NAND2_X1 U16659 ( .A1(n20462), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13236) );
  AOI21_X1 U16660 ( .B1(n13236), .B2(n20885), .A(n20881), .ZN(n13226) );
  INV_X1 U16661 ( .A(n13236), .ZN(n13225) );
  NAND2_X1 U16662 ( .A1(n13225), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20728) );
  AOI22_X1 U16663 ( .A1(n13247), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13226), .B2(n20728), .ZN(n13227) );
  NOR2_X1 U16664 ( .A1(n14094), .A2(n13231), .ZN(n13232) );
  NAND2_X1 U16665 ( .A1(n13256), .A2(n13232), .ZN(n16219) );
  OAI21_X1 U16666 ( .B1(n13256), .B2(n13232), .A(n16219), .ZN(n14035) );
  INV_X1 U16667 ( .A(n14035), .ZN(n13253) );
  NOR2_X1 U16668 ( .A1(n14094), .A2(n13233), .ZN(n13241) );
  INV_X1 U16669 ( .A(n20462), .ZN(n13234) );
  NAND2_X1 U16670 ( .A1(n13234), .A2(n20894), .ZN(n13235) );
  NAND2_X1 U16671 ( .A1(n13236), .A2(n13235), .ZN(n20381) );
  NOR2_X1 U16672 ( .A1(n20381), .A2(n20881), .ZN(n13237) );
  AOI21_X1 U16673 ( .B1(n13247), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13237), .ZN(n13238) );
  NAND2_X1 U16674 ( .A1(n13239), .A2(n13238), .ZN(n13240) );
  NAND2_X1 U16675 ( .A1(n13240), .A2(n13241), .ZN(n13252) );
  NAND2_X1 U16676 ( .A1(n13247), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13242) );
  NAND2_X1 U16677 ( .A1(n17256), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20525) );
  NAND2_X1 U16678 ( .A1(n20679), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20555) );
  NAND2_X1 U16679 ( .A1(n20525), .A2(n20555), .ZN(n20434) );
  NAND2_X1 U16680 ( .A1(n20434), .A2(n20906), .ZN(n20557) );
  NAND2_X1 U16681 ( .A1(n13242), .A2(n20557), .ZN(n13243) );
  NOR2_X1 U16682 ( .A1(n20881), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13246) );
  INV_X1 U16683 ( .A(n13249), .ZN(n13250) );
  NAND2_X1 U16684 ( .A1(n13253), .A2(n14034), .ZN(n14033) );
  NAND2_X1 U16685 ( .A1(n13254), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13255) );
  NAND4_X1 U16686 ( .A1(n16401), .A2(n13258), .A3(n13257), .A4(n16392), .ZN(
        n13262) );
  NAND2_X1 U16687 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16391) );
  NAND2_X1 U16688 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13259) );
  NOR2_X1 U16689 ( .A1(n16391), .A2(n13259), .ZN(n13260) );
  NAND3_X1 U16690 ( .A1(n16409), .A2(n16394), .A3(n13260), .ZN(n13261) );
  NOR3_X1 U16691 ( .A1(n14094), .A2(n13262), .A3(n13261), .ZN(n13263) );
  INV_X1 U16692 ( .A(n16375), .ZN(n13277) );
  AOI22_X1 U16693 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13269) );
  NAND2_X1 U16694 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13265) );
  AOI22_X1 U16695 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13264) );
  AND2_X1 U16696 ( .A1(n13265), .A2(n13264), .ZN(n13268) );
  AOI22_X1 U16697 ( .A1(n13389), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13390), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16698 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13266) );
  NAND4_X1 U16699 ( .A1(n13269), .A2(n13268), .A3(n13267), .A4(n13266), .ZN(
        n13275) );
  AOI22_X1 U16700 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13397), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U16701 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U16702 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U16703 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13270) );
  NAND4_X1 U16704 ( .A1(n13273), .A2(n13272), .A3(n13271), .A4(n13270), .ZN(
        n13274) );
  NOR2_X1 U16705 ( .A1(n13275), .A2(n13274), .ZN(n16377) );
  AOI22_X1 U16706 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11395), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13283) );
  NAND2_X1 U16707 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13279) );
  AOI22_X1 U16708 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13278) );
  AND2_X1 U16709 ( .A1(n13279), .A2(n13278), .ZN(n13282) );
  AOI22_X1 U16710 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13390), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16711 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13280) );
  NAND4_X1 U16712 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13289) );
  AOI22_X1 U16713 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16714 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U16715 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13285) );
  NAND2_X1 U16716 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13284) );
  NAND4_X1 U16717 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13288) );
  NOR2_X1 U16718 ( .A1(n13289), .A2(n13288), .ZN(n16372) );
  INV_X1 U16719 ( .A(n16372), .ZN(n13290) );
  AOI22_X1 U16720 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11395), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U16721 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13292) );
  AOI22_X1 U16722 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13291) );
  AND2_X1 U16723 ( .A1(n13292), .A2(n13291), .ZN(n13295) );
  AOI22_X1 U16724 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13390), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U16725 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13293) );
  NAND4_X1 U16726 ( .A1(n13296), .A2(n13295), .A3(n13294), .A4(n13293), .ZN(
        n13302) );
  AOI22_X1 U16727 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16728 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U16729 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13298) );
  NAND2_X1 U16730 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13297) );
  NAND4_X1 U16731 ( .A1(n13300), .A2(n13299), .A3(n13298), .A4(n13297), .ZN(
        n13301) );
  NOR2_X1 U16732 ( .A1(n13302), .A2(n13301), .ZN(n16367) );
  OAI22_X1 U16733 ( .A1(n13322), .A2(n13303), .B1(n13320), .B2(n13458), .ZN(
        n13307) );
  INV_X1 U16734 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13305) );
  INV_X1 U16735 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13304) );
  OAI22_X1 U16736 ( .A1(n13305), .A2(n13324), .B1(n14041), .B2(n13304), .ZN(
        n13306) );
  NOR2_X1 U16737 ( .A1(n13307), .A2(n13306), .ZN(n13319) );
  NAND2_X1 U16738 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16739 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13310) );
  NAND2_X1 U16740 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13309) );
  AOI22_X1 U16741 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13308) );
  AND4_X1 U16742 ( .A1(n13311), .A2(n13310), .A3(n13309), .A4(n13308), .ZN(
        n13318) );
  AOI22_X1 U16743 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16744 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U16745 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13314) );
  NAND2_X1 U16746 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13313) );
  NAND2_X1 U16747 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13312) );
  AND4_X1 U16748 ( .A1(n13315), .A2(n13314), .A3(n13313), .A4(n13312), .ZN(
        n13316) );
  NAND4_X1 U16749 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n16363) );
  INV_X1 U16750 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13321) );
  INV_X1 U16751 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13485) );
  OAI22_X1 U16752 ( .A1(n13322), .A2(n13321), .B1(n13320), .B2(n13485), .ZN(
        n13327) );
  INV_X1 U16753 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13325) );
  OAI22_X1 U16754 ( .A1(n13325), .A2(n13324), .B1(n14041), .B2(n13323), .ZN(
        n13326) );
  NOR2_X1 U16755 ( .A1(n13327), .A2(n13326), .ZN(n13339) );
  NAND2_X1 U16756 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13331) );
  NAND2_X1 U16757 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13330) );
  NAND2_X1 U16758 ( .A1(n10736), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13329) );
  AOI22_X1 U16759 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13328) );
  AND4_X1 U16760 ( .A1(n13331), .A2(n13330), .A3(n13329), .A4(n13328), .ZN(
        n13338) );
  AOI22_X1 U16761 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U16762 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U16763 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13334) );
  NAND2_X1 U16764 ( .A1(n13397), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13333) );
  NAND2_X1 U16765 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13332) );
  AND4_X1 U16766 ( .A1(n13335), .A2(n13334), .A3(n13333), .A4(n13332), .ZN(
        n13336) );
  NAND4_X1 U16767 ( .A1(n13339), .A2(n13338), .A3(n13337), .A4(n13336), .ZN(
        n16359) );
  AOI22_X1 U16768 ( .A1(n11395), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U16769 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13341) );
  AOI22_X1 U16770 ( .A1(n10758), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13386), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13340) );
  AND2_X1 U16771 ( .A1(n13341), .A2(n13340), .ZN(n13344) );
  AOI22_X1 U16772 ( .A1(n13389), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13390), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16773 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13342) );
  NAND4_X1 U16774 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13351) );
  AOI22_X1 U16775 ( .A1(n10743), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13397), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U16776 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U16777 ( .A1(n13400), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U16778 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13346) );
  NAND4_X1 U16779 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13350) );
  NOR2_X1 U16780 ( .A1(n13351), .A2(n13350), .ZN(n16354) );
  AOI22_X1 U16781 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11395), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13358) );
  NAND2_X1 U16782 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13354) );
  AOI22_X1 U16783 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13353) );
  AND2_X1 U16784 ( .A1(n13354), .A2(n13353), .ZN(n13357) );
  AOI22_X1 U16785 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n13390), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13356) );
  AOI22_X1 U16786 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13355) );
  NAND4_X1 U16787 ( .A1(n13358), .A2(n13357), .A3(n13356), .A4(n13355), .ZN(
        n13364) );
  AOI22_X1 U16788 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U16789 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U16790 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U16791 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13359) );
  NAND4_X1 U16792 ( .A1(n13362), .A2(n13361), .A3(n13360), .A4(n13359), .ZN(
        n13363) );
  AOI22_X1 U16793 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13567), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16794 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13554), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U16795 ( .A1(n13413), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13374) );
  INV_X1 U16797 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13371) );
  INV_X1 U16798 ( .A(n13366), .ZN(n13562) );
  INV_X1 U16799 ( .A(n13562), .ZN(n17154) );
  NAND2_X1 U16800 ( .A1(n17154), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13370) );
  INV_X1 U16801 ( .A(n13367), .ZN(n13369) );
  NAND2_X1 U16802 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13368) );
  OAI211_X1 U16803 ( .C1(n10503), .C2(n13371), .A(n13370), .B(n13535), .ZN(
        n13372) );
  INV_X1 U16804 ( .A(n13372), .ZN(n13373) );
  NAND4_X1 U16805 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13385) );
  AOI22_X1 U16806 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13383) );
  INV_X1 U16807 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n20412) );
  INV_X1 U16808 ( .A(n13554), .ZN(n13560) );
  INV_X1 U16809 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13377) );
  OR2_X1 U16810 ( .A1(n13560), .A2(n13377), .ZN(n13378) );
  OAI211_X1 U16811 ( .C1(n13365), .C2(n20412), .A(n13558), .B(n13378), .ZN(
        n13379) );
  INV_X1 U16812 ( .A(n13379), .ZN(n13382) );
  AOI22_X1 U16813 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U16814 ( .A1(n13413), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13380) );
  NAND4_X1 U16815 ( .A1(n13383), .A2(n13382), .A3(n13381), .A4(n13380), .ZN(
        n13384) );
  NAND2_X1 U16816 ( .A1(n13385), .A2(n13384), .ZN(n13434) );
  NOR2_X1 U16817 ( .A1(n16324), .A2(n13434), .ZN(n13407) );
  AOI22_X1 U16818 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11395), .B1(
        n10736), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U16819 ( .A1(n10773), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13388) );
  AOI22_X1 U16820 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13386), .B1(
        n10758), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13387) );
  AND2_X1 U16821 ( .A1(n13388), .A2(n13387), .ZN(n13395) );
  AOI22_X1 U16822 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13390), .B1(
        n13389), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U16823 ( .A1(n13392), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13391), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13393) );
  NAND4_X1 U16824 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        n13406) );
  AOI22_X1 U16825 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13397), .B1(
        n10743), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U16826 ( .A1(n10802), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13398), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16827 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13400), .B1(
        n13399), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13402) );
  NAND2_X1 U16828 ( .A1(n10765), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13401) );
  NAND4_X1 U16829 ( .A1(n13404), .A2(n13403), .A3(n13402), .A4(n13401), .ZN(
        n13405) );
  NOR2_X1 U16830 ( .A1(n13406), .A2(n13405), .ZN(n13428) );
  XNOR2_X1 U16831 ( .A(n13407), .B(n13428), .ZN(n13432) );
  INV_X1 U16832 ( .A(n13434), .ZN(n13429) );
  NAND2_X1 U16833 ( .A1(n16324), .A2(n13429), .ZN(n16346) );
  NOR2_X2 U16834 ( .A1(n16343), .A2(n16346), .ZN(n16344) );
  AOI22_X1 U16835 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13417) );
  INV_X1 U16836 ( .A(n9624), .ZN(n13564) );
  OR2_X1 U16837 ( .A1(n13560), .A2(n13410), .ZN(n13411) );
  OAI211_X1 U16838 ( .C1(n13564), .C2(n17198), .A(n13558), .B(n13411), .ZN(
        n13412) );
  INV_X1 U16839 ( .A(n13412), .ZN(n13416) );
  AOI22_X1 U16840 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U16841 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U16842 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13427) );
  AOI22_X1 U16843 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13425) );
  OR2_X1 U16844 ( .A1(n13560), .A2(n13418), .ZN(n13419) );
  OAI211_X1 U16845 ( .C1(n13564), .C2(n13420), .A(n13535), .B(n13419), .ZN(
        n13421) );
  INV_X1 U16846 ( .A(n13421), .ZN(n13424) );
  AOI22_X1 U16847 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U16848 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13422) );
  NAND4_X1 U16849 ( .A1(n13425), .A2(n13424), .A3(n13423), .A4(n13422), .ZN(
        n13426) );
  AND2_X1 U16850 ( .A1(n13427), .A2(n13426), .ZN(n13433) );
  INV_X1 U16851 ( .A(n13428), .ZN(n13430) );
  AND2_X1 U16852 ( .A1(n13430), .A2(n13429), .ZN(n13431) );
  NAND2_X1 U16853 ( .A1(n13431), .A2(n13433), .ZN(n13436) );
  OAI211_X1 U16854 ( .C1(n13433), .C2(n13431), .A(n13473), .B(n13436), .ZN(
        n16338) );
  NAND2_X1 U16855 ( .A1(n16324), .A2(n13433), .ZN(n16340) );
  INV_X1 U16856 ( .A(n13436), .ZN(n13454) );
  AOI22_X1 U16857 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9617), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U16858 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U16859 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13442) );
  INV_X1 U16860 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13439) );
  INV_X1 U16861 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13437) );
  OR2_X1 U16862 ( .A1(n13560), .A2(n13437), .ZN(n13438) );
  OAI211_X1 U16863 ( .C1(n10707), .C2(n13439), .A(n13438), .B(n13558), .ZN(
        n13440) );
  INV_X1 U16864 ( .A(n13440), .ZN(n13441) );
  NAND4_X1 U16865 ( .A1(n13444), .A2(n13443), .A3(n13442), .A4(n13441), .ZN(
        n13453) );
  AOI22_X1 U16866 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13451) );
  INV_X1 U16867 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13446) );
  INV_X1 U16868 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17242) );
  OR2_X1 U16869 ( .A1(n13560), .A2(n17242), .ZN(n13445) );
  OAI211_X1 U16870 ( .C1(n13365), .C2(n13446), .A(n13535), .B(n13445), .ZN(
        n13447) );
  INV_X1 U16871 ( .A(n13447), .ZN(n13450) );
  AOI22_X1 U16872 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U16873 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13448) );
  NAND4_X1 U16874 ( .A1(n13451), .A2(n13450), .A3(n13449), .A4(n13448), .ZN(
        n13452) );
  AND2_X1 U16875 ( .A1(n13453), .A2(n13452), .ZN(n13477) );
  NAND2_X1 U16876 ( .A1(n13454), .A2(n13477), .ZN(n13455) );
  OAI211_X1 U16877 ( .C1(n13454), .C2(n13477), .A(n13473), .B(n13455), .ZN(
        n13475) );
  INV_X1 U16878 ( .A(n13455), .ZN(n13474) );
  AOI22_X1 U16879 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13463) );
  OR2_X1 U16880 ( .A1(n13560), .A2(n13456), .ZN(n13457) );
  OAI211_X1 U16881 ( .C1(n13564), .C2(n13458), .A(n13558), .B(n13457), .ZN(
        n13459) );
  INV_X1 U16882 ( .A(n13459), .ZN(n13462) );
  AOI22_X1 U16883 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U16884 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13460) );
  NAND4_X1 U16885 ( .A1(n13463), .A2(n13462), .A3(n13461), .A4(n13460), .ZN(
        n13472) );
  AOI22_X1 U16886 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13470) );
  OR2_X1 U16887 ( .A1(n13560), .A2(n17245), .ZN(n13464) );
  OAI211_X1 U16888 ( .C1(n13564), .C2(n13465), .A(n13535), .B(n13464), .ZN(
        n13466) );
  INV_X1 U16889 ( .A(n13466), .ZN(n13469) );
  AOI22_X1 U16890 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16891 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U16892 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  AND2_X1 U16893 ( .A1(n13472), .A2(n13471), .ZN(n16323) );
  NAND2_X1 U16894 ( .A1(n13474), .A2(n16323), .ZN(n13503) );
  OAI211_X1 U16895 ( .C1(n13474), .C2(n16323), .A(n13503), .B(n13473), .ZN(
        n16325) );
  XNOR2_X1 U16896 ( .A(n13476), .B(n10451), .ZN(n16321) );
  INV_X1 U16897 ( .A(n13477), .ZN(n13478) );
  NOR2_X1 U16898 ( .A1(n11309), .A2(n13478), .ZN(n16333) );
  NAND2_X1 U16899 ( .A1(n16321), .A2(n13479), .ZN(n13480) );
  INV_X1 U16900 ( .A(n10503), .ZN(n13551) );
  AOI22_X1 U16901 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13490) );
  INV_X1 U16902 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13483) );
  OR2_X1 U16903 ( .A1(n13560), .A2(n13483), .ZN(n13484) );
  OAI211_X1 U16904 ( .C1(n13564), .C2(n13485), .A(n13558), .B(n13484), .ZN(
        n13486) );
  INV_X1 U16905 ( .A(n13486), .ZN(n13489) );
  AOI22_X1 U16906 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U16907 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13487) );
  NAND4_X1 U16908 ( .A1(n13490), .A2(n13489), .A3(n13488), .A4(n13487), .ZN(
        n13500) );
  AOI22_X1 U16909 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13498) );
  INV_X1 U16910 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13491) );
  OR2_X1 U16911 ( .A1(n13560), .A2(n13491), .ZN(n13492) );
  OAI211_X1 U16912 ( .C1(n13564), .C2(n13493), .A(n13535), .B(n13492), .ZN(
        n13494) );
  INV_X1 U16913 ( .A(n13494), .ZN(n13497) );
  AOI22_X1 U16914 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U16915 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13495) );
  NAND4_X1 U16916 ( .A1(n13498), .A2(n13497), .A3(n13496), .A4(n13495), .ZN(
        n13499) );
  AND2_X1 U16917 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  INV_X1 U16918 ( .A(n13501), .ZN(n13506) );
  INV_X1 U16919 ( .A(n13503), .ZN(n13502) );
  NOR2_X1 U16920 ( .A1(n11297), .A2(n13506), .ZN(n16317) );
  AOI22_X1 U16921 ( .A1(n9609), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13514) );
  OR2_X1 U16922 ( .A1(n13560), .A2(n13507), .ZN(n13508) );
  OAI211_X1 U16923 ( .C1(n13564), .C2(n13509), .A(n13558), .B(n13508), .ZN(
        n13510) );
  INV_X1 U16924 ( .A(n13510), .ZN(n13513) );
  AOI22_X1 U16925 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U16926 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13511) );
  NAND4_X1 U16927 ( .A1(n13514), .A2(n13513), .A3(n13512), .A4(n13511), .ZN(
        n13524) );
  AOI22_X1 U16928 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13522) );
  OR2_X1 U16929 ( .A1(n13560), .A2(n13515), .ZN(n13516) );
  OAI211_X1 U16930 ( .C1(n13564), .C2(n13517), .A(n13535), .B(n13516), .ZN(
        n13518) );
  INV_X1 U16931 ( .A(n13518), .ZN(n13521) );
  AOI22_X1 U16932 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U16933 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13519) );
  NAND4_X1 U16934 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13523) );
  NAND2_X1 U16935 ( .A1(n13524), .A2(n13523), .ZN(n13545) );
  AOI22_X1 U16936 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9609), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U16937 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U16938 ( .A1(n13570), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13530) );
  INV_X1 U16939 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13527) );
  OR2_X1 U16940 ( .A1(n13560), .A2(n13525), .ZN(n13526) );
  OAI211_X1 U16941 ( .C1(n13365), .C2(n13527), .A(n13558), .B(n13526), .ZN(
        n13528) );
  INV_X1 U16942 ( .A(n13528), .ZN(n13529) );
  NAND4_X1 U16943 ( .A1(n13532), .A2(n13531), .A3(n13530), .A4(n13529), .ZN(
        n13543) );
  AOI22_X1 U16944 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13571), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U16945 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U16946 ( .A1(n13570), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17154), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13539) );
  INV_X1 U16947 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13536) );
  OR2_X1 U16948 ( .A1(n13560), .A2(n13533), .ZN(n13534) );
  OAI211_X1 U16949 ( .C1(n13564), .C2(n13536), .A(n13535), .B(n13534), .ZN(
        n13537) );
  INV_X1 U16950 ( .A(n13537), .ZN(n13538) );
  NAND4_X1 U16951 ( .A1(n13541), .A2(n13540), .A3(n13539), .A4(n13538), .ZN(
        n13542) );
  NAND2_X1 U16952 ( .A1(n13543), .A2(n13542), .ZN(n13548) );
  INV_X1 U16953 ( .A(n13545), .ZN(n16311) );
  NAND2_X1 U16954 ( .A1(n11309), .A2(n16311), .ZN(n13546) );
  OR2_X1 U16955 ( .A1(n16309), .A2(n13546), .ZN(n13547) );
  NOR2_X1 U16956 ( .A1(n13547), .A2(n13548), .ZN(n13549) );
  AOI21_X1 U16957 ( .B1(n13548), .B2(n13547), .A(n13549), .ZN(n16304) );
  NAND2_X1 U16958 ( .A1(n16305), .A2(n16304), .ZN(n16306) );
  INV_X1 U16959 ( .A(n13549), .ZN(n13550) );
  NAND2_X1 U16960 ( .A1(n16306), .A2(n13550), .ZN(n13579) );
  AOI22_X1 U16961 ( .A1(n13567), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13571), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U16962 ( .A1(n9617), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U16963 ( .A1(n13553), .A2(n13552), .ZN(n13577) );
  INV_X1 U16964 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13557) );
  AOI22_X1 U16965 ( .A1(n9624), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13556) );
  AOI21_X1 U16966 ( .B1(n13554), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13558), .ZN(n13555) );
  OAI211_X1 U16967 ( .C1(n13562), .C2(n13557), .A(n13556), .B(n13555), .ZN(
        n13576) );
  INV_X1 U16968 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13559) );
  OAI21_X1 U16969 ( .B1(n13560), .B2(n13559), .A(n13558), .ZN(n13566) );
  INV_X1 U16970 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13561) );
  OAI22_X1 U16971 ( .A1(n13564), .A2(n13563), .B1(n13562), .B2(n13561), .ZN(
        n13565) );
  AOI211_X1 U16972 ( .C1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n13567), .A(
        n13566), .B(n13565), .ZN(n13574) );
  AOI22_X1 U16973 ( .A1(n9616), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13551), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13573) );
  AOI22_X1 U16974 ( .A1(n13571), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13570), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13572) );
  NAND3_X1 U16975 ( .A1(n13574), .A2(n13573), .A3(n13572), .ZN(n13575) );
  OAI21_X1 U16976 ( .B1(n13577), .B2(n13576), .A(n13575), .ZN(n13578) );
  XNOR2_X1 U16977 ( .A(n13579), .B(n13578), .ZN(n13601) );
  NAND2_X1 U16978 ( .A1(n11221), .A2(n20917), .ZN(n13614) );
  OAI22_X1 U16979 ( .A1(n17266), .A2(n14043), .B1(n13616), .B2(n13614), .ZN(
        n13639) );
  INV_X1 U16980 ( .A(n13580), .ZN(n13581) );
  NOR2_X1 U16981 ( .A1(n11307), .A2(n20133), .ZN(n20128) );
  NAND2_X1 U16982 ( .A1(n13601), .A2(n20128), .ZN(n13600) );
  NOR4_X1 U16983 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13587) );
  NOR4_X1 U16984 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13586) );
  NOR4_X1 U16985 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13585) );
  NOR4_X1 U16986 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13584) );
  AND4_X1 U16987 ( .A1(n13587), .A2(n13586), .A3(n13585), .A4(n13584), .ZN(
        n13592) );
  NOR4_X1 U16988 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13590) );
  NOR4_X1 U16989 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13589) );
  NOR4_X1 U16990 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13588) );
  AND4_X1 U16991 ( .A1(n13590), .A2(n13589), .A3(n13588), .A4(n20812), .ZN(
        n13591) );
  NAND2_X1 U16992 ( .A1(n13592), .A2(n13591), .ZN(n13593) );
  INV_X1 U16993 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n13596) );
  MUX2_X1 U16994 ( .A(BUF2_REG_14__SCAN_IN), .B(BUF1_REG_14__SCAN_IN), .S(
        n17185), .Z(n14352) );
  AOI22_X1 U16995 ( .A1(n20114), .A2(n14352), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20133), .ZN(n13595) );
  OAI21_X1 U16996 ( .B1(n16513), .B2(n13596), .A(n13595), .ZN(n13597) );
  AOI21_X1 U16997 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n20116), .A(n13597), .ZN(
        n13598) );
  NAND2_X1 U16998 ( .A1(n13600), .A2(n10471), .ZN(P2_U2889) );
  NAND2_X1 U16999 ( .A1(n16418), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13603) );
  INV_X1 U17000 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20896) );
  NOR2_X1 U17001 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n20896), .ZN(n13605) );
  NOR4_X1 U17002 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13604) );
  NAND4_X1 U17003 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13605), .A3(n13604), .A4(
        n20861), .ZN(n13608) );
  INV_X1 U17004 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21460) );
  NOR3_X1 U17005 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21460), .ZN(n13607) );
  NOR4_X1 U17006 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13606) );
  NAND4_X1 U17007 ( .A1(n14974), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13607), .A4(
        n13606), .ZN(U214) );
  NOR2_X1 U17008 ( .A1(n17186), .A2(n13608), .ZN(n17708) );
  NAND2_X1 U17009 ( .A1(n17708), .A2(U214), .ZN(U212) );
  NAND2_X1 U17010 ( .A1(n20917), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U17011 ( .B1(n20050), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17289), 
        .ZN(n13609) );
  AOI21_X1 U17012 ( .B1(n13609), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13610) );
  NOR2_X1 U17013 ( .A1(n17115), .A2(n20912), .ZN(n17675) );
  NOR2_X1 U17014 ( .A1(n13610), .A2(n17675), .ZN(P2_U3178) );
  NOR2_X1 U17015 ( .A1(n11243), .A2(n17677), .ZN(n13675) );
  NAND2_X1 U17016 ( .A1(n13675), .A2(n13611), .ZN(n16303) );
  INV_X1 U17017 ( .A(n16303), .ZN(n13613) );
  INV_X1 U17018 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13612) );
  OAI211_X1 U17019 ( .C1(n13613), .C2(n13612), .A(n13621), .B(n13668), .ZN(
        P2_U2814) );
  INV_X1 U17020 ( .A(n13614), .ZN(n13615) );
  NOR3_X1 U17021 ( .A1(n13616), .A2(n13615), .A3(n13640), .ZN(n17273) );
  NOR2_X1 U17022 ( .A1(n17273), .A2(n17677), .ZN(n20897) );
  OAI21_X1 U17023 ( .B1(n20897), .B2(n13618), .A(n13617), .ZN(P2_U2819) );
  INV_X1 U17024 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13619) );
  OAI22_X1 U17025 ( .A1(n13620), .A2(n13619), .B1(n20912), .B2(n13621), .ZN(
        P2_U2816) );
  INV_X1 U17026 ( .A(n13621), .ZN(n13622) );
  OAI21_X1 U17027 ( .B1(n13622), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20908), 
        .ZN(n13623) );
  OAI21_X1 U17028 ( .B1(n20915), .B2(n20908), .A(n13623), .ZN(P2_U3612) );
  AND2_X1 U17029 ( .A1(n13657), .A2(n12614), .ZN(n13650) );
  NAND2_X1 U17030 ( .A1(n13650), .A2(n13624), .ZN(n14535) );
  AND2_X1 U17031 ( .A1(n21285), .A2(n13625), .ZN(n14732) );
  AOI21_X1 U17032 ( .B1(n14535), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14732), 
        .ZN(n13626) );
  NAND2_X1 U17033 ( .A1(n14536), .A2(n13626), .ZN(P1_U2801) );
  INV_X1 U17034 ( .A(n13627), .ZN(n16291) );
  NOR2_X1 U17035 ( .A1(n16291), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13629) );
  NOR2_X1 U17036 ( .A1(n13629), .A2(n13628), .ZN(n17660) );
  OAI21_X1 U17037 ( .B1(n13631), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13630), .ZN(n17664) );
  NAND2_X1 U17038 ( .A1(n20179), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n17662) );
  OAI21_X1 U17039 ( .B1(n16773), .B2(n17664), .A(n17662), .ZN(n13632) );
  AOI21_X1 U17040 ( .B1(n20196), .B2(n17660), .A(n13632), .ZN(n13635) );
  OAI21_X1 U17041 ( .B1(n20204), .B2(n13633), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13634) );
  OAI211_X1 U17042 ( .C1(n20194), .C2(n13666), .A(n13635), .B(n13634), .ZN(
        P2_U3014) );
  NAND2_X1 U17043 ( .A1(n13637), .A2(n13636), .ZN(n13638) );
  NOR2_X1 U17044 ( .A1(n13639), .A2(n13638), .ZN(n13642) );
  INV_X1 U17045 ( .A(n11243), .ZN(n13648) );
  NAND3_X1 U17046 ( .A1(n13676), .A2(n13648), .A3(n13640), .ZN(n13641) );
  NAND2_X1 U17047 ( .A1(n13642), .A2(n13641), .ZN(n17253) );
  NAND2_X1 U17048 ( .A1(n17253), .A2(n13643), .ZN(n13646) );
  NAND2_X1 U17049 ( .A1(n20912), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17294) );
  INV_X1 U17050 ( .A(n17294), .ZN(n13644) );
  AOI21_X1 U17051 ( .B1(n17675), .B2(P2_FLUSH_REG_SCAN_IN), .A(n13644), .ZN(
        n13645) );
  AND2_X1 U17052 ( .A1(n17149), .A2(n17288), .ZN(n17169) );
  INV_X1 U17053 ( .A(n17169), .ZN(n13649) );
  NAND3_X1 U17054 ( .A1(n13648), .A2(n16324), .A3(n13647), .ZN(n17274) );
  OAI22_X1 U17055 ( .A1(n13649), .A2(n17274), .B1(n10937), .B2(n17149), .ZN(
        P2_U3595) );
  INV_X1 U17056 ( .A(n11674), .ZN(n13651) );
  OAI22_X1 U17057 ( .A1(n13851), .A2(n9625), .B1(n13651), .B2(n13650), .ZN(
        n20928) );
  NOR3_X1 U17058 ( .A1(n9625), .A2(n13829), .A3(n17543), .ZN(n13652) );
  NOR2_X1 U17059 ( .A1(n13652), .A2(n21467), .ZN(n21469) );
  NOR2_X1 U17060 ( .A1(n20928), .A2(n21469), .ZN(n17513) );
  NOR2_X1 U17061 ( .A1(n17513), .A2(n20927), .ZN(n20934) );
  INV_X1 U17062 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13662) );
  OAI21_X1 U17063 ( .B1(n14541), .B2(n13654), .A(n13653), .ZN(n13655) );
  MUX2_X1 U17064 ( .A(n14220), .B(n13655), .S(n17532), .Z(n13659) );
  INV_X1 U17065 ( .A(n12614), .ZN(n13656) );
  NOR2_X1 U17066 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  OAI21_X1 U17067 ( .B1(n13659), .B2(n13658), .A(n14317), .ZN(n17515) );
  INV_X1 U17068 ( .A(n17515), .ZN(n13660) );
  NAND2_X1 U17069 ( .A1(n20934), .A2(n13660), .ZN(n13661) );
  OAI21_X1 U17070 ( .B1(n20934), .B2(n13662), .A(n13661), .ZN(P1_U3484) );
  NAND2_X1 U17071 ( .A1(n11309), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13664) );
  MUX2_X1 U17072 ( .A(n10628), .B(n13666), .S(n20112), .Z(n13667) );
  OAI21_X1 U17073 ( .B1(n17220), .B2(n20101), .A(n13667), .ZN(P2_U2887) );
  NOR2_X1 U17074 ( .A1(n13668), .A2(n20910), .ZN(n13669) );
  INV_X1 U17075 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13674) );
  INV_X1 U17076 ( .A(n13783), .ZN(n13673) );
  INV_X1 U17077 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14438) );
  NOR2_X1 U17078 ( .A1(n17186), .A2(n14438), .ZN(n13671) );
  AOI21_X1 U17079 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n17186), .A(n13671), .ZN(
        n14478) );
  INV_X1 U17080 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13672) );
  OAI222_X1 U17081 ( .A1(n13743), .A2(n13674), .B1(n13673), .B2(n14478), .C1(
        n13672), .C2(n13762), .ZN(P2_U2982) );
  INV_X1 U17082 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U17083 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  INV_X1 U17084 ( .A(n20794), .ZN(n20911) );
  INV_X1 U17085 ( .A(n20178), .ZN(n13681) );
  NAND2_X1 U17086 ( .A1(n13681), .A2(n13680), .ZN(n13705) );
  INV_X1 U17087 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13752) );
  INV_X1 U17088 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n13682) );
  OAI222_X1 U17089 ( .A1(n13683), .A2(n20145), .B1(n13705), .B2(n13752), .C1(
        n20909), .C2(n13682), .ZN(P2_U2921) );
  INV_X1 U17090 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13685) );
  INV_X1 U17091 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13763) );
  INV_X1 U17092 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13684) );
  OAI222_X1 U17093 ( .A1(n13685), .A2(n20145), .B1(n13705), .B2(n13763), .C1(
        n20909), .C2(n13684), .ZN(P2_U2923) );
  INV_X1 U17094 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13687) );
  INV_X1 U17095 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13736) );
  INV_X1 U17096 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13686) );
  OAI222_X1 U17097 ( .A1(n13687), .A2(n20145), .B1(n13705), .B2(n13736), .C1(
        n20909), .C2(n13686), .ZN(P2_U2931) );
  INV_X1 U17098 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13689) );
  INV_X1 U17099 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13759) );
  INV_X1 U17100 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13688) );
  OAI222_X1 U17101 ( .A1(n13689), .A2(n20145), .B1(n13705), .B2(n13759), .C1(
        n20909), .C2(n13688), .ZN(P2_U2929) );
  INV_X1 U17102 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13691) );
  INV_X1 U17103 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13742) );
  INV_X1 U17104 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13690) );
  OAI222_X1 U17105 ( .A1(n13691), .A2(n20145), .B1(n13705), .B2(n13742), .C1(
        n20909), .C2(n13690), .ZN(P2_U2935) );
  INV_X1 U17106 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13693) );
  INV_X1 U17107 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13739) );
  INV_X1 U17108 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13692) );
  OAI222_X1 U17109 ( .A1(n13693), .A2(n20145), .B1(n13705), .B2(n13739), .C1(
        n20909), .C2(n13692), .ZN(P2_U2933) );
  INV_X1 U17110 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13695) );
  INV_X1 U17111 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13694) );
  OAI222_X1 U17112 ( .A1(n13695), .A2(n20145), .B1(n13705), .B2(n16494), .C1(
        n20909), .C2(n13694), .ZN(P2_U2932) );
  INV_X1 U17113 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13697) );
  INV_X1 U17114 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13755) );
  INV_X1 U17115 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13696) );
  OAI222_X1 U17116 ( .A1(n13697), .A2(n20145), .B1(n13705), .B2(n13755), .C1(
        n20909), .C2(n13696), .ZN(P2_U2925) );
  INV_X1 U17117 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16480) );
  INV_X1 U17118 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13698) );
  OAI222_X1 U17119 ( .A1(n13705), .A2(n16480), .B1(n20145), .B2(n17789), .C1(
        n20909), .C2(n13698), .ZN(P2_U2930) );
  INV_X1 U17120 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13700) );
  INV_X1 U17121 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n17795) );
  OAI222_X1 U17122 ( .A1(n13705), .A2(n13700), .B1(n20145), .B2(n17795), .C1(
        n20909), .C2(n13699), .ZN(P2_U2924) );
  NOR2_X1 U17123 ( .A1(n20243), .A2(n16418), .ZN(n13703) );
  AOI21_X1 U17124 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16418), .A(n13703), .ZN(
        n13704) );
  OAI21_X1 U17125 ( .B1(n20251), .B2(n20101), .A(n13704), .ZN(P2_U2886) );
  INV_X1 U17126 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13707) );
  INV_X1 U17127 ( .A(n13705), .ZN(n13714) );
  AOI22_X1 U17128 ( .A1(n13714), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n20175), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13706) );
  OAI21_X1 U17129 ( .B1(n20145), .B2(n13707), .A(n13706), .ZN(P2_U2928) );
  INV_X1 U17130 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U17131 ( .A1(n13714), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n20175), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U17132 ( .B1(n20145), .B2(n13709), .A(n13708), .ZN(P2_U2926) );
  INV_X1 U17133 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U17134 ( .A1(n13714), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n20175), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13710) );
  OAI21_X1 U17135 ( .B1(n20145), .B2(n13711), .A(n13710), .ZN(P2_U2934) );
  INV_X1 U17136 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17137 ( .A1(n13714), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n20175), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U17138 ( .B1(n20145), .B2(n13713), .A(n13712), .ZN(P2_U2927) );
  INV_X1 U17139 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U17140 ( .A1(n13714), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n20175), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13715) );
  OAI21_X1 U17141 ( .B1(n20145), .B2(n13716), .A(n13715), .ZN(P2_U2922) );
  INV_X1 U17142 ( .A(n17168), .ZN(n20221) );
  INV_X1 U17143 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n16263) );
  MUX2_X1 U17144 ( .A(n20221), .B(n16263), .S(n16418), .Z(n13720) );
  OAI21_X1 U17145 ( .B1(n20889), .B2(n20101), .A(n13720), .ZN(P2_U2885) );
  INV_X1 U17146 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13726) );
  INV_X1 U17147 ( .A(n15501), .ZN(n13721) );
  NAND2_X1 U17148 ( .A1(n13721), .A2(n17543), .ZN(n13831) );
  AND2_X1 U17149 ( .A1(n14436), .A2(n17543), .ZN(n13722) );
  NAND2_X1 U17150 ( .A1(n12603), .A2(n13722), .ZN(n17523) );
  AND2_X1 U17151 ( .A1(n13831), .A2(n17523), .ZN(n13723) );
  NAND2_X1 U17152 ( .A1(n21369), .A2(n17632), .ZN(n21466) );
  NOR2_X4 U17153 ( .A1(n21044), .A2(n21067), .ZN(n21055) );
  AOI22_X1 U17154 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13725) );
  OAI21_X1 U17155 ( .B1(n13726), .B2(n14163), .A(n13725), .ZN(P1_U2910) );
  INV_X1 U17156 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U17157 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13727) );
  OAI21_X1 U17158 ( .B1(n13728), .B2(n14163), .A(n13727), .ZN(P1_U2908) );
  INV_X1 U17159 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U17160 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13729) );
  OAI21_X1 U17161 ( .B1(n13730), .B2(n14163), .A(n13729), .ZN(P1_U2911) );
  INV_X1 U17162 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13732) );
  AOI22_X1 U17163 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17164 ( .B1(n13732), .B2(n14163), .A(n13731), .ZN(P1_U2907) );
  NAND2_X1 U17165 ( .A1(n13801), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13735) );
  NAND2_X1 U17166 ( .A1(n17186), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U17167 ( .A1(n17185), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13733) );
  AND2_X1 U17168 ( .A1(n13734), .A2(n13733), .ZN(n20132) );
  NAND2_X1 U17169 ( .A1(n13783), .A2(n17210), .ZN(n13764) );
  OAI211_X1 U17170 ( .C1(n13736), .C2(n13762), .A(n13735), .B(n13764), .ZN(
        P2_U2956) );
  NAND2_X1 U17171 ( .A1(n13801), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13738) );
  INV_X1 U17172 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19433) );
  NAND2_X1 U17173 ( .A1(n17185), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13737) );
  OAI21_X1 U17174 ( .B1(n17185), .B2(n19433), .A(n13737), .ZN(n17238) );
  NAND2_X1 U17175 ( .A1(n13783), .A2(n17238), .ZN(n13775) );
  OAI211_X1 U17176 ( .C1(n13739), .C2(n13762), .A(n13738), .B(n13775), .ZN(
        P2_U2954) );
  NAND2_X1 U17177 ( .A1(n13801), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13741) );
  NOR2_X1 U17178 ( .A1(n17185), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13740) );
  AOI21_X1 U17179 ( .B1(n17185), .B2(n12880), .A(n13740), .ZN(n20113) );
  NAND2_X1 U17180 ( .A1(n13783), .A2(n20113), .ZN(n13746) );
  OAI211_X1 U17181 ( .C1(n13742), .C2(n13762), .A(n13741), .B(n13746), .ZN(
        P2_U2952) );
  INV_X1 U17182 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20152) );
  INV_X2 U17183 ( .A(n13743), .ZN(n13801) );
  NAND2_X1 U17184 ( .A1(n13801), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13745) );
  INV_X1 U17185 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18721) );
  NAND2_X1 U17186 ( .A1(n17185), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13744) );
  OAI21_X1 U17187 ( .B1(n17185), .B2(n18721), .A(n13744), .ZN(n16433) );
  NAND2_X1 U17188 ( .A1(n13783), .A2(n16433), .ZN(n13760) );
  OAI211_X1 U17189 ( .C1(n20152), .C2(n13762), .A(n13745), .B(n13760), .ZN(
        P2_U2979) );
  NAND2_X1 U17190 ( .A1(n13801), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13747) );
  OAI211_X1 U17191 ( .C1(n11299), .C2(n13762), .A(n13747), .B(n13746), .ZN(
        P2_U2967) );
  INV_X1 U17192 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20156) );
  NAND2_X1 U17193 ( .A1(n13801), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13748) );
  MUX2_X1 U17194 ( .A(BUF2_REG_10__SCAN_IN), .B(BUF1_REG_10__SCAN_IN), .S(
        n17185), .Z(n16447) );
  NAND2_X1 U17195 ( .A1(n13783), .A2(n16447), .ZN(n13753) );
  OAI211_X1 U17196 ( .C1(n20156), .C2(n13762), .A(n13748), .B(n13753), .ZN(
        P2_U2977) );
  INV_X1 U17197 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20148) );
  NAND2_X1 U17198 ( .A1(n13801), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U17199 ( .A1(n13783), .A2(n14352), .ZN(n13750) );
  OAI211_X1 U17200 ( .C1(n20148), .C2(n13762), .A(n13749), .B(n13750), .ZN(
        P2_U2981) );
  NAND2_X1 U17201 ( .A1(n13801), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13751) );
  OAI211_X1 U17202 ( .C1(n13752), .C2(n13762), .A(n13751), .B(n13750), .ZN(
        P2_U2966) );
  NAND2_X1 U17203 ( .A1(n13801), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13754) );
  OAI211_X1 U17204 ( .C1(n13755), .C2(n13762), .A(n13754), .B(n13753), .ZN(
        P2_U2962) );
  NAND2_X1 U17205 ( .A1(n13801), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13758) );
  INV_X1 U17206 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U17207 ( .A1(n17185), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13756) );
  OAI21_X1 U17208 ( .B1(n17185), .B2(n13757), .A(n13756), .ZN(n20278) );
  NAND2_X1 U17209 ( .A1(n13783), .A2(n20278), .ZN(n13772) );
  OAI211_X1 U17210 ( .C1(n13759), .C2(n13762), .A(n13758), .B(n13772), .ZN(
        P2_U2958) );
  NAND2_X1 U17211 ( .A1(n13801), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13761) );
  OAI211_X1 U17212 ( .C1(n13763), .C2(n13762), .A(n13761), .B(n13760), .ZN(
        P2_U2964) );
  AOI22_X1 U17213 ( .A1(n13801), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13791), .ZN(n13765) );
  NAND2_X1 U17214 ( .A1(n13765), .A2(n13764), .ZN(P2_U2971) );
  AOI22_X1 U17215 ( .A1(n13801), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n13791), .ZN(n13767) );
  INV_X1 U17216 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17755) );
  NAND2_X1 U17217 ( .A1(n17185), .A2(n17755), .ZN(n13766) );
  OAI21_X1 U17218 ( .B1(n17185), .B2(BUF2_REG_5__SCAN_IN), .A(n13766), .ZN(
        n20271) );
  INV_X1 U17219 ( .A(n20271), .ZN(n16521) );
  NAND2_X1 U17220 ( .A1(n13783), .A2(n16521), .ZN(n13795) );
  NAND2_X1 U17221 ( .A1(n13767), .A2(n13795), .ZN(P2_U2972) );
  AOI22_X1 U17222 ( .A1(n13801), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13791), .ZN(n13770) );
  INV_X1 U17223 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17759) );
  NAND2_X1 U17224 ( .A1(n17185), .A2(n17759), .ZN(n13768) );
  OAI21_X1 U17225 ( .B1(n17185), .B2(BUF2_REG_3__SCAN_IN), .A(n13768), .ZN(
        n20143) );
  INV_X1 U17226 ( .A(n20143), .ZN(n13769) );
  NAND2_X1 U17227 ( .A1(n13783), .A2(n13769), .ZN(n13802) );
  NAND2_X1 U17228 ( .A1(n13770), .A2(n13802), .ZN(P2_U2970) );
  AOI22_X1 U17229 ( .A1(n13801), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13794), .ZN(n13771) );
  MUX2_X1 U17230 ( .A(BUF2_REG_13__SCAN_IN), .B(BUF1_REG_13__SCAN_IN), .S(
        n17185), .Z(n16426) );
  NAND2_X1 U17231 ( .A1(n13783), .A2(n16426), .ZN(n13785) );
  NAND2_X1 U17232 ( .A1(n13771), .A2(n13785), .ZN(P2_U2965) );
  AOI22_X1 U17233 ( .A1(n13801), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n13794), .ZN(n13773) );
  NAND2_X1 U17234 ( .A1(n13773), .A2(n13772), .ZN(P2_U2973) );
  AOI22_X1 U17235 ( .A1(n13801), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n13794), .ZN(n13774) );
  MUX2_X1 U17236 ( .A(BUF2_REG_8__SCAN_IN), .B(BUF1_REG_8__SCAN_IN), .S(n17185), .Z(n16460) );
  NAND2_X1 U17237 ( .A1(n13783), .A2(n16460), .ZN(n13792) );
  NAND2_X1 U17238 ( .A1(n13774), .A2(n13792), .ZN(P2_U2975) );
  AOI22_X1 U17239 ( .A1(n13801), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n13794), .ZN(n13776) );
  NAND2_X1 U17240 ( .A1(n13776), .A2(n13775), .ZN(P2_U2969) );
  AOI22_X1 U17241 ( .A1(n13801), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n13794), .ZN(n13779) );
  NAND2_X1 U17242 ( .A1(n17186), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U17243 ( .A1(n17185), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13777) );
  AND2_X1 U17244 ( .A1(n13778), .A2(n13777), .ZN(n17192) );
  INV_X1 U17245 ( .A(n17192), .ZN(n16510) );
  NAND2_X1 U17246 ( .A1(n13783), .A2(n16510), .ZN(n13799) );
  NAND2_X1 U17247 ( .A1(n13779), .A2(n13799), .ZN(P2_U2968) );
  AOI22_X1 U17248 ( .A1(n13801), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13794), .ZN(n13780) );
  MUX2_X1 U17249 ( .A(BUF2_REG_11__SCAN_IN), .B(BUF1_REG_11__SCAN_IN), .S(
        n17185), .Z(n16440) );
  NAND2_X1 U17250 ( .A1(n13783), .A2(n16440), .ZN(n13797) );
  NAND2_X1 U17251 ( .A1(n13780), .A2(n13797), .ZN(P2_U2978) );
  AOI22_X1 U17252 ( .A1(n13801), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13794), .ZN(n13781) );
  MUX2_X1 U17253 ( .A(BUF2_REG_9__SCAN_IN), .B(BUF1_REG_9__SCAN_IN), .S(n17185), .Z(n16454) );
  NAND2_X1 U17254 ( .A1(n13783), .A2(n16454), .ZN(n13787) );
  NAND2_X1 U17255 ( .A1(n13781), .A2(n13787), .ZN(P2_U2976) );
  AOI22_X1 U17256 ( .A1(n13801), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n13794), .ZN(n13784) );
  INV_X1 U17257 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19452) );
  NAND2_X1 U17258 ( .A1(n17185), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U17259 ( .B1(n17185), .B2(n19452), .A(n13782), .ZN(n20284) );
  NAND2_X1 U17260 ( .A1(n13783), .A2(n20284), .ZN(n13789) );
  NAND2_X1 U17261 ( .A1(n13784), .A2(n13789), .ZN(P2_U2974) );
  AOI22_X1 U17262 ( .A1(n13801), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13794), .ZN(n13786) );
  NAND2_X1 U17263 ( .A1(n13786), .A2(n13785), .ZN(P2_U2980) );
  AOI22_X1 U17264 ( .A1(n13801), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13791), .ZN(n13788) );
  NAND2_X1 U17265 ( .A1(n13788), .A2(n13787), .ZN(P2_U2961) );
  AOI22_X1 U17266 ( .A1(n13801), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n13791), .ZN(n13790) );
  NAND2_X1 U17267 ( .A1(n13790), .A2(n13789), .ZN(P2_U2959) );
  AOI22_X1 U17268 ( .A1(n13801), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n13791), .ZN(n13793) );
  NAND2_X1 U17269 ( .A1(n13793), .A2(n13792), .ZN(P2_U2960) );
  AOI22_X1 U17270 ( .A1(n13801), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n13794), .ZN(n13796) );
  NAND2_X1 U17271 ( .A1(n13796), .A2(n13795), .ZN(P2_U2957) );
  AOI22_X1 U17272 ( .A1(n13801), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13794), .ZN(n13798) );
  NAND2_X1 U17273 ( .A1(n13798), .A2(n13797), .ZN(P2_U2963) );
  AOI22_X1 U17274 ( .A1(n13801), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n13794), .ZN(n13800) );
  NAND2_X1 U17275 ( .A1(n13800), .A2(n13799), .ZN(P2_U2953) );
  AOI22_X1 U17276 ( .A1(n13801), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n13794), .ZN(n13803) );
  NAND2_X1 U17277 ( .A1(n13803), .A2(n13802), .ZN(P2_U2955) );
  NOR2_X1 U17278 ( .A1(n13804), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13806) );
  OAI211_X1 U17279 ( .C1(n15559), .C2(n13807), .A(n13806), .B(n13805), .ZN(
        n13809) );
  NAND2_X1 U17280 ( .A1(n13809), .A2(n13808), .ZN(n13822) );
  OAI21_X1 U17281 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17600), .A(
        n21129), .ZN(n21144) );
  INV_X1 U17282 ( .A(n15434), .ZN(n15362) );
  NAND3_X1 U17283 ( .A1(n15342), .A2(n17600), .A3(n12748), .ZN(n13810) );
  OAI21_X1 U17284 ( .B1(n21144), .B2(n15362), .A(n13810), .ZN(n13816) );
  INV_X2 U17285 ( .A(n17622), .ZN(n21142) );
  INV_X1 U17286 ( .A(n13811), .ZN(n13813) );
  OR2_X1 U17287 ( .A1(n14580), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13812) );
  AND2_X1 U17288 ( .A1(n13813), .A2(n13812), .ZN(n14910) );
  INV_X1 U17289 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13814) );
  NOR2_X1 U17290 ( .A1(n15176), .A2(n13814), .ZN(n13826) );
  AOI21_X1 U17291 ( .B1(n21142), .B2(n14910), .A(n13826), .ZN(n13815) );
  OAI211_X1 U17292 ( .C1(n13822), .C2(n15482), .A(n13816), .B(n13815), .ZN(
        P1_U3031) );
  INV_X1 U17293 ( .A(n14910), .ZN(n13821) );
  OAI21_X1 U17294 ( .B1(n13819), .B2(n13818), .A(n13817), .ZN(n13820) );
  INV_X1 U17295 ( .A(n13820), .ZN(n14917) );
  OAI222_X1 U17296 ( .A1(n13821), .A2(n14960), .B1(n12630), .B2(n21035), .C1(
        n14963), .C2(n14917), .ZN(P1_U2872) );
  INV_X1 U17297 ( .A(n13822), .ZN(n13827) );
  INV_X1 U17298 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13823) );
  AOI21_X1 U17299 ( .B1(n15249), .B2(n13824), .A(n13823), .ZN(n13825) );
  AOI211_X1 U17300 ( .C1(n13827), .C2(n21102), .A(n13826), .B(n13825), .ZN(
        n13828) );
  OAI21_X1 U17301 ( .B1(n14917), .B2(n15264), .A(n13828), .ZN(P1_U2999) );
  OAI21_X1 U17302 ( .B1(n17543), .B2(n13829), .A(n12603), .ZN(n13830) );
  AOI21_X1 U17303 ( .B1(n13831), .B2(n13830), .A(n21467), .ZN(n13832) );
  MUX2_X1 U17304 ( .A(n13832), .B(n14220), .S(n17532), .Z(n13837) );
  NOR2_X1 U17305 ( .A1(n14885), .A2(n14309), .ZN(n13833) );
  OR2_X1 U17306 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  OR3_X1 U17307 ( .A1(n13837), .A2(n13836), .A3(n13835), .ZN(n14246) );
  INV_X1 U17308 ( .A(n14246), .ZN(n17501) );
  INV_X1 U17309 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20933) );
  NAND2_X1 U17310 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17632), .ZN(n17635) );
  OAI22_X1 U17311 ( .A1(n17501), .A2(n20927), .B1(n20933), .B2(n17635), .ZN(
        n13840) );
  AOI21_X1 U17312 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21369), .A(n13840), 
        .ZN(n15524) );
  INV_X1 U17313 ( .A(n15524), .ZN(n15516) );
  INV_X1 U17314 ( .A(n14392), .ZN(n14292) );
  XNOR2_X1 U17315 ( .A(n13838), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20994) );
  INV_X1 U17316 ( .A(n13849), .ZN(n13839) );
  AND2_X1 U17317 ( .A1(n20994), .A2(n13839), .ZN(n14247) );
  NAND3_X1 U17318 ( .A1(n14247), .A2(n15504), .A3(n13840), .ZN(n13841) );
  OAI21_X1 U17319 ( .B1(n11850), .B2(n15516), .A(n13841), .ZN(P1_U3468) );
  INV_X1 U17320 ( .A(n12603), .ZN(n13845) );
  INV_X1 U17321 ( .A(n13842), .ZN(n13844) );
  NAND3_X1 U17322 ( .A1(n13845), .A2(n13844), .A3(n13843), .ZN(n13846) );
  NOR2_X1 U17323 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  AND2_X1 U17324 ( .A1(n13849), .A2(n13848), .ZN(n14242) );
  INV_X1 U17325 ( .A(n14242), .ZN(n15503) );
  NOR2_X1 U17326 ( .A1(n15500), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13850) );
  AOI21_X1 U17327 ( .B1(n14290), .B2(n15503), .A(n13850), .ZN(n17500) );
  OAI21_X1 U17328 ( .B1(n17500), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n13625), 
        .ZN(n13852) );
  NOR2_X1 U17329 ( .A1(n13625), .A2(n12748), .ZN(n15506) );
  INV_X1 U17330 ( .A(n15506), .ZN(n15513) );
  INV_X1 U17331 ( .A(n15520), .ZN(n15508) );
  AOI22_X1 U17332 ( .A1(n13852), .A2(n15513), .B1(n15508), .B2(n12356), .ZN(
        n13854) );
  NOR2_X1 U17333 ( .A1(n15501), .A2(n12356), .ZN(n17498) );
  AOI22_X1 U17334 ( .A1(n17498), .A2(n15504), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15524), .ZN(n13853) );
  OAI21_X1 U17335 ( .B1(n13854), .B2(n15524), .A(n13853), .ZN(P1_U3474) );
  AOI22_X1 U17336 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13858) );
  AOI22_X1 U17337 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U17338 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17339 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13855) );
  NAND4_X1 U17340 ( .A1(n13858), .A2(n13857), .A3(n13856), .A4(n13855), .ZN(
        n13866) );
  AOI22_X1 U17341 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17342 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13863) );
  INV_X2 U17343 ( .A(n17436), .ZN(n18324) );
  AOI22_X1 U17344 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U17345 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13861) );
  NAND4_X1 U17346 ( .A1(n13864), .A2(n13863), .A3(n13862), .A4(n13861), .ZN(
        n13865) );
  AOI22_X1 U17347 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17348 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U17349 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U17350 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U17351 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13878) );
  AOI22_X1 U17352 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17353 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U17354 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17355 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13873) );
  NAND4_X1 U17356 ( .A1(n13876), .A2(n13875), .A3(n13874), .A4(n13873), .ZN(
        n13877) );
  AOI22_X1 U17357 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17358 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17359 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17360 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17361 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U17362 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17363 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U17364 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13883) );
  INV_X1 U17365 ( .A(n13996), .ZN(n14090) );
  AOI22_X1 U17366 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U17367 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U17368 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13860), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U17369 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U17370 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17371 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13893) );
  AOI22_X1 U17372 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13892) );
  AOI22_X1 U17373 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13891) );
  AOI22_X1 U17374 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17375 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17376 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17377 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13895) );
  NAND4_X1 U17378 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        n13904) );
  AOI22_X1 U17379 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17380 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9599), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17381 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17382 ( .A1(n18427), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13899) );
  NAND4_X1 U17383 ( .A1(n13902), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13903) );
  AOI22_X1 U17384 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17385 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17386 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17387 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13906) );
  NAND4_X1 U17388 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13915) );
  AOI22_X1 U17389 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17390 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17391 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17392 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13910) );
  NAND4_X1 U17393 ( .A1(n13913), .A2(n13912), .A3(n13911), .A4(n13910), .ZN(
        n13914) );
  INV_X1 U17394 ( .A(n14006), .ZN(n18606) );
  AOI22_X1 U17395 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17396 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17397 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13917) );
  AOI22_X1 U17398 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13916) );
  NAND4_X1 U17399 ( .A1(n13919), .A2(n13918), .A3(n13917), .A4(n13916), .ZN(
        n13926) );
  AOI22_X1 U17400 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13924) );
  AOI22_X1 U17401 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U17402 ( .A1(n13069), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U17403 ( .A1(n13860), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13921) );
  NAND4_X1 U17404 ( .A1(n13924), .A2(n13923), .A3(n13922), .A4(n13921), .ZN(
        n13925) );
  NAND2_X1 U17405 ( .A1(n13940), .A2(n14017), .ZN(n13938) );
  AOI22_X1 U17406 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17407 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17408 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17409 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13927) );
  NAND4_X1 U17410 ( .A1(n13930), .A2(n13929), .A3(n13928), .A4(n13927), .ZN(
        n13936) );
  AOI22_X1 U17411 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17412 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17413 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13932) );
  AOI22_X1 U17414 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13931) );
  NAND4_X1 U17415 ( .A1(n13934), .A2(n13933), .A3(n13932), .A4(n13931), .ZN(
        n13935) );
  NAND2_X1 U17416 ( .A1(n13937), .A2(n14024), .ZN(n17332) );
  XNOR2_X1 U17417 ( .A(n17386), .B(n17332), .ZN(n17337) );
  XOR2_X1 U17418 ( .A(n13937), .B(n14024), .Z(n13953) );
  XNOR2_X1 U17419 ( .A(n18598), .B(n13938), .ZN(n13939) );
  XOR2_X1 U17420 ( .A(n19346), .B(n13939), .Z(n19037) );
  XOR2_X1 U17421 ( .A(n13940), .B(n14017), .Z(n13950) );
  OR2_X1 U17422 ( .A1(n19367), .A2(n13941), .ZN(n13948) );
  XOR2_X1 U17423 ( .A(n19367), .B(n13941), .Z(n19065) );
  NAND2_X1 U17424 ( .A1(n18611), .A2(n13996), .ZN(n14005) );
  OAI21_X1 U17425 ( .B1(n14005), .B2(n19094), .A(n13942), .ZN(n13946) );
  NAND2_X1 U17426 ( .A1(n13946), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13947) );
  AOI21_X1 U17427 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18611), .A(
        n13905), .ZN(n13944) );
  INV_X1 U17428 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19396) );
  NOR2_X1 U17429 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18611), .ZN(
        n13943) );
  AOI221_X1 U17430 ( .B1(n13905), .B2(n18611), .C1(n13944), .C2(n19396), .A(
        n13943), .ZN(n19074) );
  INV_X1 U17431 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13945) );
  XNOR2_X1 U17432 ( .A(n13946), .B(n13945), .ZN(n19073) );
  NAND2_X1 U17433 ( .A1(n19074), .A2(n19073), .ZN(n19075) );
  NAND2_X1 U17434 ( .A1(n13947), .A2(n19075), .ZN(n19064) );
  NAND2_X1 U17435 ( .A1(n19065), .A2(n19064), .ZN(n19063) );
  NAND2_X1 U17436 ( .A1(n13950), .A2(n13949), .ZN(n13951) );
  NAND2_X1 U17437 ( .A1(n13953), .A2(n13954), .ZN(n13955) );
  AOI21_X1 U17438 ( .B1(n17337), .B2(n17336), .A(n17334), .ZN(n13956) );
  XOR2_X1 U17439 ( .A(n13956), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19021) );
  INV_X1 U17440 ( .A(n19021), .ZN(n14032) );
  NAND2_X1 U17441 ( .A1(n13958), .A2(n13957), .ZN(n20041) );
  NOR2_X1 U17442 ( .A1(n19442), .A2(n18476), .ZN(n14067) );
  NAND3_X1 U17443 ( .A1(n13963), .A2(n13972), .A3(n14067), .ZN(n14060) );
  NAND2_X2 U17444 ( .A1(n13964), .A2(n13959), .ZN(n19224) );
  NAND2_X1 U17445 ( .A1(n14057), .A2(n13960), .ZN(n13962) );
  OAI21_X1 U17446 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n14070) );
  AOI21_X2 U17447 ( .B1(n14069), .B2(n13964), .A(n14070), .ZN(n19314) );
  INV_X1 U17448 ( .A(n13965), .ZN(n13966) );
  NAND2_X1 U17449 ( .A1(n13967), .A2(n13966), .ZN(n13970) );
  AOI211_X1 U17450 ( .C1(n17806), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        n14063) );
  XNOR2_X1 U17451 ( .A(n19430), .B(n13985), .ZN(n13995) );
  OAI21_X1 U17452 ( .B1(n20027), .B2(n13995), .A(n20023), .ZN(n17813) );
  OR3_X1 U17453 ( .A1(n13972), .A2(n13971), .A3(n17813), .ZN(n13989) );
  AND2_X1 U17454 ( .A1(n14104), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13973) );
  NOR2_X1 U17455 ( .A1(n13974), .A2(n13973), .ZN(n13982) );
  AND2_X1 U17456 ( .A1(n13982), .A2(n13975), .ZN(n13978) );
  NAND2_X1 U17457 ( .A1(n13977), .A2(n13976), .ZN(n13983) );
  AOI21_X1 U17458 ( .B1(n19442), .B2(n13980), .A(n19879), .ZN(n13981) );
  INV_X1 U17459 ( .A(n13981), .ZN(n13988) );
  NAND2_X1 U17460 ( .A1(n13983), .A2(n13982), .ZN(n13984) );
  NOR3_X1 U17461 ( .A1(n19430), .A2(n19449), .A3(n13985), .ZN(n13986) );
  NAND2_X1 U17462 ( .A1(n19873), .A2(n13986), .ZN(n13987) );
  NAND4_X1 U17463 ( .A1(n14063), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13990) );
  AND2_X1 U17464 ( .A1(n19878), .A2(n19397), .ZN(n19389) );
  INV_X1 U17465 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17333) );
  INV_X1 U17466 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19337) );
  NOR2_X1 U17467 ( .A1(n17333), .A2(n19337), .ZN(n13992) );
  INV_X1 U17468 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19354) );
  INV_X1 U17469 ( .A(n19314), .ZN(n19277) );
  NOR2_X1 U17470 ( .A1(n19224), .A2(n19277), .ZN(n19369) );
  INV_X1 U17471 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17358) );
  NOR2_X1 U17472 ( .A1(n13945), .A2(n17358), .ZN(n13993) );
  OAI21_X1 U17473 ( .B1(n19396), .B2(n17358), .A(n13945), .ZN(n19376) );
  INV_X1 U17474 ( .A(n19376), .ZN(n17360) );
  NOR2_X1 U17475 ( .A1(n19314), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19371) );
  AOI211_X1 U17476 ( .C1(n19880), .C2(n17360), .A(n19371), .B(n19367), .ZN(
        n13991) );
  OAI21_X1 U17477 ( .B1(n19369), .B2(n13993), .A(n13991), .ZN(n19364) );
  NOR3_X1 U17478 ( .A1(n19346), .A2(n19354), .A3(n19364), .ZN(n19333) );
  OR2_X1 U17479 ( .A1(n19227), .A2(n19390), .ZN(n19385) );
  AOI21_X1 U17480 ( .B1(n13992), .B2(n19333), .A(n19385), .ZN(n19327) );
  AOI21_X1 U17481 ( .B1(n19277), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n19224), .ZN(n17364) );
  INV_X1 U17482 ( .A(n17364), .ZN(n19372) );
  AOI22_X1 U17483 ( .A1(n19880), .A2(n19376), .B1(n19372), .B2(n13993), .ZN(
        n19359) );
  NOR3_X1 U17484 ( .A1(n19346), .A2(n19367), .A3(n19354), .ZN(n19338) );
  NAND2_X1 U17485 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19338), .ZN(
        n13994) );
  OAI21_X1 U17486 ( .B1(n19359), .B2(n13994), .A(n17333), .ZN(n14030) );
  NAND2_X2 U17487 ( .A1(n19227), .A2(n13995), .ZN(n19875) );
  INV_X1 U17488 ( .A(n18611), .ZN(n13997) );
  NAND2_X1 U17489 ( .A1(n13997), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13998) );
  INV_X1 U17490 ( .A(n13999), .ZN(n14000) );
  NAND2_X1 U17491 ( .A1(n14000), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14001) );
  NAND2_X1 U17492 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  XNOR2_X1 U17493 ( .A(n14005), .B(n14006), .ZN(n19066) );
  NAND2_X1 U17494 ( .A1(n14003), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14004) );
  INV_X1 U17495 ( .A(n14005), .ZN(n14007) );
  NAND2_X1 U17496 ( .A1(n14007), .A2(n14006), .ZN(n14011) );
  INV_X1 U17497 ( .A(n14017), .ZN(n18601) );
  XNOR2_X1 U17498 ( .A(n14011), .B(n18601), .ZN(n19053) );
  INV_X1 U17499 ( .A(n19053), .ZN(n14008) );
  NAND2_X1 U17500 ( .A1(n14008), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14009) );
  NAND2_X1 U17501 ( .A1(n14010), .A2(n14009), .ZN(n19042) );
  NAND2_X1 U17502 ( .A1(n14019), .A2(n14017), .ZN(n14012) );
  XNOR2_X1 U17503 ( .A(n14012), .B(n18598), .ZN(n19040) );
  NAND2_X1 U17504 ( .A1(n19040), .A2(n19346), .ZN(n14013) );
  INV_X1 U17505 ( .A(n19040), .ZN(n14014) );
  NAND2_X1 U17506 ( .A1(n14014), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14015) );
  XNOR2_X1 U17507 ( .A(n14023), .B(n18594), .ZN(n14020) );
  XNOR2_X1 U17508 ( .A(n14020), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19028) );
  INV_X1 U17509 ( .A(n14020), .ZN(n14021) );
  NAND2_X1 U17510 ( .A1(n14021), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14022) );
  OAI21_X1 U17511 ( .B1(n14023), .B2(n18594), .A(n18591), .ZN(n14027) );
  NAND2_X1 U17512 ( .A1(n14027), .A2(n19006), .ZN(n17297) );
  XNOR2_X1 U17513 ( .A(n17296), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19018) );
  AOI22_X1 U17514 ( .A1(n19392), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19402), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n14028) );
  OAI21_X1 U17515 ( .B1(n19404), .B2(n19018), .A(n14028), .ZN(n14029) );
  AOI21_X1 U17516 ( .B1(n19327), .B2(n14030), .A(n14029), .ZN(n14031) );
  OAI21_X1 U17517 ( .B1(n14032), .B2(n19406), .A(n14031), .ZN(P3_U2855) );
  NAND2_X1 U17518 ( .A1(n14036), .A2(n14035), .ZN(n14037) );
  MUX2_X1 U17519 ( .A(n17649), .B(n16255), .S(n16418), .Z(n14038) );
  OAI21_X1 U17520 ( .B1(n17184), .B2(n20101), .A(n14038), .ZN(P2_U2884) );
  NAND3_X1 U17521 ( .A1(n20876), .A2(n17668), .A3(n17149), .ZN(n14055) );
  INV_X1 U17522 ( .A(n17127), .ZN(n17167) );
  NAND2_X1 U17523 ( .A1(n9615), .A2(n17167), .ZN(n14053) );
  NAND2_X1 U17524 ( .A1(n14040), .A2(n11260), .ZN(n17156) );
  OAI21_X1 U17525 ( .B1(n17154), .B2(n14056), .A(n14041), .ZN(n14051) );
  NAND2_X1 U17526 ( .A1(n14043), .A2(n14042), .ZN(n17163) );
  NOR2_X1 U17527 ( .A1(n14044), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17155) );
  INV_X1 U17528 ( .A(n17155), .ZN(n14045) );
  XNOR2_X1 U17529 ( .A(n14045), .B(n14056), .ZN(n14046) );
  NAND2_X1 U17530 ( .A1(n17163), .A2(n14046), .ZN(n14049) );
  OAI211_X1 U17531 ( .C1(n10694), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17161), .B(n14047), .ZN(n14048) );
  NAND2_X1 U17532 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  AOI21_X1 U17533 ( .B1(n17156), .B2(n14051), .A(n14050), .ZN(n14052) );
  NAND2_X1 U17534 ( .A1(n14053), .A2(n14052), .ZN(n17249) );
  NAND2_X1 U17535 ( .A1(n17249), .A2(n17169), .ZN(n14054) );
  OAI211_X1 U17536 ( .C1(n17149), .C2(n14056), .A(n14055), .B(n14054), .ZN(
        P2_U3596) );
  NAND2_X1 U17537 ( .A1(n19876), .A2(n20023), .ZN(n14064) );
  NAND2_X1 U17538 ( .A1(n19430), .A2(n17814), .ZN(n19899) );
  INV_X1 U17539 ( .A(n19899), .ZN(n14061) );
  OAI21_X1 U17540 ( .B1(n14064), .B2(n18619), .A(n14063), .ZN(n14065) );
  NOR3_X1 U17541 ( .A1(n14087), .A2(n14085), .A3(n14065), .ZN(n19894) );
  INV_X1 U17542 ( .A(n19894), .ZN(n19884) );
  NOR2_X1 U17543 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20009), .ZN(n19425) );
  INV_X1 U17544 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19408) );
  NAND3_X1 U17545 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n20007)
         );
  NOR2_X1 U17546 ( .A1(n19408), .A2(n20007), .ZN(n14066) );
  INV_X1 U17547 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17368) );
  OAI22_X1 U17548 ( .A1(n17368), .A2(n17358), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14138) );
  INV_X1 U17549 ( .A(n14138), .ZN(n14075) );
  NOR2_X1 U17550 ( .A1(n19895), .A2(n19396), .ZN(n14137) );
  NOR2_X1 U17551 ( .A1(n14132), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14118) );
  INV_X1 U17552 ( .A(n14118), .ZN(n14121) );
  NAND2_X1 U17553 ( .A1(n14119), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14126) );
  NAND2_X1 U17554 ( .A1(n14121), .A2(n14126), .ZN(n18160) );
  OAI21_X1 U17555 ( .B1(n19314), .B2(n14104), .A(n19398), .ZN(n14120) );
  INV_X1 U17556 ( .A(n14120), .ZN(n14136) );
  NOR2_X1 U17557 ( .A1(n14136), .A2(n14143), .ZN(n14072) );
  AOI21_X1 U17558 ( .B1(n14067), .B2(n14069), .A(n14070), .ZN(n14068) );
  OR2_X1 U17559 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14068), .ZN(
        n14116) );
  NOR3_X1 U17560 ( .A1(n14070), .A2(n14069), .A3(n19224), .ZN(n14117) );
  AOI21_X1 U17561 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14116), .A(
        n14117), .ZN(n14071) );
  MUX2_X1 U17562 ( .A(n14072), .B(n14071), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n14073) );
  AOI21_X1 U17563 ( .B1(n19880), .B2(n18160), .A(n14073), .ZN(n19863) );
  INV_X1 U17564 ( .A(n20040), .ZN(n14522) );
  INV_X1 U17565 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U17566 ( .A1(n14519), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n14526) );
  OAI22_X1 U17567 ( .A1(n19863), .A2(n14522), .B1(n14526), .B2(n18160), .ZN(
        n14074) );
  AOI21_X1 U17568 ( .B1(n14075), .B2(n14137), .A(n14074), .ZN(n14076) );
  INV_X1 U17569 ( .A(n14523), .ZN(n14139) );
  AOI22_X1 U17570 ( .A1(n14523), .A2(n14077), .B1(n14076), .B2(n14139), .ZN(
        P3_U3288) );
  OAI21_X1 U17571 ( .B1(n14079), .B2(n14078), .A(n14198), .ZN(n14909) );
  INV_X1 U17572 ( .A(n14909), .ZN(n14114) );
  XNOR2_X1 U17573 ( .A(n14907), .B(n14579), .ZN(n21139) );
  OAI22_X1 U17574 ( .A1(n14960), .A2(n21139), .B1(n14899), .B2(n21035), .ZN(
        n14080) );
  AOI21_X1 U17575 ( .B1(n14114), .B2(n21031), .A(n14080), .ZN(n14081) );
  INV_X1 U17576 ( .A(n14081), .ZN(P1_U2871) );
  NAND2_X1 U17577 ( .A1(n11662), .A2(n14317), .ZN(n14082) );
  MUX2_X1 U17578 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n14974), .Z(
        n15007) );
  INV_X1 U17579 ( .A(n15007), .ZN(n14303) );
  INV_X1 U17580 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21070) );
  OAI222_X1 U17581 ( .A1(n15033), .A2(n14303), .B1(n15031), .B2(n14917), .C1(
        n21070), .C2(n15029), .ZN(P1_U2904) );
  INV_X1 U17582 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21066) );
  MUX2_X1 U17583 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n14974), .Z(
        n15001) );
  INV_X1 U17584 ( .A(n15001), .ZN(n14313) );
  OAI222_X1 U17585 ( .A1(n14909), .A2(n15031), .B1(n15029), .B2(n21066), .C1(
        n15033), .C2(n14313), .ZN(P1_U2903) );
  NAND2_X1 U17586 ( .A1(n14088), .A2(n9967), .ZN(n18610) );
  AND2_X1 U17587 ( .A1(n18518), .A2(n9967), .ZN(n18576) );
  NAND3_X1 U17588 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(n9967), .ZN(n18614) );
  NOR2_X1 U17589 ( .A1(n18518), .A2(n18614), .ZN(n14089) );
  AOI21_X1 U17590 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18615), .A(n14089), .ZN(
        n14091) );
  NAND2_X1 U17591 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n14089), .ZN(n18604) );
  INV_X1 U17592 ( .A(n18604), .ZN(n18605) );
  OAI222_X1 U17593 ( .A1(n19433), .A2(n18610), .B1(n14091), .B2(n18605), .C1(
        n18607), .C2(n14090), .ZN(P3_U2733) );
  NOR2_X1 U17594 ( .A1(n14094), .A2(n14093), .ZN(n16220) );
  XNOR2_X1 U17595 ( .A(n16217), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14102) );
  AND2_X1 U17596 ( .A1(n14097), .A2(n14098), .ZN(n14099) );
  NOR2_X1 U17597 ( .A1(n14096), .A2(n14099), .ZN(n17640) );
  NOR2_X1 U17598 ( .A1(n20112), .A2(n10961), .ZN(n14100) );
  AOI21_X1 U17599 ( .B1(n17640), .B2(n20112), .A(n14100), .ZN(n14101) );
  OAI21_X1 U17600 ( .B1(n14102), .B2(n20101), .A(n14101), .ZN(P2_U2882) );
  INV_X1 U17601 ( .A(n14526), .ZN(n19896) );
  NAND2_X1 U17602 ( .A1(n19896), .A2(n14104), .ZN(n14108) );
  NOR2_X1 U17603 ( .A1(n14103), .A2(n19277), .ZN(n14135) );
  MUX2_X1 U17604 ( .A(n19398), .B(n14135), .S(n14104), .Z(n19865) );
  NAND2_X1 U17605 ( .A1(n19396), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n14105) );
  OAI211_X1 U17606 ( .C1(n19865), .C2(n14522), .A(n14139), .B(n14105), .ZN(
        n14106) );
  OAI21_X1 U17607 ( .B1(n14139), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n14106), .ZN(n14107) );
  OAI21_X1 U17608 ( .B1(n14523), .B2(n14108), .A(n14107), .ZN(P3_U3290) );
  OAI21_X1 U17609 ( .B1(n14110), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14109), .ZN(n21143) );
  INV_X1 U17610 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14111) );
  NOR2_X1 U17611 ( .A1(n15176), .A2(n14111), .ZN(n21140) );
  AOI21_X1 U17612 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n21140), .ZN(n14112) );
  OAI21_X1 U17613 ( .B1(n21106), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14112), .ZN(n14113) );
  AOI21_X1 U17614 ( .B1(n14114), .B2(n21101), .A(n14113), .ZN(n14115) );
  OAI21_X1 U17615 ( .B1(n20932), .B2(n21143), .A(n14115), .ZN(P1_U2998) );
  OAI211_X1 U17616 ( .C1(n14117), .C2(n14119), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14116), .ZN(n14122) );
  NOR2_X1 U17617 ( .A1(n14122), .A2(n14118), .ZN(n14125) );
  AOI21_X1 U17618 ( .B1(n14120), .B2(n14119), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14124) );
  NAND3_X1 U17619 ( .A1(n14122), .A2(n19880), .A3(n14121), .ZN(n14123) );
  OAI21_X1 U17620 ( .B1(n14125), .B2(n14124), .A(n14123), .ZN(n19885) );
  NAND2_X1 U17621 ( .A1(n14126), .A2(n14130), .ZN(n14127) );
  NAND2_X1 U17622 ( .A1(n17438), .A2(n14127), .ZN(n18146) );
  OAI21_X1 U17623 ( .B1(n14526), .B2(n18146), .A(n14139), .ZN(n14128) );
  AOI21_X1 U17624 ( .B1(n19885), .B2(n20040), .A(n14128), .ZN(n14129) );
  AOI21_X1 U17625 ( .B1(n14523), .B2(n14130), .A(n14129), .ZN(P3_U3285) );
  INV_X1 U17626 ( .A(n14131), .ZN(n14134) );
  INV_X1 U17627 ( .A(n14132), .ZN(n14133) );
  NAND2_X1 U17628 ( .A1(n14134), .A2(n14133), .ZN(n18178) );
  OAI22_X1 U17629 ( .A1(n14136), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14135), .B2(n18178), .ZN(n19869) );
  NAND2_X1 U17630 ( .A1(n14138), .A2(n14137), .ZN(n14140) );
  OAI211_X1 U17631 ( .C1(n18178), .C2(n14526), .A(n14140), .B(n14139), .ZN(
        n14141) );
  AOI21_X1 U17632 ( .B1(n19869), .B2(n20040), .A(n14141), .ZN(n14142) );
  AOI21_X1 U17633 ( .B1(n14523), .B2(n14143), .A(n14142), .ZN(P3_U3289) );
  AOI22_X1 U17634 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14144) );
  OAI21_X1 U17635 ( .B1(n12227), .B2(n14163), .A(n14144), .ZN(P1_U2912) );
  INV_X1 U17636 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U17637 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14145) );
  OAI21_X1 U17638 ( .B1(n14146), .B2(n14163), .A(n14145), .ZN(P1_U2916) );
  INV_X1 U17639 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U17640 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17641 ( .B1(n14148), .B2(n14163), .A(n14147), .ZN(P1_U2915) );
  INV_X1 U17642 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U17643 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U17644 ( .B1(n14150), .B2(n14163), .A(n14149), .ZN(P1_U2913) );
  INV_X1 U17645 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14152) );
  AOI22_X1 U17646 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U17647 ( .B1(n14152), .B2(n14163), .A(n14151), .ZN(P1_U2918) );
  INV_X1 U17648 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17649 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14153) );
  OAI21_X1 U17650 ( .B1(n14154), .B2(n14163), .A(n14153), .ZN(P1_U2917) );
  INV_X1 U17651 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U17652 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14155) );
  OAI21_X1 U17653 ( .B1(n14156), .B2(n14163), .A(n14155), .ZN(P1_U2919) );
  INV_X1 U17654 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17655 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14157) );
  OAI21_X1 U17656 ( .B1(n14158), .B2(n14163), .A(n14157), .ZN(P1_U2920) );
  AOI22_X1 U17657 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14159) );
  OAI21_X1 U17658 ( .B1(n12345), .B2(n14163), .A(n14159), .ZN(P1_U2906) );
  INV_X1 U17659 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U17660 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14160) );
  OAI21_X1 U17661 ( .B1(n14161), .B2(n14163), .A(n14160), .ZN(P1_U2914) );
  INV_X1 U17662 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U17663 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14162) );
  OAI21_X1 U17664 ( .B1(n14164), .B2(n14163), .A(n14162), .ZN(P1_U2909) );
  INV_X1 U17665 ( .A(n20113), .ZN(n14171) );
  OAI21_X1 U17666 ( .B1(n14167), .B2(n14166), .A(n11316), .ZN(n17656) );
  INV_X1 U17667 ( .A(n17656), .ZN(n16293) );
  NOR2_X1 U17668 ( .A1(n17220), .A2(n17656), .ZN(n14189) );
  INV_X1 U17669 ( .A(n14189), .ZN(n14168) );
  OAI211_X1 U17670 ( .C1(n17219), .C2(n16293), .A(n14168), .B(n20128), .ZN(
        n14170) );
  AOI22_X1 U17671 ( .A1(n20134), .A2(n16293), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n20133), .ZN(n14169) );
  OAI211_X1 U17672 ( .C1(n20142), .C2(n14171), .A(n14170), .B(n14169), .ZN(
        P2_U2919) );
  OR2_X1 U17673 ( .A1(n14173), .A2(n14172), .ZN(n14174) );
  NAND2_X1 U17674 ( .A1(n14175), .A2(n14174), .ZN(n14183) );
  XOR2_X1 U17675 ( .A(n14183), .B(n20889), .Z(n14182) );
  OAI21_X1 U17676 ( .B1(n14178), .B2(n14177), .A(n14176), .ZN(n20237) );
  INV_X1 U17677 ( .A(n20237), .ZN(n16284) );
  NAND2_X1 U17678 ( .A1(n20251), .A2(n16284), .ZN(n14179) );
  OAI21_X1 U17679 ( .B1(n20251), .B2(n16284), .A(n14179), .ZN(n14188) );
  NOR2_X1 U17680 ( .A1(n14188), .A2(n14189), .ZN(n14187) );
  INV_X1 U17681 ( .A(n14179), .ZN(n14180) );
  NOR2_X1 U17682 ( .A1(n14187), .A2(n14180), .ZN(n14181) );
  NOR2_X1 U17683 ( .A1(n14181), .A2(n14182), .ZN(n16519) );
  AOI21_X1 U17684 ( .B1(n14182), .B2(n14181), .A(n16519), .ZN(n14186) );
  INV_X1 U17685 ( .A(n14183), .ZN(n20887) );
  INV_X1 U17686 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20172) );
  OAI22_X1 U17687 ( .A1(n16517), .A2(n20887), .B1(n16495), .B2(n20172), .ZN(
        n14184) );
  AOI21_X1 U17688 ( .B1(n17238), .B2(n16522), .A(n14184), .ZN(n14185) );
  OAI21_X1 U17689 ( .B1(n14186), .B2(n20138), .A(n14185), .ZN(P2_U2917) );
  AOI21_X1 U17690 ( .B1(n14189), .B2(n14188), .A(n14187), .ZN(n14192) );
  INV_X1 U17691 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20174) );
  OAI22_X1 U17692 ( .A1(n16517), .A2(n16284), .B1(n16495), .B2(n20174), .ZN(
        n14190) );
  AOI21_X1 U17693 ( .B1(n16522), .B2(n16510), .A(n14190), .ZN(n14191) );
  OAI21_X1 U17694 ( .B1(n14192), .B2(n20138), .A(n14191), .ZN(P2_U2918) );
  OAI21_X1 U17695 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n21128) );
  INV_X1 U17696 ( .A(n14196), .ZN(n14197) );
  AOI21_X1 U17697 ( .B1(n14199), .B2(n14198), .A(n14197), .ZN(n21025) );
  AOI22_X1 U17698 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21133), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14200) );
  OAI21_X1 U17699 ( .B1(n21106), .B2(n21015), .A(n14200), .ZN(n14201) );
  AOI21_X1 U17700 ( .B1(n21025), .B2(n21101), .A(n14201), .ZN(n14202) );
  OAI21_X1 U17701 ( .B1(n20932), .B2(n21128), .A(n14202), .ZN(P1_U2997) );
  XOR2_X1 U17702 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(n16414), .Z(n14207)
         );
  NOR2_X1 U17703 ( .A1(n14096), .A2(n14204), .ZN(n14205) );
  OR2_X1 U17704 ( .A1(n14203), .A2(n14205), .ZN(n20088) );
  INV_X1 U17705 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n20071) );
  MUX2_X1 U17706 ( .A(n20088), .B(n20071), .S(n16418), .Z(n14206) );
  OAI21_X1 U17707 ( .B1(n14207), .B2(n20101), .A(n14206), .ZN(P2_U2881) );
  INV_X1 U17708 ( .A(n21025), .ZN(n14211) );
  INV_X1 U17709 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21064) );
  MUX2_X1 U17710 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n14974), .Z(
        n14998) );
  INV_X1 U17711 ( .A(n14998), .ZN(n14308) );
  OAI222_X1 U17712 ( .A1(n14211), .A2(n15031), .B1(n15029), .B2(n21064), .C1(
        n15033), .C2(n14308), .ZN(P1_U2902) );
  NAND2_X1 U17713 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U17714 ( .A1(n14429), .A2(n14210), .ZN(n21012) );
  INV_X1 U17715 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14212) );
  OAI222_X1 U17716 ( .A1(n21012), .A2(n14960), .B1(n14212), .B2(n21035), .C1(
        n14211), .C2(n14963), .ZN(P1_U2870) );
  INV_X1 U17717 ( .A(n15531), .ZN(n14894) );
  MUX2_X1 U17718 ( .A(n14215), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14214), .Z(n14217) );
  NOR2_X1 U17719 ( .A1(n14217), .A2(n14216), .ZN(n14230) );
  INV_X1 U17720 ( .A(n14218), .ZN(n14219) );
  OR2_X1 U17721 ( .A1(n14220), .A2(n14219), .ZN(n14240) );
  XNOR2_X1 U17722 ( .A(n14221), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14228) );
  NOR2_X1 U17723 ( .A1(n15500), .A2(n14222), .ZN(n14236) );
  NOR2_X1 U17724 ( .A1(n14214), .A2(n11823), .ZN(n14225) );
  NOR2_X1 U17725 ( .A1(n14225), .A2(n14224), .ZN(n14226) );
  NAND2_X1 U17726 ( .A1(n11733), .A2(n14226), .ZN(n15519) );
  NAND3_X1 U17727 ( .A1(n14236), .A2(n9625), .A3(n15519), .ZN(n14227) );
  OAI21_X1 U17728 ( .B1(n15501), .B2(n14228), .A(n14227), .ZN(n14229) );
  AOI21_X1 U17729 ( .B1(n14230), .B2(n14240), .A(n14229), .ZN(n14231) );
  OAI21_X1 U17730 ( .B1(n14894), .B2(n14242), .A(n14231), .ZN(n15518) );
  MUX2_X1 U17731 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15518), .S(
        n14246), .Z(n17509) );
  NOR2_X1 U17732 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13625), .ZN(n14248) );
  AOI22_X1 U17733 ( .A1(n17509), .A2(n13625), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14248), .ZN(n14244) );
  XNOR2_X1 U17734 ( .A(n14214), .B(n14233), .ZN(n14234) );
  INV_X1 U17735 ( .A(n14234), .ZN(n15515) );
  XNOR2_X1 U17736 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14238) );
  NAND3_X1 U17737 ( .A1(n14236), .A2(n9625), .A3(n14234), .ZN(n14237) );
  OAI21_X1 U17738 ( .B1(n15501), .B2(n14238), .A(n14237), .ZN(n14239) );
  AOI21_X1 U17739 ( .B1(n14240), .B2(n15515), .A(n14239), .ZN(n14241) );
  OAI21_X1 U17740 ( .B1(n14232), .B2(n14242), .A(n14241), .ZN(n15511) );
  MUX2_X1 U17741 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15511), .S(
        n14246), .Z(n17508) );
  AOI22_X1 U17742 ( .A1(n14248), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17508), .B2(n13625), .ZN(n14243) );
  NOR2_X1 U17743 ( .A1(n14244), .A2(n14243), .ZN(n17520) );
  INV_X1 U17744 ( .A(n14245), .ZN(n15499) );
  NAND2_X1 U17745 ( .A1(n17520), .A2(n15499), .ZN(n14252) );
  MUX2_X1 U17746 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n14247), .S(
        n14246), .Z(n14250) );
  AND2_X1 U17747 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14248), .ZN(
        n14249) );
  AOI21_X1 U17748 ( .B1(n14250), .B2(n13625), .A(n14249), .ZN(n17518) );
  AND3_X1 U17749 ( .A1(n14252), .A2(n17518), .A3(n20933), .ZN(n14251) );
  AND3_X1 U17750 ( .A1(n14252), .A2(n17518), .A3(n17632), .ZN(n17529) );
  INV_X1 U17751 ( .A(n14290), .ZN(n14913) );
  NAND2_X1 U17752 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n17636), .ZN(n14340) );
  INV_X1 U17753 ( .A(n14340), .ZN(n15495) );
  OAI22_X1 U17754 ( .A1(n15559), .A2(n21311), .B1(n14913), .B2(n15495), .ZN(
        n14253) );
  OAI21_X1 U17755 ( .B1(n17529), .B2(n14253), .A(n21153), .ZN(n14254) );
  OAI21_X1 U17756 ( .B1(n21153), .B2(n21307), .A(n14254), .ZN(P1_U3478) );
  INV_X1 U17757 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n21062) );
  MUX2_X1 U17758 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n14974), .Z(
        n14994) );
  INV_X1 U17759 ( .A(n14994), .ZN(n14298) );
  OAI222_X1 U17760 ( .A1(n14898), .A2(n15031), .B1(n15029), .B2(n21062), .C1(
        n15033), .C2(n14298), .ZN(P1_U2901) );
  INV_X1 U17761 ( .A(n14431), .ZN(n14256) );
  XNOR2_X1 U17762 ( .A(n14429), .B(n14256), .ZN(n21114) );
  OAI222_X1 U17763 ( .A1(n14963), .A2(n14898), .B1(n14257), .B2(n21035), .C1(
        n14960), .C2(n21114), .ZN(P1_U2869) );
  NAND2_X1 U17764 ( .A1(n14259), .A2(n14260), .ZN(n14261) );
  AND2_X1 U17765 ( .A1(n14267), .A2(n14261), .ZN(n16998) );
  INV_X1 U17766 ( .A(n16998), .ZN(n16159) );
  AOI22_X1 U17767 ( .A1(n16522), .A2(n16447), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20133), .ZN(n14262) );
  OAI21_X1 U17768 ( .B1(n16159), .B2(n16525), .A(n14262), .ZN(P2_U2909) );
  OR2_X1 U17769 ( .A1(n14263), .A2(n14264), .ZN(n14265) );
  AND2_X1 U17770 ( .A1(n10355), .A2(n14265), .ZN(n16981) );
  INV_X1 U17771 ( .A(n16981), .ZN(n16132) );
  AOI22_X1 U17772 ( .A1(n16522), .A2(n16433), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n20133), .ZN(n14266) );
  OAI21_X1 U17773 ( .B1(n16132), .B2(n16525), .A(n14266), .ZN(P2_U2907) );
  AOI21_X1 U17774 ( .B1(n14268), .B2(n14267), .A(n14263), .ZN(n16992) );
  INV_X1 U17775 ( .A(n16992), .ZN(n14270) );
  INV_X1 U17776 ( .A(n16440), .ZN(n14269) );
  INV_X1 U17777 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20154) );
  OAI222_X1 U17778 ( .A1(n14270), .A2(n16525), .B1(n14269), .B2(n20142), .C1(
        n20154), .C2(n16495), .ZN(P2_U2908) );
  NAND2_X1 U17779 ( .A1(n14272), .A2(n14273), .ZN(n14274) );
  NAND2_X1 U17780 ( .A1(n14277), .A2(n14274), .ZN(n17023) );
  INV_X1 U17781 ( .A(n16460), .ZN(n14275) );
  INV_X1 U17782 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20160) );
  OAI222_X1 U17783 ( .A1(n17023), .A2(n16525), .B1(n14275), .B2(n20142), .C1(
        n20160), .C2(n16495), .ZN(P2_U2911) );
  NAND2_X1 U17784 ( .A1(n14277), .A2(n14276), .ZN(n14278) );
  AND2_X1 U17785 ( .A1(n14259), .A2(n14278), .ZN(n17018) );
  INV_X1 U17786 ( .A(n17018), .ZN(n14280) );
  INV_X1 U17787 ( .A(n16454), .ZN(n14279) );
  INV_X1 U17788 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20158) );
  OAI222_X1 U17789 ( .A1(n14280), .A2(n16525), .B1(n14279), .B2(n20142), .C1(
        n20158), .C2(n16495), .ZN(P2_U2910) );
  NAND2_X1 U17790 ( .A1(n10355), .A2(n14282), .ZN(n14283) );
  NAND2_X1 U17791 ( .A1(n14281), .A2(n14283), .ZN(n16967) );
  INV_X1 U17792 ( .A(n16426), .ZN(n14284) );
  INV_X1 U17793 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20150) );
  OAI222_X1 U17794 ( .A1(n16967), .A2(n16525), .B1(n14284), .B2(n20142), .C1(
        n20150), .C2(n16495), .ZN(P2_U2906) );
  NAND2_X1 U17795 ( .A1(n15603), .A2(n21285), .ZN(n14359) );
  INV_X1 U17796 ( .A(n14359), .ZN(n14286) );
  AOI21_X1 U17797 ( .B1(n15803), .B2(n14286), .A(n14289), .ZN(n14288) );
  INV_X1 U17798 ( .A(n21315), .ZN(n14287) );
  INV_X1 U17799 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14297) );
  MUX2_X1 U17800 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n14974), .Z(
        n14991) );
  INV_X1 U17801 ( .A(n14991), .ZN(n14390) );
  INV_X1 U17802 ( .A(n14289), .ZN(n15801) );
  NAND2_X1 U17803 ( .A1(n14291), .A2(n14290), .ZN(n14393) );
  OR2_X1 U17804 ( .A1(n14232), .A2(n14292), .ZN(n15763) );
  INV_X1 U17805 ( .A(n15763), .ZN(n15804) );
  NAND2_X1 U17806 ( .A1(n15804), .A2(n21285), .ZN(n21308) );
  OAI222_X1 U17807 ( .A1(n21311), .A2(n14293), .B1(n15801), .B2(n11775), .C1(
        n14393), .C2(n21308), .ZN(n14327) );
  INV_X1 U17808 ( .A(n14293), .ZN(n14326) );
  NAND2_X1 U17809 ( .A1(n14294), .A2(n14324), .ZN(n15699) );
  AOI22_X1 U17810 ( .A1(n21341), .A2(n14327), .B1(n14326), .B2(n21340), .ZN(
        n14296) );
  NAND2_X1 U17811 ( .A1(n15560), .A2(n15559), .ZN(n15562) );
  INV_X1 U17812 ( .A(n14974), .ZN(n14440) );
  AOI22_X1 U17813 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14328), .B1(DATAI_28_), 
        .B2(n14329), .ZN(n21345) );
  INV_X1 U17814 ( .A(n21345), .ZN(n21227) );
  AOI22_X1 U17815 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n14328), .B1(DATAI_20_), 
        .B2(n14329), .ZN(n21230) );
  INV_X1 U17816 ( .A(n21230), .ZN(n21342) );
  AOI22_X1 U17817 ( .A1(n15833), .A2(n21227), .B1(n21164), .B2(n21342), .ZN(
        n14295) );
  OAI211_X1 U17818 ( .C1(n14333), .C2(n14297), .A(n14296), .B(n14295), .ZN(
        P1_U3157) );
  INV_X1 U17819 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14302) );
  NAND2_X1 U17820 ( .A1(n14299), .A2(n14324), .ZN(n15695) );
  AOI22_X1 U17821 ( .A1(n21335), .A2(n14327), .B1(n14326), .B2(n21334), .ZN(
        n14301) );
  AOI22_X1 U17822 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14328), .B1(DATAI_27_), 
        .B2(n14329), .ZN(n21339) );
  INV_X1 U17823 ( .A(n21339), .ZN(n21223) );
  AOI22_X1 U17824 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n14328), .B1(DATAI_19_), 
        .B2(n14329), .ZN(n21226) );
  INV_X1 U17825 ( .A(n21226), .ZN(n21336) );
  AOI22_X1 U17826 ( .A1(n15833), .A2(n21223), .B1(n21164), .B2(n21336), .ZN(
        n14300) );
  OAI211_X1 U17827 ( .C1(n14333), .C2(n14302), .A(n14301), .B(n14300), .ZN(
        P1_U3156) );
  INV_X1 U17828 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U17829 ( .A1(n14304), .A2(n14324), .ZN(n15683) );
  AOI22_X1 U17830 ( .A1(n21314), .A2(n14327), .B1(n14326), .B2(n21313), .ZN(
        n14306) );
  AOI22_X1 U17831 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n14328), .B1(DATAI_24_), 
        .B2(n14329), .ZN(n21321) );
  INV_X1 U17832 ( .A(n21321), .ZN(n21211) );
  AOI22_X1 U17833 ( .A1(DATAI_16_), .A2(n14329), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n14328), .ZN(n21214) );
  INV_X1 U17834 ( .A(n21214), .ZN(n21318) );
  AOI22_X1 U17835 ( .A1(n15833), .A2(n21211), .B1(n21164), .B2(n21318), .ZN(
        n14305) );
  OAI211_X1 U17836 ( .C1(n14333), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        P1_U3153) );
  INV_X1 U17837 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17838 ( .A1(n14309), .A2(n14324), .ZN(n15691) );
  AOI22_X1 U17839 ( .A1(n21329), .A2(n14327), .B1(n14326), .B2(n21328), .ZN(
        n14311) );
  AOI22_X1 U17840 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14328), .B1(DATAI_26_), 
        .B2(n14329), .ZN(n21333) );
  INV_X1 U17841 ( .A(n21333), .ZN(n21219) );
  AOI22_X1 U17842 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n14328), .B1(DATAI_18_), 
        .B2(n14329), .ZN(n21222) );
  INV_X1 U17843 ( .A(n21222), .ZN(n21330) );
  AOI22_X1 U17844 ( .A1(n15833), .A2(n21219), .B1(n21164), .B2(n21330), .ZN(
        n14310) );
  OAI211_X1 U17845 ( .C1(n14333), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        P1_U3155) );
  INV_X1 U17846 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U17847 ( .A1(n14542), .A2(n14324), .ZN(n15687) );
  AOI22_X1 U17848 ( .A1(n21323), .A2(n14327), .B1(n14326), .B2(n21322), .ZN(
        n14315) );
  AOI22_X1 U17849 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14328), .B1(DATAI_25_), 
        .B2(n14329), .ZN(n21327) );
  INV_X1 U17850 ( .A(n21327), .ZN(n21215) );
  AOI22_X1 U17851 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n14328), .B1(DATAI_17_), 
        .B2(n14329), .ZN(n21218) );
  INV_X1 U17852 ( .A(n21218), .ZN(n21324) );
  AOI22_X1 U17853 ( .A1(n15833), .A2(n21215), .B1(n21164), .B2(n21324), .ZN(
        n14314) );
  OAI211_X1 U17854 ( .C1(n14333), .C2(n14316), .A(n14315), .B(n14314), .ZN(
        P1_U3154) );
  INV_X1 U17855 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14320) );
  MUX2_X1 U17856 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n14974), .Z(
        n14980) );
  INV_X1 U17857 ( .A(n14980), .ZN(n14496) );
  NAND2_X1 U17858 ( .A1(n14317), .A2(n14324), .ZN(n15712) );
  AOI22_X1 U17859 ( .A1(n21361), .A2(n14327), .B1(n14326), .B2(n21359), .ZN(
        n14319) );
  AOI22_X1 U17860 ( .A1(DATAI_31_), .A2(n14329), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n14328), .ZN(n21368) );
  INV_X1 U17861 ( .A(n21368), .ZN(n21241) );
  AOI22_X1 U17862 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n14328), .B1(DATAI_23_), 
        .B2(n14329), .ZN(n21246) );
  INV_X1 U17863 ( .A(n21246), .ZN(n21362) );
  AOI22_X1 U17864 ( .A1(n15833), .A2(n21241), .B1(n21164), .B2(n21362), .ZN(
        n14318) );
  OAI211_X1 U17865 ( .C1(n14333), .C2(n14320), .A(n14319), .B(n14318), .ZN(
        P1_U3160) );
  INV_X1 U17866 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14323) );
  MUX2_X1 U17867 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n14974), .Z(
        n14987) );
  INV_X1 U17868 ( .A(n14987), .ZN(n14490) );
  NAND2_X1 U17869 ( .A1(n14568), .A2(n14324), .ZN(n15703) );
  AOI22_X1 U17870 ( .A1(n21347), .A2(n14327), .B1(n14326), .B2(n21346), .ZN(
        n14322) );
  AOI22_X1 U17871 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14328), .B1(DATAI_29_), 
        .B2(n14329), .ZN(n21351) );
  INV_X1 U17872 ( .A(n21351), .ZN(n21231) );
  AOI22_X1 U17873 ( .A1(DATAI_21_), .A2(n14329), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n14328), .ZN(n21234) );
  INV_X1 U17874 ( .A(n21234), .ZN(n21348) );
  AOI22_X1 U17875 ( .A1(n15833), .A2(n21231), .B1(n21164), .B2(n21348), .ZN(
        n14321) );
  OAI211_X1 U17876 ( .C1(n14333), .C2(n14323), .A(n14322), .B(n14321), .ZN(
        P1_U3158) );
  INV_X1 U17877 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14332) );
  MUX2_X1 U17878 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n14974), .Z(
        n14984) );
  INV_X1 U17879 ( .A(n14984), .ZN(n15032) );
  NAND2_X1 U17880 ( .A1(n14325), .A2(n14324), .ZN(n15707) );
  AOI22_X1 U17881 ( .A1(n21353), .A2(n14327), .B1(n14326), .B2(n21352), .ZN(
        n14331) );
  AOI22_X1 U17882 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14328), .B1(DATAI_30_), 
        .B2(n14329), .ZN(n21357) );
  INV_X1 U17883 ( .A(n21357), .ZN(n21235) );
  AOI22_X1 U17884 ( .A1(DATAI_22_), .A2(n14329), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n14328), .ZN(n21238) );
  INV_X1 U17885 ( .A(n21238), .ZN(n21354) );
  AOI22_X1 U17886 ( .A1(n15833), .A2(n21235), .B1(n21164), .B2(n21354), .ZN(
        n14330) );
  OAI211_X1 U17887 ( .C1(n14333), .C2(n14332), .A(n14331), .B(n14330), .ZN(
        P1_U3159) );
  NAND2_X1 U17888 ( .A1(n9891), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21281) );
  NOR2_X1 U17889 ( .A1(n21281), .A2(n21311), .ZN(n14334) );
  AND2_X1 U17890 ( .A1(n15803), .A2(n14334), .ZN(n21316) );
  INV_X1 U17891 ( .A(n14285), .ZN(n14335) );
  AOI21_X1 U17892 ( .B1(n15526), .B2(n21204), .A(n15719), .ZN(n14338) );
  NAND2_X1 U17893 ( .A1(n21250), .A2(n15603), .ZN(n14398) );
  AOI21_X1 U17894 ( .B1(n14338), .B2(n14398), .A(n21311), .ZN(n14339) );
  AOI211_X1 U17895 ( .C1(n14340), .C2(n15531), .A(n21316), .B(n14339), .ZN(
        n14343) );
  INV_X1 U17896 ( .A(n21153), .ZN(n14342) );
  NAND2_X1 U17897 ( .A1(n14342), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14341) );
  OAI21_X1 U17898 ( .B1(n14343), .B2(n14342), .A(n14341), .ZN(P1_U3475) );
  INV_X1 U17899 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20164) );
  XNOR2_X1 U17900 ( .A(n14344), .B(n14345), .ZN(n20078) );
  INV_X1 U17901 ( .A(n20278), .ZN(n14346) );
  OAI222_X1 U17902 ( .A1(n20164), .A2(n16495), .B1(n20078), .B2(n16525), .C1(
        n20142), .C2(n14346), .ZN(P2_U2913) );
  INV_X1 U17903 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20162) );
  OAI21_X1 U17904 ( .B1(n14348), .B2(n14347), .A(n14272), .ZN(n17044) );
  INV_X1 U17905 ( .A(n20284), .ZN(n14349) );
  OAI222_X1 U17906 ( .A1(n20162), .A2(n16495), .B1(n17044), .B2(n16525), .C1(
        n20142), .C2(n14349), .ZN(P2_U2912) );
  AOI21_X1 U17907 ( .B1(n14351), .B2(n14281), .A(n14350), .ZN(n16952) );
  INV_X1 U17908 ( .A(n16952), .ZN(n14354) );
  AOI22_X1 U17909 ( .A1(n16522), .A2(n14352), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20133), .ZN(n14353) );
  OAI21_X1 U17910 ( .B1(n14354), .B2(n16525), .A(n14353), .ZN(P2_U2905) );
  NAND2_X1 U17911 ( .A1(n15531), .A2(n14232), .ZN(n21276) );
  INV_X1 U17912 ( .A(n14355), .ZN(n15599) );
  NAND2_X1 U17913 ( .A1(n15599), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14381) );
  OAI21_X1 U17914 ( .B1(n21276), .B2(n14393), .A(n14381), .ZN(n14357) );
  NOR3_X1 U17915 ( .A1(n17510), .A2(n14356), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15724) );
  AOI22_X1 U17916 ( .A1(n14357), .A2(n21285), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15724), .ZN(n14382) );
  OAI22_X1 U17917 ( .A1(n15827), .A2(n14382), .B1(n15703), .B2(n14381), .ZN(
        n14358) );
  AOI21_X1 U17918 ( .B1(n15795), .B2(n21348), .A(n14358), .ZN(n14362) );
  INV_X1 U17919 ( .A(n15719), .ZN(n21282) );
  NOR2_X1 U17920 ( .A1(n21282), .A2(n14359), .ZN(n14360) );
  NAND2_X1 U17921 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14361) );
  OAI211_X1 U17922 ( .C1(n21351), .C2(n15757), .A(n14362), .B(n14361), .ZN(
        P1_U3126) );
  OAI22_X1 U17923 ( .A1(n15830), .A2(n14382), .B1(n15707), .B2(n14381), .ZN(
        n14363) );
  AOI21_X1 U17924 ( .B1(n15795), .B2(n21354), .A(n14363), .ZN(n14365) );
  NAND2_X1 U17925 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14364) );
  OAI211_X1 U17926 ( .C1(n21357), .C2(n15757), .A(n14365), .B(n14364), .ZN(
        P1_U3127) );
  OAI22_X1 U17927 ( .A1(n15818), .A2(n14382), .B1(n15691), .B2(n14381), .ZN(
        n14366) );
  AOI21_X1 U17928 ( .B1(n15795), .B2(n21330), .A(n14366), .ZN(n14368) );
  NAND2_X1 U17929 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14367) );
  OAI211_X1 U17930 ( .C1(n21333), .C2(n15757), .A(n14368), .B(n14367), .ZN(
        P1_U3123) );
  OAI22_X1 U17931 ( .A1(n15815), .A2(n14382), .B1(n15687), .B2(n14381), .ZN(
        n14369) );
  AOI21_X1 U17932 ( .B1(n15795), .B2(n21324), .A(n14369), .ZN(n14371) );
  NAND2_X1 U17933 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14370) );
  OAI211_X1 U17934 ( .C1(n21327), .C2(n15757), .A(n14371), .B(n14370), .ZN(
        P1_U3122) );
  OAI22_X1 U17935 ( .A1(n15837), .A2(n14382), .B1(n15712), .B2(n14381), .ZN(
        n14372) );
  AOI21_X1 U17936 ( .B1(n15795), .B2(n21362), .A(n14372), .ZN(n14374) );
  NAND2_X1 U17937 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14373) );
  OAI211_X1 U17938 ( .C1(n21368), .C2(n15757), .A(n14374), .B(n14373), .ZN(
        P1_U3128) );
  OAI22_X1 U17939 ( .A1(n15821), .A2(n14382), .B1(n15695), .B2(n14381), .ZN(
        n14375) );
  AOI21_X1 U17940 ( .B1(n15795), .B2(n21336), .A(n14375), .ZN(n14377) );
  NAND2_X1 U17941 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14376) );
  OAI211_X1 U17942 ( .C1(n21339), .C2(n15757), .A(n14377), .B(n14376), .ZN(
        P1_U3124) );
  OAI22_X1 U17943 ( .A1(n15812), .A2(n14382), .B1(n15683), .B2(n14381), .ZN(
        n14378) );
  AOI21_X1 U17944 ( .B1(n15795), .B2(n21318), .A(n14378), .ZN(n14380) );
  NAND2_X1 U17945 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14379) );
  OAI211_X1 U17946 ( .C1(n21321), .C2(n15757), .A(n14380), .B(n14379), .ZN(
        P1_U3121) );
  OAI22_X1 U17947 ( .A1(n15824), .A2(n14382), .B1(n15699), .B2(n14381), .ZN(
        n14383) );
  AOI21_X1 U17948 ( .B1(n15795), .B2(n21342), .A(n14383), .ZN(n14386) );
  NAND2_X1 U17949 ( .A1(n14384), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14385) );
  OAI211_X1 U17950 ( .C1(n21345), .C2(n15757), .A(n14386), .B(n14385), .ZN(
        P1_U3125) );
  NAND2_X1 U17951 ( .A1(n14388), .A2(n14387), .ZN(n14389) );
  AND2_X1 U17952 ( .A1(n14484), .A2(n14389), .ZN(n21100) );
  INV_X1 U17953 ( .A(n21100), .ZN(n14391) );
  INV_X1 U17954 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21060) );
  OAI222_X1 U17955 ( .A1(n15031), .A2(n14391), .B1(n15029), .B2(n21060), .C1(
        n15033), .C2(n14390), .ZN(P1_U2900) );
  NOR2_X1 U17956 ( .A1(n14232), .A2(n14392), .ZN(n21248) );
  INV_X1 U17957 ( .A(n14393), .ZN(n15601) );
  INV_X1 U17958 ( .A(n14394), .ZN(n14422) );
  AOI21_X1 U17959 ( .B1(n21248), .B2(n15601), .A(n14422), .ZN(n14399) );
  INV_X1 U17960 ( .A(n14399), .ZN(n14395) );
  NOR2_X1 U17961 ( .A1(n14395), .A2(n21311), .ZN(n14397) );
  OAI21_X1 U17962 ( .B1(n21285), .B2(n11804), .A(n21315), .ZN(n14396) );
  INV_X1 U17963 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14403) );
  OAI22_X1 U17964 ( .A1(n14399), .A2(n21311), .B1(n15641), .B2(n11775), .ZN(
        n14423) );
  AOI22_X1 U17965 ( .A1(n21347), .A2(n14423), .B1(n14422), .B2(n21346), .ZN(
        n14402) );
  AOI22_X1 U17966 ( .A1(n14424), .A2(n21231), .B1(n15716), .B2(n21348), .ZN(
        n14401) );
  OAI211_X1 U17967 ( .C1(n14428), .C2(n14403), .A(n14402), .B(n14401), .ZN(
        P1_U3094) );
  INV_X1 U17968 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U17969 ( .A1(n21353), .A2(n14423), .B1(n14422), .B2(n21352), .ZN(
        n14405) );
  AOI22_X1 U17970 ( .A1(n14424), .A2(n21235), .B1(n15716), .B2(n21354), .ZN(
        n14404) );
  OAI211_X1 U17971 ( .C1(n14428), .C2(n14406), .A(n14405), .B(n14404), .ZN(
        P1_U3095) );
  INV_X1 U17972 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17973 ( .A1(n21361), .A2(n14423), .B1(n14422), .B2(n21359), .ZN(
        n14408) );
  AOI22_X1 U17974 ( .A1(n14424), .A2(n21241), .B1(n15716), .B2(n21362), .ZN(
        n14407) );
  OAI211_X1 U17975 ( .C1(n14428), .C2(n14409), .A(n14408), .B(n14407), .ZN(
        P1_U3096) );
  INV_X1 U17976 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17977 ( .A1(n21314), .A2(n14423), .B1(n14422), .B2(n21313), .ZN(
        n14411) );
  AOI22_X1 U17978 ( .A1(n14424), .A2(n21211), .B1(n15716), .B2(n21318), .ZN(
        n14410) );
  OAI211_X1 U17979 ( .C1(n14428), .C2(n14412), .A(n14411), .B(n14410), .ZN(
        P1_U3089) );
  INV_X1 U17980 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14415) );
  AOI22_X1 U17981 ( .A1(n21341), .A2(n14423), .B1(n14422), .B2(n21340), .ZN(
        n14414) );
  AOI22_X1 U17982 ( .A1(n14424), .A2(n21227), .B1(n15716), .B2(n21342), .ZN(
        n14413) );
  OAI211_X1 U17983 ( .C1(n14428), .C2(n14415), .A(n14414), .B(n14413), .ZN(
        P1_U3093) );
  INV_X1 U17984 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17985 ( .A1(n21329), .A2(n14423), .B1(n14422), .B2(n21328), .ZN(
        n14417) );
  AOI22_X1 U17986 ( .A1(n14424), .A2(n21219), .B1(n15716), .B2(n21330), .ZN(
        n14416) );
  OAI211_X1 U17987 ( .C1(n14428), .C2(n14418), .A(n14417), .B(n14416), .ZN(
        P1_U3091) );
  INV_X1 U17988 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U17989 ( .A1(n21335), .A2(n14423), .B1(n14422), .B2(n21334), .ZN(
        n14420) );
  AOI22_X1 U17990 ( .A1(n14424), .A2(n21223), .B1(n15716), .B2(n21336), .ZN(
        n14419) );
  OAI211_X1 U17991 ( .C1(n14428), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        P1_U3092) );
  INV_X1 U17992 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17993 ( .A1(n21323), .A2(n14423), .B1(n14422), .B2(n21322), .ZN(
        n14426) );
  AOI22_X1 U17994 ( .A1(n14424), .A2(n21215), .B1(n15716), .B2(n21324), .ZN(
        n14425) );
  OAI211_X1 U17995 ( .C1(n14428), .C2(n14427), .A(n14426), .B(n14425), .ZN(
        P1_U3090) );
  INV_X1 U17996 ( .A(n14429), .ZN(n14432) );
  AOI21_X1 U17997 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14433) );
  OR2_X1 U17998 ( .A1(n14433), .A2(n14487), .ZN(n21003) );
  OAI22_X1 U17999 ( .A1(n14960), .A2(n21003), .B1(n21007), .B2(n21035), .ZN(
        n14434) );
  AOI21_X1 U18000 ( .B1(n21100), .B2(n21031), .A(n14434), .ZN(n14435) );
  INV_X1 U18001 ( .A(n14435), .ZN(P1_U2868) );
  NOR2_X1 U18002 ( .A1(n14436), .A2(n21389), .ZN(n14437) );
  INV_X2 U18003 ( .A(n14444), .ZN(n21090) );
  INV_X1 U18004 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n21037) );
  NOR2_X2 U18005 ( .A1(n21090), .A2(n14546), .ZN(n21080) );
  INV_X1 U18006 ( .A(n21080), .ZN(n14442) );
  NOR2_X1 U18007 ( .A1(n14440), .A2(n14438), .ZN(n14439) );
  AOI21_X1 U18008 ( .B1(DATAI_15_), .B2(n14440), .A(n14439), .ZN(n15012) );
  INV_X1 U18009 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14441) );
  OAI222_X1 U18010 ( .A1(n14443), .A2(n21037), .B1(n14442), .B2(n15012), .C1(
        n14441), .C2(n14444), .ZN(P1_U2967) );
  AOI22_X1 U18011 ( .A1(n21091), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n21090), .ZN(n14445) );
  NAND2_X1 U18012 ( .A1(n21080), .A2(n15007), .ZN(n14462) );
  NAND2_X1 U18013 ( .A1(n14445), .A2(n14462), .ZN(P1_U2952) );
  AOI22_X1 U18014 ( .A1(n21091), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n21090), .ZN(n14446) );
  NAND2_X1 U18015 ( .A1(n21080), .A2(n15001), .ZN(n14460) );
  NAND2_X1 U18016 ( .A1(n14446), .A2(n14460), .ZN(P1_U2953) );
  AOI22_X1 U18017 ( .A1(n21091), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n21090), .ZN(n14447) );
  MUX2_X1 U18018 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14974), .Z(
        n15025) );
  NAND2_X1 U18019 ( .A1(n21080), .A2(n15025), .ZN(n14456) );
  NAND2_X1 U18020 ( .A1(n14447), .A2(n14456), .ZN(P1_U2945) );
  AOI22_X1 U18021 ( .A1(n21091), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n21090), .ZN(n14448) );
  NAND2_X1 U18022 ( .A1(n21080), .A2(n14980), .ZN(n14464) );
  NAND2_X1 U18023 ( .A1(n14448), .A2(n14464), .ZN(P1_U2944) );
  AOI22_X1 U18024 ( .A1(n21091), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n21090), .ZN(n14449) );
  NAND2_X1 U18025 ( .A1(n21080), .A2(n14984), .ZN(n14471) );
  NAND2_X1 U18026 ( .A1(n14449), .A2(n14471), .ZN(P1_U2943) );
  AOI22_X1 U18027 ( .A1(n21091), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n21090), .ZN(n14450) );
  NAND2_X1 U18028 ( .A1(n21080), .A2(n14987), .ZN(n14468) );
  NAND2_X1 U18029 ( .A1(n14450), .A2(n14468), .ZN(P1_U2942) );
  AOI22_X1 U18030 ( .A1(n21091), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n21090), .ZN(n14451) );
  NAND2_X1 U18031 ( .A1(n21080), .A2(n14991), .ZN(n14454) );
  NAND2_X1 U18032 ( .A1(n14451), .A2(n14454), .ZN(P1_U2941) );
  AOI22_X1 U18033 ( .A1(n21091), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n21090), .ZN(n14452) );
  NAND2_X1 U18034 ( .A1(n21080), .A2(n14994), .ZN(n14466) );
  NAND2_X1 U18035 ( .A1(n14452), .A2(n14466), .ZN(P1_U2955) );
  AOI22_X1 U18036 ( .A1(n21091), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n21090), .ZN(n14453) );
  NAND2_X1 U18037 ( .A1(n21080), .A2(n14998), .ZN(n14458) );
  NAND2_X1 U18038 ( .A1(n14453), .A2(n14458), .ZN(P1_U2954) );
  AOI22_X1 U18039 ( .A1(n21091), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n21090), .ZN(n14455) );
  NAND2_X1 U18040 ( .A1(n14455), .A2(n14454), .ZN(P1_U2956) );
  AOI22_X1 U18041 ( .A1(n21091), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n21090), .ZN(n14457) );
  NAND2_X1 U18042 ( .A1(n14457), .A2(n14456), .ZN(P1_U2960) );
  AOI22_X1 U18043 ( .A1(n21091), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21090), .ZN(n14459) );
  NAND2_X1 U18044 ( .A1(n14459), .A2(n14458), .ZN(P1_U2939) );
  AOI22_X1 U18045 ( .A1(n21091), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n21090), .ZN(n14461) );
  NAND2_X1 U18046 ( .A1(n14461), .A2(n14460), .ZN(P1_U2938) );
  AOI22_X1 U18047 ( .A1(n21091), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n21090), .ZN(n14463) );
  NAND2_X1 U18048 ( .A1(n14463), .A2(n14462), .ZN(P1_U2937) );
  AOI22_X1 U18049 ( .A1(n21091), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n21090), .ZN(n14465) );
  NAND2_X1 U18050 ( .A1(n14465), .A2(n14464), .ZN(P1_U2959) );
  AOI22_X1 U18051 ( .A1(n21091), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n21090), .ZN(n14467) );
  NAND2_X1 U18052 ( .A1(n14467), .A2(n14466), .ZN(P1_U2940) );
  AOI22_X1 U18053 ( .A1(n21091), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n21090), .ZN(n14469) );
  NAND2_X1 U18054 ( .A1(n14469), .A2(n14468), .ZN(P1_U2957) );
  AOI22_X1 U18055 ( .A1(n21091), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n21090), .ZN(n14470) );
  MUX2_X1 U18056 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14974), .Z(
        n15016) );
  NAND2_X1 U18057 ( .A1(n21080), .A2(n15016), .ZN(n14473) );
  NAND2_X1 U18058 ( .A1(n14470), .A2(n14473), .ZN(P1_U2949) );
  AOI22_X1 U18059 ( .A1(n21091), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n21090), .ZN(n14472) );
  NAND2_X1 U18060 ( .A1(n14472), .A2(n14471), .ZN(P1_U2958) );
  AOI22_X1 U18061 ( .A1(n21091), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n21090), .ZN(n14474) );
  NAND2_X1 U18062 ( .A1(n14474), .A2(n14473), .ZN(P1_U2964) );
  NOR2_X1 U18063 ( .A1(n14350), .A2(n14476), .ZN(n14477) );
  OR2_X1 U18064 ( .A1(n14475), .A2(n14477), .ZN(n16934) );
  OAI222_X1 U18065 ( .A1(n16934), .A2(n16525), .B1(n16495), .B2(n13672), .C1(
        n14478), .C2(n20142), .ZN(P2_U2904) );
  XNOR2_X1 U18066 ( .A(n21096), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14480) );
  NOR2_X1 U18067 ( .A1(n14480), .A2(n10175), .ZN(n21095) );
  AOI21_X1 U18068 ( .B1(n14480), .B2(n10175), .A(n21095), .ZN(n21118) );
  NAND2_X1 U18069 ( .A1(n21118), .A2(n21102), .ZN(n14483) );
  AND2_X1 U18070 ( .A1(n21133), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n21115) );
  NOR2_X1 U18071 ( .A1(n21106), .A2(n14890), .ZN(n14481) );
  AOI211_X1 U18072 ( .C1(n21094), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n21115), .B(n14481), .ZN(n14482) );
  OAI211_X1 U18073 ( .C1(n15264), .C2(n14898), .A(n14483), .B(n14482), .ZN(
        P1_U2996) );
  OAI21_X1 U18074 ( .B1(n9600), .B2(n9887), .A(n15027), .ZN(n17582) );
  INV_X1 U18075 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14489) );
  NOR2_X1 U18076 ( .A1(n14487), .A2(n14486), .ZN(n14488) );
  OR2_X1 U18077 ( .A1(n17612), .A2(n14488), .ZN(n17621) );
  OAI222_X1 U18078 ( .A1(n17582), .A2(n14963), .B1(n21035), .B2(n14489), .C1(
        n17621), .C2(n14960), .ZN(P1_U2867) );
  OAI222_X1 U18079 ( .A1(n15031), .A2(n17582), .B1(n15029), .B2(n11875), .C1(
        n15033), .C2(n14490), .ZN(P1_U2899) );
  OAI21_X1 U18080 ( .B1(n14493), .B2(n14492), .A(n14491), .ZN(n20973) );
  XNOR2_X1 U18081 ( .A(n14494), .B(n14862), .ZN(n20977) );
  AOI22_X1 U18082 ( .A1(n21030), .A2(n20977), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14961), .ZN(n14495) );
  OAI21_X1 U18083 ( .B1(n20973), .B2(n14963), .A(n14495), .ZN(P1_U2865) );
  INV_X1 U18084 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n21054) );
  OAI222_X1 U18085 ( .A1(n15031), .A2(n20973), .B1(n15029), .B2(n21054), .C1(
        n15033), .C2(n14496), .ZN(P1_U2897) );
  INV_X1 U18086 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n14498) );
  NAND2_X1 U18087 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18462) );
  NOR2_X1 U18088 ( .A1(n9829), .A2(n18462), .ZN(n18452) );
  NAND3_X1 U18089 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18452), .ZN(n18450) );
  NAND3_X1 U18090 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n18438) );
  INV_X1 U18091 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n14499) );
  NOR2_X1 U18092 ( .A1(n18518), .A2(n18470), .ZN(n18451) );
  NOR4_X1 U18093 ( .A1(n14499), .A2(n18442), .A3(n18450), .A4(n18473), .ZN(
        n18445) );
  AOI21_X1 U18094 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18445), .A(
        P3_EBX_REG_8__SCAN_IN), .ZN(n14500) );
  NOR2_X1 U18095 ( .A1(n18436), .A2(n14500), .ZN(n14512) );
  AOI22_X1 U18096 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U18097 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U18098 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U18099 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14501) );
  NAND4_X1 U18100 ( .A1(n14504), .A2(n14503), .A3(n14502), .A4(n14501), .ZN(
        n14510) );
  AOI22_X1 U18101 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14508) );
  AOI22_X1 U18102 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U18103 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U18104 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14505) );
  NAND4_X1 U18105 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        n14509) );
  NOR2_X1 U18106 ( .A1(n14510), .A2(n14509), .ZN(n18588) );
  INV_X1 U18107 ( .A(n18588), .ZN(n14511) );
  MUX2_X1 U18108 ( .A(n14512), .B(n14511), .S(n18471), .Z(P3_U2695) );
  INV_X1 U18109 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18320) );
  INV_X1 U18110 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18017) );
  NAND4_X1 U18111 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n14513) );
  NOR3_X1 U18112 ( .A1(n18450), .A2(n18438), .A3(n14513), .ZN(n18376) );
  NAND2_X1 U18113 ( .A1(n18468), .A2(n18376), .ZN(n18377) );
  NAND2_X1 U18114 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18362), .ZN(n18361) );
  NAND4_X1 U18115 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17392)
         );
  AND2_X1 U18116 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17393) );
  NAND3_X1 U18117 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17393), .ZN(n18222) );
  NOR4_X1 U18118 ( .A1(n14514), .A2(n18278), .A3(n17392), .A4(n18222), .ZN(
        n18216) );
  NAND2_X1 U18119 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18216), .ZN(n14515) );
  NOR2_X1 U18120 ( .A1(n18518), .A2(n14515), .ZN(n14517) );
  NAND2_X1 U18121 ( .A1(n18458), .A2(n14515), .ZN(n18217) );
  INV_X1 U18122 ( .A(n18217), .ZN(n14516) );
  MUX2_X1 U18123 ( .A(n14517), .B(n14516), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NAND2_X1 U18124 ( .A1(n14518), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14520) );
  NAND2_X1 U18125 ( .A1(n14520), .A2(n14519), .ZN(n14525) );
  NAND2_X1 U18126 ( .A1(n14521), .A2(n14525), .ZN(n19856) );
  NOR2_X1 U18127 ( .A1(n14522), .A2(n19856), .ZN(n14524) );
  MUX2_X1 U18128 ( .A(n14524), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n14523), .Z(P3_U3284) );
  OR2_X1 U18129 ( .A1(n13868), .A2(n14525), .ZN(n19409) );
  NOR2_X1 U18130 ( .A1(n19409), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(n14527) );
  OAI21_X1 U18131 ( .B1(n14527), .B2(n20007), .A(n19523), .ZN(n19419) );
  INV_X1 U18132 ( .A(n19419), .ZN(n14528) );
  OAI21_X1 U18133 ( .B1(n20039), .B2(n19895), .A(n20009), .ZN(n20025) );
  NOR2_X1 U18134 ( .A1(n19895), .A2(n17812), .ZN(n19004) );
  NOR2_X1 U18135 ( .A1(n20025), .A2(n19004), .ZN(n19412) );
  AOI21_X1 U18136 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19412), .ZN(n19413) );
  NOR2_X1 U18137 ( .A1(n14528), .A2(n19413), .ZN(n14530) );
  INV_X1 U18138 ( .A(n19756), .ZN(n19414) );
  NOR2_X1 U18139 ( .A1(n20009), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19458) );
  OR2_X1 U18140 ( .A1(n19458), .A2(n14528), .ZN(n19411) );
  OR2_X1 U18141 ( .A1(n19414), .A2(n19411), .ZN(n14529) );
  MUX2_X1 U18142 ( .A(n14530), .B(n14529), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U18143 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14587) );
  XNOR2_X2 U18144 ( .A(n14534), .B(n14587), .ZN(n15040) );
  NAND2_X1 U18145 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21468), .ZN(n17534) );
  AND2_X1 U18146 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21369), .ZN(n14537) );
  NAND2_X1 U18147 ( .A1(n14538), .A2(n14537), .ZN(n14539) );
  OAI211_X1 U18148 ( .C1(n17534), .C2(n21369), .A(n15176), .B(n14539), .ZN(
        n14540) );
  NAND2_X1 U18149 ( .A1(n14884), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14560) );
  OR2_X1 U18150 ( .A1(n14886), .A2(n14541), .ZN(n14544) );
  AND2_X1 U18151 ( .A1(n14542), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U18152 ( .A1(n21389), .A2(n21204), .ZN(n17522) );
  NAND2_X1 U18153 ( .A1(n14547), .A2(n17522), .ZN(n14543) );
  NOR2_X4 U18154 ( .A1(n14544), .A2(n14543), .ZN(n21013) );
  AOI21_X1 U18155 ( .B1(n14546), .B2(n14545), .A(n17522), .ZN(n14549) );
  NOR2_X1 U18156 ( .A1(n14549), .A2(n14547), .ZN(n14548) );
  INV_X1 U18157 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14574) );
  INV_X1 U18158 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21399) );
  NAND3_X1 U18159 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n21000) );
  NOR2_X1 U18160 ( .A1(n21399), .A2(n21000), .ZN(n14874) );
  INV_X1 U18161 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21406) );
  NAND2_X1 U18162 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20968) );
  NOR2_X1 U18163 ( .A1(n21406), .A2(n20968), .ZN(n14860) );
  NAND3_X1 U18164 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14874), .A3(n14860), 
        .ZN(n14819) );
  NAND2_X1 U18165 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14818) );
  INV_X1 U18166 ( .A(n14818), .ZN(n17550) );
  AND4_X1 U18167 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_14__SCAN_IN), .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U18168 ( .A1(n17550), .A2(n14551), .ZN(n14552) );
  NOR2_X1 U18169 ( .A1(n14819), .A2(n14552), .ZN(n14731) );
  INV_X1 U18170 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15175) );
  INV_X1 U18171 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15187) );
  NOR2_X1 U18172 ( .A1(n15175), .A2(n15187), .ZN(n14779) );
  AND2_X1 U18173 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14779), .ZN(n14730) );
  AND3_X1 U18174 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(n14730), .ZN(n14553) );
  AND2_X1 U18175 ( .A1(n14731), .A2(n14553), .ZN(n14718) );
  AND2_X1 U18176 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14554) );
  AND2_X1 U18177 ( .A1(n14718), .A2(n14554), .ZN(n14691) );
  NAND3_X1 U18178 ( .A1(n14691), .A2(P1_REIP_REG_23__SCAN_IN), .A3(
        P1_REIP_REG_22__SCAN_IN), .ZN(n14668) );
  INV_X1 U18179 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15089) );
  NOR3_X1 U18180 ( .A1(n14668), .A2(n21429), .A3(n15089), .ZN(n14642) );
  INV_X1 U18181 ( .A(n14642), .ZN(n14555) );
  INV_X1 U18182 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15080) );
  NOR3_X1 U18183 ( .A1(n20970), .A2(n14555), .A3(n15080), .ZN(n14624) );
  NAND2_X1 U18184 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14557) );
  INV_X1 U18185 ( .A(n14557), .ZN(n14556) );
  NAND2_X1 U18186 ( .A1(n14624), .A2(n14556), .ZN(n14603) );
  INV_X1 U18187 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21437) );
  NOR2_X1 U18188 ( .A1(n14603), .A2(n21437), .ZN(n14559) );
  AND2_X1 U18189 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14585) );
  NAND2_X1 U18190 ( .A1(n20970), .A2(n14884), .ZN(n14915) );
  INV_X1 U18191 ( .A(n14915), .ZN(n14558) );
  NOR2_X1 U18192 ( .A1(n20970), .A2(n14642), .ZN(n14655) );
  INV_X1 U18193 ( .A(n14884), .ZN(n14902) );
  NOR2_X1 U18194 ( .A1(n14655), .A2(n14902), .ZN(n14654) );
  OAI21_X1 U18195 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n20970), .A(n14654), 
        .ZN(n14641) );
  AOI21_X1 U18196 ( .B1(n14915), .B2(n14557), .A(n14641), .ZN(n14616) );
  OAI21_X1 U18197 ( .B1(n14585), .B2(n14558), .A(n14616), .ZN(n14590) );
  OAI21_X1 U18198 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14559), .A(n14590), 
        .ZN(n14564) );
  INV_X1 U18199 ( .A(n14560), .ZN(n14561) );
  AOI22_X1 U18200 ( .A1(n21018), .A2(n14562), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21016), .ZN(n14563) );
  OAI211_X1 U18201 ( .C1(n21006), .C2(n14574), .A(n14564), .B(n14563), .ZN(
        n14565) );
  AOI21_X1 U18202 ( .B1(n14573), .B2(n21013), .A(n14565), .ZN(n14566) );
  OAI21_X1 U18203 ( .B1(n14531), .B2(n20974), .A(n14566), .ZN(P1_U2810) );
  AOI22_X1 U18204 ( .A1(n15005), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15022), .ZN(n14572) );
  NOR3_X1 U18205 ( .A1(n15022), .A2(n14569), .A3(n14568), .ZN(n14570) );
  MUX2_X1 U18206 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14974), .Z(
        n21079) );
  AOI22_X1 U18207 ( .A1(n15008), .A2(n21079), .B1(n15006), .B2(DATAI_30_), 
        .ZN(n14571) );
  OAI211_X1 U18208 ( .C1(n14531), .C2(n15031), .A(n14572), .B(n14571), .ZN(
        P1_U2874) );
  INV_X1 U18209 ( .A(n14573), .ZN(n14575) );
  OAI222_X1 U18210 ( .A1(n14960), .A2(n14575), .B1(n14574), .B2(n21035), .C1(
        n14531), .C2(n14963), .ZN(P1_U2842) );
  OR2_X1 U18211 ( .A1(n14732), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14578) );
  NAND2_X1 U18212 ( .A1(n14872), .A2(n14576), .ZN(n14577) );
  MUX2_X1 U18213 ( .A(n14578), .B(n14577), .S(n21462), .Z(P1_U3487) );
  AOI22_X1 U18214 ( .A1(n14580), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14579), .ZN(n14582) );
  XNOR2_X1 U18215 ( .A(n14582), .B(n14581), .ZN(n14584) );
  OR2_X1 U18216 ( .A1(n14582), .A2(n10323), .ZN(n14583) );
  MUX2_X1 U18217 ( .A(n14584), .B(n14583), .S(n14593), .Z(n15265) );
  NAND2_X1 U18218 ( .A1(n15042), .A2(n20989), .ZN(n14592) );
  INV_X1 U18219 ( .A(n14585), .ZN(n14586) );
  NOR3_X1 U18220 ( .A1(n14603), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14586), 
        .ZN(n14589) );
  INV_X1 U18221 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14919) );
  OAI22_X1 U18222 ( .A1(n21006), .A2(n14919), .B1(n14587), .B2(n20980), .ZN(
        n14588) );
  AOI211_X1 U18223 ( .C1(n14590), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14589), 
        .B(n14588), .ZN(n14591) );
  OAI211_X1 U18224 ( .C1(n15265), .C2(n14888), .A(n14592), .B(n14591), .ZN(
        P1_U2809) );
  OAI21_X1 U18225 ( .B1(n14611), .B2(n14594), .A(n14593), .ZN(n15273) );
  INV_X1 U18226 ( .A(n14595), .ZN(n14599) );
  INV_X1 U18227 ( .A(n14596), .ZN(n14598) );
  NAND2_X1 U18228 ( .A1(n15051), .A2(n20989), .ZN(n14607) );
  INV_X1 U18229 ( .A(n14616), .ZN(n14605) );
  INV_X1 U18230 ( .A(n15049), .ZN(n14600) );
  AOI22_X1 U18231 ( .A1(n21018), .A2(n14600), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21016), .ZN(n14602) );
  NAND2_X1 U18232 ( .A1(n21014), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14601) );
  OAI211_X1 U18233 ( .C1(n14603), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14602), 
        .B(n14601), .ZN(n14604) );
  AOI21_X1 U18234 ( .B1(n14605), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14604), 
        .ZN(n14606) );
  OAI211_X1 U18235 ( .C1(n15273), .C2(n14888), .A(n14607), .B(n14606), .ZN(
        P1_U2811) );
  NOR2_X1 U18236 ( .A1(n14608), .A2(n14609), .ZN(n14610) );
  AOI21_X1 U18237 ( .B1(n14613), .B2(n14612), .A(n14596), .ZN(n15066) );
  NAND2_X1 U18238 ( .A1(n15066), .A2(n20989), .ZN(n14620) );
  OAI22_X1 U18239 ( .A1(n20983), .A2(n15064), .B1(n14614), .B2(n20980), .ZN(
        n14618) );
  AOI21_X1 U18240 ( .B1(n14624), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14615) );
  NOR2_X1 U18241 ( .A1(n14616), .A2(n14615), .ZN(n14617) );
  AOI211_X1 U18242 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n21014), .A(n14618), .B(
        n14617), .ZN(n14619) );
  OAI211_X1 U18243 ( .C1(n15287), .C2(n14888), .A(n14620), .B(n14619), .ZN(
        P1_U2812) );
  AND2_X1 U18244 ( .A1(n14686), .A2(n14688), .ZN(n14622) );
  OAI21_X1 U18245 ( .B1(n14635), .B2(n14623), .A(n14612), .ZN(n15071) );
  INV_X1 U18246 ( .A(n14624), .ZN(n14628) );
  OAI22_X1 U18247 ( .A1(n20983), .A2(n15073), .B1(n14625), .B2(n20980), .ZN(
        n14626) );
  AOI21_X1 U18248 ( .B1(n21014), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14626), .ZN(
        n14627) );
  OAI21_X1 U18249 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14628), .A(n14627), 
        .ZN(n14632) );
  NOR2_X1 U18250 ( .A1(n14640), .A2(n14629), .ZN(n14630) );
  OR2_X1 U18251 ( .A1(n14608), .A2(n14630), .ZN(n15292) );
  NOR2_X1 U18252 ( .A1(n15292), .A2(n14888), .ZN(n14631) );
  OAI21_X1 U18253 ( .B1(n15071), .B2(n20974), .A(n14633), .ZN(P1_U2813) );
  INV_X1 U18254 ( .A(n14635), .ZN(n14636) );
  AND2_X1 U18255 ( .A1(n14653), .A2(n14638), .ZN(n14639) );
  NOR2_X1 U18256 ( .A1(n14640), .A2(n14639), .ZN(n15308) );
  INV_X1 U18257 ( .A(n14641), .ZN(n14647) );
  AOI21_X1 U18258 ( .B1(n21002), .B2(n14642), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14646) );
  INV_X1 U18259 ( .A(n15082), .ZN(n14643) );
  AOI22_X1 U18260 ( .A1(n21018), .A2(n14643), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21016), .ZN(n14645) );
  NAND2_X1 U18261 ( .A1(n21014), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14644) );
  OAI211_X1 U18262 ( .C1(n14647), .C2(n14646), .A(n14645), .B(n14644), .ZN(
        n14648) );
  AOI21_X1 U18263 ( .B1(n15308), .B2(n21013), .A(n14648), .ZN(n14649) );
  OAI21_X1 U18264 ( .B1(n15079), .B2(n20974), .A(n14649), .ZN(P1_U2814) );
  NAND2_X1 U18265 ( .A1(n14673), .A2(n14651), .ZN(n14652) );
  NAND2_X1 U18266 ( .A1(n14653), .A2(n14652), .ZN(n14924) );
  INV_X1 U18267 ( .A(n14924), .ZN(n15318) );
  NOR2_X1 U18268 ( .A1(n14654), .A2(n21429), .ZN(n14661) );
  INV_X1 U18269 ( .A(n14668), .ZN(n14667) );
  NAND3_X1 U18270 ( .A1(n14655), .A2(n14667), .A3(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14659) );
  INV_X1 U18271 ( .A(n14656), .ZN(n14657) );
  AOI22_X1 U18272 ( .A1(n21018), .A2(n14657), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21016), .ZN(n14658) );
  OAI211_X1 U18273 ( .C1(n14925), .C2(n21006), .A(n14659), .B(n14658), .ZN(
        n14660) );
  AOI211_X1 U18274 ( .C1(n15318), .C2(n21013), .A(n14661), .B(n14660), .ZN(
        n14662) );
  OAI21_X1 U18275 ( .B1(n14650), .B2(n20974), .A(n14662), .ZN(P1_U2815) );
  OAI21_X1 U18276 ( .B1(n20970), .B2(n14667), .A(n14884), .ZN(n14679) );
  NOR3_X1 U18277 ( .A1(n20970), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14668), 
        .ZN(n14672) );
  INV_X1 U18278 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14670) );
  AOI22_X1 U18279 ( .A1(n21018), .A2(n15088), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21016), .ZN(n14669) );
  OAI21_X1 U18280 ( .B1(n21006), .B2(n14670), .A(n14669), .ZN(n14671) );
  AOI211_X1 U18281 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14679), .A(n14672), 
        .B(n14671), .ZN(n14678) );
  INV_X1 U18282 ( .A(n14673), .ZN(n14674) );
  AOI21_X1 U18283 ( .B1(n14676), .B2(n14675), .A(n14674), .ZN(n15327) );
  NAND2_X1 U18284 ( .A1(n15327), .A2(n21013), .ZN(n14677) );
  OAI211_X1 U18285 ( .C1(n14979), .C2(n20974), .A(n14678), .B(n14677), .ZN(
        P1_U2816) );
  INV_X1 U18286 ( .A(n15100), .ZN(n14983) );
  INV_X1 U18287 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14683) );
  AND3_X1 U18288 ( .A1(n21002), .A2(n14691), .A3(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14680) );
  OAI21_X1 U18289 ( .B1(n14680), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14679), 
        .ZN(n14682) );
  AOI22_X1 U18290 ( .A1(n21018), .A2(n15096), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21016), .ZN(n14681) );
  OAI211_X1 U18291 ( .C1(n14683), .C2(n21006), .A(n14682), .B(n14681), .ZN(
        n14684) );
  AOI21_X1 U18292 ( .B1(n15335), .B2(n21013), .A(n14684), .ZN(n14685) );
  OAI21_X1 U18293 ( .B1(n14983), .B2(n20974), .A(n14685), .ZN(P1_U2817) );
  OAI21_X1 U18294 ( .B1(n14701), .B2(n14688), .A(n14687), .ZN(n15105) );
  INV_X1 U18295 ( .A(n14718), .ZN(n14703) );
  INV_X1 U18296 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21423) );
  OAI21_X1 U18297 ( .B1(n14703), .B2(n21423), .A(n21002), .ZN(n14689) );
  NAND2_X1 U18298 ( .A1(n14689), .A2(n14884), .ZN(n14717) );
  INV_X1 U18299 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U18300 ( .A1(n21018), .A2(n15106), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21016), .ZN(n14693) );
  NAND2_X1 U18301 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14690) );
  OAI211_X1 U18302 ( .C1(n14691), .C2(P1_REIP_REG_22__SCAN_IN), .A(n21002), 
        .B(n14690), .ZN(n14692) );
  OAI211_X1 U18303 ( .C1(n14927), .C2(n21006), .A(n14693), .B(n14692), .ZN(
        n14698) );
  INV_X1 U18304 ( .A(n12860), .ZN(n14694) );
  OAI21_X1 U18305 ( .B1(n14696), .B2(n14695), .A(n14694), .ZN(n15348) );
  NOR2_X1 U18306 ( .A1(n15348), .A2(n14888), .ZN(n14697) );
  AOI211_X1 U18307 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14717), .A(n14698), 
        .B(n14697), .ZN(n14699) );
  OAI21_X1 U18308 ( .B1(n15105), .B2(n20974), .A(n14699), .ZN(P1_U2818) );
  NOR2_X1 U18309 ( .A1(n10480), .A2(n14700), .ZN(n14702) );
  NOR2_X1 U18310 ( .A1(n14702), .A2(n14701), .ZN(n15126) );
  INV_X1 U18311 ( .A(n15126), .ZN(n14990) );
  NOR4_X1 U18312 ( .A1(n20970), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14703), 
        .A4(n21423), .ZN(n14708) );
  INV_X1 U18313 ( .A(n15124), .ZN(n14704) );
  AOI22_X1 U18314 ( .A1(n21018), .A2(n14704), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21016), .ZN(n14705) );
  OAI21_X1 U18315 ( .B1(n21006), .B2(n14706), .A(n14705), .ZN(n14707) );
  AOI211_X1 U18316 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n14717), .A(n14708), 
        .B(n14707), .ZN(n14711) );
  XOR2_X1 U18317 ( .A(n14709), .B(n14716), .Z(n15357) );
  NAND2_X1 U18318 ( .A1(n15357), .A2(n21013), .ZN(n14710) );
  OAI211_X1 U18319 ( .C1(n14990), .C2(n20974), .A(n14711), .B(n14710), .ZN(
        P1_U2819) );
  XNOR2_X1 U18320 ( .A(n14727), .B(n14713), .ZN(n15131) );
  NAND2_X1 U18321 ( .A1(n14725), .A2(n14714), .ZN(n14715) );
  AND2_X1 U18322 ( .A1(n14716), .A2(n14715), .ZN(n15371) );
  INV_X1 U18323 ( .A(n14717), .ZN(n14722) );
  AOI21_X1 U18324 ( .B1(n21002), .B2(n14718), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14721) );
  AOI22_X1 U18325 ( .A1(n21018), .A2(n15134), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21016), .ZN(n14720) );
  NAND2_X1 U18326 ( .A1(n21014), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n14719) );
  OAI211_X1 U18327 ( .C1(n14722), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        n14723) );
  AOI21_X1 U18328 ( .B1(n15371), .B2(n21013), .A(n14723), .ZN(n14724) );
  OAI21_X1 U18329 ( .B1(n15131), .B2(n20974), .A(n14724), .ZN(P1_U2820) );
  OAI21_X1 U18330 ( .B1(n14750), .B2(n14726), .A(n14725), .ZN(n15374) );
  AOI21_X1 U18331 ( .B1(n14728), .B2(n14740), .A(n14712), .ZN(n15144) );
  NAND2_X1 U18332 ( .A1(n15144), .A2(n20989), .ZN(n14739) );
  INV_X1 U18333 ( .A(n14731), .ZN(n14729) );
  AOI21_X1 U18334 ( .B1(n21002), .B2(n14729), .A(n14902), .ZN(n17552) );
  OAI21_X1 U18335 ( .B1(n14730), .B2(n20970), .A(n17552), .ZN(n14762) );
  INV_X1 U18336 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14930) );
  NOR2_X1 U18337 ( .A1(n21006), .A2(n14930), .ZN(n14737) );
  XOR2_X1 U18338 ( .A(P1_REIP_REG_18__SCAN_IN), .B(P1_REIP_REG_19__SCAN_IN), 
        .Z(n14733) );
  INV_X1 U18339 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21418) );
  NAND2_X1 U18340 ( .A1(n21002), .A2(n14731), .ZN(n14799) );
  INV_X1 U18341 ( .A(n14799), .ZN(n14781) );
  NAND2_X1 U18342 ( .A1(n14781), .A2(n14779), .ZN(n14764) );
  NOR2_X1 U18343 ( .A1(n21418), .A2(n14764), .ZN(n14745) );
  NAND2_X1 U18344 ( .A1(n14884), .A2(n14732), .ZN(n20998) );
  INV_X1 U18345 ( .A(n20998), .ZN(n20952) );
  AOI21_X1 U18346 ( .B1(n14733), .B2(n14745), .A(n20952), .ZN(n14735) );
  NAND2_X1 U18347 ( .A1(n21016), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14734) );
  OAI211_X1 U18348 ( .C1(n20983), .C2(n15142), .A(n14735), .B(n14734), .ZN(
        n14736) );
  AOI211_X1 U18349 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n14762), .A(n14737), 
        .B(n14736), .ZN(n14738) );
  OAI211_X1 U18350 ( .C1(n15374), .C2(n14888), .A(n14739), .B(n14738), .ZN(
        P1_U2821) );
  OAI21_X1 U18351 ( .B1(n14756), .B2(n14741), .A(n14740), .ZN(n15147) );
  INV_X1 U18352 ( .A(n14742), .ZN(n15150) );
  INV_X1 U18353 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15148) );
  INV_X1 U18354 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14743) );
  NOR2_X1 U18355 ( .A1(n20980), .A2(n14743), .ZN(n14744) );
  AOI211_X1 U18356 ( .C1(n14745), .C2(n15148), .A(n20952), .B(n14744), .ZN(
        n14747) );
  NAND2_X1 U18357 ( .A1(n21014), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14746) );
  OAI211_X1 U18358 ( .C1(n20983), .C2(n15150), .A(n14747), .B(n14746), .ZN(
        n14748) );
  AOI21_X1 U18359 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n14762), .A(n14748), 
        .ZN(n14754) );
  INV_X1 U18360 ( .A(n14767), .ZN(n14749) );
  NAND2_X1 U18361 ( .A1(n14776), .A2(n14749), .ZN(n14751) );
  AOI21_X1 U18362 ( .B1(n14752), .B2(n14751), .A(n14750), .ZN(n15391) );
  NAND2_X1 U18363 ( .A1(n15391), .A2(n21013), .ZN(n14753) );
  OAI211_X1 U18364 ( .C1(n15147), .C2(n20974), .A(n14754), .B(n14753), .ZN(
        P1_U2822) );
  INV_X1 U18365 ( .A(n14755), .ZN(n14758) );
  INV_X1 U18366 ( .A(n14771), .ZN(n14757) );
  AOI21_X1 U18367 ( .B1(n14758), .B2(n14757), .A(n14756), .ZN(n15166) );
  INV_X1 U18368 ( .A(n15166), .ZN(n15004) );
  INV_X1 U18369 ( .A(n15164), .ZN(n14759) );
  NAND2_X1 U18370 ( .A1(n21018), .A2(n14759), .ZN(n14760) );
  OAI211_X1 U18371 ( .C1(n20980), .C2(n14761), .A(n14760), .B(n20998), .ZN(
        n14766) );
  INV_X1 U18372 ( .A(n14762), .ZN(n14763) );
  AOI21_X1 U18373 ( .B1(n21418), .B2(n14764), .A(n14763), .ZN(n14765) );
  AOI211_X1 U18374 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n21014), .A(n14766), .B(
        n14765), .ZN(n14769) );
  XNOR2_X1 U18375 ( .A(n14776), .B(n14767), .ZN(n15400) );
  NAND2_X1 U18376 ( .A1(n15400), .A2(n21013), .ZN(n14768) );
  OAI211_X1 U18377 ( .C1(n15004), .C2(n20974), .A(n14769), .B(n14768), .ZN(
        P1_U2823) );
  AOI21_X1 U18378 ( .B1(n14772), .B2(n10086), .A(n14771), .ZN(n15180) );
  INV_X1 U18379 ( .A(n15180), .ZN(n15011) );
  AND2_X1 U18380 ( .A1(n14802), .A2(n14774), .ZN(n14775) );
  NOR2_X1 U18381 ( .A1(n14776), .A2(n14775), .ZN(n15407) );
  NAND2_X1 U18382 ( .A1(n21018), .A2(n15179), .ZN(n14777) );
  OAI211_X1 U18383 ( .C1(n20980), .C2(n15177), .A(n14777), .B(n20998), .ZN(
        n14778) );
  AOI21_X1 U18384 ( .B1(n21014), .B2(P1_EBX_REG_16__SCAN_IN), .A(n14778), .ZN(
        n14783) );
  INV_X1 U18385 ( .A(n14779), .ZN(n14780) );
  OAI211_X1 U18386 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14781), .B(n14780), .ZN(n14782) );
  OAI211_X1 U18387 ( .C1(n17552), .C2(n15175), .A(n14783), .B(n14782), .ZN(
        n14784) );
  AOI21_X1 U18388 ( .B1(n15407), .B2(n21013), .A(n14784), .ZN(n14785) );
  OAI21_X1 U18389 ( .B1(n15011), .B2(n20974), .A(n14785), .ZN(P1_U2824) );
  INV_X1 U18390 ( .A(n14786), .ZN(n14807) );
  INV_X1 U18391 ( .A(n14808), .ZN(n14788) );
  INV_X1 U18392 ( .A(n14809), .ZN(n14945) );
  OR2_X1 U18393 ( .A1(n14848), .A2(n14945), .ZN(n14787) );
  NAND2_X1 U18394 ( .A1(n14788), .A2(n14787), .ZN(n14790) );
  AND2_X1 U18395 ( .A1(n14811), .A2(n14810), .ZN(n14789) );
  NAND2_X1 U18396 ( .A1(n14790), .A2(n14789), .ZN(n14936) );
  INV_X1 U18397 ( .A(n14791), .ZN(n14935) );
  INV_X1 U18398 ( .A(n14938), .ZN(n14793) );
  OAI21_X1 U18399 ( .B1(n14793), .B2(n14792), .A(n10086), .ZN(n15186) );
  INV_X1 U18400 ( .A(n17552), .ZN(n14805) );
  INV_X1 U18401 ( .A(n15189), .ZN(n14794) );
  NAND2_X1 U18402 ( .A1(n9627), .A2(n14794), .ZN(n14795) );
  OAI211_X1 U18403 ( .C1(n20980), .C2(n14796), .A(n14795), .B(n20998), .ZN(
        n14797) );
  AOI21_X1 U18404 ( .B1(n21014), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14797), .ZN(
        n14798) );
  OAI21_X1 U18405 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n14799), .A(n14798), 
        .ZN(n14804) );
  NAND2_X1 U18406 ( .A1(n14941), .A2(n14800), .ZN(n14801) );
  NAND2_X1 U18407 ( .A1(n14802), .A2(n14801), .ZN(n15416) );
  NOR2_X1 U18408 ( .A1(n15416), .A2(n14888), .ZN(n14803) );
  AOI211_X1 U18409 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n14805), .A(n14804), 
        .B(n14803), .ZN(n14806) );
  OAI21_X1 U18410 ( .B1(n15186), .B2(n20974), .A(n14806), .ZN(P1_U2825) );
  AOI21_X1 U18411 ( .B1(n14807), .B2(n14848), .A(n14808), .ZN(n14946) );
  AOI21_X1 U18412 ( .B1(n14946), .B2(n14809), .A(n14808), .ZN(n14833) );
  INV_X1 U18413 ( .A(n14810), .ZN(n14832) );
  NOR2_X1 U18414 ( .A1(n14833), .A2(n14832), .ZN(n14831) );
  INV_X1 U18415 ( .A(n15212), .ZN(n14829) );
  AND2_X1 U18416 ( .A1(n14839), .A2(n14812), .ZN(n14813) );
  OR2_X1 U18417 ( .A1(n14813), .A2(n14940), .ZN(n15440) );
  OAI22_X1 U18418 ( .A1(n15440), .A2(n14888), .B1(n14814), .B2(n21006), .ZN(
        n14815) );
  INV_X1 U18419 ( .A(n14815), .ZN(n14816) );
  OAI211_X1 U18420 ( .C1(n20980), .C2(n14817), .A(n14816), .B(n20998), .ZN(
        n14828) );
  NOR2_X1 U18421 ( .A1(n20970), .A2(n14819), .ZN(n20957) );
  NAND3_X1 U18422 ( .A1(n20957), .A2(P1_REIP_REG_9__SCAN_IN), .A3(
        P1_REIP_REG_10__SCAN_IN), .ZN(n17569) );
  NOR2_X1 U18423 ( .A1(n14818), .A2(n17569), .ZN(n14826) );
  INV_X1 U18424 ( .A(n14819), .ZN(n14820) );
  NAND2_X1 U18425 ( .A1(n14884), .A2(n14820), .ZN(n14821) );
  AND2_X1 U18426 ( .A1(n14915), .A2(n14821), .ZN(n20958) );
  INV_X1 U18427 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21410) );
  INV_X1 U18428 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20956) );
  OR2_X1 U18429 ( .A1(n21410), .A2(n20956), .ZN(n14822) );
  AND2_X1 U18430 ( .A1(n14915), .A2(n14822), .ZN(n14823) );
  NOR2_X1 U18431 ( .A1(n20970), .A2(n17550), .ZN(n14824) );
  NOR2_X1 U18432 ( .A1(n17565), .A2(n14824), .ZN(n14845) );
  INV_X1 U18433 ( .A(n14845), .ZN(n14825) );
  MUX2_X1 U18434 ( .A(n14826), .B(n14825), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14827) );
  AOI211_X1 U18435 ( .C1(n21018), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14830) );
  OAI21_X1 U18436 ( .B1(n15209), .B2(n20974), .A(n14830), .ZN(P1_U2827) );
  INV_X1 U18437 ( .A(n17569), .ZN(n17551) );
  AOI21_X1 U18438 ( .B1(n17551), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U18439 ( .A1(n15221), .A2(n20989), .ZN(n14843) );
  INV_X1 U18440 ( .A(n15219), .ZN(n14834) );
  NAND2_X1 U18441 ( .A1(n21018), .A2(n14834), .ZN(n14835) );
  OAI211_X1 U18442 ( .C1(n20980), .C2(n14836), .A(n14835), .B(n20998), .ZN(
        n14841) );
  NAND2_X1 U18443 ( .A1(n14950), .A2(n14837), .ZN(n14838) );
  NAND2_X1 U18444 ( .A1(n14839), .A2(n14838), .ZN(n15454) );
  NOR2_X1 U18445 ( .A1(n14888), .A2(n15454), .ZN(n14840) );
  AOI211_X1 U18446 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n21014), .A(n14841), .B(
        n14840), .ZN(n14842) );
  OAI211_X1 U18447 ( .C1(n14845), .C2(n14844), .A(n14843), .B(n14842), .ZN(
        P1_U2828) );
  OAI21_X1 U18448 ( .B1(n14847), .B2(n14849), .A(n14848), .ZN(n15239) );
  NAND2_X1 U18449 ( .A1(n21014), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14850) );
  OAI211_X1 U18450 ( .C1(n20983), .C2(n15241), .A(n20998), .B(n14850), .ZN(
        n14856) );
  NAND2_X1 U18451 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20957), .ZN(n14854) );
  OR2_X1 U18452 ( .A1(n14957), .A2(n14851), .ZN(n14852) );
  AND2_X1 U18453 ( .A1(n14948), .A2(n14852), .ZN(n15474) );
  AOI22_X1 U18454 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n21016), .B1(
        n21013), .B2(n15474), .ZN(n14853) );
  OAI21_X1 U18455 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n14854), .A(n14853), 
        .ZN(n14855) );
  AOI211_X1 U18456 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n17565), .A(n14856), 
        .B(n14855), .ZN(n14857) );
  OAI21_X1 U18457 ( .B1(n15239), .B2(n20974), .A(n14857), .ZN(P1_U2830) );
  INV_X1 U18458 ( .A(n14491), .ZN(n14859) );
  OAI21_X1 U18459 ( .B1(n14859), .B2(n10481), .A(n14955), .ZN(n15263) );
  NAND3_X1 U18460 ( .A1(n21002), .A2(n14874), .A3(n14860), .ZN(n14867) );
  INV_X1 U18461 ( .A(n14494), .ZN(n14863) );
  AOI21_X1 U18462 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(n14865) );
  INV_X1 U18463 ( .A(n14958), .ZN(n14864) );
  NOR2_X1 U18464 ( .A1(n14865), .A2(n14864), .ZN(n17596) );
  AOI22_X1 U18465 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n21016), .B1(
        n21013), .B2(n17596), .ZN(n14866) );
  OAI211_X1 U18466 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n14867), .A(n14866), .B(
        n20998), .ZN(n14868) );
  AOI21_X1 U18467 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20958), .A(n14868), .ZN(
        n14871) );
  INV_X1 U18468 ( .A(n15259), .ZN(n14869) );
  AOI22_X1 U18469 ( .A1(n21014), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n21018), .B2(
        n14869), .ZN(n14870) );
  OAI211_X1 U18470 ( .C1(n15263), .C2(n20974), .A(n14871), .B(n14870), .ZN(
        P1_U2832) );
  OR2_X1 U18471 ( .A1(n14886), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U18472 ( .A1(n20974), .A2(n14873), .ZN(n21024) );
  OAI21_X1 U18473 ( .B1(n14874), .B2(n20970), .A(n14884), .ZN(n20972) );
  INV_X1 U18474 ( .A(n20972), .ZN(n21011) );
  NAND2_X1 U18475 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21011), .ZN(n20985) );
  INV_X1 U18476 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n17620) );
  NAND2_X1 U18477 ( .A1(n21002), .A2(n14874), .ZN(n20963) );
  NAND2_X1 U18478 ( .A1(n17620), .A2(n20963), .ZN(n14875) );
  NAND2_X1 U18479 ( .A1(n20985), .A2(n14875), .ZN(n14882) );
  INV_X1 U18480 ( .A(n17590), .ZN(n14876) );
  AND2_X1 U18481 ( .A1(n21018), .A2(n14876), .ZN(n14880) );
  NOR2_X1 U18482 ( .A1(n21006), .A2(n14489), .ZN(n14879) );
  OAI22_X1 U18483 ( .A1(n14877), .A2(n20980), .B1(n14888), .B2(n17621), .ZN(
        n14878) );
  NOR4_X1 U18484 ( .A1(n14880), .A2(n14879), .A3(n20952), .A4(n14878), .ZN(
        n14881) );
  OAI211_X1 U18485 ( .C1(n14918), .C2(n17582), .A(n14882), .B(n14881), .ZN(
        P1_U2835) );
  NAND2_X1 U18486 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14883) );
  NAND2_X1 U18487 ( .A1(n21002), .A2(n14883), .ZN(n21028) );
  AND2_X1 U18488 ( .A1(n21028), .A2(n14884), .ZN(n21021) );
  INV_X1 U18489 ( .A(n21021), .ZN(n14896) );
  OR2_X1 U18490 ( .A1(n14886), .A2(n14885), .ZN(n21020) );
  INV_X1 U18491 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21401) );
  NAND4_X1 U18492 ( .A1(n21002), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n21401), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n14887) );
  OAI21_X1 U18493 ( .B1(n14888), .B2(n21114), .A(n14887), .ZN(n14892) );
  OAI22_X1 U18494 ( .A1(n20983), .A2(n14890), .B1(n14889), .B2(n20980), .ZN(
        n14891) );
  OAI21_X1 U18495 ( .B1(n14894), .B2(n21020), .A(n14893), .ZN(n14895) );
  AOI21_X1 U18496 ( .B1(n14896), .B2(P1_REIP_REG_3__SCAN_IN), .A(n14895), .ZN(
        n14897) );
  OAI21_X1 U18497 ( .B1(n14918), .B2(n14898), .A(n14897), .ZN(P1_U2837) );
  INV_X1 U18498 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14899) );
  OAI22_X1 U18499 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20970), .B1(n21006), 
        .B2(n14899), .ZN(n14906) );
  INV_X1 U18500 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U18501 ( .A1(n21018), .A2(n14901), .ZN(n14904) );
  AOI22_X1 U18502 ( .A1(n21016), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14902), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14903) );
  OAI211_X1 U18503 ( .C1(n21020), .C2(n21206), .A(n14904), .B(n14903), .ZN(
        n14905) );
  AOI211_X1 U18504 ( .C1(n21013), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14908) );
  OAI21_X1 U18505 ( .B1(n14918), .B2(n14909), .A(n14908), .ZN(P1_U2839) );
  AOI22_X1 U18506 ( .A1(n21014), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n21013), .B2(
        n14910), .ZN(n14912) );
  OAI21_X1 U18507 ( .B1(n21018), .B2(n21016), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14911) );
  OAI211_X1 U18508 ( .C1(n21020), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14914) );
  AOI21_X1 U18509 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n14915), .A(n14914), .ZN(
        n14916) );
  OAI21_X1 U18510 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(P1_U2840) );
  OAI22_X1 U18511 ( .A1(n15265), .A2(n14960), .B1(n21035), .B2(n14919), .ZN(
        P1_U2841) );
  INV_X1 U18512 ( .A(n15051), .ZN(n14966) );
  OAI222_X1 U18513 ( .A1(n14966), .A2(n14963), .B1(n14920), .B2(n21035), .C1(
        n15273), .C2(n14960), .ZN(P1_U2843) );
  INV_X1 U18514 ( .A(n15066), .ZN(n14969) );
  OAI222_X1 U18515 ( .A1(n14963), .A2(n14969), .B1(n14921), .B2(n21035), .C1(
        n15287), .C2(n14960), .ZN(P1_U2844) );
  INV_X1 U18516 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14922) );
  OAI222_X1 U18517 ( .A1(n14963), .A2(n15071), .B1(n14922), .B2(n21035), .C1(
        n15292), .C2(n14960), .ZN(P1_U2845) );
  AOI22_X1 U18518 ( .A1(n15308), .A2(n21030), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14961), .ZN(n14923) );
  OAI21_X1 U18519 ( .B1(n15079), .B2(n14963), .A(n14923), .ZN(P1_U2846) );
  OAI222_X1 U18520 ( .A1(n14650), .A2(n14963), .B1(n14925), .B2(n21035), .C1(
        n14924), .C2(n14960), .ZN(P1_U2847) );
  AOI22_X1 U18521 ( .A1(n15327), .A2(n21030), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14961), .ZN(n14926) );
  OAI21_X1 U18522 ( .B1(n14979), .B2(n14963), .A(n14926), .ZN(P1_U2848) );
  OAI222_X1 U18523 ( .A1(n15105), .A2(n14963), .B1(n14927), .B2(n21035), .C1(
        n15348), .C2(n14960), .ZN(P1_U2850) );
  AOI22_X1 U18524 ( .A1(n15357), .A2(n21030), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14961), .ZN(n14928) );
  OAI21_X1 U18525 ( .B1(n14990), .B2(n14963), .A(n14928), .ZN(P1_U2851) );
  AOI22_X1 U18526 ( .A1(n15371), .A2(n21030), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14961), .ZN(n14929) );
  OAI21_X1 U18527 ( .B1(n15131), .B2(n14963), .A(n14929), .ZN(P1_U2852) );
  INV_X1 U18528 ( .A(n15144), .ZN(n14997) );
  OAI222_X1 U18529 ( .A1(n14997), .A2(n14963), .B1(n14930), .B2(n21035), .C1(
        n15374), .C2(n14960), .ZN(P1_U2853) );
  AOI22_X1 U18530 ( .A1(n15391), .A2(n21030), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14961), .ZN(n14931) );
  OAI21_X1 U18531 ( .B1(n15147), .B2(n14963), .A(n14931), .ZN(P1_U2854) );
  AOI22_X1 U18532 ( .A1(n15400), .A2(n21030), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14961), .ZN(n14932) );
  OAI21_X1 U18533 ( .B1(n15004), .B2(n14963), .A(n14932), .ZN(P1_U2855) );
  AOI22_X1 U18534 ( .A1(n15407), .A2(n21030), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14961), .ZN(n14933) );
  OAI21_X1 U18535 ( .B1(n15011), .B2(n14963), .A(n14933), .ZN(P1_U2856) );
  OAI222_X1 U18536 ( .A1(n15186), .A2(n14963), .B1(n14934), .B2(n21035), .C1(
        n15416), .C2(n14960), .ZN(P1_U2857) );
  NAND2_X1 U18537 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  OR2_X1 U18538 ( .A1(n14940), .A2(n14939), .ZN(n14942) );
  AND2_X1 U18539 ( .A1(n14942), .A2(n14941), .ZN(n17549) );
  AOI22_X1 U18540 ( .A1(n17549), .A2(n21030), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14961), .ZN(n14943) );
  OAI21_X1 U18541 ( .B1(n15014), .B2(n14963), .A(n14943), .ZN(P1_U2858) );
  OAI222_X1 U18542 ( .A1(n15209), .A2(n14963), .B1(n21035), .B2(n14814), .C1(
        n15440), .C2(n14960), .ZN(P1_U2859) );
  INV_X1 U18543 ( .A(n15221), .ZN(n15018) );
  INV_X1 U18544 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14944) );
  OAI222_X1 U18545 ( .A1(n15018), .A2(n14963), .B1(n14944), .B2(n21035), .C1(
        n15454), .C2(n14960), .ZN(P1_U2860) );
  XNOR2_X1 U18546 ( .A(n14946), .B(n14945), .ZN(n17566) );
  NAND2_X1 U18547 ( .A1(n17566), .A2(n21031), .ZN(n14952) );
  NAND2_X1 U18548 ( .A1(n14948), .A2(n14947), .ZN(n14949) );
  AND2_X1 U18549 ( .A1(n14950), .A2(n14949), .ZN(n17564) );
  NAND2_X1 U18550 ( .A1(n17564), .A2(n21030), .ZN(n14951) );
  OAI211_X1 U18551 ( .C1(n14953), .C2(n21035), .A(n14952), .B(n14951), .ZN(
        P1_U2861) );
  AOI22_X1 U18552 ( .A1(n15474), .A2(n21030), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14961), .ZN(n14954) );
  OAI21_X1 U18553 ( .B1(n15239), .B2(n14963), .A(n14954), .ZN(P1_U2862) );
  AOI21_X1 U18554 ( .B1(n14956), .B2(n14955), .A(n14847), .ZN(n20959) );
  INV_X1 U18555 ( .A(n20959), .ZN(n15254) );
  AOI21_X1 U18556 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n20950) );
  INV_X1 U18557 ( .A(n20950), .ZN(n15485) );
  OAI222_X1 U18558 ( .A1(n15254), .A2(n14963), .B1(n20954), .B2(n21035), .C1(
        n15485), .C2(n14960), .ZN(P1_U2863) );
  AOI22_X1 U18559 ( .A1(n17596), .A2(n21030), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14961), .ZN(n14962) );
  OAI21_X1 U18560 ( .B1(n15263), .B2(n14963), .A(n14962), .ZN(P1_U2864) );
  AOI22_X1 U18561 ( .A1(n15005), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15022), .ZN(n14965) );
  MUX2_X1 U18562 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14974), .Z(
        n21077) );
  AOI22_X1 U18563 ( .A1(n15008), .A2(n21077), .B1(n15006), .B2(DATAI_29_), 
        .ZN(n14964) );
  OAI211_X1 U18564 ( .C1(n14966), .C2(n15031), .A(n14965), .B(n14964), .ZN(
        P1_U2875) );
  AOI22_X1 U18565 ( .A1(n15005), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15022), .ZN(n14968) );
  AOI22_X1 U18566 ( .A1(n15008), .A2(n15016), .B1(n15006), .B2(DATAI_28_), 
        .ZN(n14967) );
  OAI211_X1 U18567 ( .C1(n14969), .C2(n15031), .A(n14968), .B(n14967), .ZN(
        P1_U2876) );
  AOI22_X1 U18568 ( .A1(n15005), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15022), .ZN(n14971) );
  MUX2_X1 U18569 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14974), .Z(
        n21075) );
  AOI22_X1 U18570 ( .A1(n15008), .A2(n21075), .B1(n15006), .B2(DATAI_27_), 
        .ZN(n14970) );
  OAI211_X1 U18571 ( .C1(n15071), .C2(n15031), .A(n14971), .B(n14970), .ZN(
        P1_U2877) );
  AOI22_X1 U18572 ( .A1(n15005), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15022), .ZN(n14973) );
  MUX2_X1 U18573 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14974), .Z(
        n21073) );
  AOI22_X1 U18574 ( .A1(n15008), .A2(n21073), .B1(n15006), .B2(DATAI_26_), 
        .ZN(n14972) );
  OAI211_X1 U18575 ( .C1(n15079), .C2(n15031), .A(n14973), .B(n14972), .ZN(
        P1_U2878) );
  AOI22_X1 U18576 ( .A1(n15005), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15022), .ZN(n14976) );
  MUX2_X1 U18577 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14974), .Z(
        n21071) );
  AOI22_X1 U18578 ( .A1(n15008), .A2(n21071), .B1(n15006), .B2(DATAI_25_), 
        .ZN(n14975) );
  OAI211_X1 U18579 ( .C1(n14650), .C2(n15031), .A(n14976), .B(n14975), .ZN(
        P1_U2879) );
  AOI22_X1 U18580 ( .A1(n15005), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15022), .ZN(n14978) );
  AOI22_X1 U18581 ( .A1(n15008), .A2(n15025), .B1(n15006), .B2(DATAI_24_), 
        .ZN(n14977) );
  OAI211_X1 U18582 ( .C1(n14979), .C2(n15031), .A(n14978), .B(n14977), .ZN(
        P1_U2880) );
  AOI22_X1 U18583 ( .A1(n15005), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15022), .ZN(n14982) );
  AOI22_X1 U18584 ( .A1(n15008), .A2(n14980), .B1(n15006), .B2(DATAI_23_), 
        .ZN(n14981) );
  OAI211_X1 U18585 ( .C1(n14983), .C2(n15031), .A(n14982), .B(n14981), .ZN(
        P1_U2881) );
  AOI22_X1 U18586 ( .A1(n15005), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15022), .ZN(n14986) );
  AOI22_X1 U18587 ( .A1(n15008), .A2(n14984), .B1(n15006), .B2(DATAI_22_), 
        .ZN(n14985) );
  OAI211_X1 U18588 ( .C1(n15105), .C2(n15031), .A(n14986), .B(n14985), .ZN(
        P1_U2882) );
  AOI22_X1 U18589 ( .A1(n15005), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15022), .ZN(n14989) );
  AOI22_X1 U18590 ( .A1(n15008), .A2(n14987), .B1(n15006), .B2(DATAI_21_), 
        .ZN(n14988) );
  OAI211_X1 U18591 ( .C1(n14990), .C2(n15031), .A(n14989), .B(n14988), .ZN(
        P1_U2883) );
  AOI22_X1 U18592 ( .A1(n15005), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15022), .ZN(n14993) );
  AOI22_X1 U18593 ( .A1(n15008), .A2(n14991), .B1(n15006), .B2(DATAI_20_), 
        .ZN(n14992) );
  OAI211_X1 U18594 ( .C1(n15131), .C2(n15031), .A(n14993), .B(n14992), .ZN(
        P1_U2884) );
  AOI22_X1 U18595 ( .A1(n15005), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15022), .ZN(n14996) );
  AOI22_X1 U18596 ( .A1(n15008), .A2(n14994), .B1(n15006), .B2(DATAI_19_), 
        .ZN(n14995) );
  OAI211_X1 U18597 ( .C1(n14997), .C2(n15031), .A(n14996), .B(n14995), .ZN(
        P1_U2885) );
  AOI22_X1 U18598 ( .A1(n15005), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15022), .ZN(n15000) );
  AOI22_X1 U18599 ( .A1(n15008), .A2(n14998), .B1(n15006), .B2(DATAI_18_), 
        .ZN(n14999) );
  OAI211_X1 U18600 ( .C1(n15147), .C2(n15031), .A(n15000), .B(n14999), .ZN(
        P1_U2886) );
  AOI22_X1 U18601 ( .A1(n15005), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n15022), .ZN(n15003) );
  AOI22_X1 U18602 ( .A1(n15008), .A2(n15001), .B1(n15006), .B2(DATAI_17_), 
        .ZN(n15002) );
  OAI211_X1 U18603 ( .C1(n15004), .C2(n15031), .A(n15003), .B(n15002), .ZN(
        P1_U2887) );
  AOI22_X1 U18604 ( .A1(n15005), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15022), .ZN(n15010) );
  AOI22_X1 U18605 ( .A1(n15008), .A2(n15007), .B1(n15006), .B2(DATAI_16_), 
        .ZN(n15009) );
  OAI211_X1 U18606 ( .C1(n15011), .C2(n15031), .A(n15010), .B(n15009), .ZN(
        P1_U2888) );
  OAI222_X1 U18607 ( .A1(n15031), .A2(n15186), .B1(n15033), .B2(n15012), .C1(
        n21037), .C2(n15029), .ZN(P1_U2889) );
  AOI22_X1 U18608 ( .A1(n15023), .A2(n21079), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15022), .ZN(n15013) );
  OAI21_X1 U18609 ( .B1(n15014), .B2(n15031), .A(n15013), .ZN(P1_U2890) );
  AOI22_X1 U18610 ( .A1(n15023), .A2(n21077), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15022), .ZN(n15015) );
  OAI21_X1 U18611 ( .B1(n15209), .B2(n15031), .A(n15015), .ZN(P1_U2891) );
  INV_X1 U18612 ( .A(n15016), .ZN(n15017) );
  OAI222_X1 U18613 ( .A1(n15018), .A2(n15031), .B1(n21043), .B2(n15029), .C1(
        n15033), .C2(n15017), .ZN(P1_U2892) );
  INV_X1 U18614 ( .A(n17566), .ZN(n15020) );
  AOI22_X1 U18615 ( .A1(n15023), .A2(n21075), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15022), .ZN(n15019) );
  OAI21_X1 U18616 ( .B1(n15020), .B2(n15031), .A(n15019), .ZN(P1_U2893) );
  AOI22_X1 U18617 ( .A1(n15023), .A2(n21073), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15022), .ZN(n15021) );
  OAI21_X1 U18618 ( .B1(n15239), .B2(n15031), .A(n15021), .ZN(P1_U2894) );
  AOI22_X1 U18619 ( .A1(n15023), .A2(n21071), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15022), .ZN(n15024) );
  OAI21_X1 U18620 ( .B1(n15254), .B2(n15031), .A(n15024), .ZN(P1_U2895) );
  INV_X1 U18621 ( .A(n15025), .ZN(n15026) );
  OAI222_X1 U18622 ( .A1(n15031), .A2(n15263), .B1(n15029), .B2(n21052), .C1(
        n15033), .C2(n15026), .ZN(P1_U2896) );
  XOR2_X1 U18623 ( .A(n15028), .B(n15027), .Z(n21032) );
  INV_X1 U18624 ( .A(n21032), .ZN(n15030) );
  OAI222_X1 U18625 ( .A1(n15033), .A2(n15032), .B1(n15031), .B2(n15030), .C1(
        n21057), .C2(n15029), .ZN(P1_U2898) );
  INV_X1 U18626 ( .A(n15034), .ZN(n15035) );
  NAND2_X1 U18627 ( .A1(n15035), .A2(n10334), .ZN(n15037) );
  NAND2_X1 U18628 ( .A1(n21133), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U18629 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15039) );
  OAI211_X1 U18630 ( .C1(n15040), .C2(n21106), .A(n15268), .B(n15039), .ZN(
        n15041) );
  NAND2_X1 U18631 ( .A1(n15045), .A2(n15044), .ZN(n15046) );
  XNOR2_X1 U18632 ( .A(n15047), .B(n15046), .ZN(n15282) );
  NOR2_X1 U18633 ( .A1(n15176), .A2(n21437), .ZN(n15274) );
  AOI21_X1 U18634 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15274), .ZN(n15048) );
  OAI21_X1 U18635 ( .B1(n21106), .B2(n15049), .A(n15048), .ZN(n15050) );
  AOI21_X1 U18636 ( .B1(n15051), .B2(n21101), .A(n15050), .ZN(n15052) );
  OAI21_X1 U18637 ( .B1(n20932), .B2(n15282), .A(n15052), .ZN(P1_U2970) );
  INV_X1 U18638 ( .A(n15053), .ZN(n15054) );
  MUX2_X1 U18639 ( .A(n15054), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15227), .Z(n15059) );
  NAND2_X1 U18640 ( .A1(n15303), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15057) );
  INV_X1 U18641 ( .A(n15055), .ZN(n15056) );
  OAI21_X1 U18642 ( .B1(n12991), .B2(n15057), .A(n15056), .ZN(n15058) );
  NAND2_X1 U18643 ( .A1(n15059), .A2(n15058), .ZN(n15061) );
  XNOR2_X1 U18644 ( .A(n15061), .B(n15060), .ZN(n15291) );
  INV_X1 U18645 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n15062) );
  NOR2_X1 U18646 ( .A1(n15176), .A2(n15062), .ZN(n15286) );
  AOI21_X1 U18647 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15286), .ZN(n15063) );
  OAI21_X1 U18648 ( .B1(n21106), .B2(n15064), .A(n15063), .ZN(n15065) );
  AOI21_X1 U18649 ( .B1(n15066), .B2(n21101), .A(n15065), .ZN(n15067) );
  OAI21_X1 U18650 ( .B1(n20932), .B2(n15291), .A(n15067), .ZN(P1_U2971) );
  MUX2_X1 U18651 ( .A(n15069), .B(n15068), .S(n10334), .Z(n15070) );
  XNOR2_X1 U18652 ( .A(n15070), .B(n15297), .ZN(n15302) );
  INV_X1 U18653 ( .A(n15071), .ZN(n15075) );
  INV_X1 U18654 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21434) );
  NOR2_X1 U18655 ( .A1(n15176), .A2(n21434), .ZN(n15294) );
  AOI21_X1 U18656 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15294), .ZN(n15072) );
  OAI21_X1 U18657 ( .B1(n21106), .B2(n15073), .A(n15072), .ZN(n15074) );
  AOI21_X1 U18658 ( .B1(n15075), .B2(n21101), .A(n15074), .ZN(n15076) );
  OAI21_X1 U18659 ( .B1(n20932), .B2(n15302), .A(n15076), .ZN(P1_U2972) );
  OAI211_X1 U18660 ( .C1(n10334), .C2(n15303), .A(n15077), .B(n15084), .ZN(
        n15078) );
  XOR2_X1 U18661 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15078), .Z(
        n15310) );
  NOR2_X1 U18662 ( .A1(n15176), .A2(n15080), .ZN(n15307) );
  AOI21_X1 U18663 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15307), .ZN(n15081) );
  OAI21_X1 U18664 ( .B1(n21106), .B2(n15082), .A(n15081), .ZN(n15083) );
  XNOR2_X1 U18665 ( .A(n15245), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15095) );
  NAND3_X1 U18666 ( .A1(n15085), .A2(n15095), .A3(n15084), .ZN(n15087) );
  XNOR2_X1 U18667 ( .A(n15087), .B(n15086), .ZN(n15330) );
  INV_X1 U18668 ( .A(n15088), .ZN(n15091) );
  NOR2_X1 U18669 ( .A1(n15176), .A2(n15089), .ZN(n15325) );
  AOI21_X1 U18670 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15325), .ZN(n15090) );
  OAI21_X1 U18671 ( .B1(n21106), .B2(n15091), .A(n15090), .ZN(n15092) );
  AOI21_X1 U18672 ( .B1(n15093), .B2(n21101), .A(n15092), .ZN(n15094) );
  OAI21_X1 U18673 ( .B1(n20932), .B2(n15330), .A(n15094), .ZN(P1_U2975) );
  XNOR2_X1 U18674 ( .A(n9923), .B(n15095), .ZN(n15338) );
  INV_X1 U18675 ( .A(n15096), .ZN(n15098) );
  INV_X1 U18676 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21427) );
  NOR2_X1 U18677 ( .A1(n15176), .A2(n21427), .ZN(n15333) );
  AOI21_X1 U18678 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15333), .ZN(n15097) );
  OAI21_X1 U18679 ( .B1(n21106), .B2(n15098), .A(n15097), .ZN(n15099) );
  AOI21_X1 U18680 ( .B1(n15100), .B2(n21101), .A(n15099), .ZN(n15101) );
  OAI21_X1 U18681 ( .B1(n15338), .B2(n20932), .A(n15101), .ZN(P1_U2976) );
  NAND2_X1 U18682 ( .A1(n15102), .A2(n15103), .ZN(n15104) );
  XOR2_X1 U18683 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15104), .Z(
        n15352) );
  INV_X1 U18684 ( .A(n15105), .ZN(n15111) );
  INV_X1 U18685 ( .A(n15106), .ZN(n15109) );
  INV_X1 U18686 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U18687 ( .A1(n15176), .A2(n15107), .ZN(n15347) );
  AOI21_X1 U18688 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15347), .ZN(n15108) );
  OAI21_X1 U18689 ( .B1(n21106), .B2(n15109), .A(n15108), .ZN(n15110) );
  AOI21_X1 U18690 ( .B1(n15111), .B2(n21101), .A(n15110), .ZN(n15112) );
  OAI21_X1 U18691 ( .B1(n20932), .B2(n15352), .A(n15112), .ZN(P1_U2977) );
  OR2_X1 U18692 ( .A1(n15245), .A2(n15113), .ZN(n15114) );
  AND2_X1 U18693 ( .A1(n15115), .A2(n15114), .ZN(n15140) );
  NOR2_X1 U18694 ( .A1(n15245), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15138) );
  INV_X1 U18695 ( .A(n15116), .ZN(n15118) );
  INV_X1 U18696 ( .A(n15146), .ZN(n15117) );
  NAND2_X1 U18697 ( .A1(n15227), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15136) );
  AOI21_X1 U18698 ( .B1(n15140), .B2(n15138), .A(n15119), .ZN(n15129) );
  NOR2_X1 U18699 ( .A1(n15129), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15128) );
  AOI22_X1 U18700 ( .A1(n15128), .A2(n10334), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15119), .ZN(n15121) );
  XNOR2_X1 U18701 ( .A(n15121), .B(n15120), .ZN(n15360) );
  INV_X1 U18702 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U18703 ( .A1(n15176), .A2(n15122), .ZN(n15355) );
  AOI21_X1 U18704 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15355), .ZN(n15123) );
  OAI21_X1 U18705 ( .B1(n21106), .B2(n15124), .A(n15123), .ZN(n15125) );
  AOI21_X1 U18706 ( .B1(n15126), .B2(n21101), .A(n15125), .ZN(n15127) );
  OAI21_X1 U18707 ( .B1(n15360), .B2(n20932), .A(n15127), .ZN(P1_U2978) );
  AOI21_X1 U18708 ( .B1(n15129), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15128), .ZN(n15373) );
  OR2_X1 U18709 ( .A1(n15176), .A2(n21423), .ZN(n15367) );
  OAI21_X1 U18710 ( .B1(n15249), .B2(n15130), .A(n15367), .ZN(n15133) );
  NOR2_X1 U18711 ( .A1(n15131), .A2(n15264), .ZN(n15132) );
  AOI211_X1 U18712 ( .C1(n15251), .C2(n15134), .A(n15133), .B(n15132), .ZN(
        n15135) );
  OAI21_X1 U18713 ( .B1(n15373), .B2(n20932), .A(n15135), .ZN(P1_U2979) );
  INV_X1 U18714 ( .A(n15136), .ZN(n15137) );
  NOR2_X1 U18715 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  XNOR2_X1 U18716 ( .A(n15140), .B(n15139), .ZN(n15382) );
  INV_X1 U18717 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21420) );
  NOR2_X1 U18718 ( .A1(n15176), .A2(n21420), .ZN(n15375) );
  AOI21_X1 U18719 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15375), .ZN(n15141) );
  OAI21_X1 U18720 ( .B1(n21106), .B2(n15142), .A(n15141), .ZN(n15143) );
  AOI21_X1 U18721 ( .B1(n15144), .B2(n21101), .A(n15143), .ZN(n15145) );
  OAI21_X1 U18722 ( .B1(n20932), .B2(n15382), .A(n15145), .ZN(P1_U2980) );
  XNOR2_X1 U18723 ( .A(n15116), .B(n15146), .ZN(n15394) );
  INV_X1 U18724 ( .A(n15147), .ZN(n15152) );
  NOR2_X1 U18725 ( .A1(n15176), .A2(n15148), .ZN(n15390) );
  AOI21_X1 U18726 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15390), .ZN(n15149) );
  OAI21_X1 U18727 ( .B1(n21106), .B2(n15150), .A(n15149), .ZN(n15151) );
  AOI21_X1 U18728 ( .B1(n15152), .B2(n21101), .A(n15151), .ZN(n15153) );
  OAI21_X1 U18729 ( .B1(n15394), .B2(n20932), .A(n15153), .ZN(P1_U2981) );
  INV_X1 U18730 ( .A(n15155), .ZN(n15156) );
  NAND2_X1 U18731 ( .A1(n15154), .A2(n15156), .ZN(n15196) );
  OAI21_X1 U18732 ( .B1(n15196), .B2(n15158), .A(n15157), .ZN(n15161) );
  NAND2_X1 U18733 ( .A1(n15161), .A2(n15159), .ZN(n15160) );
  MUX2_X1 U18734 ( .A(n15161), .B(n15160), .S(n10334), .Z(n15162) );
  XNOR2_X1 U18735 ( .A(n15162), .B(n15395), .ZN(n15403) );
  NOR2_X1 U18736 ( .A1(n15176), .A2(n21418), .ZN(n15397) );
  AOI21_X1 U18737 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15397), .ZN(n15163) );
  OAI21_X1 U18738 ( .B1(n21106), .B2(n15164), .A(n15163), .ZN(n15165) );
  AOI21_X1 U18739 ( .B1(n15166), .B2(n21101), .A(n15165), .ZN(n15167) );
  OAI21_X1 U18740 ( .B1(n20932), .B2(n15403), .A(n15167), .ZN(P1_U2982) );
  OAI21_X1 U18741 ( .B1(n15154), .B2(n15168), .A(n10476), .ZN(n15185) );
  INV_X1 U18742 ( .A(n15169), .ZN(n15170) );
  NAND2_X1 U18743 ( .A1(n15170), .A2(n15171), .ZN(n15184) );
  NOR2_X1 U18744 ( .A1(n15185), .A2(n15184), .ZN(n15183) );
  INV_X1 U18745 ( .A(n15171), .ZN(n15172) );
  NOR2_X1 U18746 ( .A1(n15183), .A2(n15172), .ZN(n15174) );
  XNOR2_X1 U18747 ( .A(n15174), .B(n15173), .ZN(n15413) );
  NOR2_X1 U18748 ( .A1(n15176), .A2(n15175), .ZN(n15406) );
  NOR2_X1 U18749 ( .A1(n15249), .A2(n15177), .ZN(n15178) );
  AOI211_X1 U18750 ( .C1(n15251), .C2(n15179), .A(n15406), .B(n15178), .ZN(
        n15182) );
  NAND2_X1 U18751 ( .A1(n15180), .A2(n21101), .ZN(n15181) );
  OAI211_X1 U18752 ( .C1(n15413), .C2(n20932), .A(n15182), .B(n15181), .ZN(
        P1_U2983) );
  AOI21_X1 U18753 ( .B1(n15185), .B2(n15184), .A(n15183), .ZN(n15421) );
  INV_X1 U18754 ( .A(n15186), .ZN(n15191) );
  NOR2_X1 U18755 ( .A1(n15176), .A2(n15187), .ZN(n15414) );
  AOI21_X1 U18756 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15414), .ZN(n15188) );
  OAI21_X1 U18757 ( .B1(n21106), .B2(n15189), .A(n15188), .ZN(n15190) );
  AOI21_X1 U18758 ( .B1(n15191), .B2(n21101), .A(n15190), .ZN(n15192) );
  OAI21_X1 U18759 ( .B1(n15421), .B2(n20932), .A(n15192), .ZN(P1_U2984) );
  AND2_X1 U18760 ( .A1(n15227), .A2(n15193), .ZN(n15204) );
  INV_X1 U18761 ( .A(n12586), .ZN(n15194) );
  AOI21_X1 U18762 ( .B1(n15196), .B2(n15195), .A(n15194), .ZN(n15198) );
  XNOR2_X1 U18763 ( .A(n10334), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15197) );
  XNOR2_X1 U18764 ( .A(n15198), .B(n15197), .ZN(n15431) );
  INV_X1 U18765 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n17553) );
  NOR2_X1 U18766 ( .A1(n15176), .A2(n17553), .ZN(n15422) );
  AOI21_X1 U18767 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15422), .ZN(n15199) );
  OAI21_X1 U18768 ( .B1(n21106), .B2(n17547), .A(n15199), .ZN(n15200) );
  AOI21_X1 U18769 ( .B1(n17556), .B2(n21101), .A(n15200), .ZN(n15201) );
  OAI21_X1 U18770 ( .B1(n15431), .B2(n20932), .A(n15201), .ZN(P1_U2985) );
  INV_X1 U18771 ( .A(n15202), .ZN(n15203) );
  OAI22_X1 U18772 ( .A1(n15154), .A2(n15204), .B1(n15203), .B2(n15245), .ZN(
        n15216) );
  INV_X1 U18773 ( .A(n15206), .ZN(n15205) );
  OAI21_X1 U18774 ( .B1(n15245), .B2(n15449), .A(n15205), .ZN(n15215) );
  NOR2_X1 U18775 ( .A1(n15216), .A2(n15215), .ZN(n15214) );
  NOR2_X1 U18776 ( .A1(n15214), .A2(n15206), .ZN(n15207) );
  XOR2_X1 U18777 ( .A(n15208), .B(n15207), .Z(n15446) );
  INV_X1 U18778 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15210) );
  NOR2_X1 U18779 ( .A1(n15176), .A2(n15210), .ZN(n15432) );
  AOI21_X1 U18780 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15432), .ZN(n15211) );
  OAI21_X1 U18781 ( .B1(n21106), .B2(n15212), .A(n15211), .ZN(n15213) );
  AOI21_X1 U18782 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15458) );
  INV_X1 U18783 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15217) );
  NOR2_X1 U18784 ( .A1(n15176), .A2(n15217), .ZN(n15451) );
  AOI21_X1 U18785 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15451), .ZN(n15218) );
  OAI21_X1 U18786 ( .B1(n21106), .B2(n15219), .A(n15218), .ZN(n15220) );
  AOI21_X1 U18787 ( .B1(n15221), .B2(n21101), .A(n15220), .ZN(n15222) );
  OAI21_X1 U18788 ( .B1(n15458), .B2(n20932), .A(n15222), .ZN(P1_U2987) );
  INV_X1 U18789 ( .A(n15223), .ZN(n15225) );
  NOR2_X1 U18790 ( .A1(n10334), .A2(n15224), .ZN(n15256) );
  AOI21_X1 U18791 ( .B1(n15225), .B2(n15255), .A(n15256), .ZN(n15226) );
  AOI21_X1 U18792 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15223), .A(
        n15226), .ZN(n15247) );
  NAND2_X1 U18793 ( .A1(n15247), .A2(n15491), .ZN(n15234) );
  NOR3_X1 U18794 ( .A1(n15234), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15227), .ZN(n15238) );
  NOR3_X1 U18795 ( .A1(n15154), .A2(n10334), .A3(n15478), .ZN(n15228) );
  NOR2_X1 U18796 ( .A1(n15238), .A2(n15228), .ZN(n15229) );
  XNOR2_X1 U18797 ( .A(n15229), .B(n15459), .ZN(n15466) );
  INV_X1 U18798 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15230) );
  NOR2_X1 U18799 ( .A1(n15176), .A2(n15230), .ZN(n15462) );
  AOI21_X1 U18800 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15462), .ZN(n15231) );
  OAI21_X1 U18801 ( .B1(n21106), .B2(n17562), .A(n15231), .ZN(n15232) );
  AOI21_X1 U18802 ( .B1(n17566), .B2(n21101), .A(n15232), .ZN(n15233) );
  OAI21_X1 U18803 ( .B1(n15466), .B2(n20932), .A(n15233), .ZN(P1_U2988) );
  XNOR2_X1 U18804 ( .A(n15154), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15236) );
  AND2_X1 U18805 ( .A1(n15234), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15235) );
  MUX2_X1 U18806 ( .A(n15236), .B(n15235), .S(n10334), .Z(n15237) );
  NOR2_X1 U18807 ( .A1(n15238), .A2(n15237), .ZN(n15481) );
  INV_X1 U18808 ( .A(n15239), .ZN(n15243) );
  NOR2_X1 U18809 ( .A1(n15176), .A2(n21410), .ZN(n15473) );
  AOI21_X1 U18810 ( .B1(n21094), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15473), .ZN(n15240) );
  OAI21_X1 U18811 ( .B1(n21106), .B2(n15241), .A(n15240), .ZN(n15242) );
  AOI21_X1 U18812 ( .B1(n15243), .B2(n21101), .A(n15242), .ZN(n15244) );
  OAI21_X1 U18813 ( .B1(n15481), .B2(n20932), .A(n15244), .ZN(P1_U2989) );
  XNOR2_X1 U18814 ( .A(n15245), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15246) );
  XNOR2_X1 U18815 ( .A(n15247), .B(n15246), .ZN(n15483) );
  NAND2_X1 U18816 ( .A1(n15483), .A2(n21102), .ZN(n15253) );
  NOR2_X1 U18817 ( .A1(n15176), .A2(n20956), .ZN(n15487) );
  NOR2_X1 U18818 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  AOI211_X1 U18819 ( .C1(n15251), .C2(n20951), .A(n15487), .B(n15250), .ZN(
        n15252) );
  OAI211_X1 U18820 ( .C1(n15264), .C2(n15254), .A(n15253), .B(n15252), .ZN(
        P1_U2990) );
  XNOR2_X1 U18821 ( .A(n15256), .B(n15255), .ZN(n15257) );
  XNOR2_X1 U18822 ( .A(n15223), .B(n15257), .ZN(n17602) );
  NAND2_X1 U18823 ( .A1(n17602), .A2(n21102), .ZN(n15262) );
  INV_X1 U18824 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15258) );
  NOR2_X1 U18825 ( .A1(n15176), .A2(n15258), .ZN(n17595) );
  NOR2_X1 U18826 ( .A1(n21106), .A2(n15259), .ZN(n15260) );
  AOI211_X1 U18827 ( .C1(n21094), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17595), .B(n15260), .ZN(n15261) );
  OAI211_X1 U18828 ( .C1(n15264), .C2(n15263), .A(n15262), .B(n15261), .ZN(
        P1_U2991) );
  INV_X1 U18829 ( .A(n15265), .ZN(n15271) );
  NAND3_X1 U18830 ( .A1(n9931), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15269) );
  INV_X1 U18831 ( .A(n15273), .ZN(n15280) );
  INV_X1 U18832 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15277) );
  AOI21_X1 U18833 ( .B1(n15275), .B2(n15277), .A(n15274), .ZN(n15276) );
  OAI21_X1 U18834 ( .B1(n15278), .B2(n15277), .A(n15276), .ZN(n15279) );
  AOI21_X1 U18835 ( .B1(n15280), .B2(n21142), .A(n15279), .ZN(n15281) );
  OAI21_X1 U18836 ( .B1(n15282), .B2(n15482), .A(n15281), .ZN(P1_U3002) );
  INV_X1 U18837 ( .A(n15295), .ZN(n15284) );
  XNOR2_X1 U18838 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15283) );
  NOR2_X1 U18839 ( .A1(n15284), .A2(n15283), .ZN(n15285) );
  AOI211_X1 U18840 ( .C1(n15293), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15286), .B(n15285), .ZN(n15290) );
  INV_X1 U18841 ( .A(n15287), .ZN(n15288) );
  NAND2_X1 U18842 ( .A1(n15288), .A2(n21142), .ZN(n15289) );
  OAI211_X1 U18843 ( .C1(n15291), .C2(n15482), .A(n15290), .B(n15289), .ZN(
        P1_U3003) );
  INV_X1 U18844 ( .A(n15292), .ZN(n15300) );
  INV_X1 U18845 ( .A(n15293), .ZN(n15298) );
  AOI21_X1 U18846 ( .B1(n15295), .B2(n15297), .A(n15294), .ZN(n15296) );
  OAI21_X1 U18847 ( .B1(n15298), .B2(n15297), .A(n15296), .ZN(n15299) );
  AOI21_X1 U18848 ( .B1(n15300), .B2(n21142), .A(n15299), .ZN(n15301) );
  OAI21_X1 U18849 ( .B1(n15302), .B2(n15482), .A(n15301), .ZN(P1_U3004) );
  INV_X1 U18850 ( .A(n15331), .ZN(n15311) );
  AOI21_X1 U18851 ( .B1(n15311), .B2(n15303), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15304) );
  NOR2_X1 U18852 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  AOI211_X1 U18853 ( .C1(n15308), .C2(n21142), .A(n15307), .B(n15306), .ZN(
        n15309) );
  OAI21_X1 U18854 ( .B1(n15310), .B2(n15482), .A(n15309), .ZN(P1_U3005) );
  NAND3_X1 U18855 ( .A1(n15311), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15314) );
  INV_X1 U18856 ( .A(n15312), .ZN(n15313) );
  AOI21_X1 U18857 ( .B1(n15315), .B2(n15314), .A(n15313), .ZN(n15316) );
  AOI211_X1 U18858 ( .C1(n15318), .C2(n21142), .A(n15317), .B(n15316), .ZN(
        n15319) );
  OAI21_X1 U18859 ( .B1(n15320), .B2(n15482), .A(n15319), .ZN(P1_U3006) );
  OAI21_X1 U18860 ( .B1(n15322), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15321), .ZN(n15326) );
  NOR3_X1 U18861 ( .A1(n15331), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15323), .ZN(n15324) );
  AOI211_X1 U18862 ( .C1(n15326), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15325), .B(n15324), .ZN(n15329) );
  NAND2_X1 U18863 ( .A1(n15327), .A2(n21142), .ZN(n15328) );
  OAI211_X1 U18864 ( .C1(n15330), .C2(n15482), .A(n15329), .B(n15328), .ZN(
        P1_U3007) );
  NOR2_X1 U18865 ( .A1(n15331), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15332) );
  AOI211_X1 U18866 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15334), .A(
        n15333), .B(n15332), .ZN(n15337) );
  NAND2_X1 U18867 ( .A1(n15335), .A2(n21142), .ZN(n15336) );
  OAI211_X1 U18868 ( .C1(n15338), .C2(n15482), .A(n15337), .B(n15336), .ZN(
        P1_U3008) );
  INV_X1 U18869 ( .A(n15339), .ZN(n15356) );
  NAND2_X1 U18870 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15442), .ZN(
        n15341) );
  NAND2_X1 U18871 ( .A1(n15450), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15340) );
  OAI22_X1 U18872 ( .A1(n15342), .A2(n15341), .B1(n17600), .B2(n15340), .ZN(
        n15437) );
  AND2_X1 U18873 ( .A1(n15437), .A2(n15343), .ZN(n15363) );
  AOI21_X1 U18874 ( .B1(n15362), .B2(n15344), .A(n15363), .ZN(n15378) );
  XNOR2_X1 U18875 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15345) );
  NOR3_X1 U18876 ( .A1(n15378), .A2(n15353), .A3(n15345), .ZN(n15346) );
  AOI211_X1 U18877 ( .C1(n15356), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15347), .B(n15346), .ZN(n15351) );
  INV_X1 U18878 ( .A(n15348), .ZN(n15349) );
  NAND2_X1 U18879 ( .A1(n15349), .A2(n21142), .ZN(n15350) );
  OAI211_X1 U18880 ( .C1(n15352), .C2(n15482), .A(n15351), .B(n15350), .ZN(
        P1_U3009) );
  NOR3_X1 U18881 ( .A1(n15378), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15353), .ZN(n15354) );
  AOI211_X1 U18882 ( .C1(n15356), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15355), .B(n15354), .ZN(n15359) );
  NAND2_X1 U18883 ( .A1(n15357), .A2(n21142), .ZN(n15358) );
  OAI211_X1 U18884 ( .C1(n15360), .C2(n15482), .A(n15359), .B(n15358), .ZN(
        P1_U3010) );
  OAI21_X1 U18885 ( .B1(n15363), .B2(n15362), .A(n15361), .ZN(n15365) );
  INV_X1 U18886 ( .A(n15376), .ZN(n15364) );
  AOI21_X1 U18887 ( .B1(n15365), .B2(n15364), .A(n15366), .ZN(n15370) );
  NAND2_X1 U18888 ( .A1(n15366), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15368) );
  OAI21_X1 U18889 ( .B1(n15378), .B2(n15368), .A(n15367), .ZN(n15369) );
  AOI211_X1 U18890 ( .C1(n15371), .C2(n21142), .A(n15370), .B(n15369), .ZN(
        n15372) );
  OAI21_X1 U18891 ( .B1(n15373), .B2(n15482), .A(n15372), .ZN(P1_U3011) );
  INV_X1 U18892 ( .A(n15374), .ZN(n15380) );
  AOI21_X1 U18893 ( .B1(n15376), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15375), .ZN(n15377) );
  OAI21_X1 U18894 ( .B1(n15378), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15377), .ZN(n15379) );
  AOI21_X1 U18895 ( .B1(n15380), .B2(n21142), .A(n15379), .ZN(n15381) );
  OAI21_X1 U18896 ( .B1(n15382), .B2(n15482), .A(n15381), .ZN(P1_U3012) );
  NAND2_X1 U18897 ( .A1(n15468), .A2(n15383), .ZN(n15386) );
  INV_X1 U18898 ( .A(n15424), .ZN(n15384) );
  NAND2_X1 U18899 ( .A1(n21127), .A2(n15384), .ZN(n15385) );
  OAI21_X1 U18900 ( .B1(n17601), .B2(n15387), .A(n15428), .ZN(n15398) );
  INV_X1 U18901 ( .A(n15410), .ZN(n15404) );
  NOR3_X1 U18902 ( .A1(n15404), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15388), .ZN(n15389) );
  AOI211_X1 U18903 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15398), .A(
        n15390), .B(n15389), .ZN(n15393) );
  NAND2_X1 U18904 ( .A1(n15391), .A2(n21142), .ZN(n15392) );
  OAI211_X1 U18905 ( .C1(n15394), .C2(n15482), .A(n15393), .B(n15392), .ZN(
        P1_U3013) );
  NAND3_X1 U18906 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15396) );
  OAI21_X1 U18907 ( .B1(n15404), .B2(n15396), .A(n15395), .ZN(n15399) );
  AOI21_X1 U18908 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(n15402) );
  NAND2_X1 U18909 ( .A1(n15400), .A2(n21142), .ZN(n15401) );
  OAI211_X1 U18910 ( .C1(n15403), .C2(n15482), .A(n15402), .B(n15401), .ZN(
        P1_U3014) );
  NOR4_X1 U18911 ( .A1(n15404), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15427), .A4(n15408), .ZN(n15405) );
  AOI211_X1 U18912 ( .C1(n21142), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15412) );
  AND2_X1 U18913 ( .A1(n15408), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15409) );
  AND2_X1 U18914 ( .A1(n15410), .A2(n15409), .ZN(n15418) );
  OAI21_X1 U18915 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17601), .A(
        n15428), .ZN(n15419) );
  OAI21_X1 U18916 ( .B1(n15418), .B2(n15419), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15411) );
  OAI211_X1 U18917 ( .C1(n15413), .C2(n15482), .A(n15412), .B(n15411), .ZN(
        P1_U3015) );
  INV_X1 U18918 ( .A(n15414), .ZN(n15415) );
  OAI21_X1 U18919 ( .B1(n15416), .B2(n17622), .A(n15415), .ZN(n15417) );
  AOI211_X1 U18920 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15419), .A(
        n15418), .B(n15417), .ZN(n15420) );
  OAI21_X1 U18921 ( .B1(n15421), .B2(n15482), .A(n15420), .ZN(P1_U3016) );
  AOI21_X1 U18922 ( .B1(n17549), .B2(n21142), .A(n15422), .ZN(n15426) );
  NAND3_X1 U18923 ( .A1(n17591), .A2(n15424), .A3(n15427), .ZN(n15425) );
  OAI211_X1 U18924 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15429) );
  INV_X1 U18925 ( .A(n15429), .ZN(n15430) );
  OAI21_X1 U18926 ( .B1(n15431), .B2(n15482), .A(n15430), .ZN(P1_U3017) );
  INV_X1 U18927 ( .A(n15432), .ZN(n15439) );
  INV_X1 U18928 ( .A(n15442), .ZN(n15433) );
  NOR2_X1 U18929 ( .A1(n15434), .A2(n15433), .ZN(n15436) );
  OAI21_X1 U18930 ( .B1(n15437), .B2(n15436), .A(n15435), .ZN(n15438) );
  OAI211_X1 U18931 ( .C1(n15440), .C2(n17622), .A(n15439), .B(n15438), .ZN(
        n15441) );
  INV_X1 U18932 ( .A(n15441), .ZN(n15445) );
  OAI21_X1 U18933 ( .B1(n15450), .B2(n17600), .A(n21129), .ZN(n15447) );
  OAI22_X1 U18934 ( .A1(n21130), .A2(n15442), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17600), .ZN(n15443) );
  OAI21_X1 U18935 ( .B1(n15447), .B2(n15443), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15444) );
  OAI211_X1 U18936 ( .C1(n15446), .C2(n15482), .A(n15445), .B(n15444), .ZN(
        P1_U3018) );
  AOI21_X1 U18937 ( .B1(n15448), .B2(n15468), .A(n15447), .ZN(n15460) );
  OAI21_X1 U18938 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21134), .A(
        n15460), .ZN(n15456) );
  NAND3_X1 U18939 ( .A1(n17591), .A2(n15450), .A3(n15449), .ZN(n15453) );
  INV_X1 U18940 ( .A(n15451), .ZN(n15452) );
  OAI211_X1 U18941 ( .C1(n17622), .C2(n15454), .A(n15453), .B(n15452), .ZN(
        n15455) );
  AOI21_X1 U18942 ( .B1(n15456), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15455), .ZN(n15457) );
  OAI21_X1 U18943 ( .B1(n15458), .B2(n15482), .A(n15457), .ZN(P1_U3019) );
  NOR2_X1 U18944 ( .A1(n15460), .A2(n15459), .ZN(n15461) );
  AOI211_X1 U18945 ( .C1(n21142), .C2(n17564), .A(n15462), .B(n15461), .ZN(
        n15465) );
  NOR3_X1 U18946 ( .A1(n15491), .A2(n15478), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15463) );
  NAND3_X1 U18947 ( .A1(n17591), .A2(n15484), .A3(n15463), .ZN(n15464) );
  OAI211_X1 U18948 ( .C1(n15466), .C2(n15482), .A(n15465), .B(n15464), .ZN(
        P1_U3020) );
  NAND2_X1 U18949 ( .A1(n15468), .A2(n15467), .ZN(n15469) );
  NAND2_X1 U18950 ( .A1(n15469), .A2(n21129), .ZN(n17598) );
  INV_X1 U18951 ( .A(n15484), .ZN(n15470) );
  OR2_X1 U18952 ( .A1(n17598), .A2(n15470), .ZN(n15472) );
  NAND2_X1 U18953 ( .A1(n15472), .A2(n15471), .ZN(n15492) );
  AOI21_X1 U18954 ( .B1(n21142), .B2(n15474), .A(n15473), .ZN(n15477) );
  XNOR2_X1 U18955 ( .A(n15491), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15475) );
  NAND3_X1 U18956 ( .A1(n17591), .A2(n15484), .A3(n15475), .ZN(n15476) );
  OAI211_X1 U18957 ( .C1(n15492), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15479) );
  INV_X1 U18958 ( .A(n15479), .ZN(n15480) );
  OAI21_X1 U18959 ( .B1(n15481), .B2(n15482), .A(n15480), .ZN(P1_U3021) );
  NAND2_X1 U18960 ( .A1(n15483), .A2(n21145), .ZN(n15490) );
  AND2_X1 U18961 ( .A1(n17591), .A2(n15484), .ZN(n15488) );
  NOR2_X1 U18962 ( .A1(n15485), .A2(n17622), .ZN(n15486) );
  AOI211_X1 U18963 ( .C1(n15488), .C2(n15491), .A(n15487), .B(n15486), .ZN(
        n15489) );
  OAI211_X1 U18964 ( .C1(n15492), .C2(n15491), .A(n15490), .B(n15489), .ZN(
        P1_U3022) );
  OAI21_X1 U18965 ( .B1(n15560), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21285), 
        .ZN(n15493) );
  OAI22_X1 U18966 ( .A1(n15493), .A2(n15603), .B1(n21206), .B2(n15495), .ZN(
        n15494) );
  MUX2_X1 U18967 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15494), .S(
        n21153), .Z(P1_U3477) );
  XNOR2_X1 U18968 ( .A(n14285), .B(n15603), .ZN(n15496) );
  OAI22_X1 U18969 ( .A1(n15496), .A2(n21311), .B1(n14232), .B2(n15495), .ZN(
        n15497) );
  MUX2_X1 U18970 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15497), .S(
        n21153), .Z(P1_U3476) );
  INV_X1 U18971 ( .A(n14214), .ZN(n15498) );
  NAND2_X1 U18972 ( .A1(n15499), .A2(n15498), .ZN(n15505) );
  OAI22_X1 U18973 ( .A1(n15501), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15505), .B2(n15500), .ZN(n15502) );
  AOI21_X1 U18974 ( .B1(n15805), .B2(n15503), .A(n15502), .ZN(n17502) );
  INV_X1 U18975 ( .A(n15504), .ZN(n15522) );
  INV_X1 U18976 ( .A(n15505), .ZN(n15507) );
  INV_X1 U18977 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21149) );
  AOI22_X1 U18978 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21149), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n9931), .ZN(n15514) );
  AOI22_X1 U18979 ( .A1(n15508), .A2(n15507), .B1(n15514), .B2(n15506), .ZN(
        n15509) );
  OAI21_X1 U18980 ( .B1(n17502), .B2(n15522), .A(n15509), .ZN(n15510) );
  MUX2_X1 U18981 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15510), .S(
        n15516), .Z(P1_U3473) );
  INV_X1 U18982 ( .A(n15511), .ZN(n15512) );
  OAI222_X1 U18983 ( .A1(n15520), .A2(n15515), .B1(n15514), .B2(n15513), .C1(
        n15522), .C2(n15512), .ZN(n15517) );
  MUX2_X1 U18984 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15517), .S(
        n15516), .Z(P1_U3472) );
  INV_X1 U18985 ( .A(n15518), .ZN(n15523) );
  INV_X1 U18986 ( .A(n15519), .ZN(n15521) );
  OAI22_X1 U18987 ( .A1(n15523), .A2(n15522), .B1(n15521), .B2(n15520), .ZN(
        n15525) );
  MUX2_X1 U18988 ( .A(n15525), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15524), .Z(P1_U3469) );
  INV_X1 U18989 ( .A(n21199), .ZN(n15528) );
  OAI21_X1 U18990 ( .B1(n21155), .B2(n21164), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15529) );
  NAND2_X1 U18991 ( .A1(n15529), .A2(n21285), .ZN(n15541) );
  INV_X1 U18992 ( .A(n15541), .ZN(n15536) );
  INV_X1 U18993 ( .A(n14232), .ZN(n15530) );
  OR2_X1 U18994 ( .A1(n15531), .A2(n15530), .ZN(n21170) );
  NOR3_X1 U18995 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21177) );
  INV_X1 U18996 ( .A(n21177), .ZN(n21173) );
  NOR2_X1 U18997 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21173), .ZN(
        n21163) );
  INV_X1 U18998 ( .A(n15681), .ZN(n15532) );
  NAND2_X1 U18999 ( .A1(n15532), .A2(n15722), .ZN(n21201) );
  NAND2_X1 U19000 ( .A1(n21201), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15534) );
  NAND2_X1 U19001 ( .A1(n15538), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21202) );
  NAND2_X1 U19002 ( .A1(n15533), .A2(n21202), .ZN(n15729) );
  INV_X1 U19003 ( .A(n15729), .ZN(n15679) );
  OAI211_X1 U19004 ( .C1(n21163), .C2(n17636), .A(n15534), .B(n15679), .ZN(
        n15535) );
  INV_X1 U19005 ( .A(n21164), .ZN(n15554) );
  INV_X1 U19006 ( .A(n21163), .ZN(n15553) );
  OAI22_X1 U19007 ( .A1(n15554), .A2(n21321), .B1(n15553), .B2(n15683), .ZN(
        n15537) );
  AOI21_X1 U19008 ( .B1(n21155), .B2(n21318), .A(n15537), .ZN(n15543) );
  NOR2_X1 U19009 ( .A1(n15538), .A2(n11775), .ZN(n15723) );
  INV_X1 U19010 ( .A(n15723), .ZN(n15539) );
  NAND2_X1 U19011 ( .A1(n21165), .A2(n21314), .ZN(n15542) );
  OAI211_X1 U19012 ( .C1(n21158), .C2(n15544), .A(n15543), .B(n15542), .ZN(
        P1_U3033) );
  INV_X1 U19013 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15548) );
  OAI22_X1 U19014 ( .A1(n15554), .A2(n21333), .B1(n15553), .B2(n15691), .ZN(
        n15545) );
  AOI21_X1 U19015 ( .B1(n21155), .B2(n21330), .A(n15545), .ZN(n15547) );
  NAND2_X1 U19016 ( .A1(n21165), .A2(n21329), .ZN(n15546) );
  OAI211_X1 U19017 ( .C1(n21158), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        P1_U3035) );
  INV_X1 U19018 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15552) );
  OAI22_X1 U19019 ( .A1(n15554), .A2(n21339), .B1(n15553), .B2(n15695), .ZN(
        n15549) );
  AOI21_X1 U19020 ( .B1(n21155), .B2(n21336), .A(n15549), .ZN(n15551) );
  NAND2_X1 U19021 ( .A1(n21165), .A2(n21335), .ZN(n15550) );
  OAI211_X1 U19022 ( .C1(n21158), .C2(n15552), .A(n15551), .B(n15550), .ZN(
        P1_U3036) );
  INV_X1 U19023 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15558) );
  OAI22_X1 U19024 ( .A1(n15554), .A2(n21345), .B1(n15553), .B2(n15699), .ZN(
        n15555) );
  AOI21_X1 U19025 ( .B1(n21155), .B2(n21342), .A(n15555), .ZN(n15557) );
  NAND2_X1 U19026 ( .A1(n21165), .A2(n21341), .ZN(n15556) );
  OAI211_X1 U19027 ( .C1(n21158), .C2(n15558), .A(n15557), .B(n15556), .ZN(
        P1_U3037) );
  INV_X1 U19028 ( .A(n15802), .ZN(n15561) );
  NAND3_X1 U19029 ( .A1(n15564), .A2(n15635), .A3(n21285), .ZN(n15563) );
  NAND2_X1 U19030 ( .A1(n21285), .A2(n21204), .ZN(n15720) );
  NAND2_X1 U19031 ( .A1(n15563), .A2(n15720), .ZN(n15568) );
  NOR2_X1 U19032 ( .A1(n21170), .A2(n21206), .ZN(n15565) );
  OR2_X1 U19033 ( .A1(n15722), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15566) );
  INV_X1 U19034 ( .A(n15566), .ZN(n15640) );
  NAND3_X1 U19035 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17510), .A3(
        n21203), .ZN(n15608) );
  NOR2_X1 U19036 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15608), .ZN(
        n15592) );
  INV_X1 U19037 ( .A(n15565), .ZN(n15567) );
  AND2_X1 U19038 ( .A1(n15566), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15644) );
  AOI211_X1 U19039 ( .C1(n15568), .C2(n15567), .A(n15729), .B(n15644), .ZN(
        n15569) );
  OAI21_X1 U19040 ( .B1(n15592), .B2(n17636), .A(n15569), .ZN(n15591) );
  AOI22_X1 U19041 ( .A1(n21313), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n15591), .ZN(n15570) );
  OAI21_X1 U19042 ( .B1(n15635), .B2(n21214), .A(n15570), .ZN(n15571) );
  AOI21_X1 U19043 ( .B1(n21194), .B2(n21211), .A(n15571), .ZN(n15572) );
  OAI21_X1 U19044 ( .B1(n15812), .B2(n15596), .A(n15572), .ZN(P1_U3049) );
  AOI22_X1 U19045 ( .A1(n21322), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n15591), .ZN(n15573) );
  OAI21_X1 U19046 ( .B1(n15635), .B2(n21218), .A(n15573), .ZN(n15574) );
  AOI21_X1 U19047 ( .B1(n21194), .B2(n21215), .A(n15574), .ZN(n15575) );
  OAI21_X1 U19048 ( .B1(n15815), .B2(n15596), .A(n15575), .ZN(P1_U3050) );
  AOI22_X1 U19049 ( .A1(n21328), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n15591), .ZN(n15576) );
  OAI21_X1 U19050 ( .B1(n15635), .B2(n21222), .A(n15576), .ZN(n15577) );
  AOI21_X1 U19051 ( .B1(n21194), .B2(n21219), .A(n15577), .ZN(n15578) );
  OAI21_X1 U19052 ( .B1(n15818), .B2(n15596), .A(n15578), .ZN(P1_U3051) );
  AOI22_X1 U19053 ( .A1(n21334), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n15591), .ZN(n15579) );
  OAI21_X1 U19054 ( .B1(n15635), .B2(n21226), .A(n15579), .ZN(n15580) );
  AOI21_X1 U19055 ( .B1(n21194), .B2(n21223), .A(n15580), .ZN(n15581) );
  OAI21_X1 U19056 ( .B1(n15821), .B2(n15596), .A(n15581), .ZN(P1_U3052) );
  AOI22_X1 U19057 ( .A1(n21340), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n15591), .ZN(n15582) );
  OAI21_X1 U19058 ( .B1(n15635), .B2(n21230), .A(n15582), .ZN(n15583) );
  AOI21_X1 U19059 ( .B1(n21194), .B2(n21227), .A(n15583), .ZN(n15584) );
  OAI21_X1 U19060 ( .B1(n15824), .B2(n15596), .A(n15584), .ZN(P1_U3053) );
  AOI22_X1 U19061 ( .A1(n21346), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n15591), .ZN(n15585) );
  OAI21_X1 U19062 ( .B1(n15635), .B2(n21234), .A(n15585), .ZN(n15586) );
  AOI21_X1 U19063 ( .B1(n21194), .B2(n21231), .A(n15586), .ZN(n15587) );
  OAI21_X1 U19064 ( .B1(n15827), .B2(n15596), .A(n15587), .ZN(P1_U3054) );
  AOI22_X1 U19065 ( .A1(n21352), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n15591), .ZN(n15588) );
  OAI21_X1 U19066 ( .B1(n15635), .B2(n21238), .A(n15588), .ZN(n15589) );
  AOI21_X1 U19067 ( .B1(n21194), .B2(n21235), .A(n15589), .ZN(n15590) );
  OAI21_X1 U19068 ( .B1(n15830), .B2(n15596), .A(n15590), .ZN(P1_U3055) );
  AOI22_X1 U19069 ( .A1(n21359), .A2(n15592), .B1(
        P1_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n15591), .ZN(n15593) );
  OAI21_X1 U19070 ( .B1(n15635), .B2(n21246), .A(n15593), .ZN(n15594) );
  AOI21_X1 U19071 ( .B1(n21194), .B2(n21241), .A(n15594), .ZN(n15595) );
  OAI21_X1 U19072 ( .B1(n15837), .B2(n15596), .A(n15595), .ZN(P1_U3056) );
  INV_X1 U19073 ( .A(n21175), .ZN(n15598) );
  INV_X1 U19074 ( .A(n21170), .ZN(n15602) );
  NAND2_X1 U19075 ( .A1(n15599), .A2(n17510), .ZN(n15634) );
  INV_X1 U19076 ( .A(n15634), .ZN(n15600) );
  AOI21_X1 U19077 ( .B1(n15602), .B2(n15601), .A(n15600), .ZN(n15610) );
  INV_X1 U19078 ( .A(n15603), .ZN(n15604) );
  OR2_X1 U19079 ( .A1(n21175), .A2(n15604), .ZN(n15605) );
  AOI22_X1 U19080 ( .A1(n15610), .A2(n15607), .B1(n21311), .B2(n15608), .ZN(
        n15606) );
  NAND2_X1 U19081 ( .A1(n21315), .A2(n15606), .ZN(n15633) );
  INV_X1 U19082 ( .A(n15607), .ZN(n15609) );
  AOI22_X1 U19083 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n15633), .B1(
        n21314), .B2(n15632), .ZN(n15613) );
  OAI22_X1 U19084 ( .A1(n15635), .A2(n21321), .B1(n15634), .B2(n15683), .ZN(
        n15611) );
  INV_X1 U19085 ( .A(n15611), .ZN(n15612) );
  OAI211_X1 U19086 ( .C1(n21214), .C2(n21210), .A(n15613), .B(n15612), .ZN(
        P1_U3057) );
  AOI22_X1 U19087 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n15633), .B1(
        n21323), .B2(n15632), .ZN(n15616) );
  OAI22_X1 U19088 ( .A1(n15635), .A2(n21327), .B1(n15634), .B2(n15687), .ZN(
        n15614) );
  INV_X1 U19089 ( .A(n15614), .ZN(n15615) );
  OAI211_X1 U19090 ( .C1(n21218), .C2(n21210), .A(n15616), .B(n15615), .ZN(
        P1_U3058) );
  AOI22_X1 U19091 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n15633), .B1(
        n21329), .B2(n15632), .ZN(n15619) );
  OAI22_X1 U19092 ( .A1(n15635), .A2(n21333), .B1(n15634), .B2(n15691), .ZN(
        n15617) );
  INV_X1 U19093 ( .A(n15617), .ZN(n15618) );
  OAI211_X1 U19094 ( .C1(n21222), .C2(n21210), .A(n15619), .B(n15618), .ZN(
        P1_U3059) );
  AOI22_X1 U19095 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n15633), .B1(
        n21335), .B2(n15632), .ZN(n15622) );
  OAI22_X1 U19096 ( .A1(n15635), .A2(n21339), .B1(n15634), .B2(n15695), .ZN(
        n15620) );
  INV_X1 U19097 ( .A(n15620), .ZN(n15621) );
  OAI211_X1 U19098 ( .C1(n21226), .C2(n21210), .A(n15622), .B(n15621), .ZN(
        P1_U3060) );
  AOI22_X1 U19099 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n15633), .B1(
        n21341), .B2(n15632), .ZN(n15625) );
  OAI22_X1 U19100 ( .A1(n15635), .A2(n21345), .B1(n15634), .B2(n15699), .ZN(
        n15623) );
  INV_X1 U19101 ( .A(n15623), .ZN(n15624) );
  OAI211_X1 U19102 ( .C1(n21230), .C2(n21210), .A(n15625), .B(n15624), .ZN(
        P1_U3061) );
  AOI22_X1 U19103 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n15633), .B1(
        n21347), .B2(n15632), .ZN(n15628) );
  OAI22_X1 U19104 ( .A1(n15635), .A2(n21351), .B1(n15634), .B2(n15703), .ZN(
        n15626) );
  INV_X1 U19105 ( .A(n15626), .ZN(n15627) );
  OAI211_X1 U19106 ( .C1(n21234), .C2(n21210), .A(n15628), .B(n15627), .ZN(
        P1_U3062) );
  AOI22_X1 U19107 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n15633), .B1(
        n21353), .B2(n15632), .ZN(n15631) );
  OAI22_X1 U19108 ( .A1(n15635), .A2(n21357), .B1(n15634), .B2(n15707), .ZN(
        n15629) );
  INV_X1 U19109 ( .A(n15629), .ZN(n15630) );
  OAI211_X1 U19110 ( .C1(n21238), .C2(n21210), .A(n15631), .B(n15630), .ZN(
        P1_U3063) );
  AOI22_X1 U19111 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n15633), .B1(
        n21361), .B2(n15632), .ZN(n15638) );
  OAI22_X1 U19112 ( .A1(n15635), .A2(n21368), .B1(n15634), .B2(n15712), .ZN(
        n15636) );
  INV_X1 U19113 ( .A(n15636), .ZN(n15637) );
  OAI211_X1 U19114 ( .C1(n21246), .C2(n21210), .A(n15638), .B(n15637), .ZN(
        P1_U3064) );
  NAND2_X1 U19115 ( .A1(n15672), .A2(n21285), .ZN(n15639) );
  OAI21_X1 U19116 ( .B1(n15639), .B2(n21271), .A(n15720), .ZN(n15646) );
  AND2_X1 U19117 ( .A1(n21248), .A2(n15805), .ZN(n15643) );
  INV_X1 U19118 ( .A(n21202), .ZN(n15798) );
  NOR2_X1 U19119 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15641), .ZN(
        n15670) );
  NOR2_X1 U19120 ( .A1(n15642), .A2(n15723), .ZN(n21208) );
  INV_X1 U19121 ( .A(n15643), .ZN(n15645) );
  AOI21_X1 U19122 ( .B1(n15646), .B2(n15645), .A(n15644), .ZN(n15647) );
  OAI211_X1 U19123 ( .C1(n15670), .C2(n17636), .A(n21208), .B(n15647), .ZN(
        n15669) );
  AOI22_X1 U19124 ( .A1(n21313), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n15669), .ZN(n15648) );
  OAI21_X1 U19125 ( .B1(n15672), .B2(n21214), .A(n15648), .ZN(n15649) );
  AOI21_X1 U19126 ( .B1(n21271), .B2(n21211), .A(n15649), .ZN(n15650) );
  OAI21_X1 U19127 ( .B1(n15812), .B2(n15675), .A(n15650), .ZN(P1_U3081) );
  AOI22_X1 U19128 ( .A1(n21322), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n15669), .ZN(n15651) );
  OAI21_X1 U19129 ( .B1(n15672), .B2(n21218), .A(n15651), .ZN(n15652) );
  AOI21_X1 U19130 ( .B1(n21271), .B2(n21215), .A(n15652), .ZN(n15653) );
  OAI21_X1 U19131 ( .B1(n15815), .B2(n15675), .A(n15653), .ZN(P1_U3082) );
  AOI22_X1 U19132 ( .A1(n21328), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n15669), .ZN(n15654) );
  OAI21_X1 U19133 ( .B1(n15672), .B2(n21222), .A(n15654), .ZN(n15655) );
  AOI21_X1 U19134 ( .B1(n21271), .B2(n21219), .A(n15655), .ZN(n15656) );
  OAI21_X1 U19135 ( .B1(n15818), .B2(n15675), .A(n15656), .ZN(P1_U3083) );
  AOI22_X1 U19136 ( .A1(n21334), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n15669), .ZN(n15657) );
  OAI21_X1 U19137 ( .B1(n15672), .B2(n21226), .A(n15657), .ZN(n15658) );
  AOI21_X1 U19138 ( .B1(n21271), .B2(n21223), .A(n15658), .ZN(n15659) );
  OAI21_X1 U19139 ( .B1(n15821), .B2(n15675), .A(n15659), .ZN(P1_U3084) );
  AOI22_X1 U19140 ( .A1(n21340), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n15669), .ZN(n15660) );
  OAI21_X1 U19141 ( .B1(n15672), .B2(n21230), .A(n15660), .ZN(n15661) );
  AOI21_X1 U19142 ( .B1(n21271), .B2(n21227), .A(n15661), .ZN(n15662) );
  OAI21_X1 U19143 ( .B1(n15824), .B2(n15675), .A(n15662), .ZN(P1_U3085) );
  AOI22_X1 U19144 ( .A1(n21346), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n15669), .ZN(n15663) );
  OAI21_X1 U19145 ( .B1(n15672), .B2(n21234), .A(n15663), .ZN(n15664) );
  AOI21_X1 U19146 ( .B1(n21271), .B2(n21231), .A(n15664), .ZN(n15665) );
  OAI21_X1 U19147 ( .B1(n15827), .B2(n15675), .A(n15665), .ZN(P1_U3086) );
  AOI22_X1 U19148 ( .A1(n21352), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n15669), .ZN(n15666) );
  OAI21_X1 U19149 ( .B1(n15672), .B2(n21238), .A(n15666), .ZN(n15667) );
  AOI21_X1 U19150 ( .B1(n21271), .B2(n21235), .A(n15667), .ZN(n15668) );
  OAI21_X1 U19151 ( .B1(n15830), .B2(n15675), .A(n15668), .ZN(P1_U3087) );
  AOI22_X1 U19152 ( .A1(n21359), .A2(n15670), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n15669), .ZN(n15671) );
  OAI21_X1 U19153 ( .B1(n15672), .B2(n21246), .A(n15671), .ZN(n15673) );
  AOI21_X1 U19154 ( .B1(n21271), .B2(n21241), .A(n15673), .ZN(n15674) );
  OAI21_X1 U19155 ( .B1(n15837), .B2(n15675), .A(n15674), .ZN(P1_U3088) );
  NOR3_X1 U19156 ( .A1(n17510), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21284) );
  INV_X1 U19157 ( .A(n21284), .ZN(n21279) );
  NOR2_X1 U19158 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21279), .ZN(
        n15680) );
  INV_X1 U19159 ( .A(n15716), .ZN(n15676) );
  AOI21_X1 U19160 ( .B1(n15676), .B2(n21306), .A(n21204), .ZN(n15677) );
  INV_X1 U19161 ( .A(n15680), .ZN(n15713) );
  OAI21_X1 U19162 ( .B1(n21276), .B2(n15805), .A(n15713), .ZN(n15682) );
  NAND2_X1 U19163 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n15686) );
  AND2_X1 U19164 ( .A1(n15681), .A2(n15722), .ZN(n15765) );
  AOI22_X1 U19165 ( .A1(n15682), .A2(n21285), .B1(n15765), .B2(n15723), .ZN(
        n15714) );
  OAI22_X1 U19166 ( .A1(n15812), .A2(n15714), .B1(n15683), .B2(n15713), .ZN(
        n15684) );
  AOI21_X1 U19167 ( .B1(n15716), .B2(n21211), .A(n15684), .ZN(n15685) );
  OAI211_X1 U19168 ( .C1(n21214), .C2(n21306), .A(n15686), .B(n15685), .ZN(
        P1_U3097) );
  NAND2_X1 U19169 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15690) );
  OAI22_X1 U19170 ( .A1(n15815), .A2(n15714), .B1(n15713), .B2(n15687), .ZN(
        n15688) );
  AOI21_X1 U19171 ( .B1(n15716), .B2(n21215), .A(n15688), .ZN(n15689) );
  OAI211_X1 U19172 ( .C1(n21218), .C2(n21306), .A(n15690), .B(n15689), .ZN(
        P1_U3098) );
  NAND2_X1 U19173 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n15694) );
  OAI22_X1 U19174 ( .A1(n15818), .A2(n15714), .B1(n15713), .B2(n15691), .ZN(
        n15692) );
  AOI21_X1 U19175 ( .B1(n15716), .B2(n21219), .A(n15692), .ZN(n15693) );
  OAI211_X1 U19176 ( .C1(n21222), .C2(n21306), .A(n15694), .B(n15693), .ZN(
        P1_U3099) );
  NAND2_X1 U19177 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15698) );
  OAI22_X1 U19178 ( .A1(n15821), .A2(n15714), .B1(n15713), .B2(n15695), .ZN(
        n15696) );
  AOI21_X1 U19179 ( .B1(n15716), .B2(n21223), .A(n15696), .ZN(n15697) );
  OAI211_X1 U19180 ( .C1(n21226), .C2(n21306), .A(n15698), .B(n15697), .ZN(
        P1_U3100) );
  NAND2_X1 U19181 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15702) );
  OAI22_X1 U19182 ( .A1(n15824), .A2(n15714), .B1(n15713), .B2(n15699), .ZN(
        n15700) );
  AOI21_X1 U19183 ( .B1(n15716), .B2(n21227), .A(n15700), .ZN(n15701) );
  OAI211_X1 U19184 ( .C1(n21230), .C2(n21306), .A(n15702), .B(n15701), .ZN(
        P1_U3101) );
  NAND2_X1 U19185 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15706) );
  OAI22_X1 U19186 ( .A1(n15827), .A2(n15714), .B1(n15713), .B2(n15703), .ZN(
        n15704) );
  AOI21_X1 U19187 ( .B1(n15716), .B2(n21231), .A(n15704), .ZN(n15705) );
  OAI211_X1 U19188 ( .C1(n21234), .C2(n21306), .A(n15706), .B(n15705), .ZN(
        P1_U3102) );
  NAND2_X1 U19189 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15710) );
  OAI22_X1 U19190 ( .A1(n15830), .A2(n15714), .B1(n15713), .B2(n15707), .ZN(
        n15708) );
  AOI21_X1 U19191 ( .B1(n15716), .B2(n21235), .A(n15708), .ZN(n15709) );
  OAI211_X1 U19192 ( .C1(n21238), .C2(n21306), .A(n15710), .B(n15709), .ZN(
        P1_U3103) );
  NAND2_X1 U19193 ( .A1(n15711), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n15718) );
  OAI22_X1 U19194 ( .A1(n15837), .A2(n15714), .B1(n15713), .B2(n15712), .ZN(
        n15715) );
  AOI21_X1 U19195 ( .B1(n15716), .B2(n21241), .A(n15715), .ZN(n15717) );
  OAI211_X1 U19196 ( .C1(n21246), .C2(n21306), .A(n15718), .B(n15717), .ZN(
        P1_U3104) );
  NAND2_X1 U19197 ( .A1(n15757), .A2(n21285), .ZN(n15721) );
  OAI21_X1 U19198 ( .B1(n15721), .B2(n21302), .A(n15720), .ZN(n15731) );
  NOR2_X1 U19199 ( .A1(n21276), .A2(n21206), .ZN(n15726) );
  OR2_X1 U19200 ( .A1(n15722), .A2(n17510), .ZN(n15727) );
  INV_X1 U19201 ( .A(n15727), .ZN(n15799) );
  INV_X1 U19202 ( .A(n15724), .ZN(n15725) );
  NOR2_X1 U19203 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15725), .ZN(
        n15755) );
  INV_X1 U19204 ( .A(n15726), .ZN(n15730) );
  NAND2_X1 U19205 ( .A1(n15727), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15808) );
  INV_X1 U19206 ( .A(n15808), .ZN(n15728) );
  AOI211_X1 U19207 ( .C1(n15731), .C2(n15730), .A(n15729), .B(n15728), .ZN(
        n15732) );
  OAI21_X1 U19208 ( .B1(n15755), .B2(n17636), .A(n15732), .ZN(n15754) );
  AOI22_X1 U19209 ( .A1(n21313), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__0__SCAN_IN), .B2(n15754), .ZN(n15733) );
  OAI21_X1 U19210 ( .B1(n15757), .B2(n21214), .A(n15733), .ZN(n15734) );
  AOI21_X1 U19211 ( .B1(n21302), .B2(n21211), .A(n15734), .ZN(n15735) );
  OAI21_X1 U19212 ( .B1(n15812), .B2(n15760), .A(n15735), .ZN(P1_U3113) );
  AOI22_X1 U19213 ( .A1(n21322), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n15754), .ZN(n15736) );
  OAI21_X1 U19214 ( .B1(n15757), .B2(n21218), .A(n15736), .ZN(n15737) );
  AOI21_X1 U19215 ( .B1(n21302), .B2(n21215), .A(n15737), .ZN(n15738) );
  OAI21_X1 U19216 ( .B1(n15815), .B2(n15760), .A(n15738), .ZN(P1_U3114) );
  AOI22_X1 U19217 ( .A1(n21328), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n15754), .ZN(n15739) );
  OAI21_X1 U19218 ( .B1(n15757), .B2(n21222), .A(n15739), .ZN(n15740) );
  AOI21_X1 U19219 ( .B1(n21302), .B2(n21219), .A(n15740), .ZN(n15741) );
  OAI21_X1 U19220 ( .B1(n15818), .B2(n15760), .A(n15741), .ZN(P1_U3115) );
  AOI22_X1 U19221 ( .A1(n21334), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n15754), .ZN(n15742) );
  OAI21_X1 U19222 ( .B1(n15757), .B2(n21226), .A(n15742), .ZN(n15743) );
  AOI21_X1 U19223 ( .B1(n21302), .B2(n21223), .A(n15743), .ZN(n15744) );
  OAI21_X1 U19224 ( .B1(n15821), .B2(n15760), .A(n15744), .ZN(P1_U3116) );
  AOI22_X1 U19225 ( .A1(n21340), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n15754), .ZN(n15745) );
  OAI21_X1 U19226 ( .B1(n15757), .B2(n21230), .A(n15745), .ZN(n15746) );
  AOI21_X1 U19227 ( .B1(n21302), .B2(n21227), .A(n15746), .ZN(n15747) );
  OAI21_X1 U19228 ( .B1(n15824), .B2(n15760), .A(n15747), .ZN(P1_U3117) );
  AOI22_X1 U19229 ( .A1(n21346), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(n15754), .ZN(n15748) );
  OAI21_X1 U19230 ( .B1(n15757), .B2(n21234), .A(n15748), .ZN(n15749) );
  AOI21_X1 U19231 ( .B1(n21302), .B2(n21231), .A(n15749), .ZN(n15750) );
  OAI21_X1 U19232 ( .B1(n15827), .B2(n15760), .A(n15750), .ZN(P1_U3118) );
  AOI22_X1 U19233 ( .A1(n21352), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n15754), .ZN(n15751) );
  OAI21_X1 U19234 ( .B1(n15757), .B2(n21238), .A(n15751), .ZN(n15752) );
  AOI21_X1 U19235 ( .B1(n21302), .B2(n21235), .A(n15752), .ZN(n15753) );
  OAI21_X1 U19236 ( .B1(n15830), .B2(n15760), .A(n15753), .ZN(P1_U3119) );
  AOI22_X1 U19237 ( .A1(n21359), .A2(n15755), .B1(
        P1_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n15754), .ZN(n15756) );
  OAI21_X1 U19238 ( .B1(n15757), .B2(n21246), .A(n15756), .ZN(n15758) );
  AOI21_X1 U19239 ( .B1(n21302), .B2(n21241), .A(n15758), .ZN(n15759) );
  OAI21_X1 U19240 ( .B1(n15837), .B2(n15760), .A(n15759), .ZN(P1_U3120) );
  INV_X1 U19241 ( .A(n21367), .ZN(n15761) );
  OAI21_X1 U19242 ( .B1(n15795), .B2(n15761), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15762) );
  NOR2_X1 U19243 ( .A1(n15763), .A2(n15805), .ZN(n15764) );
  NOR3_X1 U19244 ( .A1(n21203), .A2(n17510), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21317) );
  INV_X1 U19245 ( .A(n21317), .ZN(n21310) );
  NOR2_X1 U19246 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21310), .ZN(
        n15792) );
  INV_X1 U19247 ( .A(n15764), .ZN(n15767) );
  NOR2_X1 U19248 ( .A1(n15765), .A2(n11775), .ZN(n15766) );
  AOI21_X1 U19249 ( .B1(n15768), .B2(n15767), .A(n15766), .ZN(n15769) );
  OAI211_X1 U19250 ( .C1(n15792), .C2(n17636), .A(n21208), .B(n15769), .ZN(
        n15791) );
  AOI22_X1 U19251 ( .A1(n21313), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n15791), .ZN(n15770) );
  OAI21_X1 U19252 ( .B1(n21367), .B2(n21214), .A(n15770), .ZN(n15771) );
  AOI21_X1 U19253 ( .B1(n15795), .B2(n21211), .A(n15771), .ZN(n15772) );
  OAI21_X1 U19254 ( .B1(n15812), .B2(n15797), .A(n15772), .ZN(P1_U3129) );
  AOI22_X1 U19255 ( .A1(n21322), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15791), .ZN(n15773) );
  OAI21_X1 U19256 ( .B1(n21367), .B2(n21218), .A(n15773), .ZN(n15774) );
  AOI21_X1 U19257 ( .B1(n15795), .B2(n21215), .A(n15774), .ZN(n15775) );
  OAI21_X1 U19258 ( .B1(n15815), .B2(n15797), .A(n15775), .ZN(P1_U3130) );
  AOI22_X1 U19259 ( .A1(n21328), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n15791), .ZN(n15776) );
  OAI21_X1 U19260 ( .B1(n21367), .B2(n21222), .A(n15776), .ZN(n15777) );
  AOI21_X1 U19261 ( .B1(n15795), .B2(n21219), .A(n15777), .ZN(n15778) );
  OAI21_X1 U19262 ( .B1(n15818), .B2(n15797), .A(n15778), .ZN(P1_U3131) );
  AOI22_X1 U19263 ( .A1(n21334), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n15791), .ZN(n15779) );
  OAI21_X1 U19264 ( .B1(n21367), .B2(n21226), .A(n15779), .ZN(n15780) );
  AOI21_X1 U19265 ( .B1(n15795), .B2(n21223), .A(n15780), .ZN(n15781) );
  OAI21_X1 U19266 ( .B1(n15821), .B2(n15797), .A(n15781), .ZN(P1_U3132) );
  AOI22_X1 U19267 ( .A1(n21340), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n15791), .ZN(n15782) );
  OAI21_X1 U19268 ( .B1(n21367), .B2(n21230), .A(n15782), .ZN(n15783) );
  AOI21_X1 U19269 ( .B1(n15795), .B2(n21227), .A(n15783), .ZN(n15784) );
  OAI21_X1 U19270 ( .B1(n15824), .B2(n15797), .A(n15784), .ZN(P1_U3133) );
  AOI22_X1 U19271 ( .A1(n21346), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n15791), .ZN(n15785) );
  OAI21_X1 U19272 ( .B1(n21367), .B2(n21234), .A(n15785), .ZN(n15786) );
  AOI21_X1 U19273 ( .B1(n15795), .B2(n21231), .A(n15786), .ZN(n15787) );
  OAI21_X1 U19274 ( .B1(n15827), .B2(n15797), .A(n15787), .ZN(P1_U3134) );
  AOI22_X1 U19275 ( .A1(n21352), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n15791), .ZN(n15788) );
  OAI21_X1 U19276 ( .B1(n21367), .B2(n21238), .A(n15788), .ZN(n15789) );
  AOI21_X1 U19277 ( .B1(n15795), .B2(n21235), .A(n15789), .ZN(n15790) );
  OAI21_X1 U19278 ( .B1(n15830), .B2(n15797), .A(n15790), .ZN(P1_U3135) );
  AOI22_X1 U19279 ( .A1(n21359), .A2(n15792), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n15791), .ZN(n15793) );
  OAI21_X1 U19280 ( .B1(n21367), .B2(n21246), .A(n15793), .ZN(n15794) );
  AOI21_X1 U19281 ( .B1(n15795), .B2(n21241), .A(n15794), .ZN(n15796) );
  OAI21_X1 U19282 ( .B1(n15837), .B2(n15797), .A(n15796), .ZN(P1_U3136) );
  INV_X1 U19283 ( .A(n21308), .ZN(n15800) );
  AOI22_X1 U19284 ( .A1(n15800), .A2(n15805), .B1(n15799), .B2(n15798), .ZN(
        n15836) );
  NOR2_X1 U19285 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15801), .ZN(
        n15832) );
  OAI21_X1 U19286 ( .B1(n21363), .B2(n15833), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15807) );
  NAND2_X1 U19287 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  AOI21_X1 U19288 ( .B1(n15807), .B2(n15806), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15809) );
  AOI22_X1 U19289 ( .A1(n21313), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n15831), .ZN(n15811) );
  AOI22_X1 U19290 ( .A1(n21363), .A2(n21211), .B1(n15833), .B2(n21318), .ZN(
        n15810) );
  OAI211_X1 U19291 ( .C1(n15812), .C2(n15836), .A(n15811), .B(n15810), .ZN(
        P1_U3145) );
  AOI22_X1 U19292 ( .A1(n21322), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n15831), .ZN(n15814) );
  AOI22_X1 U19293 ( .A1(n21363), .A2(n21215), .B1(n15833), .B2(n21324), .ZN(
        n15813) );
  OAI211_X1 U19294 ( .C1(n15815), .C2(n15836), .A(n15814), .B(n15813), .ZN(
        P1_U3146) );
  AOI22_X1 U19295 ( .A1(n21328), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n15831), .ZN(n15817) );
  AOI22_X1 U19296 ( .A1(n21363), .A2(n21219), .B1(n15833), .B2(n21330), .ZN(
        n15816) );
  OAI211_X1 U19297 ( .C1(n15818), .C2(n15836), .A(n15817), .B(n15816), .ZN(
        P1_U3147) );
  AOI22_X1 U19298 ( .A1(n21334), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n15831), .ZN(n15820) );
  AOI22_X1 U19299 ( .A1(n21363), .A2(n21223), .B1(n15833), .B2(n21336), .ZN(
        n15819) );
  OAI211_X1 U19300 ( .C1(n15821), .C2(n15836), .A(n15820), .B(n15819), .ZN(
        P1_U3148) );
  AOI22_X1 U19301 ( .A1(n21340), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n15831), .ZN(n15823) );
  AOI22_X1 U19302 ( .A1(n21363), .A2(n21227), .B1(n15833), .B2(n21342), .ZN(
        n15822) );
  OAI211_X1 U19303 ( .C1(n15824), .C2(n15836), .A(n15823), .B(n15822), .ZN(
        P1_U3149) );
  AOI22_X1 U19304 ( .A1(n21346), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__5__SCAN_IN), .B2(n15831), .ZN(n15826) );
  AOI22_X1 U19305 ( .A1(n21363), .A2(n21231), .B1(n15833), .B2(n21348), .ZN(
        n15825) );
  OAI211_X1 U19306 ( .C1(n15827), .C2(n15836), .A(n15826), .B(n15825), .ZN(
        P1_U3150) );
  AOI22_X1 U19307 ( .A1(n21352), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n15831), .ZN(n15829) );
  AOI22_X1 U19308 ( .A1(n21363), .A2(n21235), .B1(n15833), .B2(n21354), .ZN(
        n15828) );
  OAI211_X1 U19309 ( .C1(n15830), .C2(n15836), .A(n15829), .B(n15828), .ZN(
        P1_U3151) );
  AOI22_X1 U19310 ( .A1(n21359), .A2(n15832), .B1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n15831), .ZN(n15835) );
  AOI22_X1 U19311 ( .A1(n21363), .A2(n21241), .B1(n15833), .B2(n21362), .ZN(
        n15834) );
  OAI211_X1 U19312 ( .C1(n15837), .C2(n15836), .A(n15835), .B(n15834), .ZN(
        P1_U3152) );
  NAND3_X1 U19313 ( .A1(n13794), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n15838), 
        .ZN(n15839) );
  OAI21_X1 U19314 ( .B1(n16262), .B2(n20858), .A(n15839), .ZN(n15843) );
  INV_X2 U19315 ( .A(n16274), .ZN(n20083) );
  NOR3_X1 U19316 ( .A1(n15841), .A2(n15840), .A3(n16297), .ZN(n15842) );
  AOI211_X1 U19317 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n16275), .A(
        n15843), .B(n15842), .ZN(n15844) );
  OAI21_X1 U19318 ( .B1(n15845), .B2(n20073), .A(n15844), .ZN(n15846) );
  AOI21_X1 U19319 ( .B1(n16530), .B2(n16301), .A(n15846), .ZN(n15847) );
  OAI21_X1 U19320 ( .B1(n16424), .B2(n20077), .A(n15847), .ZN(P2_U2824) );
  AOI21_X1 U19321 ( .B1(n15849), .B2(n9655), .A(n15848), .ZN(n16783) );
  INV_X1 U19322 ( .A(n16783), .ZN(n16432) );
  OR2_X1 U19323 ( .A1(n13202), .A2(n15850), .ZN(n15851) );
  NAND2_X1 U19324 ( .A1(n15852), .A2(n15851), .ZN(n16781) );
  AOI21_X1 U19325 ( .B1(n15855), .B2(n20083), .A(n16282), .ZN(n15859) );
  INV_X1 U19326 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15853) );
  OAI22_X1 U19327 ( .A1(n20072), .A2(n15853), .B1(n20853), .B2(n16262), .ZN(
        n15857) );
  INV_X1 U19328 ( .A(n16538), .ZN(n15854) );
  NOR3_X1 U19329 ( .A1(n15855), .A2(n15854), .A3(n16297), .ZN(n15856) );
  AOI211_X1 U19330 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15857), .B(n15856), .ZN(n15858) );
  OAI21_X1 U19331 ( .B1(n16432), .B2(n20077), .A(n15864), .ZN(P2_U2826) );
  NAND2_X1 U19332 ( .A1(n15865), .A2(n15866), .ZN(n15867) );
  INV_X1 U19333 ( .A(n16796), .ZN(n15881) );
  OAI22_X1 U19334 ( .A1(n20072), .A2(n15869), .B1(n15868), .B2(n16262), .ZN(
        n15871) );
  INV_X1 U19335 ( .A(n15872), .ZN(n15889) );
  NOR3_X1 U19336 ( .A1(n15889), .A2(n15873), .A3(n16297), .ZN(n15870) );
  AOI211_X1 U19337 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15871), .B(n15870), .ZN(n15876) );
  NOR2_X1 U19338 ( .A1(n15872), .A2(n16274), .ZN(n15874) );
  OAI21_X1 U19339 ( .B1(n15874), .B2(n16282), .A(n15873), .ZN(n15875) );
  OAI211_X1 U19340 ( .C1(n15877), .C2(n20073), .A(n15876), .B(n15875), .ZN(
        n15878) );
  AOI21_X1 U19341 ( .B1(n15879), .B2(n15862), .A(n15878), .ZN(n15880) );
  OAI21_X1 U19342 ( .B1(n15881), .B2(n20077), .A(n15880), .ZN(P2_U2827) );
  OR2_X1 U19343 ( .A1(n15882), .A2(n15883), .ZN(n15884) );
  NAND2_X1 U19344 ( .A1(n15865), .A2(n15884), .ZN(n16810) );
  XNOR2_X1 U19345 ( .A(n15886), .B(n15885), .ZN(n16318) );
  INV_X1 U19346 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15887) );
  OAI22_X1 U19347 ( .A1(n20072), .A2(n15887), .B1(n20851), .B2(n16262), .ZN(
        n15892) );
  OAI21_X1 U19348 ( .B1(n15888), .B2(n16549), .A(n20083), .ZN(n15890) );
  AOI21_X1 U19349 ( .B1(n16288), .B2(n15890), .A(n15889), .ZN(n15891) );
  AOI211_X1 U19350 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15892), .B(n15891), .ZN(n15893) );
  OAI21_X1 U19351 ( .B1(n15894), .B2(n20073), .A(n15893), .ZN(n15895) );
  AOI21_X1 U19352 ( .B1(n16808), .B2(n16301), .A(n15895), .ZN(n15896) );
  OAI21_X1 U19353 ( .B1(n16810), .B2(n20077), .A(n15896), .ZN(P2_U2828) );
  AOI21_X1 U19354 ( .B1(n15898), .B2(n15913), .A(n15882), .ZN(n16822) );
  INV_X1 U19355 ( .A(n16822), .ZN(n15911) );
  INV_X1 U19356 ( .A(n15899), .ZN(n15900) );
  AOI211_X1 U19357 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n15900), .A(n20073), .B(
        n11543), .ZN(n15909) );
  INV_X1 U19358 ( .A(n16262), .ZN(n20076) );
  AOI22_X1 U19359 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16275), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n20076), .ZN(n15907) );
  NOR2_X1 U19360 ( .A1(n20080), .A2(n10223), .ZN(n15903) );
  OAI21_X1 U19361 ( .B1(n15904), .B2(n15903), .A(n20083), .ZN(n15902) );
  AOI21_X1 U19362 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(n15905) );
  INV_X1 U19363 ( .A(n15905), .ZN(n15906) );
  OAI211_X1 U19364 ( .C1(n20072), .C2(n16330), .A(n15907), .B(n15906), .ZN(
        n15908) );
  AOI211_X1 U19365 ( .C1(n16329), .C2(n15862), .A(n15909), .B(n15908), .ZN(
        n15910) );
  OAI21_X1 U19366 ( .B1(n15911), .B2(n20077), .A(n15910), .ZN(P2_U2829) );
  AOI21_X1 U19367 ( .B1(n15914), .B2(n15912), .A(n15897), .ZN(n16835) );
  INV_X1 U19368 ( .A(n16835), .ZN(n15929) );
  OAI21_X1 U19369 ( .B1(n15915), .B2(n15916), .A(n11159), .ZN(n16832) );
  INV_X1 U19370 ( .A(n16832), .ZN(n15927) );
  INV_X1 U19371 ( .A(n15917), .ZN(n15925) );
  INV_X1 U19372 ( .A(n15918), .ZN(n15919) );
  NOR2_X1 U19373 ( .A1(n20080), .A2(n15919), .ZN(n15921) );
  OAI21_X1 U19374 ( .B1(n16560), .B2(n15921), .A(n20083), .ZN(n15920) );
  AOI21_X1 U19375 ( .B1(n16560), .B2(n15921), .A(n15920), .ZN(n15923) );
  INV_X1 U19376 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20846) );
  OAI22_X1 U19377 ( .A1(n16557), .A2(n20092), .B1(n20846), .B2(n16262), .ZN(
        n15922) );
  AOI211_X1 U19378 ( .C1(n16292), .C2(P2_EBX_REG_25__SCAN_IN), .A(n15923), .B(
        n15922), .ZN(n15924) );
  OAI21_X1 U19379 ( .B1(n15925), .B2(n20073), .A(n15924), .ZN(n15926) );
  AOI21_X1 U19380 ( .B1(n15927), .B2(n16301), .A(n15926), .ZN(n15928) );
  OAI21_X1 U19381 ( .B1(n15929), .B2(n20077), .A(n15928), .ZN(P2_U2830) );
  OAI21_X1 U19382 ( .B1(n15930), .B2(n15931), .A(n15912), .ZN(n16848) );
  NOR2_X1 U19383 ( .A1(n15932), .A2(n15933), .ZN(n15934) );
  OR2_X1 U19384 ( .A1(n15915), .A2(n15934), .ZN(n16570) );
  INV_X1 U19385 ( .A(n16570), .ZN(n16846) );
  AOI21_X1 U19386 ( .B1(n20083), .B2(n15936), .A(n16282), .ZN(n15942) );
  XOR2_X1 U19387 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n9682), .Z(n15935) );
  NAND2_X1 U19388 ( .A1(n15935), .A2(n16290), .ZN(n15940) );
  INV_X1 U19389 ( .A(n15941), .ZN(n16568) );
  NOR3_X1 U19390 ( .A1(n16297), .A2(n16568), .A3(n15936), .ZN(n15938) );
  OAI22_X1 U19391 ( .A1(n20072), .A2(n11088), .B1(n20844), .B2(n16262), .ZN(
        n15937) );
  AOI211_X1 U19392 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15938), .B(n15937), .ZN(n15939) );
  OAI211_X1 U19393 ( .C1(n15942), .C2(n15941), .A(n15940), .B(n15939), .ZN(
        n15943) );
  AOI21_X1 U19394 ( .B1(n16846), .B2(n16301), .A(n15943), .ZN(n15944) );
  OAI21_X1 U19395 ( .B1(n16848), .B2(n20077), .A(n15944), .ZN(P2_U2831) );
  NOR2_X1 U19396 ( .A1(n15945), .A2(n15946), .ZN(n15947) );
  OR2_X1 U19397 ( .A1(n15930), .A2(n15947), .ZN(n16853) );
  INV_X1 U19398 ( .A(n15948), .ZN(n15969) );
  AND2_X1 U19399 ( .A1(n15969), .A2(n15949), .ZN(n15950) );
  OR2_X1 U19400 ( .A1(n15950), .A2(n15932), .ZN(n16859) );
  INV_X1 U19401 ( .A(n16859), .ZN(n15960) );
  OAI21_X1 U19402 ( .B1(n15952), .B2(n15951), .A(n16273), .ZN(n15953) );
  XNOR2_X1 U19403 ( .A(n15953), .B(n9737), .ZN(n15956) );
  AOI22_X1 U19404 ( .A1(n16292), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n20076), .ZN(n15954) );
  OAI21_X1 U19405 ( .B1(n16576), .B2(n20092), .A(n15954), .ZN(n15955) );
  AOI21_X1 U19406 ( .B1(n20083), .B2(n15956), .A(n15955), .ZN(n15957) );
  OAI21_X1 U19407 ( .B1(n15958), .B2(n20073), .A(n15957), .ZN(n15959) );
  AOI21_X1 U19408 ( .B1(n15960), .B2(n16301), .A(n15959), .ZN(n15961) );
  OAI21_X1 U19409 ( .B1(n16853), .B2(n20077), .A(n15961), .ZN(P2_U2832) );
  INV_X1 U19410 ( .A(n15945), .ZN(n15965) );
  NAND2_X1 U19411 ( .A1(n15962), .A2(n15963), .ZN(n15964) );
  NAND2_X1 U19412 ( .A1(n15965), .A2(n15964), .ZN(n16870) );
  NAND2_X1 U19413 ( .A1(n15987), .A2(n15967), .ZN(n15968) );
  NAND2_X1 U19414 ( .A1(n15969), .A2(n15968), .ZN(n16869) );
  INV_X1 U19415 ( .A(n16869), .ZN(n15981) );
  INV_X1 U19416 ( .A(n16607), .ZN(n15972) );
  NOR2_X1 U19417 ( .A1(n20080), .A2(n15970), .ZN(n15989) );
  INV_X1 U19418 ( .A(n15989), .ZN(n15971) );
  OAI21_X1 U19419 ( .B1(n20080), .B2(n15972), .A(n15971), .ZN(n15974) );
  OAI21_X1 U19420 ( .B1(n16590), .B2(n15974), .A(n20083), .ZN(n15973) );
  AOI21_X1 U19421 ( .B1(n16590), .B2(n15974), .A(n15973), .ZN(n15977) );
  OAI22_X1 U19422 ( .A1(n20072), .A2(n15975), .B1(n16589), .B2(n16262), .ZN(
        n15976) );
  AOI211_X1 U19423 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15977), .B(n15976), .ZN(n15978) );
  OAI21_X1 U19424 ( .B1(n15979), .B2(n20073), .A(n15978), .ZN(n15980) );
  AOI21_X1 U19425 ( .B1(n15981), .B2(n16301), .A(n15980), .ZN(n15982) );
  OAI21_X1 U19426 ( .B1(n16870), .B2(n20077), .A(n15982), .ZN(P2_U2833) );
  NAND2_X1 U19427 ( .A1(n12462), .A2(n15983), .ZN(n15984) );
  NAND2_X1 U19428 ( .A1(n15962), .A2(n15984), .ZN(n16876) );
  OR2_X1 U19429 ( .A1(n12457), .A2(n15985), .ZN(n15986) );
  NAND2_X1 U19430 ( .A1(n15987), .A2(n15986), .ZN(n16883) );
  INV_X1 U19431 ( .A(n16883), .ZN(n15995) );
  OAI21_X1 U19432 ( .B1(n16607), .B2(n15989), .A(n20083), .ZN(n15988) );
  AOI21_X1 U19433 ( .B1(n16607), .B2(n15989), .A(n15988), .ZN(n15991) );
  INV_X1 U19434 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20839) );
  OAI22_X1 U19435 ( .A1(n16605), .A2(n20092), .B1(n20839), .B2(n16262), .ZN(
        n15990) );
  AOI211_X1 U19436 ( .C1(n16292), .C2(P2_EBX_REG_21__SCAN_IN), .A(n15991), .B(
        n15990), .ZN(n15992) );
  OAI21_X1 U19437 ( .B1(n15993), .B2(n20073), .A(n15992), .ZN(n15994) );
  AOI21_X1 U19438 ( .B1(n15995), .B2(n16301), .A(n15994), .ZN(n15996) );
  OAI21_X1 U19439 ( .B1(n16876), .B2(n20077), .A(n15996), .ZN(P2_U2834) );
  NOR2_X1 U19440 ( .A1(n16361), .A2(n20087), .ZN(n16009) );
  AND2_X1 U19441 ( .A1(n15997), .A2(n16290), .ZN(n16008) );
  NAND2_X1 U19442 ( .A1(n16005), .A2(n20083), .ZN(n15998) );
  AOI21_X1 U19443 ( .B1(n15998), .B2(n16288), .A(n15999), .ZN(n16007) );
  NAND2_X1 U19444 ( .A1(n16250), .A2(n15999), .ZN(n16004) );
  OAI22_X1 U19445 ( .A1(n20072), .A2(n16360), .B1(n16000), .B2(n16262), .ZN(
        n16001) );
  INV_X1 U19446 ( .A(n16001), .ZN(n16003) );
  NAND2_X1 U19447 ( .A1(n16275), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16002) );
  OAI211_X1 U19448 ( .C1(n16005), .C2(n16004), .A(n16003), .B(n16002), .ZN(
        n16006) );
  NOR4_X1 U19449 ( .A1(n16009), .A2(n16008), .A3(n16007), .A4(n16006), .ZN(
        n16010) );
  OAI21_X1 U19450 ( .B1(n16493), .B2(n20077), .A(n16010), .ZN(P2_U2835) );
  NOR2_X1 U19451 ( .A1(n16028), .A2(n16011), .ZN(n16012) );
  OR2_X1 U19452 ( .A1(n12459), .A2(n16012), .ZN(n16894) );
  AND2_X1 U19453 ( .A1(n16013), .A2(n16014), .ZN(n16015) );
  NOR2_X1 U19454 ( .A1(n12463), .A2(n16015), .ZN(n16888) );
  NAND2_X1 U19455 ( .A1(n16888), .A2(n16294), .ZN(n16027) );
  INV_X1 U19456 ( .A(n16016), .ZN(n16025) );
  AOI21_X1 U19457 ( .B1(n16017), .B2(n20083), .A(n16282), .ZN(n16023) );
  NAND2_X1 U19458 ( .A1(n16292), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16018) );
  OAI211_X1 U19459 ( .C1(n20836), .C2(n16262), .A(n16018), .B(n20207), .ZN(
        n16019) );
  AOI21_X1 U19460 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16275), .A(
        n16019), .ZN(n16022) );
  NAND3_X1 U19461 ( .A1(n16617), .A2(n16250), .A3(n16020), .ZN(n16021) );
  OAI211_X1 U19462 ( .C1(n16023), .C2(n16617), .A(n16022), .B(n16021), .ZN(
        n16024) );
  AOI21_X1 U19463 ( .B1(n16025), .B2(n16290), .A(n16024), .ZN(n16026) );
  OAI211_X1 U19464 ( .C1(n16894), .C2(n20087), .A(n16027), .B(n16026), .ZN(
        P2_U2836) );
  AOI21_X1 U19465 ( .B1(n16029), .B2(n16043), .A(n16028), .ZN(n16629) );
  INV_X1 U19466 ( .A(n16629), .ZN(n16905) );
  NOR3_X1 U19467 ( .A1(n10228), .A2(n9738), .A3(n16297), .ZN(n16035) );
  AOI21_X1 U19468 ( .B1(n20083), .B2(n9738), .A(n16282), .ZN(n16033) );
  NAND2_X1 U19469 ( .A1(n16292), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16030) );
  OAI211_X1 U19470 ( .C1(n20834), .C2(n16262), .A(n16030), .B(n20207), .ZN(
        n16031) );
  AOI21_X1 U19471 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16275), .A(
        n16031), .ZN(n16032) );
  OAI21_X1 U19472 ( .B1(n16625), .B2(n16033), .A(n16032), .ZN(n16034) );
  AOI211_X1 U19473 ( .C1(n16036), .C2(n16290), .A(n16035), .B(n16034), .ZN(
        n16041) );
  INV_X1 U19474 ( .A(n16013), .ZN(n16038) );
  AOI21_X1 U19475 ( .B1(n16039), .B2(n16037), .A(n16038), .ZN(n16907) );
  NAND2_X1 U19476 ( .A1(n16907), .A2(n16294), .ZN(n16040) );
  OAI211_X1 U19477 ( .C1(n16905), .C2(n20087), .A(n16041), .B(n16040), .ZN(
        P2_U2837) );
  INV_X1 U19478 ( .A(n16042), .ZN(n16044) );
  OAI21_X1 U19479 ( .B1(n9657), .B2(n16044), .A(n16043), .ZN(n16917) );
  INV_X1 U19480 ( .A(n16037), .ZN(n16046) );
  AOI21_X1 U19481 ( .B1(n16047), .B2(n16045), .A(n16046), .ZN(n16920) );
  NAND2_X1 U19482 ( .A1(n16920), .A2(n16294), .ZN(n16058) );
  OAI21_X1 U19483 ( .B1(n16048), .B2(n16274), .A(n16288), .ZN(n16056) );
  INV_X1 U19484 ( .A(n16638), .ZN(n16049) );
  NAND3_X1 U19485 ( .A1(n16049), .A2(n16250), .A3(n16048), .ZN(n16052) );
  OAI21_X1 U19486 ( .B1(n16262), .B2(n20832), .A(n20207), .ZN(n16050) );
  AOI21_X1 U19487 ( .B1(n16292), .B2(P2_EBX_REG_17__SCAN_IN), .A(n16050), .ZN(
        n16051) );
  OAI211_X1 U19488 ( .C1(n20092), .C2(n16635), .A(n16052), .B(n16051), .ZN(
        n16055) );
  NOR2_X1 U19489 ( .A1(n16053), .A2(n20073), .ZN(n16054) );
  AOI211_X1 U19490 ( .C1(n16638), .C2(n16056), .A(n16055), .B(n16054), .ZN(
        n16057) );
  OAI211_X1 U19491 ( .C1(n20087), .C2(n16917), .A(n16058), .B(n16057), .ZN(
        P2_U2838) );
  OAI21_X1 U19492 ( .B1(n14475), .B2(n16059), .A(n16045), .ZN(n20117) );
  AOI21_X1 U19493 ( .B1(n16061), .B2(n16060), .A(n9657), .ZN(n16926) );
  NAND2_X1 U19494 ( .A1(n16926), .A2(n16301), .ZN(n16074) );
  NAND2_X1 U19495 ( .A1(n16065), .A2(n20083), .ZN(n16062) );
  NAND2_X1 U19496 ( .A1(n16062), .A2(n16288), .ZN(n16063) );
  NAND2_X1 U19497 ( .A1(n16063), .A2(n10227), .ZN(n16070) );
  OAI21_X1 U19498 ( .B1(n16262), .B2(n16643), .A(n20207), .ZN(n16064) );
  AOI21_X1 U19499 ( .B1(n16292), .B2(P2_EBX_REG_16__SCAN_IN), .A(n16064), .ZN(
        n16069) );
  INV_X1 U19500 ( .A(n16065), .ZN(n16066) );
  NAND3_X1 U19501 ( .A1(n16066), .A2(n16250), .A3(n16645), .ZN(n16068) );
  NAND2_X1 U19502 ( .A1(n16275), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16067) );
  NAND4_X1 U19503 ( .A1(n16070), .A2(n16069), .A3(n16068), .A4(n16067), .ZN(
        n16071) );
  AOI21_X1 U19504 ( .B1(n16072), .B2(n16290), .A(n16071), .ZN(n16073) );
  OAI211_X1 U19505 ( .C1(n20077), .C2(n20117), .A(n16074), .B(n16073), .ZN(
        P2_U2839) );
  OAI21_X1 U19506 ( .B1(n16075), .B2(n16076), .A(n16060), .ZN(n16939) );
  INV_X1 U19507 ( .A(n16939), .ZN(n16656) );
  NOR2_X1 U19508 ( .A1(n16077), .A2(n20080), .ZN(n16078) );
  XNOR2_X1 U19509 ( .A(n16078), .B(n16654), .ZN(n16082) );
  AOI21_X1 U19510 ( .B1(n20076), .B2(P2_REIP_REG_15__SCAN_IN), .A(n20179), 
        .ZN(n16080) );
  NAND2_X1 U19511 ( .A1(n16275), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16079) );
  OAI211_X1 U19512 ( .C1(n20072), .C2(n11031), .A(n16080), .B(n16079), .ZN(
        n16081) );
  AOI21_X1 U19513 ( .B1(n16082), .B2(n20083), .A(n16081), .ZN(n16083) );
  OAI21_X1 U19514 ( .B1(n16084), .B2(n20073), .A(n16083), .ZN(n16085) );
  AOI21_X1 U19515 ( .B1(n16656), .B2(n16301), .A(n16085), .ZN(n16086) );
  OAI21_X1 U19516 ( .B1(n16934), .B2(n20077), .A(n16086), .ZN(P2_U2840) );
  NOR2_X1 U19517 ( .A1(n16087), .A2(n16088), .ZN(n16089) );
  OR2_X1 U19518 ( .A1(n16075), .A2(n16089), .ZN(n16948) );
  NAND2_X1 U19519 ( .A1(n16952), .A2(n16294), .ZN(n16099) );
  NOR2_X1 U19520 ( .A1(n16090), .A2(n20080), .ZN(n16104) );
  XNOR2_X1 U19521 ( .A(n16104), .B(n16664), .ZN(n16097) );
  OAI21_X1 U19522 ( .B1(n16262), .B2(n20827), .A(n20207), .ZN(n16091) );
  AOI21_X1 U19523 ( .B1(n16292), .B2(P2_EBX_REG_14__SCAN_IN), .A(n16091), .ZN(
        n16092) );
  OAI21_X1 U19524 ( .B1(n16093), .B2(n20092), .A(n16092), .ZN(n16096) );
  NOR2_X1 U19525 ( .A1(n16094), .A2(n20073), .ZN(n16095) );
  AOI211_X1 U19526 ( .C1(n20083), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        n16098) );
  OAI211_X1 U19527 ( .C1(n20087), .C2(n16948), .A(n16099), .B(n16098), .ZN(
        P2_U2841) );
  AOI21_X1 U19528 ( .B1(n16101), .B2(n16100), .A(n16087), .ZN(n16965) );
  INV_X1 U19529 ( .A(n16102), .ZN(n16110) );
  INV_X1 U19530 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n16398) );
  OR2_X1 U19531 ( .A1(n16262), .A2(n16675), .ZN(n16103) );
  OAI211_X1 U19532 ( .C1(n20072), .C2(n16398), .A(n20207), .B(n16103), .ZN(
        n16108) );
  OAI211_X1 U19533 ( .C1(n16105), .C2(n16678), .A(n16104), .B(n20083), .ZN(
        n16106) );
  OAI21_X1 U19534 ( .B1(n16288), .B2(n16678), .A(n16106), .ZN(n16107) );
  AOI211_X1 U19535 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16275), .A(
        n16108), .B(n16107), .ZN(n16109) );
  OAI21_X1 U19536 ( .B1(n16110), .B2(n20073), .A(n16109), .ZN(n16111) );
  AOI21_X1 U19537 ( .B1(n16965), .B2(n16301), .A(n16111), .ZN(n16112) );
  OAI21_X1 U19538 ( .B1(n20077), .B2(n16967), .A(n16112), .ZN(P2_U2842) );
  INV_X1 U19539 ( .A(n16100), .ZN(n16114) );
  AOI21_X1 U19540 ( .B1(n16115), .B2(n16113), .A(n16114), .ZN(n20095) );
  INV_X1 U19541 ( .A(n20095), .ZN(n16116) );
  NOR2_X1 U19542 ( .A1(n16116), .A2(n20087), .ZN(n16130) );
  NAND2_X1 U19543 ( .A1(n20083), .A2(n16118), .ZN(n16117) );
  AOI21_X1 U19544 ( .B1(n16288), .B2(n16117), .A(n16687), .ZN(n16129) );
  INV_X1 U19545 ( .A(n16118), .ZN(n16119) );
  NAND2_X1 U19546 ( .A1(n16687), .A2(n16119), .ZN(n16120) );
  NOR2_X1 U19547 ( .A1(n16297), .A2(n16120), .ZN(n16128) );
  INV_X1 U19548 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n20098) );
  INV_X1 U19549 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16121) );
  OAI22_X1 U19550 ( .A1(n16122), .A2(n20073), .B1(n16121), .B2(n20092), .ZN(
        n16123) );
  INV_X1 U19551 ( .A(n16123), .ZN(n16124) );
  OAI21_X1 U19552 ( .B1(n20072), .B2(n20098), .A(n16124), .ZN(n16125) );
  INV_X1 U19553 ( .A(n16125), .ZN(n16126) );
  OAI211_X1 U19554 ( .C1(n16262), .C2(n16685), .A(n20207), .B(n16126), .ZN(
        n16127) );
  NOR4_X1 U19555 ( .A1(n16130), .A2(n16129), .A3(n16128), .A4(n16127), .ZN(
        n16131) );
  OAI21_X1 U19556 ( .B1(n16132), .B2(n20077), .A(n16131), .ZN(P2_U2843) );
  OR2_X1 U19557 ( .A1(n16147), .A2(n16133), .ZN(n16134) );
  NAND2_X1 U19558 ( .A1(n16113), .A2(n16134), .ZN(n16711) );
  NAND2_X1 U19559 ( .A1(n16992), .A2(n16294), .ZN(n16144) );
  OAI21_X1 U19560 ( .B1(n16274), .B2(n16136), .A(n16288), .ZN(n16142) );
  INV_X1 U19561 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16706) );
  OAI21_X1 U19562 ( .B1(n16262), .B2(n16706), .A(n20207), .ZN(n16135) );
  AOI21_X1 U19563 ( .B1(n16292), .B2(P2_EBX_REG_11__SCAN_IN), .A(n16135), .ZN(
        n16138) );
  NAND3_X1 U19564 ( .A1(n16250), .A2(n10232), .A3(n16136), .ZN(n16137) );
  OAI211_X1 U19565 ( .C1(n20092), .C2(n16707), .A(n16138), .B(n16137), .ZN(
        n16141) );
  NOR2_X1 U19566 ( .A1(n16139), .A2(n20073), .ZN(n16140) );
  AOI211_X1 U19567 ( .C1(n16709), .C2(n16142), .A(n16141), .B(n16140), .ZN(
        n16143) );
  OAI211_X1 U19568 ( .C1(n20087), .C2(n16711), .A(n16144), .B(n16143), .ZN(
        P2_U2844) );
  AND2_X1 U19569 ( .A1(n16163), .A2(n16145), .ZN(n16146) );
  NOR2_X1 U19570 ( .A1(n16147), .A2(n16146), .ZN(n20105) );
  AOI21_X1 U19571 ( .B1(n20083), .B2(n16152), .A(n16282), .ZN(n16156) );
  INV_X1 U19572 ( .A(n16148), .ZN(n16149) );
  AOI22_X1 U19573 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16275), .B1(
        n16149), .B2(n16290), .ZN(n16150) );
  OAI21_X1 U19574 ( .B1(n20072), .B2(n20107), .A(n16150), .ZN(n16151) );
  AOI211_X1 U19575 ( .C1(n20076), .C2(P2_REIP_REG_10__SCAN_IN), .A(n20179), 
        .B(n16151), .ZN(n16155) );
  INV_X1 U19576 ( .A(n16152), .ZN(n16153) );
  NAND3_X1 U19577 ( .A1(n16250), .A2(n16724), .A3(n16153), .ZN(n16154) );
  OAI211_X1 U19578 ( .C1(n16156), .C2(n16724), .A(n16155), .B(n16154), .ZN(
        n16157) );
  AOI21_X1 U19579 ( .B1(n20105), .B2(n16301), .A(n16157), .ZN(n16158) );
  OAI21_X1 U19580 ( .B1(n20077), .B2(n16159), .A(n16158), .ZN(P2_U2845) );
  NAND2_X1 U19581 ( .A1(n16160), .A2(n16161), .ZN(n16162) );
  NAND2_X1 U19582 ( .A1(n16163), .A2(n16162), .ZN(n17012) );
  NAND2_X1 U19583 ( .A1(n17018), .A2(n16294), .ZN(n16175) );
  INV_X1 U19584 ( .A(n16167), .ZN(n16164) );
  AOI21_X1 U19585 ( .B1(n20083), .B2(n16164), .A(n16282), .ZN(n16171) );
  INV_X1 U19586 ( .A(n16735), .ZN(n16170) );
  OAI21_X1 U19587 ( .B1(n20821), .B2(n16262), .A(n20207), .ZN(n16166) );
  NOR2_X1 U19588 ( .A1(n20072), .A2(n10376), .ZN(n16165) );
  AOI211_X1 U19589 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16166), .B(n16165), .ZN(n16169) );
  NAND3_X1 U19590 ( .A1(n16250), .A2(n16170), .A3(n16167), .ZN(n16168) );
  OAI211_X1 U19591 ( .C1(n16171), .C2(n16170), .A(n16169), .B(n16168), .ZN(
        n16172) );
  AOI21_X1 U19592 ( .B1(n16173), .B2(n16290), .A(n16172), .ZN(n16174) );
  OAI211_X1 U19593 ( .C1(n17012), .C2(n20087), .A(n16175), .B(n16174), .ZN(
        P2_U2846) );
  NAND2_X1 U19594 ( .A1(n16176), .A2(n16177), .ZN(n16178) );
  NAND2_X1 U19595 ( .A1(n16160), .A2(n16178), .ZN(n17029) );
  INV_X1 U19596 ( .A(n17029), .ZN(n16747) );
  NOR2_X1 U19597 ( .A1(n16179), .A2(n20073), .ZN(n16188) );
  AOI21_X1 U19598 ( .B1(n20083), .B2(n16182), .A(n16282), .ZN(n16186) );
  OAI21_X1 U19599 ( .B1(n20819), .B2(n16262), .A(n20207), .ZN(n16181) );
  INV_X1 U19600 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n16410) );
  NOR2_X1 U19601 ( .A1(n20072), .A2(n16410), .ZN(n16180) );
  AOI211_X1 U19602 ( .C1(n16275), .C2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16181), .B(n16180), .ZN(n16185) );
  INV_X1 U19603 ( .A(n16182), .ZN(n16183) );
  NAND3_X1 U19604 ( .A1(n16250), .A2(n16745), .A3(n16183), .ZN(n16184) );
  OAI211_X1 U19605 ( .C1(n16186), .C2(n16745), .A(n16185), .B(n16184), .ZN(
        n16187) );
  AOI211_X1 U19606 ( .C1(n16747), .C2(n15862), .A(n16188), .B(n16187), .ZN(
        n16189) );
  OAI21_X1 U19607 ( .B1(n20077), .B2(n17023), .A(n16189), .ZN(P2_U2847) );
  OR2_X1 U19608 ( .A1(n14203), .A2(n16190), .ZN(n16191) );
  NAND2_X1 U19609 ( .A1(n16176), .A2(n16191), .ZN(n16764) );
  INV_X1 U19610 ( .A(n16764), .ZN(n17039) );
  INV_X1 U19611 ( .A(n16196), .ZN(n16192) );
  AOI21_X1 U19612 ( .B1(n20083), .B2(n16192), .A(n16282), .ZN(n16200) );
  INV_X1 U19613 ( .A(n16762), .ZN(n16199) );
  AOI22_X1 U19614 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16275), .B1(
        n16290), .B2(n16193), .ZN(n16194) );
  OAI211_X1 U19615 ( .C1(n20817), .C2(n16262), .A(n16194), .B(n20207), .ZN(
        n16195) );
  AOI21_X1 U19616 ( .B1(n16292), .B2(P2_EBX_REG_7__SCAN_IN), .A(n16195), .ZN(
        n16198) );
  NAND3_X1 U19617 ( .A1(n16250), .A2(n16196), .A3(n16199), .ZN(n16197) );
  OAI211_X1 U19618 ( .C1(n16200), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        n16201) );
  AOI21_X1 U19619 ( .B1(n17039), .B2(n16301), .A(n16201), .ZN(n16202) );
  OAI21_X1 U19620 ( .B1(n20077), .B2(n17044), .A(n16202), .ZN(P2_U2848) );
  OR2_X1 U19621 ( .A1(n16204), .A2(n16203), .ZN(n16205) );
  NAND2_X1 U19622 ( .A1(n16206), .A2(n16205), .ZN(n17077) );
  OAI21_X1 U19623 ( .B1(n11346), .B2(n16262), .A(n20207), .ZN(n16215) );
  OAI21_X1 U19624 ( .B1(n16208), .B2(n16274), .A(n16288), .ZN(n16212) );
  INV_X1 U19625 ( .A(n17638), .ZN(n16207) );
  NAND3_X1 U19626 ( .A1(n16250), .A2(n16208), .A3(n16207), .ZN(n16210) );
  NAND2_X1 U19627 ( .A1(n16275), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16209) );
  OAI211_X1 U19628 ( .C1(n20072), .C2(n10961), .A(n16210), .B(n16209), .ZN(
        n16211) );
  AOI21_X1 U19629 ( .B1(n17638), .B2(n16212), .A(n16211), .ZN(n16213) );
  OAI21_X1 U19630 ( .B1(n17067), .B2(n20073), .A(n16213), .ZN(n16214) );
  AOI211_X1 U19631 ( .C1(n17640), .C2(n15862), .A(n16215), .B(n16214), .ZN(
        n16216) );
  OAI21_X1 U19632 ( .B1(n20077), .B2(n17077), .A(n16216), .ZN(P2_U2850) );
  INV_X1 U19633 ( .A(n16217), .ZN(n16223) );
  INV_X1 U19634 ( .A(n16220), .ZN(n16221) );
  NAND3_X1 U19635 ( .A1(n16218), .A2(n16219), .A3(n16221), .ZN(n16222) );
  NAND2_X1 U19636 ( .A1(n16223), .A2(n16222), .ZN(n20126) );
  XNOR2_X1 U19637 ( .A(n16224), .B(n16225), .ZN(n20124) );
  NAND2_X1 U19638 ( .A1(n16227), .A2(n16226), .ZN(n16228) );
  AND2_X1 U19639 ( .A1(n14097), .A2(n16228), .ZN(n20181) );
  NAND2_X1 U19640 ( .A1(n20181), .A2(n16301), .ZN(n16242) );
  OAI21_X1 U19641 ( .B1(n16262), .B2(n11104), .A(n20207), .ZN(n16229) );
  AOI21_X1 U19642 ( .B1(n16292), .B2(P2_EBX_REG_4__SCAN_IN), .A(n16229), .ZN(
        n16238) );
  INV_X1 U19643 ( .A(n16232), .ZN(n16230) );
  NOR2_X1 U19644 ( .A1(n16274), .A2(n16230), .ZN(n16231) );
  INV_X1 U19645 ( .A(n20185), .ZN(n16233) );
  OAI21_X1 U19646 ( .B1(n16282), .B2(n16231), .A(n16233), .ZN(n16237) );
  NOR2_X1 U19647 ( .A1(n16233), .A2(n16232), .ZN(n16234) );
  NAND2_X1 U19648 ( .A1(n16250), .A2(n16234), .ZN(n16236) );
  NAND2_X1 U19649 ( .A1(n16275), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16235) );
  NAND4_X1 U19650 ( .A1(n16238), .A2(n16237), .A3(n16236), .A4(n16235), .ZN(
        n16240) );
  NOR2_X1 U19651 ( .A1(n17082), .A2(n20073), .ZN(n16239) );
  NOR2_X1 U19652 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  OAI211_X1 U19653 ( .C1(n20124), .C2(n20077), .A(n16242), .B(n16241), .ZN(
        n16243) );
  INV_X1 U19654 ( .A(n16243), .ZN(n16244) );
  OAI21_X1 U19655 ( .B1(n20126), .B2(n16303), .A(n16244), .ZN(P2_U2851) );
  NAND2_X1 U19656 ( .A1(n16246), .A2(n16245), .ZN(n16247) );
  AND2_X1 U19657 ( .A1(n16224), .A2(n16247), .ZN(n20878) );
  NOR2_X1 U19658 ( .A1(n16248), .A2(n20073), .ZN(n16257) );
  INV_X1 U19659 ( .A(n17645), .ZN(n16249) );
  NAND3_X1 U19660 ( .A1(n16250), .A2(n16251), .A3(n16249), .ZN(n16254) );
  NOR2_X1 U19661 ( .A1(n16251), .A2(n16274), .ZN(n16252) );
  OAI21_X1 U19662 ( .B1(n16282), .B2(n16252), .A(n17645), .ZN(n16253) );
  OAI211_X1 U19663 ( .C1(n20072), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        n16256) );
  AOI211_X1 U19664 ( .C1(n20878), .C2(n16294), .A(n16257), .B(n16256), .ZN(
        n16260) );
  INV_X1 U19665 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20811) );
  OAI22_X1 U19666 ( .A1(n17655), .A2(n20092), .B1(n20811), .B2(n16262), .ZN(
        n16258) );
  AOI21_X1 U19667 ( .B1(n16301), .B2(n9615), .A(n16258), .ZN(n16259) );
  OAI211_X1 U19668 ( .C1(n17184), .C2(n16303), .A(n16260), .B(n16259), .ZN(
        P2_U2852) );
  AOI21_X1 U19669 ( .B1(n20083), .B2(n16271), .A(n16282), .ZN(n16267) );
  INV_X1 U19670 ( .A(n20200), .ZN(n16261) );
  NOR3_X1 U19671 ( .A1(n16297), .A2(n16271), .A3(n16261), .ZN(n16265) );
  OAI22_X1 U19672 ( .A1(n20072), .A2(n16263), .B1(n20809), .B2(n16262), .ZN(
        n16264) );
  OAI21_X1 U19673 ( .B1(n20889), .B2(n16303), .A(n16268), .ZN(P2_U2853) );
  AND2_X1 U19674 ( .A1(n16269), .A2(n16289), .ZN(n16270) );
  NOR2_X1 U19675 ( .A1(n16271), .A2(n16270), .ZN(n16272) );
  NAND2_X1 U19676 ( .A1(n16273), .A2(n16272), .ZN(n17144) );
  NOR2_X1 U19677 ( .A1(n17144), .A2(n16274), .ZN(n16281) );
  INV_X1 U19678 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n16279) );
  AOI22_X1 U19679 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16275), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n20076), .ZN(n16278) );
  NAND2_X1 U19680 ( .A1(n16290), .A2(n16276), .ZN(n16277) );
  OAI211_X1 U19681 ( .C1(n20072), .C2(n16279), .A(n16278), .B(n16277), .ZN(
        n16280) );
  AOI211_X1 U19682 ( .C1(n20208), .C2(n16282), .A(n16281), .B(n16280), .ZN(
        n16283) );
  OAI21_X1 U19683 ( .B1(n16284), .B2(n20077), .A(n16283), .ZN(n16285) );
  AOI21_X1 U19684 ( .B1(n20214), .B2(n16301), .A(n16285), .ZN(n16286) );
  OAI21_X1 U19685 ( .B1(n20251), .B2(n16303), .A(n16286), .ZN(P2_U2854) );
  INV_X1 U19686 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16287) );
  AOI21_X1 U19687 ( .B1(n20092), .B2(n16288), .A(n16287), .ZN(n16299) );
  INV_X1 U19688 ( .A(n16289), .ZN(n17126) );
  AOI22_X1 U19689 ( .A1(n16292), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n16291), .B2(
        n16290), .ZN(n16296) );
  AOI22_X1 U19690 ( .A1(n16294), .A2(n16293), .B1(n20076), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n16295) );
  OAI211_X1 U19691 ( .C1(n16297), .C2(n17126), .A(n16296), .B(n16295), .ZN(
        n16298) );
  AOI211_X1 U19692 ( .C1(n16301), .C2(n16300), .A(n16299), .B(n16298), .ZN(
        n16302) );
  OAI21_X1 U19693 ( .B1(n17220), .B2(n16303), .A(n16302), .ZN(P2_U2855) );
  OR2_X1 U19694 ( .A1(n16305), .A2(n16304), .ZN(n16425) );
  NAND3_X1 U19695 ( .A1(n16425), .A2(n16306), .A3(n20108), .ZN(n16308) );
  NAND2_X1 U19696 ( .A1(n16418), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16307) );
  OAI211_X1 U19697 ( .C1(n16418), .C2(n16781), .A(n16308), .B(n16307), .ZN(
        P2_U2858) );
  NAND2_X1 U19698 ( .A1(n16310), .A2(n16309), .ZN(n16312) );
  XNOR2_X1 U19699 ( .A(n16312), .B(n16311), .ZN(n16439) );
  NOR2_X1 U19700 ( .A1(n16794), .A2(n16418), .ZN(n16313) );
  AOI21_X1 U19701 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16418), .A(n16313), .ZN(
        n16314) );
  OAI21_X1 U19702 ( .B1(n16439), .B2(n20101), .A(n16314), .ZN(P2_U2859) );
  OAI21_X1 U19703 ( .B1(n16315), .B2(n16317), .A(n16316), .ZN(n16446) );
  NOR2_X1 U19704 ( .A1(n16318), .A2(n16418), .ZN(n16319) );
  AOI21_X1 U19705 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16418), .A(n16319), .ZN(
        n16320) );
  OAI21_X1 U19706 ( .B1(n16446), .B2(n20101), .A(n16320), .ZN(P2_U2860) );
  NAND2_X1 U19707 ( .A1(n16334), .A2(n16333), .ZN(n16332) );
  NAND2_X1 U19708 ( .A1(n16332), .A2(n16322), .ZN(n16328) );
  NAND2_X1 U19709 ( .A1(n16324), .A2(n16323), .ZN(n16326) );
  XOR2_X1 U19710 ( .A(n16326), .B(n16325), .Z(n16327) );
  XNOR2_X1 U19711 ( .A(n16328), .B(n16327), .ZN(n16453) );
  INV_X1 U19712 ( .A(n16329), .ZN(n16819) );
  MUX2_X1 U19713 ( .A(n16330), .B(n16819), .S(n20112), .Z(n16331) );
  OAI21_X1 U19714 ( .B1(n16453), .B2(n20101), .A(n16331), .ZN(P2_U2861) );
  OAI21_X1 U19715 ( .B1(n16334), .B2(n16333), .A(n16332), .ZN(n16459) );
  NOR2_X1 U19716 ( .A1(n16832), .A2(n16418), .ZN(n16335) );
  AOI21_X1 U19717 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16418), .A(n16335), .ZN(
        n16336) );
  OAI21_X1 U19718 ( .B1(n16459), .B2(n20101), .A(n16336), .ZN(P2_U2862) );
  AOI21_X1 U19719 ( .B1(n16337), .B2(n16338), .A(n9686), .ZN(n16339) );
  XOR2_X1 U19720 ( .A(n16340), .B(n16339), .Z(n16466) );
  NOR2_X1 U19721 ( .A1(n16570), .A2(n16418), .ZN(n16341) );
  AOI21_X1 U19722 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16418), .A(n16341), .ZN(
        n16342) );
  OAI21_X1 U19723 ( .B1(n16466), .B2(n20101), .A(n16342), .ZN(P2_U2863) );
  AOI21_X1 U19724 ( .B1(n16343), .B2(n16346), .A(n16345), .ZN(n16467) );
  NAND2_X1 U19725 ( .A1(n16467), .A2(n20108), .ZN(n16348) );
  NAND2_X1 U19726 ( .A1(n16418), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16347) );
  OAI211_X1 U19727 ( .C1(n16859), .C2(n16418), .A(n16348), .B(n16347), .ZN(
        P2_U2864) );
  AOI21_X1 U19728 ( .B1(n16350), .B2(n16349), .A(n13408), .ZN(n16477) );
  NAND2_X1 U19729 ( .A1(n16477), .A2(n20108), .ZN(n16352) );
  NAND2_X1 U19730 ( .A1(n16418), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16351) );
  OAI211_X1 U19731 ( .C1(n16869), .C2(n16418), .A(n16352), .B(n16351), .ZN(
        P2_U2865) );
  NAND2_X1 U19732 ( .A1(n16353), .A2(n16354), .ZN(n16355) );
  NAND2_X1 U19733 ( .A1(n16349), .A2(n16355), .ZN(n16486) );
  MUX2_X1 U19734 ( .A(n16883), .B(n16356), .S(n16418), .Z(n16357) );
  OAI21_X1 U19735 ( .B1(n20101), .B2(n16486), .A(n16357), .ZN(P2_U2866) );
  OAI21_X1 U19736 ( .B1(n16358), .B2(n16359), .A(n16353), .ZN(n16489) );
  MUX2_X1 U19737 ( .A(n16361), .B(n16360), .S(n16418), .Z(n16362) );
  OAI21_X1 U19738 ( .B1(n20101), .B2(n16489), .A(n16362), .ZN(P2_U2867) );
  OAI21_X1 U19739 ( .B1(n9642), .B2(n16363), .A(n10153), .ZN(n16502) );
  NOR2_X1 U19740 ( .A1(n16894), .A2(n16418), .ZN(n16364) );
  AOI21_X1 U19741 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16418), .A(n16364), .ZN(
        n16365) );
  OAI21_X1 U19742 ( .B1(n20101), .B2(n16502), .A(n16365), .ZN(P2_U2868) );
  AOI21_X1 U19743 ( .B1(n16367), .B2(n16366), .A(n9642), .ZN(n16507) );
  NAND2_X1 U19744 ( .A1(n16507), .A2(n20108), .ZN(n16369) );
  NAND2_X1 U19745 ( .A1(n16418), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16368) );
  OAI211_X1 U19746 ( .C1(n16905), .C2(n16418), .A(n16369), .B(n16368), .ZN(
        P2_U2869) );
  INV_X1 U19747 ( .A(n16366), .ZN(n16371) );
  AOI21_X1 U19748 ( .B1(n16372), .B2(n16370), .A(n16371), .ZN(n16515) );
  NAND2_X1 U19749 ( .A1(n16515), .A2(n20108), .ZN(n16374) );
  NAND2_X1 U19750 ( .A1(n16418), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n16373) );
  OAI211_X1 U19751 ( .C1(n16917), .C2(n16418), .A(n16374), .B(n16373), .ZN(
        P2_U2870) );
  NAND2_X1 U19752 ( .A1(n16376), .A2(n16377), .ZN(n16378) );
  NAND2_X1 U19753 ( .A1(n16370), .A2(n16378), .ZN(n20118) );
  NOR2_X1 U19754 ( .A1(n20112), .A2(n16379), .ZN(n16380) );
  AOI21_X1 U19755 ( .B1(n16926), .B2(n20112), .A(n16380), .ZN(n16381) );
  OAI21_X1 U19756 ( .B1(n20101), .B2(n20118), .A(n16381), .ZN(P2_U2871) );
  NAND2_X1 U19757 ( .A1(n16656), .A2(n20112), .ZN(n16385) );
  OAI211_X1 U19758 ( .C1(n16382), .C2(n16383), .A(n16376), .B(n20108), .ZN(
        n16384) );
  OAI211_X1 U19759 ( .C1(n20112), .C2(n11031), .A(n16385), .B(n16384), .ZN(
        P2_U2872) );
  AOI211_X1 U19760 ( .C1(n16387), .C2(n16386), .A(n20101), .B(n16382), .ZN(
        n16389) );
  NOR2_X1 U19761 ( .A1(n16948), .A2(n16418), .ZN(n16388) );
  AOI211_X1 U19762 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n16418), .A(n16389), .B(
        n16388), .ZN(n16390) );
  INV_X1 U19763 ( .A(n16390), .ZN(P2_U2873) );
  NAND2_X1 U19764 ( .A1(n16415), .A2(n16409), .ZN(n16406) );
  NOR2_X1 U19765 ( .A1(n16406), .A2(n16405), .ZN(n20099) );
  NAND2_X1 U19766 ( .A1(n20099), .A2(n16392), .ZN(n16399) );
  NOR2_X1 U19767 ( .A1(n16399), .A2(n16393), .ZN(n20094) );
  INV_X1 U19768 ( .A(n20094), .ZN(n16400) );
  NOR2_X1 U19769 ( .A1(n16400), .A2(n20093), .ZN(n16395) );
  OAI211_X1 U19770 ( .C1(n16395), .C2(n16394), .A(n20108), .B(n16386), .ZN(
        n16397) );
  NAND2_X1 U19771 ( .A1(n16965), .A2(n20112), .ZN(n16396) );
  OAI211_X1 U19772 ( .C1(n20112), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        P2_U2874) );
  INV_X1 U19773 ( .A(n16399), .ZN(n20100) );
  OAI211_X1 U19774 ( .C1(n20100), .C2(n16401), .A(n16400), .B(n20108), .ZN(
        n16403) );
  INV_X1 U19775 ( .A(n16711), .ZN(n16987) );
  NAND2_X1 U19776 ( .A1(n16987), .A2(n20112), .ZN(n16402) );
  OAI211_X1 U19777 ( .C1(n20112), .C2(n16404), .A(n16403), .B(n16402), .ZN(
        P2_U2876) );
  XNOR2_X1 U19778 ( .A(n16406), .B(n16405), .ZN(n16408) );
  MUX2_X1 U19779 ( .A(n17012), .B(n10376), .S(n16418), .Z(n16407) );
  OAI21_X1 U19780 ( .B1(n16408), .B2(n20101), .A(n16407), .ZN(P2_U2878) );
  XNOR2_X1 U19781 ( .A(n16415), .B(n16409), .ZN(n16412) );
  MUX2_X1 U19782 ( .A(n16410), .B(n17029), .S(n20112), .Z(n16411) );
  OAI21_X1 U19783 ( .B1(n16412), .B2(n20101), .A(n16411), .ZN(P2_U2879) );
  NOR2_X1 U19784 ( .A1(n16414), .A2(n16413), .ZN(n16417) );
  INV_X1 U19785 ( .A(n16415), .ZN(n16416) );
  OAI211_X1 U19786 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n16417), .A(
        n16416), .B(n20108), .ZN(n16421) );
  MUX2_X1 U19787 ( .A(n16764), .B(n16419), .S(n16418), .Z(n16420) );
  NAND2_X1 U19788 ( .A1(n16421), .A2(n16420), .ZN(P2_U2880) );
  AOI22_X1 U19789 ( .A1(n20116), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20133), .ZN(n16423) );
  NAND2_X1 U19790 ( .A1(n20115), .A2(BUF2_REG_31__SCAN_IN), .ZN(n16422) );
  OAI211_X1 U19791 ( .C1(n16424), .C2(n16517), .A(n16423), .B(n16422), .ZN(
        P2_U2888) );
  NAND3_X1 U19792 ( .A1(n16425), .A2(n16306), .A3(n20128), .ZN(n16431) );
  INV_X1 U19793 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16428) );
  AOI22_X1 U19794 ( .A1(n20114), .A2(n16426), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n20133), .ZN(n16427) );
  OAI21_X1 U19795 ( .B1(n16513), .B2(n16428), .A(n16427), .ZN(n16429) );
  AOI21_X1 U19796 ( .B1(n20116), .B2(BUF1_REG_29__SCAN_IN), .A(n16429), .ZN(
        n16430) );
  OAI211_X1 U19797 ( .C1(n16517), .C2(n16432), .A(n16431), .B(n16430), .ZN(
        P2_U2890) );
  NAND2_X1 U19798 ( .A1(n20116), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16436) );
  NAND2_X1 U19799 ( .A1(n20115), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19800 ( .A1(n20114), .A2(n16433), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n20133), .ZN(n16434) );
  NAND3_X1 U19801 ( .A1(n16436), .A2(n16435), .A3(n16434), .ZN(n16437) );
  AOI21_X1 U19802 ( .B1(n16796), .B2(n20134), .A(n16437), .ZN(n16438) );
  OAI21_X1 U19803 ( .B1(n16439), .B2(n20138), .A(n16438), .ZN(P2_U2891) );
  INV_X1 U19804 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19805 ( .A1(n20114), .A2(n16440), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n20133), .ZN(n16441) );
  OAI21_X1 U19806 ( .B1(n16513), .B2(n16442), .A(n16441), .ZN(n16444) );
  NOR2_X1 U19807 ( .A1(n16810), .A2(n16517), .ZN(n16443) );
  AOI211_X1 U19808 ( .C1(n20116), .C2(BUF1_REG_27__SCAN_IN), .A(n16444), .B(
        n16443), .ZN(n16445) );
  OAI21_X1 U19809 ( .B1(n16446), .B2(n20138), .A(n16445), .ZN(P2_U2892) );
  INV_X1 U19810 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16450) );
  AOI22_X1 U19811 ( .A1(n20114), .A2(n16447), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n20133), .ZN(n16449) );
  NAND2_X1 U19812 ( .A1(n20116), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16448) );
  OAI211_X1 U19813 ( .C1(n16513), .C2(n16450), .A(n16449), .B(n16448), .ZN(
        n16451) );
  AOI21_X1 U19814 ( .B1(n16822), .B2(n20134), .A(n16451), .ZN(n16452) );
  OAI21_X1 U19815 ( .B1(n16453), .B2(n20138), .A(n16452), .ZN(P2_U2893) );
  AOI22_X1 U19816 ( .A1(n20114), .A2(n16454), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n20133), .ZN(n16456) );
  NAND2_X1 U19817 ( .A1(n20116), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16455) );
  OAI211_X1 U19818 ( .C1(n16513), .C2(n19429), .A(n16456), .B(n16455), .ZN(
        n16457) );
  AOI21_X1 U19819 ( .B1(n16835), .B2(n20134), .A(n16457), .ZN(n16458) );
  OAI21_X1 U19820 ( .B1(n16459), .B2(n20138), .A(n16458), .ZN(P2_U2894) );
  INV_X1 U19821 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19822 ( .A1(n20114), .A2(n16460), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n20133), .ZN(n16461) );
  OAI21_X1 U19823 ( .B1(n16513), .B2(n16462), .A(n16461), .ZN(n16464) );
  NOR2_X1 U19824 ( .A1(n16848), .A2(n16517), .ZN(n16463) );
  AOI211_X1 U19825 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n20116), .A(n16464), .B(
        n16463), .ZN(n16465) );
  OAI21_X1 U19826 ( .B1(n16466), .B2(n20138), .A(n16465), .ZN(P2_U2895) );
  NAND2_X1 U19827 ( .A1(n16467), .A2(n20128), .ZN(n16472) );
  INV_X1 U19828 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19829 ( .A1(n20114), .A2(n20284), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n20133), .ZN(n16468) );
  OAI21_X1 U19830 ( .B1(n16513), .B2(n16469), .A(n16468), .ZN(n16470) );
  AOI21_X1 U19831 ( .B1(n20116), .B2(BUF1_REG_23__SCAN_IN), .A(n16470), .ZN(
        n16471) );
  OAI211_X1 U19832 ( .C1(n16853), .C2(n16517), .A(n16472), .B(n16471), .ZN(
        P2_U2896) );
  INV_X1 U19833 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19834 ( .A1(n20114), .A2(n20278), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n20133), .ZN(n16474) );
  NAND2_X1 U19835 ( .A1(n20116), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16473) );
  OAI211_X1 U19836 ( .C1(n16513), .C2(n16475), .A(n16474), .B(n16473), .ZN(
        n16476) );
  AOI21_X1 U19837 ( .B1(n16477), .B2(n20128), .A(n16476), .ZN(n16478) );
  OAI21_X1 U19838 ( .B1(n16870), .B2(n16517), .A(n16478), .ZN(P2_U2897) );
  INV_X1 U19839 ( .A(n16876), .ZN(n16479) );
  NAND2_X1 U19840 ( .A1(n16479), .A2(n20134), .ZN(n16485) );
  INV_X1 U19841 ( .A(n20114), .ZN(n16496) );
  OAI22_X1 U19842 ( .A1(n16496), .A2(n20271), .B1(n16495), .B2(n16480), .ZN(
        n16483) );
  INV_X1 U19843 ( .A(n20116), .ZN(n16481) );
  INV_X1 U19844 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20275) );
  NOR2_X1 U19845 ( .A1(n16481), .A2(n20275), .ZN(n16482) );
  AOI211_X1 U19846 ( .C1(n20115), .C2(BUF2_REG_21__SCAN_IN), .A(n16483), .B(
        n16482), .ZN(n16484) );
  OAI211_X1 U19847 ( .C1(n20138), .C2(n16486), .A(n16485), .B(n16484), .ZN(
        P2_U2898) );
  INV_X1 U19848 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U19849 ( .A1(n20114), .A2(n17210), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n20133), .ZN(n16487) );
  OAI21_X1 U19850 ( .B1(n16513), .B2(n16488), .A(n16487), .ZN(n16491) );
  NOR2_X1 U19851 ( .A1(n16489), .A2(n20138), .ZN(n16490) );
  AOI211_X1 U19852 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n20116), .A(n16491), .B(
        n16490), .ZN(n16492) );
  OAI21_X1 U19853 ( .B1(n16517), .B2(n16493), .A(n16492), .ZN(P2_U2899) );
  NAND2_X1 U19854 ( .A1(n16888), .A2(n20134), .ZN(n16501) );
  OAI22_X1 U19855 ( .A1(n16496), .A2(n20143), .B1(n16495), .B2(n16494), .ZN(
        n16499) );
  INV_X1 U19856 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16497) );
  NOR2_X1 U19857 ( .A1(n16513), .A2(n16497), .ZN(n16498) );
  AOI211_X1 U19858 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n20116), .A(n16499), .B(
        n16498), .ZN(n16500) );
  OAI211_X1 U19859 ( .C1(n20138), .C2(n16502), .A(n16501), .B(n16500), .ZN(
        P2_U2900) );
  INV_X1 U19860 ( .A(n16907), .ZN(n16509) );
  INV_X1 U19861 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16505) );
  AOI22_X1 U19862 ( .A1(n20114), .A2(n17238), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n20133), .ZN(n16504) );
  NAND2_X1 U19863 ( .A1(n20116), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16503) );
  OAI211_X1 U19864 ( .C1(n16513), .C2(n16505), .A(n16504), .B(n16503), .ZN(
        n16506) );
  AOI21_X1 U19865 ( .B1(n16507), .B2(n20128), .A(n16506), .ZN(n16508) );
  OAI21_X1 U19866 ( .B1(n16509), .B2(n16517), .A(n16508), .ZN(P2_U2901) );
  INV_X1 U19867 ( .A(n16920), .ZN(n16518) );
  AOI22_X1 U19868 ( .A1(n20114), .A2(n16510), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n20133), .ZN(n16512) );
  NAND2_X1 U19869 ( .A1(n20116), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16511) );
  OAI211_X1 U19870 ( .C1(n16513), .C2(n17193), .A(n16512), .B(n16511), .ZN(
        n16514) );
  AOI21_X1 U19871 ( .B1(n16515), .B2(n20128), .A(n16514), .ZN(n16516) );
  OAI21_X1 U19872 ( .B1(n16518), .B2(n16517), .A(n16516), .ZN(P2_U2902) );
  AOI21_X1 U19873 ( .B1(n20887), .B2(n20889), .A(n16519), .ZN(n20137) );
  XNOR2_X1 U19874 ( .A(n20876), .B(n20878), .ZN(n20136) );
  NOR2_X1 U19875 ( .A1(n20137), .A2(n20136), .ZN(n20135) );
  NOR2_X1 U19876 ( .A1(n20876), .A2(n20878), .ZN(n16520) );
  OAI21_X1 U19877 ( .B1(n20135), .B2(n16520), .A(n20124), .ZN(n20127) );
  INV_X1 U19878 ( .A(n20126), .ZN(n20109) );
  NAND3_X1 U19879 ( .A1(n20127), .A2(n20109), .A3(n20128), .ZN(n16524) );
  AOI22_X1 U19880 ( .A1(n16522), .A2(n16521), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n20133), .ZN(n16523) );
  OAI211_X1 U19881 ( .C1(n16525), .C2(n17077), .A(n16524), .B(n16523), .ZN(
        P2_U2914) );
  NAND2_X1 U19882 ( .A1(n20204), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16526) );
  OAI211_X1 U19883 ( .C1(n20199), .C2(n16528), .A(n16527), .B(n16526), .ZN(
        n16529) );
  NAND2_X1 U19884 ( .A1(n10218), .A2(n16534), .ZN(n16536) );
  XNOR2_X1 U19885 ( .A(n16536), .B(n16535), .ZN(n16787) );
  AOI21_X1 U19886 ( .B1(n16775), .B2(n13210), .A(n16537), .ZN(n16784) );
  NOR2_X1 U19887 ( .A1(n20207), .A2(n20853), .ZN(n16774) );
  NOR2_X1 U19888 ( .A1(n20199), .A2(n16538), .ZN(n16539) );
  AOI211_X1 U19889 ( .C1(n20204), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16774), .B(n16539), .ZN(n16540) );
  OAI21_X1 U19890 ( .B1(n16781), .B2(n20194), .A(n16540), .ZN(n16541) );
  AOI21_X1 U19891 ( .B1(n20205), .B2(n16784), .A(n16541), .ZN(n16542) );
  OAI21_X1 U19892 ( .B1(n16787), .B2(n20211), .A(n16542), .ZN(P2_U2985) );
  XNOR2_X1 U19893 ( .A(n16545), .B(n16544), .ZN(n16546) );
  NAND2_X1 U19894 ( .A1(n16546), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16801) );
  INV_X1 U19895 ( .A(n16546), .ZN(n16547) );
  NAND3_X1 U19896 ( .A1(n16801), .A2(n16800), .A3(n20196), .ZN(n16552) );
  NOR2_X1 U19897 ( .A1(n20207), .A2(n20851), .ZN(n16802) );
  AOI21_X1 U19898 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16802), .ZN(n16548) );
  OAI21_X1 U19899 ( .B1(n20199), .B2(n16549), .A(n16548), .ZN(n16550) );
  AOI21_X1 U19900 ( .B1(n16808), .B2(n20213), .A(n16550), .ZN(n16551) );
  OAI211_X1 U19901 ( .C1(n16773), .C2(n16809), .A(n16552), .B(n16551), .ZN(
        P2_U2987) );
  NAND2_X1 U19902 ( .A1(n16554), .A2(n16553), .ZN(n16555) );
  XNOR2_X1 U19903 ( .A(n16556), .B(n16555), .ZN(n16840) );
  NAND2_X1 U19904 ( .A1(n20179), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16829) );
  OAI21_X1 U19905 ( .B1(n17654), .B2(n16557), .A(n16829), .ZN(n16559) );
  NOR2_X1 U19906 ( .A1(n16832), .A2(n20194), .ZN(n16558) );
  AOI211_X1 U19907 ( .C1(n20209), .C2(n16560), .A(n16559), .B(n16558), .ZN(
        n16563) );
  INV_X1 U19908 ( .A(n16561), .ZN(n16837) );
  NAND2_X1 U19909 ( .A1(n16571), .A2(n16830), .ZN(n16836) );
  NAND3_X1 U19910 ( .A1(n16837), .A2(n20205), .A3(n16836), .ZN(n16562) );
  OAI211_X1 U19911 ( .C1(n16840), .C2(n20211), .A(n16563), .B(n16562), .ZN(
        P2_U2989) );
  XNOR2_X1 U19912 ( .A(n16564), .B(n16843), .ZN(n16565) );
  XNOR2_X1 U19913 ( .A(n16566), .B(n16565), .ZN(n16850) );
  OR2_X1 U19914 ( .A1(n20207), .A2(n20844), .ZN(n16841) );
  OAI21_X1 U19915 ( .B1(n17654), .B2(n10298), .A(n16841), .ZN(n16567) );
  AOI21_X1 U19916 ( .B1(n20209), .B2(n16568), .A(n16567), .ZN(n16569) );
  OAI21_X1 U19917 ( .B1(n16570), .B2(n20194), .A(n16569), .ZN(n16572) );
  INV_X1 U19918 ( .A(n16573), .ZN(n16574) );
  XNOR2_X1 U19919 ( .A(n16575), .B(n16574), .ZN(n16862) );
  OR2_X1 U19920 ( .A1(n20207), .A2(n20842), .ZN(n16855) );
  OAI21_X1 U19921 ( .B1(n17654), .B2(n16576), .A(n16855), .ZN(n16577) );
  AOI21_X1 U19922 ( .B1(n20209), .B2(n9737), .A(n16577), .ZN(n16578) );
  OAI21_X1 U19923 ( .B1(n16859), .B2(n20194), .A(n16578), .ZN(n16582) );
  INV_X1 U19924 ( .A(n16580), .ZN(n16581) );
  OAI21_X1 U19925 ( .B1(n16602), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n9946), .ZN(n16875) );
  NAND2_X1 U19926 ( .A1(n16586), .A2(n16585), .ZN(n16587) );
  XNOR2_X1 U19927 ( .A(n16588), .B(n16587), .ZN(n16873) );
  NOR2_X1 U19928 ( .A1(n20207), .A2(n16589), .ZN(n16866) );
  AOI21_X1 U19929 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16866), .ZN(n16592) );
  NAND2_X1 U19930 ( .A1(n20209), .A2(n16590), .ZN(n16591) );
  OAI211_X1 U19931 ( .C1(n16869), .C2(n20194), .A(n16592), .B(n16591), .ZN(
        n16593) );
  AOI21_X1 U19932 ( .B1(n20196), .B2(n16873), .A(n16593), .ZN(n16594) );
  OAI21_X1 U19933 ( .B1(n16875), .B2(n16773), .A(n16594), .ZN(P2_U2992) );
  NAND2_X1 U19934 ( .A1(n16596), .A2(n16595), .ZN(n16601) );
  XOR2_X1 U19935 ( .A(n16601), .B(n16600), .Z(n16887) );
  OR2_X1 U19936 ( .A1(n20207), .A2(n20839), .ZN(n16882) );
  OAI21_X1 U19937 ( .B1(n17654), .B2(n16605), .A(n16882), .ZN(n16606) );
  AOI21_X1 U19938 ( .B1(n20209), .B2(n16607), .A(n16606), .ZN(n16608) );
  OAI21_X1 U19939 ( .B1(n16883), .B2(n20194), .A(n16608), .ZN(n16609) );
  AOI21_X1 U19940 ( .B1(n16886), .B2(n20205), .A(n16609), .ZN(n16610) );
  OAI21_X1 U19941 ( .B1(n16887), .B2(n20211), .A(n16610), .ZN(P2_U2993) );
  INV_X1 U19942 ( .A(n16620), .ZN(n16611) );
  NOR2_X1 U19943 ( .A1(n16894), .A2(n20194), .ZN(n16619) );
  NOR2_X1 U19944 ( .A1(n20207), .A2(n20836), .ZN(n16889) );
  AOI21_X1 U19945 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16889), .ZN(n16616) );
  OAI21_X1 U19946 ( .B1(n16617), .B2(n20199), .A(n16616), .ZN(n16618) );
  NAND2_X1 U19947 ( .A1(n16621), .A2(n16620), .ZN(n16623) );
  XOR2_X1 U19948 ( .A(n16623), .B(n16622), .Z(n16908) );
  NOR2_X1 U19949 ( .A1(n20207), .A2(n20834), .ZN(n16902) );
  AOI21_X1 U19950 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16902), .ZN(n16624) );
  OAI21_X1 U19951 ( .B1(n16625), .B2(n20199), .A(n16624), .ZN(n16628) );
  OAI21_X1 U19952 ( .B1(n20211), .B2(n16908), .A(n16630), .ZN(P2_U2996) );
  NAND2_X1 U19953 ( .A1(n16632), .A2(n16631), .ZN(n16633) );
  XNOR2_X1 U19954 ( .A(n9721), .B(n16633), .ZN(n16923) );
  XNOR2_X1 U19955 ( .A(n16913), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16634) );
  NAND2_X1 U19956 ( .A1(n16634), .A2(n20205), .ZN(n16640) );
  NAND2_X1 U19957 ( .A1(n20179), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16916) );
  OAI21_X1 U19958 ( .B1(n17654), .B2(n16635), .A(n16916), .ZN(n16637) );
  NOR2_X1 U19959 ( .A1(n16917), .A2(n20194), .ZN(n16636) );
  AOI211_X1 U19960 ( .C1(n20209), .C2(n16638), .A(n16637), .B(n16636), .ZN(
        n16639) );
  OAI211_X1 U19961 ( .C1(n16923), .C2(n20211), .A(n16640), .B(n16639), .ZN(
        P2_U2997) );
  OAI211_X1 U19962 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16918), .A(
        n16913), .B(n20205), .ZN(n16648) );
  NOR2_X1 U19963 ( .A1(n20207), .A2(n16643), .ZN(n16925) );
  AOI21_X1 U19964 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16925), .ZN(n16644) );
  OAI21_X1 U19965 ( .B1(n16645), .B2(n20199), .A(n16644), .ZN(n16646) );
  AOI21_X1 U19966 ( .B1(n16926), .B2(n20213), .A(n16646), .ZN(n16647) );
  OAI211_X1 U19967 ( .C1(n16924), .C2(n20211), .A(n16648), .B(n16647), .ZN(
        P2_U2998) );
  NAND2_X1 U19968 ( .A1(n16651), .A2(n16650), .ZN(n16652) );
  XNOR2_X1 U19969 ( .A(n16649), .B(n16652), .ZN(n16945) );
  NAND2_X1 U19970 ( .A1(n16933), .A2(n20205), .ZN(n16658) );
  NOR2_X1 U19971 ( .A1(n20207), .A2(n20829), .ZN(n16935) );
  AOI21_X1 U19972 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16935), .ZN(n16653) );
  OAI21_X1 U19973 ( .B1(n20199), .B2(n16654), .A(n16653), .ZN(n16655) );
  AOI21_X1 U19974 ( .B1(n16656), .B2(n20213), .A(n16655), .ZN(n16657) );
  OAI211_X1 U19975 ( .C1(n16945), .C2(n20211), .A(n16658), .B(n16657), .ZN(
        P2_U2999) );
  OAI21_X1 U19976 ( .B1(n9603), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16659), .ZN(n16959) );
  NAND2_X1 U19977 ( .A1(n10035), .A2(n16661), .ZN(n16662) );
  XNOR2_X1 U19978 ( .A(n16663), .B(n16662), .ZN(n16957) );
  NOR2_X1 U19979 ( .A1(n20207), .A2(n20827), .ZN(n16950) );
  NOR2_X1 U19980 ( .A1(n20199), .A2(n16664), .ZN(n16665) );
  AOI211_X1 U19981 ( .C1(n20204), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16950), .B(n16665), .ZN(n16666) );
  OAI21_X1 U19982 ( .B1(n16948), .B2(n20194), .A(n16666), .ZN(n16667) );
  AOI21_X1 U19983 ( .B1(n16957), .B2(n20196), .A(n16667), .ZN(n16668) );
  OAI21_X1 U19984 ( .B1(n16959), .B2(n16773), .A(n16668), .ZN(P2_U3000) );
  NAND2_X1 U19985 ( .A1(n16671), .A2(n16670), .ZN(n16674) );
  NAND2_X1 U19986 ( .A1(n16672), .A2(n16682), .ZN(n16673) );
  XOR2_X1 U19987 ( .A(n16674), .B(n16673), .Z(n16969) );
  NAND2_X1 U19988 ( .A1(n16965), .A2(n20213), .ZN(n16677) );
  NOR2_X1 U19989 ( .A1(n20207), .A2(n16675), .ZN(n16964) );
  AOI21_X1 U19990 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16964), .ZN(n16676) );
  OAI211_X1 U19991 ( .C1(n20199), .C2(n16678), .A(n16677), .B(n16676), .ZN(
        n16679) );
  AOI21_X1 U19992 ( .B1(n16969), .B2(n20196), .A(n16679), .ZN(n16680) );
  OAI21_X1 U19993 ( .B1(n16971), .B2(n16773), .A(n16680), .ZN(P2_U3001) );
  NAND2_X1 U19994 ( .A1(n16682), .A2(n16681), .ZN(n16684) );
  XOR2_X1 U19995 ( .A(n16684), .B(n16683), .Z(n16984) );
  NAND2_X1 U19996 ( .A1(n16728), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16727) );
  INV_X1 U19997 ( .A(n16669), .ZN(n16972) );
  NAND3_X1 U19998 ( .A1(n16973), .A2(n20205), .A3(n16972), .ZN(n16690) );
  NOR2_X1 U19999 ( .A1(n20207), .A2(n16685), .ZN(n16974) );
  AOI21_X1 U20000 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16974), .ZN(n16686) );
  OAI21_X1 U20001 ( .B1(n20199), .B2(n16687), .A(n16686), .ZN(n16688) );
  AOI21_X1 U20002 ( .B1(n20095), .B2(n20213), .A(n16688), .ZN(n16689) );
  OAI211_X1 U20003 ( .C1(n16984), .C2(n20211), .A(n16690), .B(n16689), .ZN(
        P2_U3002) );
  OAI21_X1 U20004 ( .B1(n16719), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16691), .ZN(n16996) );
  XNOR2_X1 U20005 ( .A(n16693), .B(n16692), .ZN(n16768) );
  INV_X1 U20006 ( .A(n16767), .ZN(n16696) );
  INV_X1 U20007 ( .A(n16694), .ZN(n16695) );
  INV_X1 U20008 ( .A(n16697), .ZN(n16698) );
  NAND2_X1 U20009 ( .A1(n16732), .A2(n16730), .ZN(n16716) );
  INV_X1 U20010 ( .A(n16715), .ZN(n16701) );
  OAI21_X1 U20011 ( .B1(n16716), .B2(n16701), .A(n16700), .ZN(n16705) );
  NAND2_X1 U20012 ( .A1(n16703), .A2(n16702), .ZN(n16704) );
  XNOR2_X1 U20013 ( .A(n16705), .B(n16704), .ZN(n16993) );
  NOR2_X1 U20014 ( .A1(n20207), .A2(n16706), .ZN(n16986) );
  NOR2_X1 U20015 ( .A1(n17654), .A2(n16707), .ZN(n16708) );
  AOI211_X1 U20016 ( .C1(n16709), .C2(n20209), .A(n16986), .B(n16708), .ZN(
        n16710) );
  OAI21_X1 U20017 ( .B1(n16711), .B2(n20194), .A(n16710), .ZN(n16712) );
  AOI21_X1 U20018 ( .B1(n16993), .B2(n20196), .A(n16712), .ZN(n16713) );
  OAI21_X1 U20019 ( .B1(n16996), .B2(n16773), .A(n16713), .ZN(P2_U3003) );
  NAND2_X1 U20020 ( .A1(n16715), .A2(n16714), .ZN(n16718) );
  NAND2_X1 U20021 ( .A1(n16716), .A2(n16729), .ZN(n16717) );
  XOR2_X1 U20022 ( .A(n16718), .B(n16717), .Z(n17009) );
  AOI21_X1 U20023 ( .B1(n16720), .B2(n16727), .A(n16719), .ZN(n17007) );
  NAND2_X1 U20024 ( .A1(n20105), .A2(n20213), .ZN(n16723) );
  NOR2_X1 U20025 ( .A1(n20207), .A2(n16721), .ZN(n16997) );
  AOI21_X1 U20026 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16997), .ZN(n16722) );
  OAI211_X1 U20027 ( .C1(n20199), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        n16725) );
  AOI21_X1 U20028 ( .B1(n17007), .B2(n20205), .A(n16725), .ZN(n16726) );
  OAI21_X1 U20029 ( .B1(n17009), .B2(n20211), .A(n16726), .ZN(P2_U3004) );
  OAI21_X1 U20030 ( .B1(n16728), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16727), .ZN(n17022) );
  NAND2_X1 U20031 ( .A1(n16730), .A2(n16729), .ZN(n16731) );
  XNOR2_X1 U20032 ( .A(n16732), .B(n16731), .ZN(n17019) );
  NOR2_X1 U20033 ( .A1(n20207), .A2(n20821), .ZN(n17010) );
  NOR2_X1 U20034 ( .A1(n17654), .A2(n16733), .ZN(n16734) );
  AOI211_X1 U20035 ( .C1(n16735), .C2(n20209), .A(n17010), .B(n16734), .ZN(
        n16736) );
  OAI21_X1 U20036 ( .B1(n17012), .B2(n20194), .A(n16736), .ZN(n16737) );
  AOI21_X1 U20037 ( .B1(n17019), .B2(n20196), .A(n16737), .ZN(n16738) );
  OAI21_X1 U20038 ( .B1(n17022), .B2(n16773), .A(n16738), .ZN(P2_U3005) );
  NAND2_X1 U20039 ( .A1(n16740), .A2(n16739), .ZN(n16743) );
  INV_X1 U20040 ( .A(n16756), .ZN(n16741) );
  OAI21_X1 U20041 ( .B1(n16758), .B2(n16741), .A(n16757), .ZN(n16742) );
  XOR2_X1 U20042 ( .A(n16743), .B(n16742), .Z(n17036) );
  OR2_X1 U20043 ( .A1(n20207), .A2(n20819), .ZN(n17028) );
  NAND2_X1 U20044 ( .A1(n20204), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16744) );
  OAI211_X1 U20045 ( .C1(n20199), .C2(n16745), .A(n17028), .B(n16744), .ZN(
        n16746) );
  AOI21_X1 U20046 ( .B1(n16747), .B2(n20213), .A(n16746), .ZN(n16752) );
  NAND2_X1 U20047 ( .A1(n16750), .A2(n16749), .ZN(n17032) );
  NAND3_X1 U20048 ( .A1(n17033), .A2(n17032), .A3(n20205), .ZN(n16751) );
  OAI211_X1 U20049 ( .C1(n17036), .C2(n20211), .A(n16752), .B(n16751), .ZN(
        P2_U3006) );
  XNOR2_X1 U20050 ( .A(n16754), .B(n17040), .ZN(n16755) );
  XNOR2_X1 U20051 ( .A(n16753), .B(n16755), .ZN(n17048) );
  NAND2_X1 U20052 ( .A1(n16757), .A2(n16756), .ZN(n16759) );
  XOR2_X1 U20053 ( .A(n16759), .B(n16758), .Z(n17037) );
  OAI22_X1 U20054 ( .A1(n17654), .A2(n16760), .B1(n20817), .B2(n20207), .ZN(
        n16761) );
  AOI21_X1 U20055 ( .B1(n20209), .B2(n16762), .A(n16761), .ZN(n16763) );
  OAI21_X1 U20056 ( .B1(n16764), .B2(n20194), .A(n16763), .ZN(n16765) );
  AOI21_X1 U20057 ( .B1(n17037), .B2(n20196), .A(n16765), .ZN(n16766) );
  OAI21_X1 U20058 ( .B1(n16773), .B2(n17048), .A(n16766), .ZN(P2_U3007) );
  XNOR2_X1 U20059 ( .A(n16768), .B(n16767), .ZN(n17057) );
  OAI22_X1 U20060 ( .A1(n20815), .A2(n20207), .B1(n20199), .B2(n20081), .ZN(
        n16769) );
  AOI21_X1 U20061 ( .B1(n20204), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16769), .ZN(n16770) );
  OAI21_X1 U20062 ( .B1(n20088), .B2(n20194), .A(n16770), .ZN(n16771) );
  AOI21_X1 U20063 ( .B1(n17057), .B2(n20196), .A(n16771), .ZN(n16772) );
  OAI21_X1 U20064 ( .B1(n17059), .B2(n16773), .A(n16772), .ZN(P2_U3008) );
  AOI21_X1 U20065 ( .B1(n16776), .B2(n16775), .A(n16774), .ZN(n16780) );
  INV_X1 U20066 ( .A(n16789), .ZN(n16777) );
  NAND2_X1 U20067 ( .A1(n16777), .A2(n16805), .ZN(n16803) );
  NAND2_X1 U20068 ( .A1(n16806), .A2(n16803), .ZN(n16792) );
  NOR2_X1 U20069 ( .A1(n16789), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16778) );
  OAI21_X1 U20070 ( .B1(n16792), .B2(n16778), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16779) );
  OAI211_X1 U20071 ( .C1(n16781), .C2(n20242), .A(n16780), .B(n16779), .ZN(
        n16782) );
  AOI21_X1 U20072 ( .B1(n20238), .B2(n16783), .A(n16782), .ZN(n16786) );
  NAND2_X1 U20073 ( .A1(n16784), .A2(n12495), .ZN(n16785) );
  OAI211_X1 U20074 ( .C1(n16787), .C2(n20241), .A(n16786), .B(n16785), .ZN(
        P2_U3017) );
  NAND2_X1 U20075 ( .A1(n16788), .A2(n17661), .ZN(n16798) );
  NOR3_X1 U20076 ( .A1(n16789), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16805), .ZN(n16790) );
  AOI211_X1 U20077 ( .C1(n16792), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16791), .B(n16790), .ZN(n16793) );
  OAI21_X1 U20078 ( .B1(n16794), .B2(n20242), .A(n16793), .ZN(n16795) );
  AOI21_X1 U20079 ( .B1(n20238), .B2(n16796), .A(n16795), .ZN(n16797) );
  NAND3_X1 U20080 ( .A1(n16801), .A2(n16800), .A3(n17661), .ZN(n16813) );
  INV_X1 U20081 ( .A(n16802), .ZN(n16804) );
  OAI211_X1 U20082 ( .C1(n16806), .C2(n16805), .A(n16804), .B(n16803), .ZN(
        n16807) );
  AOI21_X1 U20083 ( .B1(n16808), .B2(n17090), .A(n16807), .ZN(n16812) );
  OR2_X1 U20084 ( .A1(n16810), .A2(n20227), .ZN(n16811) );
  INV_X1 U20085 ( .A(n16814), .ZN(n16827) );
  OAI211_X1 U20086 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16827), .B(n16815), .ZN(
        n16816) );
  OAI211_X1 U20087 ( .C1(n16831), .C2(n16818), .A(n16817), .B(n16816), .ZN(
        n16821) );
  NOR2_X1 U20088 ( .A1(n16819), .A2(n20242), .ZN(n16820) );
  AOI211_X1 U20089 ( .C1(n16822), .C2(n20238), .A(n16821), .B(n16820), .ZN(
        n16825) );
  OAI211_X1 U20090 ( .C1(n16826), .C2(n20241), .A(n16825), .B(n16824), .ZN(
        P2_U3020) );
  NAND2_X1 U20091 ( .A1(n16827), .A2(n16830), .ZN(n16828) );
  OAI211_X1 U20092 ( .C1(n16831), .C2(n16830), .A(n16829), .B(n16828), .ZN(
        n16834) );
  NOR2_X1 U20093 ( .A1(n16832), .A2(n20242), .ZN(n16833) );
  AOI211_X1 U20094 ( .C1(n16835), .C2(n20238), .A(n16834), .B(n16833), .ZN(
        n16839) );
  NAND3_X1 U20095 ( .A1(n16837), .A2(n12495), .A3(n16836), .ZN(n16838) );
  OAI211_X1 U20096 ( .C1(n16840), .C2(n20241), .A(n16839), .B(n16838), .ZN(
        P2_U3021) );
  OAI211_X1 U20097 ( .C1(n16844), .C2(n16843), .A(n16842), .B(n16841), .ZN(
        n16845) );
  AOI21_X1 U20098 ( .B1(n16846), .B2(n17090), .A(n16845), .ZN(n16847) );
  OAI21_X1 U20099 ( .B1(n20227), .B2(n16848), .A(n16847), .ZN(n16849) );
  AOI21_X1 U20100 ( .B1(n17661), .B2(n16850), .A(n16849), .ZN(n16851) );
  OAI21_X1 U20101 ( .B1(n20219), .B2(n16852), .A(n16851), .ZN(P2_U3022) );
  NOR2_X1 U20102 ( .A1(n16853), .A2(n20227), .ZN(n16861) );
  OAI211_X1 U20103 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16865), .B(n16854), .ZN(
        n16856) );
  NAND2_X1 U20104 ( .A1(n16856), .A2(n16855), .ZN(n16857) );
  AOI21_X1 U20105 ( .B1(n16878), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16857), .ZN(n16858) );
  OAI21_X1 U20106 ( .B1(n16859), .B2(n20242), .A(n16858), .ZN(n16860) );
  AOI211_X1 U20107 ( .C1(n17661), .C2(n16862), .A(n16861), .B(n16860), .ZN(
        n16863) );
  OAI21_X1 U20108 ( .B1(n20219), .B2(n16864), .A(n16863), .ZN(P2_U3023) );
  MUX2_X1 U20109 ( .A(n16865), .B(n16878), .S(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n16867) );
  NOR2_X1 U20110 ( .A1(n16867), .A2(n16866), .ZN(n16868) );
  OAI21_X1 U20111 ( .B1(n16869), .B2(n20242), .A(n16868), .ZN(n16872) );
  NOR2_X1 U20112 ( .A1(n16870), .A2(n20227), .ZN(n16871) );
  AOI211_X1 U20113 ( .C1(n17661), .C2(n16873), .A(n16872), .B(n16871), .ZN(
        n16874) );
  OAI21_X1 U20114 ( .B1(n16875), .B2(n20219), .A(n16874), .ZN(P2_U3024) );
  NOR2_X1 U20115 ( .A1(n16876), .A2(n20227), .ZN(n16885) );
  NAND2_X1 U20116 ( .A1(n16877), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16880) );
  INV_X1 U20117 ( .A(n16878), .ZN(n16879) );
  MUX2_X1 U20118 ( .A(n16880), .B(n16879), .S(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(n16881) );
  OAI211_X1 U20119 ( .C1(n16883), .C2(n20242), .A(n16882), .B(n16881), .ZN(
        n16884) );
  NAND2_X1 U20120 ( .A1(n16888), .A2(n20238), .ZN(n16893) );
  OR2_X1 U20121 ( .A1(n16890), .A2(n16889), .ZN(n16891) );
  AOI21_X1 U20122 ( .B1(n16903), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16891), .ZN(n16892) );
  OAI211_X1 U20123 ( .C1(n16894), .C2(n20242), .A(n16893), .B(n16892), .ZN(
        n16895) );
  AOI21_X1 U20124 ( .B1(n16896), .B2(n12495), .A(n16895), .ZN(n16897) );
  OAI21_X1 U20125 ( .B1(n20241), .B2(n16898), .A(n16897), .ZN(P2_U3027) );
  INV_X1 U20126 ( .A(n16937), .ZN(n16900) );
  NAND3_X1 U20127 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16899) );
  NOR3_X1 U20128 ( .A1(n16900), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16899), .ZN(n16901) );
  AOI211_X1 U20129 ( .C1(n16903), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16902), .B(n16901), .ZN(n16904) );
  OAI21_X1 U20130 ( .B1(n16905), .B2(n20242), .A(n16904), .ZN(n16906) );
  NAND2_X1 U20131 ( .A1(n20219), .A2(n20217), .ZN(n16912) );
  INV_X1 U20132 ( .A(n16909), .ZN(n16910) );
  AOI21_X2 U20133 ( .B1(n16913), .B2(n16912), .A(n10459), .ZN(n16932) );
  OAI21_X1 U20134 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16914), .A(
        n16932), .ZN(n16915) );
  NAND2_X1 U20135 ( .A1(n16915), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16922) );
  OAI21_X1 U20136 ( .B1(n16917), .B2(n20242), .A(n16916), .ZN(n16919) );
  OAI211_X1 U20137 ( .C1(n16923), .C2(n20241), .A(n16922), .B(n16921), .ZN(
        P2_U3029) );
  INV_X1 U20138 ( .A(n16924), .ZN(n16930) );
  AOI21_X1 U20139 ( .B1(n16926), .B2(n17090), .A(n16925), .ZN(n16927) );
  OAI21_X1 U20140 ( .B1(n20227), .B2(n20117), .A(n16927), .ZN(n16929) );
  OAI21_X1 U20141 ( .B1(n16932), .B2(n10406), .A(n16931), .ZN(P2_U3030) );
  NAND2_X1 U20142 ( .A1(n16933), .A2(n12495), .ZN(n16944) );
  NOR2_X1 U20143 ( .A1(n16934), .A2(n20227), .ZN(n16941) );
  AOI21_X1 U20144 ( .B1(n16937), .B2(n16936), .A(n16935), .ZN(n16938) );
  OAI21_X1 U20145 ( .B1(n16939), .B2(n20242), .A(n16938), .ZN(n16940) );
  AOI211_X1 U20146 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16942), .A(
        n16941), .B(n16940), .ZN(n16943) );
  OAI211_X1 U20147 ( .C1(n16945), .C2(n20241), .A(n16944), .B(n16943), .ZN(
        P2_U3031) );
  INV_X1 U20148 ( .A(n16979), .ZN(n16946) );
  AOI21_X1 U20149 ( .B1(n16975), .B2(n16947), .A(n16946), .ZN(n16960) );
  NOR2_X1 U20150 ( .A1(n16948), .A2(n20242), .ZN(n16949) );
  AOI211_X1 U20151 ( .C1(n16951), .C2(n16955), .A(n16950), .B(n16949), .ZN(
        n16954) );
  NAND2_X1 U20152 ( .A1(n16952), .A2(n20238), .ZN(n16953) );
  OAI211_X1 U20153 ( .C1(n16960), .C2(n16955), .A(n16954), .B(n16953), .ZN(
        n16956) );
  AOI21_X1 U20154 ( .B1(n16957), .B2(n17661), .A(n16956), .ZN(n16958) );
  OAI21_X1 U20155 ( .B1(n16959), .B2(n20219), .A(n16958), .ZN(P2_U3032) );
  AOI21_X1 U20156 ( .B1(n16962), .B2(n16961), .A(n16960), .ZN(n16963) );
  AOI211_X1 U20157 ( .C1(n17090), .C2(n16965), .A(n16964), .B(n16963), .ZN(
        n16966) );
  OAI21_X1 U20158 ( .B1(n20227), .B2(n16967), .A(n16966), .ZN(n16968) );
  AOI21_X1 U20159 ( .B1(n16969), .B2(n17661), .A(n16968), .ZN(n16970) );
  OAI21_X1 U20160 ( .B1(n16971), .B2(n20219), .A(n16970), .ZN(P2_U3033) );
  NAND2_X1 U20161 ( .A1(n20095), .A2(n17090), .ZN(n16977) );
  AOI21_X1 U20162 ( .B1(n16975), .B2(n16978), .A(n16974), .ZN(n16976) );
  OAI211_X1 U20163 ( .C1(n16979), .C2(n16978), .A(n16977), .B(n16976), .ZN(
        n16980) );
  AOI21_X1 U20164 ( .B1(n20238), .B2(n16981), .A(n16980), .ZN(n16982) );
  OAI211_X1 U20165 ( .C1(n16984), .C2(n20241), .A(n16983), .B(n16982), .ZN(
        P2_U3034) );
  OAI21_X1 U20166 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16985), .ZN(n16990) );
  AOI21_X1 U20167 ( .B1(n16987), .B2(n17090), .A(n16986), .ZN(n16989) );
  INV_X1 U20168 ( .A(n17015), .ZN(n17000) );
  NAND3_X1 U20169 ( .A1(n17000), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16999), .ZN(n16988) );
  OAI211_X1 U20170 ( .C1(n17001), .C2(n16990), .A(n16989), .B(n16988), .ZN(
        n16991) );
  AOI21_X1 U20171 ( .B1(n20238), .B2(n16992), .A(n16991), .ZN(n16995) );
  NAND2_X1 U20172 ( .A1(n16993), .A2(n17661), .ZN(n16994) );
  OAI211_X1 U20173 ( .C1(n16996), .C2(n20219), .A(n16995), .B(n16994), .ZN(
        P2_U3035) );
  AOI21_X1 U20174 ( .B1(n20105), .B2(n17090), .A(n16997), .ZN(n17005) );
  NAND2_X1 U20175 ( .A1(n16998), .A2(n20238), .ZN(n17004) );
  NAND3_X1 U20176 ( .A1(n17000), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16999), .ZN(n17003) );
  OR2_X1 U20177 ( .A1(n17001), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17002) );
  NAND4_X1 U20178 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17002), .ZN(
        n17006) );
  AOI21_X1 U20179 ( .B1(n17007), .B2(n12495), .A(n17006), .ZN(n17008) );
  OAI21_X1 U20180 ( .B1(n17009), .B2(n20241), .A(n17008), .ZN(P2_U3036) );
  INV_X1 U20181 ( .A(n17010), .ZN(n17011) );
  OAI21_X1 U20182 ( .B1(n17012), .B2(n20242), .A(n17011), .ZN(n17017) );
  AOI21_X1 U20183 ( .B1(n17041), .B2(n17013), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17014) );
  NOR2_X1 U20184 ( .A1(n17015), .A2(n17014), .ZN(n17016) );
  AOI211_X1 U20185 ( .C1(n20238), .C2(n17018), .A(n17017), .B(n17016), .ZN(
        n17021) );
  NAND2_X1 U20186 ( .A1(n17019), .A2(n17661), .ZN(n17020) );
  OAI211_X1 U20187 ( .C1(n17022), .C2(n20219), .A(n17021), .B(n17020), .ZN(
        P2_U3037) );
  NOR2_X1 U20188 ( .A1(n17023), .A2(n20227), .ZN(n17031) );
  NAND2_X1 U20189 ( .A1(n17024), .A2(n17040), .ZN(n17025) );
  NAND3_X1 U20190 ( .A1(n17041), .A2(n17026), .A3(n17025), .ZN(n17027) );
  OAI211_X1 U20191 ( .C1(n17029), .C2(n20242), .A(n17028), .B(n17027), .ZN(
        n17030) );
  AOI211_X1 U20192 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n17049), .A(
        n17031), .B(n17030), .ZN(n17035) );
  NAND3_X1 U20193 ( .A1(n17033), .A2(n17032), .A3(n12495), .ZN(n17034) );
  OAI211_X1 U20194 ( .C1(n17036), .C2(n20241), .A(n17035), .B(n17034), .ZN(
        P2_U3038) );
  NAND2_X1 U20195 ( .A1(n17037), .A2(n17661), .ZN(n17047) );
  NOR2_X1 U20196 ( .A1(n20817), .A2(n20207), .ZN(n17038) );
  AOI21_X1 U20197 ( .B1(n17039), .B2(n17090), .A(n17038), .ZN(n17043) );
  NAND2_X1 U20198 ( .A1(n17041), .A2(n17040), .ZN(n17042) );
  OAI211_X1 U20199 ( .C1(n20227), .C2(n17044), .A(n17043), .B(n17042), .ZN(
        n17045) );
  AOI21_X1 U20200 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17049), .A(
        n17045), .ZN(n17046) );
  OAI211_X1 U20201 ( .C1(n17048), .C2(n20219), .A(n17047), .B(n17046), .ZN(
        P2_U3039) );
  NAND2_X1 U20202 ( .A1(n17049), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17055) );
  INV_X1 U20203 ( .A(n20088), .ZN(n17053) );
  NOR2_X1 U20204 ( .A1(n20815), .A2(n20207), .ZN(n17052) );
  INV_X1 U20205 ( .A(n17070), .ZN(n17050) );
  NOR3_X1 U20206 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17050), .A3(
        n17086), .ZN(n17051) );
  AOI211_X1 U20207 ( .C1(n17053), .C2(n17090), .A(n17052), .B(n17051), .ZN(
        n17054) );
  OAI211_X1 U20208 ( .C1(n20227), .C2(n20078), .A(n17055), .B(n17054), .ZN(
        n17056) );
  AOI21_X1 U20209 ( .B1(n17057), .B2(n17661), .A(n17056), .ZN(n17058) );
  OAI21_X1 U20210 ( .B1(n17059), .B2(n20219), .A(n17058), .ZN(P2_U3040) );
  XNOR2_X1 U20211 ( .A(n17061), .B(n10478), .ZN(n17085) );
  OAI22_X1 U20212 ( .A1(n17085), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n10478), .B2(n17061), .ZN(n17066) );
  NAND2_X1 U20213 ( .A1(n17064), .A2(n17062), .ZN(n17065) );
  AOI22_X1 U20214 ( .A1(n17066), .A2(n17065), .B1(n10880), .B2(n17064), .ZN(
        n17639) );
  INV_X1 U20215 ( .A(n17639), .ZN(n17080) );
  XNOR2_X1 U20216 ( .A(n17067), .B(n17072), .ZN(n17068) );
  XNOR2_X1 U20217 ( .A(n17069), .B(n17068), .ZN(n17641) );
  NOR2_X1 U20218 ( .A1(n11346), .A2(n20207), .ZN(n17074) );
  AOI211_X1 U20219 ( .C1(n17072), .C2(n17071), .A(n17070), .B(n17086), .ZN(
        n17073) );
  AOI211_X1 U20220 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n17087), .A(
        n17074), .B(n17073), .ZN(n17076) );
  NAND2_X1 U20221 ( .A1(n17640), .A2(n17090), .ZN(n17075) );
  OAI211_X1 U20222 ( .C1(n20227), .C2(n17077), .A(n17076), .B(n17075), .ZN(
        n17078) );
  AOI21_X1 U20223 ( .B1(n17661), .B2(n17641), .A(n17078), .ZN(n17079) );
  OAI21_X1 U20224 ( .B1(n17080), .B2(n20219), .A(n17079), .ZN(P2_U3041) );
  XNOR2_X1 U20225 ( .A(n17081), .B(n17099), .ZN(n17096) );
  AOI22_X1 U20226 ( .A1(n17096), .A2(n17097), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17081), .ZN(n17084) );
  XNOR2_X1 U20227 ( .A(n17082), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17083) );
  XNOR2_X1 U20228 ( .A(n17084), .B(n17083), .ZN(n20182) );
  INV_X1 U20229 ( .A(n20182), .ZN(n17095) );
  XNOR2_X1 U20230 ( .A(n17085), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20180) );
  INV_X1 U20231 ( .A(n17086), .ZN(n17088) );
  MUX2_X1 U20232 ( .A(n17088), .B(n17087), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n17093) );
  NOR2_X1 U20233 ( .A1(n20207), .A2(n11104), .ZN(n17089) );
  AOI21_X1 U20234 ( .B1(n20181), .B2(n17090), .A(n17089), .ZN(n17091) );
  OAI21_X1 U20235 ( .B1(n20124), .B2(n20227), .A(n17091), .ZN(n17092) );
  AOI211_X1 U20236 ( .C1(n20180), .C2(n12495), .A(n17093), .B(n17092), .ZN(
        n17094) );
  OAI21_X1 U20237 ( .B1(n17095), .B2(n20241), .A(n17094), .ZN(P2_U3042) );
  XOR2_X1 U20238 ( .A(n17097), .B(n17096), .Z(n17651) );
  INV_X1 U20239 ( .A(n17651), .ZN(n17108) );
  OAI22_X1 U20240 ( .A1(n20242), .A2(n17649), .B1(n20811), .B2(n20207), .ZN(
        n17103) );
  INV_X1 U20241 ( .A(n17098), .ZN(n17101) );
  MUX2_X1 U20242 ( .A(n17101), .B(n17100), .S(n17099), .Z(n17102) );
  AOI211_X1 U20243 ( .C1(n20238), .C2(n20878), .A(n17103), .B(n17102), .ZN(
        n17107) );
  OR2_X1 U20244 ( .A1(n17105), .A2(n17104), .ZN(n17647) );
  NAND3_X1 U20245 ( .A1(n17647), .A2(n17646), .A3(n12495), .ZN(n17106) );
  OAI211_X1 U20246 ( .C1(n17108), .C2(n20241), .A(n17107), .B(n17106), .ZN(
        P2_U3043) );
  INV_X1 U20247 ( .A(n17109), .ZN(n17121) );
  INV_X1 U20248 ( .A(n17115), .ZN(n17110) );
  AOI22_X1 U20249 ( .A1(n17111), .A2(n17110), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20679), .ZN(n17112) );
  OAI21_X1 U20250 ( .B1(n17220), .B2(n17121), .A(n17112), .ZN(n17119) );
  NAND2_X1 U20251 ( .A1(n20912), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17113) );
  INV_X1 U20252 ( .A(n17675), .ZN(n17295) );
  AOI21_X1 U20253 ( .B1(n20898), .B2(n13618), .A(n17295), .ZN(n17118) );
  OR2_X1 U20254 ( .A1(n20731), .A2(n17118), .ZN(n20892) );
  MUX2_X1 U20255 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n17119), .S(
        n20892), .Z(P2_U3605) );
  NOR3_X1 U20256 ( .A1(n20251), .A2(n17121), .A3(n17120), .ZN(n17122) );
  AOI21_X1 U20257 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20237), .A(n17122), 
        .ZN(n17123) );
  OAI21_X1 U20258 ( .B1(n20871), .B2(n20868), .A(n17123), .ZN(n17124) );
  MUX2_X1 U20259 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n17124), .S(
        n20892), .Z(P2_U3604) );
  MUX2_X1 U20260 ( .A(n17126), .B(n17125), .S(n20080), .Z(n17145) );
  INV_X1 U20261 ( .A(n13663), .ZN(n17133) );
  OR2_X1 U20262 ( .A1(n13245), .A2(n17127), .ZN(n17132) );
  INV_X1 U20263 ( .A(n11213), .ZN(n17128) );
  NAND2_X1 U20264 ( .A1(n17129), .A2(n17128), .ZN(n17136) );
  MUX2_X1 U20265 ( .A(n17136), .B(n17161), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n17130) );
  INV_X1 U20266 ( .A(n17130), .ZN(n17131) );
  NAND2_X1 U20267 ( .A1(n17132), .A2(n17131), .ZN(n17250) );
  AOI222_X1 U20268 ( .A1(n17145), .A2(P2_STATE2_REG_1__SCAN_IN), .B1(n17133), 
        .B2(n17668), .C1(n17250), .C2(n17288), .ZN(n17135) );
  INV_X1 U20269 ( .A(n17149), .ZN(n17172) );
  NAND2_X1 U20270 ( .A1(n17172), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17134) );
  OAI21_X1 U20271 ( .B1(n17135), .B2(n17172), .A(n17134), .ZN(P2_U3601) );
  INV_X1 U20272 ( .A(n17668), .ZN(n17148) );
  NAND2_X1 U20273 ( .A1(n20214), .A2(n17167), .ZN(n17142) );
  OAI21_X1 U20274 ( .B1(n10709), .B2(n17137), .A(n17136), .ZN(n17140) );
  NAND2_X1 U20275 ( .A1(n17161), .A2(n17138), .ZN(n17139) );
  AND2_X1 U20276 ( .A1(n17140), .A2(n17139), .ZN(n17141) );
  NAND2_X1 U20277 ( .A1(n17142), .A2(n17141), .ZN(n17255) );
  NAND2_X1 U20278 ( .A1(n20080), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17143) );
  NAND2_X1 U20279 ( .A1(n17144), .A2(n17143), .ZN(n17151) );
  INV_X1 U20280 ( .A(n17151), .ZN(n17146) );
  NOR2_X1 U20281 ( .A1(n17145), .A2(n17290), .ZN(n17152) );
  AOI22_X1 U20282 ( .A1(n17255), .A2(n17288), .B1(n17146), .B2(n17152), .ZN(
        n17147) );
  OAI21_X1 U20283 ( .B1(n20251), .B2(n17148), .A(n17147), .ZN(n17150) );
  MUX2_X1 U20284 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17150), .S(
        n17149), .Z(P2_U3600) );
  INV_X1 U20285 ( .A(n20889), .ZN(n17153) );
  AOI22_X1 U20286 ( .A1(n17153), .A2(n17668), .B1(n17152), .B2(n17151), .ZN(
        n17173) );
  NOR2_X1 U20287 ( .A1(n17155), .A2(n17154), .ZN(n17157) );
  NAND2_X1 U20288 ( .A1(n17156), .A2(n17157), .ZN(n17165) );
  INV_X1 U20289 ( .A(n17157), .ZN(n17162) );
  INV_X1 U20290 ( .A(n17158), .ZN(n17159) );
  OAI21_X1 U20291 ( .B1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n17248), .A(
        n17159), .ZN(n17160) );
  AOI22_X1 U20292 ( .A1(n17163), .A2(n17162), .B1(n17161), .B2(n17160), .ZN(
        n17164) );
  NAND2_X1 U20293 ( .A1(n17165), .A2(n17164), .ZN(n17166) );
  AOI21_X1 U20294 ( .B1(n17168), .B2(n17167), .A(n17166), .ZN(n17247) );
  INV_X1 U20295 ( .A(n17247), .ZN(n17170) );
  AOI22_X1 U20296 ( .A1(n17170), .A2(n17169), .B1(n17172), .B2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20297 ( .B1(n17173), .B2(n17172), .A(n17171), .ZN(P2_U3599) );
  INV_X1 U20298 ( .A(n20534), .ZN(n20529) );
  NAND2_X1 U20299 ( .A1(n20464), .A2(n20529), .ZN(n17174) );
  NOR2_X1 U20300 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20349) );
  INV_X1 U20301 ( .A(n20349), .ZN(n20322) );
  NOR2_X1 U20302 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20322), .ZN(
        n20253) );
  INV_X1 U20303 ( .A(n20253), .ZN(n17182) );
  NAND2_X1 U20304 ( .A1(n17174), .A2(n17182), .ZN(n17179) );
  OR2_X1 U20305 ( .A1(n20525), .A2(n20322), .ZN(n17195) );
  INV_X1 U20306 ( .A(n17195), .ZN(n20308) );
  NAND2_X1 U20307 ( .A1(n17195), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17175) );
  OR2_X1 U20308 ( .A1(n17176), .A2(n17175), .ZN(n17180) );
  OAI211_X1 U20309 ( .C1(n20308), .C2(n11308), .A(n17180), .B(n20731), .ZN(
        n17177) );
  INV_X1 U20310 ( .A(n17177), .ZN(n17178) );
  INV_X1 U20311 ( .A(n17180), .ZN(n17181) );
  AOI211_X2 U20312 ( .C1(n20559), .C2(n17182), .A(n20463), .B(n17181), .ZN(
        n20309) );
  NAND2_X1 U20313 ( .A1(n20113), .A2(n20731), .ZN(n20691) );
  AND2_X1 U20314 ( .A1(n17183), .A2(n20287), .ZN(n20729) );
  INV_X1 U20315 ( .A(n20729), .ZN(n20631) );
  INV_X1 U20316 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17733) );
  INV_X1 U20317 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19421) );
  OAI22_X2 U20318 ( .A1(n17733), .A2(n20290), .B1(n19421), .B2(n20289), .ZN(
        n20683) );
  INV_X1 U20319 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17720) );
  OAI22_X2 U20320 ( .A1(n16462), .A2(n20289), .B1(n17720), .B2(n20290), .ZN(
        n20738) );
  AOI22_X1 U20321 ( .A1(n20342), .A2(n20683), .B1(n20310), .B2(n20738), .ZN(
        n17188) );
  OAI21_X1 U20322 ( .B1(n20631), .B2(n17195), .A(n17188), .ZN(n17189) );
  AOI21_X1 U20323 ( .B1(n20309), .B2(n20730), .A(n17189), .ZN(n17190) );
  OAI21_X1 U20324 ( .B1(n20307), .B2(n17191), .A(n17190), .ZN(P2_U3056) );
  INV_X1 U20325 ( .A(n20742), .ZN(n20642) );
  INV_X1 U20326 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n17731) );
  INV_X1 U20327 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n17193) );
  OAI22_X2 U20328 ( .A1(n17731), .A2(n20290), .B1(n17193), .B2(n20289), .ZN(
        n20692) );
  INV_X1 U20329 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17718) );
  INV_X1 U20330 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19429) );
  OAI22_X2 U20331 ( .A1(n17718), .A2(n20290), .B1(n19429), .B2(n20289), .ZN(
        n20744) );
  AOI22_X1 U20332 ( .A1(n20342), .A2(n20692), .B1(n20310), .B2(n20744), .ZN(
        n17194) );
  OAI21_X1 U20333 ( .B1(n20642), .B2(n17195), .A(n17194), .ZN(n17196) );
  AOI21_X1 U20334 ( .B1(n20309), .B2(n20743), .A(n17196), .ZN(n17197) );
  OAI21_X1 U20335 ( .B1(n20307), .B2(n17198), .A(n17197), .ZN(P2_U3057) );
  INV_X1 U20336 ( .A(n20633), .ZN(n17199) );
  NAND2_X1 U20337 ( .A1(n20464), .A2(n17199), .ZN(n17201) );
  NOR2_X1 U20338 ( .A1(n20894), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20461) );
  INV_X1 U20339 ( .A(n20461), .ZN(n20435) );
  NOR2_X1 U20340 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20435), .ZN(
        n20379) );
  INV_X1 U20341 ( .A(n20379), .ZN(n17200) );
  NAND2_X1 U20342 ( .A1(n17201), .A2(n17200), .ZN(n17204) );
  OAI21_X1 U20343 ( .B1(n10816), .B2(n20559), .A(n11308), .ZN(n17202) );
  OR2_X1 U20344 ( .A1(n20525), .A2(n20435), .ZN(n17207) );
  AOI21_X1 U20345 ( .B1(n17202), .B2(n17207), .A(n20636), .ZN(n17203) );
  NAND2_X1 U20346 ( .A1(n17204), .A2(n17203), .ZN(n20422) );
  INV_X1 U20347 ( .A(n20422), .ZN(n20432) );
  INV_X1 U20348 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17213) );
  INV_X1 U20349 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18494) );
  INV_X1 U20350 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17712) );
  OAI22_X2 U20351 ( .A1(n18494), .A2(n20289), .B1(n17712), .B2(n20290), .ZN(
        n20762) );
  INV_X1 U20352 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17725) );
  NAND2_X1 U20353 ( .A1(n17205), .A2(n20287), .ZN(n20654) );
  OAI22_X1 U20354 ( .A1(n20765), .A2(n20409), .B1(n17207), .B2(n20654), .ZN(
        n17206) );
  AOI21_X1 U20355 ( .B1(n20427), .B2(n20762), .A(n17206), .ZN(n17212) );
  NAND2_X1 U20356 ( .A1(n20379), .A2(n20906), .ZN(n17209) );
  INV_X1 U20357 ( .A(n17207), .ZN(n20426) );
  OAI21_X1 U20358 ( .B1(n10816), .B2(n20426), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17208) );
  NAND2_X1 U20359 ( .A1(n17209), .A2(n17208), .ZN(n20428) );
  NAND2_X1 U20360 ( .A1(n20428), .A2(n20761), .ZN(n17211) );
  OAI211_X1 U20361 ( .C1(n20432), .C2(n17213), .A(n17212), .B(n17211), .ZN(
        P2_U3092) );
  NAND2_X1 U20362 ( .A1(n20735), .A2(n20870), .ZN(n17214) );
  NOR2_X1 U20363 ( .A1(n20885), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20495) );
  NAND2_X1 U20364 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20495), .ZN(
        n17223) );
  NAND2_X1 U20365 ( .A1(n17214), .A2(n17223), .ZN(n17218) );
  NAND2_X1 U20366 ( .A1(n10818), .A2(n11308), .ZN(n17216) );
  NAND2_X1 U20367 ( .A1(n20462), .A2(n20495), .ZN(n17221) );
  AND2_X1 U20368 ( .A1(n17221), .A2(n20881), .ZN(n17215) );
  AOI21_X1 U20369 ( .B1(n17216), .B2(n17215), .A(n20636), .ZN(n17217) );
  NAND2_X1 U20370 ( .A1(n17218), .A2(n17217), .ZN(n20604) );
  INV_X1 U20371 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17227) );
  INV_X1 U20372 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17727) );
  INV_X1 U20373 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17714) );
  OAI22_X2 U20374 ( .A1(n16442), .A2(n20289), .B1(n17714), .B2(n20290), .ZN(
        n20756) );
  AOI22_X1 U20375 ( .A1(n20622), .A2(n20700), .B1(n20592), .B2(n20756), .ZN(
        n17226) );
  INV_X1 U20376 ( .A(n17221), .ZN(n20602) );
  OAI21_X1 U20377 ( .B1(n10818), .B2(n20602), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17222) );
  OAI21_X1 U20378 ( .B1(n17223), .B2(n20881), .A(n17222), .ZN(n20603) );
  NOR2_X2 U20379 ( .A1(n17224), .A2(n20280), .ZN(n20754) );
  AOI22_X1 U20380 ( .A1(n20603), .A2(n20755), .B1(n20754), .B2(n20602), .ZN(
        n17225) );
  OAI211_X1 U20381 ( .C1(n20595), .C2(n17227), .A(n17226), .B(n17225), .ZN(
        P2_U3139) );
  OAI21_X1 U20382 ( .B1(n20669), .B2(n20622), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17233) );
  INV_X1 U20383 ( .A(n20381), .ZN(n17234) );
  INV_X1 U20384 ( .A(n20434), .ZN(n20323) );
  NAND3_X1 U20385 ( .A1(n17234), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20323), .ZN(n17232) );
  AND2_X1 U20386 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20678) );
  AND2_X1 U20387 ( .A1(n20678), .A2(n17256), .ZN(n20638) );
  NAND2_X1 U20388 ( .A1(n20638), .A2(n20679), .ZN(n17228) );
  INV_X1 U20389 ( .A(n17228), .ZN(n20620) );
  AND2_X1 U20390 ( .A1(n17228), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17229) );
  NAND2_X1 U20391 ( .A1(n17230), .A2(n17229), .ZN(n17235) );
  OAI211_X1 U20392 ( .C1(n20620), .C2(n11308), .A(n17235), .B(n20731), .ZN(
        n17231) );
  INV_X1 U20393 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17729) );
  INV_X1 U20394 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17716) );
  OAI22_X2 U20395 ( .A1(n16450), .A2(n20289), .B1(n17716), .B2(n20290), .ZN(
        n20750) );
  AOI22_X1 U20396 ( .A1(n20669), .A2(n20696), .B1(n20622), .B2(n20750), .ZN(
        n17241) );
  NAND4_X1 U20397 ( .A1(n17234), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20323), .A4(n11308), .ZN(n17237) );
  INV_X1 U20398 ( .A(n17235), .ZN(n17236) );
  AOI22_X1 U20399 ( .A1(n20621), .A2(n20749), .B1(n20620), .B2(n20748), .ZN(
        n17240) );
  OAI211_X1 U20400 ( .C1(n20626), .C2(n17242), .A(n17241), .B(n17240), .ZN(
        P2_U3146) );
  AOI22_X1 U20401 ( .A1(n20669), .A2(n20700), .B1(n20622), .B2(n20756), .ZN(
        n17244) );
  AOI22_X1 U20402 ( .A1(n20621), .A2(n20755), .B1(n20620), .B2(n20754), .ZN(
        n17243) );
  OAI211_X1 U20403 ( .C1(n20626), .C2(n17245), .A(n17244), .B(n17243), .ZN(
        P2_U3147) );
  NAND2_X1 U20404 ( .A1(n17246), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17286) );
  MUX2_X1 U20405 ( .A(n17248), .B(n17247), .S(n17253), .Z(n17281) );
  INV_X1 U20406 ( .A(n17281), .ZN(n17258) );
  INV_X1 U20407 ( .A(n17253), .ZN(n17279) );
  MUX2_X1 U20408 ( .A(n17249), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17279), .Z(n17259) );
  NAND2_X1 U20409 ( .A1(n17255), .A2(n17256), .ZN(n17252) );
  NOR2_X1 U20410 ( .A1(n17250), .A2(n20679), .ZN(n17251) );
  NAND2_X1 U20411 ( .A1(n17252), .A2(n17251), .ZN(n17254) );
  OAI211_X1 U20412 ( .C1(n17256), .C2(n17255), .A(n17254), .B(n17253), .ZN(
        n17257) );
  AOI21_X1 U20413 ( .B1(n17281), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n17257), .ZN(n17260) );
  AOI211_X1 U20414 ( .C1(n20894), .C2(n17258), .A(n17259), .B(n17260), .ZN(
        n17262) );
  INV_X1 U20415 ( .A(n17259), .ZN(n17282) );
  INV_X1 U20416 ( .A(n17260), .ZN(n17261) );
  OAI22_X1 U20417 ( .A1(n17262), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n17282), .B2(n17261), .ZN(n17284) );
  INV_X1 U20418 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17545) );
  AOI21_X1 U20419 ( .B1(n17265), .B2(n17264), .A(n17263), .ZN(n17270) );
  MUX2_X1 U20420 ( .A(n17268), .B(n17267), .S(n17266), .Z(n17269) );
  AOI211_X1 U20421 ( .C1(n17272), .C2(n17271), .A(n17270), .B(n17269), .ZN(
        n20899) );
  OAI21_X1 U20422 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n17273), .ZN(n17277) );
  INV_X1 U20423 ( .A(n20902), .ZN(n17275) );
  NAND4_X1 U20424 ( .A1(n17277), .A2(n17276), .A3(n17275), .A4(n17274), .ZN(
        n17278) );
  AOI21_X1 U20425 ( .B1(n17279), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n17278), .ZN(n17280) );
  OAI211_X1 U20426 ( .C1(n17282), .C2(n17281), .A(n20899), .B(n17280), .ZN(
        n17283) );
  AOI21_X1 U20427 ( .B1(n17284), .B2(n17545), .A(n17283), .ZN(n17678) );
  AOI21_X1 U20428 ( .B1(n17678), .B2(n17290), .A(n20912), .ZN(n17285) );
  AOI211_X1 U20429 ( .C1(n17287), .C2(n11258), .A(n17286), .B(n17285), .ZN(
        n17672) );
  INV_X1 U20430 ( .A(n17672), .ZN(n17667) );
  INV_X1 U20431 ( .A(n17288), .ZN(n20872) );
  OAI21_X1 U20432 ( .B1(n20872), .B2(n17289), .A(n17677), .ZN(n17292) );
  NAND2_X1 U20433 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20559), .ZN(n17666) );
  AOI211_X1 U20434 ( .C1(n17667), .C2(n17666), .A(n20917), .B(n17290), .ZN(
        n17291) );
  AOI211_X1 U20435 ( .C1(n17667), .C2(n17292), .A(n20083), .B(n17291), .ZN(
        n17293) );
  INV_X1 U20436 ( .A(n17293), .ZN(P2_U3177) );
  OAI211_X1 U20437 ( .C1(n17667), .C2(n11308), .A(n17295), .B(n17294), .ZN(
        P2_U3593) );
  INV_X1 U20438 ( .A(n17297), .ZN(n17298) );
  NAND2_X1 U20439 ( .A1(n17299), .A2(n17298), .ZN(n17300) );
  INV_X2 U20440 ( .A(n18992), .ZN(n17302) );
  INV_X1 U20441 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17301) );
  INV_X1 U20442 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17303) );
  INV_X1 U20443 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17304) );
  INV_X1 U20444 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18927) );
  NAND2_X1 U20445 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19297) );
  INV_X1 U20446 ( .A(n19297), .ZN(n18972) );
  NAND2_X1 U20447 ( .A1(n18972), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19280) );
  NOR2_X1 U20448 ( .A1(n19280), .A2(n19287), .ZN(n19251) );
  NAND2_X1 U20449 ( .A1(n19251), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19249) );
  INV_X1 U20450 ( .A(n19249), .ZN(n19254) );
  NAND2_X1 U20451 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19254), .ZN(
        n19236) );
  NOR2_X1 U20452 ( .A1(n19236), .A2(n17304), .ZN(n17387) );
  AND2_X1 U20453 ( .A1(n17387), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17305) );
  MUX2_X1 U20454 ( .A(n19006), .B(n17308), .S(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(n17306) );
  AND2_X2 U20455 ( .A1(n17309), .A2(n17306), .ZN(n18879) );
  NAND2_X1 U20456 ( .A1(n18879), .A2(n19217), .ZN(n17307) );
  NAND2_X2 U20457 ( .A1(n17307), .A2(n19006), .ZN(n18804) );
  NOR2_X1 U20458 ( .A1(n19228), .A2(n19217), .ZN(n18831) );
  NAND2_X1 U20459 ( .A1(n18891), .A2(n18831), .ZN(n17310) );
  NAND2_X2 U20460 ( .A1(n18804), .A2(n17310), .ZN(n18873) );
  INV_X1 U20461 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18839) );
  INV_X1 U20462 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18864) );
  NOR2_X1 U20463 ( .A1(n18864), .A2(n19162), .ZN(n19176) );
  INV_X1 U20464 ( .A(n19176), .ZN(n18835) );
  NOR2_X1 U20465 ( .A1(n18839), .A2(n18835), .ZN(n19165) );
  AND3_X1 U20466 ( .A1(n19165), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17311) );
  NAND2_X1 U20467 ( .A1(n18831), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19164) );
  NAND2_X1 U20468 ( .A1(n19179), .A2(n19165), .ZN(n19168) );
  NOR2_X1 U20469 ( .A1(n19168), .A2(n19174), .ZN(n19121) );
  NAND2_X1 U20470 ( .A1(n19121), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18792) );
  INV_X1 U20471 ( .A(n18792), .ZN(n17312) );
  INV_X1 U20472 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18877) );
  NAND2_X1 U20473 ( .A1(n19006), .A2(n18877), .ZN(n18871) );
  NOR2_X1 U20474 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18871), .ZN(
        n17313) );
  NAND2_X1 U20475 ( .A1(n17313), .A2(n19162), .ZN(n18833) );
  NOR2_X1 U20476 ( .A1(n18833), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18816) );
  INV_X1 U20477 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19141) );
  NAND3_X1 U20478 ( .A1(n18816), .A2(n19141), .A3(n19174), .ZN(n17314) );
  NAND2_X1 U20479 ( .A1(n17315), .A2(n17314), .ZN(n17316) );
  AND2_X1 U20480 ( .A1(n18793), .A2(n19006), .ZN(n18781) );
  INV_X1 U20481 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n19110) );
  AND2_X1 U20482 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n19102) );
  NAND2_X1 U20483 ( .A1(n17319), .A2(n17318), .ZN(n18752) );
  INV_X1 U20484 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U20485 ( .A1(n19006), .A2(n18740), .ZN(n17320) );
  NOR2_X1 U20486 ( .A1(n18752), .A2(n17320), .ZN(n17490) );
  INV_X1 U20487 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17696) );
  NAND2_X1 U20488 ( .A1(n17490), .A2(n17696), .ZN(n17536) );
  NAND2_X1 U20489 ( .A1(n17536), .A2(n19006), .ZN(n17323) );
  AND2_X2 U20490 ( .A1(n17321), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17377) );
  INV_X1 U20491 ( .A(n17377), .ZN(n18751) );
  AND2_X1 U20492 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17322) );
  AOI22_X1 U20493 ( .A1(n17323), .A2(n17679), .B1(n17537), .B2(n18890), .ZN(
        n17327) );
  XNOR2_X1 U20494 ( .A(n19006), .B(n17368), .ZN(n17326) );
  NAND2_X1 U20495 ( .A1(n17368), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17352) );
  NAND3_X1 U20496 ( .A1(n17323), .A2(n17537), .A3(n17352), .ZN(n17324) );
  OAI211_X1 U20497 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17368), .A(
        n17324), .B(n17326), .ZN(n17325) );
  OAI21_X1 U20498 ( .B1(n17327), .B2(n17326), .A(n17325), .ZN(n17375) );
  NAND2_X1 U20499 ( .A1(n19878), .A2(n17328), .ZN(n17331) );
  INV_X1 U20500 ( .A(n19873), .ZN(n17329) );
  INV_X1 U20501 ( .A(n20026), .ZN(n19906) );
  NOR2_X1 U20502 ( .A1(n18591), .A2(n17332), .ZN(n17339) );
  NAND2_X1 U20503 ( .A1(n17339), .A2(n17335), .ZN(n17340) );
  NAND2_X1 U20504 ( .A1(n17337), .A2(n17336), .ZN(n17338) );
  INV_X1 U20505 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18939) );
  INV_X1 U20506 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18794) );
  NOR2_X1 U20507 ( .A1(n18792), .A2(n18794), .ZN(n19125) );
  NAND2_X1 U20508 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19125), .ZN(
        n18770) );
  NOR2_X1 U20509 ( .A1(n19110), .A2(n18770), .ZN(n18744) );
  NAND2_X1 U20510 ( .A1(n18744), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18739) );
  NOR2_X1 U20511 ( .A1(n18739), .A2(n18740), .ZN(n17376) );
  NOR2_X1 U20512 ( .A1(n17697), .A2(n17696), .ZN(n17695) );
  NAND2_X1 U20513 ( .A1(n17695), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17341) );
  XNOR2_X1 U20514 ( .A(n17341), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17373) );
  XNOR2_X1 U20515 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17350) );
  NAND2_X1 U20516 ( .A1(n9779), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17344) );
  OAI21_X4 U20517 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20025), .A(n17342), 
        .ZN(n19096) );
  AOI21_X2 U20518 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n9612), .A(
        n19801), .ZN(n18942) );
  OR2_X1 U20519 ( .A1(n17344), .A2(n18942), .ZN(n17680) );
  NOR2_X1 U20520 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18880), .ZN(
        n17701) );
  NAND2_X1 U20521 ( .A1(n19801), .A2(n17344), .ZN(n17690) );
  OAI211_X1 U20522 ( .C1(n17345), .C2(n19095), .A(n19096), .B(n17690), .ZN(
        n17691) );
  NOR2_X1 U20523 ( .A1(n17701), .A2(n17691), .ZN(n17681) );
  OR2_X1 U20524 ( .A1(n17681), .A2(n17346), .ZN(n17349) );
  NOR2_X2 U20525 ( .A1(n19083), .A2(n19004), .ZN(n19027) );
  OR2_X1 U20526 ( .A1(n19400), .A2(n19993), .ZN(n17366) );
  INV_X1 U20527 ( .A(n17366), .ZN(n17347) );
  AOI21_X1 U20528 ( .B1(n18935), .B2(n10198), .A(n17347), .ZN(n17348) );
  OAI211_X1 U20529 ( .C1(n17350), .C2(n17680), .A(n17349), .B(n17348), .ZN(
        n17356) );
  NOR2_X2 U20530 ( .A1(n17351), .A2(n10273), .ZN(n19291) );
  NAND2_X1 U20531 ( .A1(n18744), .A2(n19157), .ZN(n19104) );
  NAND3_X1 U20532 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17689) );
  INV_X1 U20533 ( .A(n17352), .ZN(n17354) );
  AOI21_X1 U20534 ( .B1(n17693), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17368), .ZN(n17353) );
  AOI21_X1 U20535 ( .B1(n17693), .B2(n17354), .A(n17353), .ZN(n17370) );
  OR2_X2 U20536 ( .A1(n19099), .A2(n17386), .ZN(n19009) );
  NOR2_X1 U20537 ( .A1(n17370), .A2(n19009), .ZN(n17355) );
  AOI211_X1 U20538 ( .C1(n17373), .C2(n19088), .A(n17356), .B(n17355), .ZN(
        n17357) );
  OAI21_X1 U20539 ( .B1(n17375), .B2(n18991), .A(n17357), .ZN(P3_U2799) );
  INV_X1 U20540 ( .A(n19385), .ZN(n19350) );
  INV_X1 U20541 ( .A(n17387), .ZN(n19210) );
  AND3_X1 U20542 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n19338), .ZN(n19328) );
  NAND2_X1 U20543 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n19328), .ZN(
        n19209) );
  OR3_X1 U20544 ( .A1(n13945), .A2(n17358), .A3(n19209), .ZN(n19250) );
  NOR2_X1 U20545 ( .A1(n19210), .A2(n19250), .ZN(n17359) );
  NAND2_X1 U20546 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17359), .ZN(
        n19221) );
  NOR2_X1 U20547 ( .A1(n18739), .A2(n19221), .ZN(n17362) );
  INV_X1 U20548 ( .A(n18744), .ZN(n19101) );
  INV_X1 U20549 ( .A(n17359), .ZN(n19161) );
  OAI21_X1 U20550 ( .B1(n19101), .B2(n19161), .A(n19224), .ZN(n17361) );
  NOR2_X1 U20551 ( .A1(n17360), .A2(n19209), .ZN(n19223) );
  NAND2_X1 U20552 ( .A1(n17387), .A2(n19223), .ZN(n19159) );
  OAI21_X1 U20553 ( .B1(n19101), .B2(n19159), .A(n19880), .ZN(n19107) );
  OAI211_X1 U20554 ( .C1(n19314), .C2(n17362), .A(n17361), .B(n19107), .ZN(
        n17380) );
  AOI22_X1 U20555 ( .A1(n19350), .A2(n17689), .B1(n19397), .B2(n17380), .ZN(
        n17542) );
  INV_X1 U20556 ( .A(n17542), .ZN(n17363) );
  AOI211_X1 U20557 ( .C1(n19350), .C2(n17679), .A(n19392), .B(n17363), .ZN(
        n17369) );
  OAI22_X1 U20558 ( .A1(n19375), .A2(n19159), .B1(n17364), .B2(n19161), .ZN(
        n19124) );
  AND2_X1 U20559 ( .A1(n19124), .A2(n17376), .ZN(n17494) );
  NAND2_X1 U20560 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n19397), .ZN(
        n17538) );
  INV_X1 U20561 ( .A(n17538), .ZN(n17365) );
  NAND4_X1 U20562 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17494), .A3(
        n17365), .A4(n17368), .ZN(n17367) );
  OAI211_X1 U20563 ( .C1(n17369), .C2(n17368), .A(n17367), .B(n17366), .ZN(
        n17372) );
  NOR2_X1 U20564 ( .A1(n19404), .A2(n17386), .ZN(n19259) );
  INV_X1 U20565 ( .A(n19259), .ZN(n19321) );
  NOR2_X1 U20566 ( .A1(n17370), .A2(n19321), .ZN(n17371) );
  AOI211_X1 U20567 ( .C1(n17373), .C2(n19389), .A(n17372), .B(n17371), .ZN(
        n17374) );
  OAI21_X1 U20568 ( .B1(n17375), .B2(n19310), .A(n17374), .ZN(P3_U2831) );
  INV_X1 U20569 ( .A(n17697), .ZN(n17384) );
  NAND2_X1 U20570 ( .A1(n17376), .A2(n19157), .ZN(n17694) );
  OAI21_X1 U20571 ( .B1(n17377), .B2(n19006), .A(n18752), .ZN(n18738) );
  XNOR2_X1 U20572 ( .A(n19006), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18737) );
  NAND2_X1 U20573 ( .A1(n18738), .A2(n18737), .ZN(n18736) );
  MUX2_X1 U20574 ( .A(n17694), .B(n18736), .S(n17386), .Z(n17379) );
  INV_X1 U20575 ( .A(n19875), .ZN(n17378) );
  NAND3_X1 U20576 ( .A1(n17379), .A2(n17378), .A3(n18754), .ZN(n17383) );
  INV_X1 U20577 ( .A(n17380), .ZN(n17381) );
  OAI21_X1 U20578 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n19269), .A(
        n17381), .ZN(n17489) );
  INV_X1 U20579 ( .A(n17489), .ZN(n17382) );
  OAI211_X1 U20580 ( .C1(n17384), .C2(n19379), .A(n17383), .B(n17382), .ZN(
        n17385) );
  AOI21_X1 U20581 ( .B1(n17385), .B2(n19400), .A(n19392), .ZN(n17391) );
  INV_X1 U20582 ( .A(n19289), .ZN(n18971) );
  OAI22_X1 U20583 ( .A1(n18971), .A2(n19379), .B1(n18969), .B2(n19290), .ZN(
        n19274) );
  AOI21_X1 U20584 ( .B1(n19274), .B2(n17387), .A(n19124), .ZN(n19169) );
  NOR2_X1 U20585 ( .A1(n19169), .A2(n19390), .ZN(n19186) );
  INV_X1 U20586 ( .A(n19186), .ZN(n19148) );
  OAI22_X1 U20587 ( .A1(n18739), .A2(n19148), .B1(n18754), .B2(n19404), .ZN(
        n17389) );
  NOR2_X1 U20588 ( .A1(n19400), .A2(n19990), .ZN(n18733) );
  NOR3_X1 U20589 ( .A1(n18752), .A2(n18737), .A3(n19310), .ZN(n17388) );
  AOI211_X1 U20590 ( .C1(n17389), .C2(n18740), .A(n18733), .B(n17388), .ZN(
        n17390) );
  OAI21_X1 U20591 ( .B1(n17391), .B2(n18740), .A(n17390), .ZN(P3_U2834) );
  NAND2_X1 U20592 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n18246), .ZN(n18235) );
  NAND2_X1 U20593 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18239), .ZN(n18229) );
  OR2_X1 U20594 ( .A1(n17867), .A2(n18229), .ZN(n17475) );
  NAND2_X1 U20595 ( .A1(n18458), .A2(n18229), .ZN(n18233) );
  OAI21_X1 U20596 ( .B1(n17393), .B2(n18473), .A(n18233), .ZN(n18224) );
  AOI22_X1 U20597 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9592), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20598 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18258), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20599 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20600 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17394) );
  NAND4_X1 U20601 ( .A1(n17397), .A2(n17396), .A3(n17395), .A4(n17394), .ZN(
        n17403) );
  AOI22_X1 U20602 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20603 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20604 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20605 ( .A1(n18426), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17398) );
  NAND4_X1 U20606 ( .A1(n17401), .A2(n17400), .A3(n17399), .A4(n17398), .ZN(
        n17402) );
  NOR2_X1 U20607 ( .A1(n17403), .A2(n17402), .ZN(n17473) );
  AOI22_X1 U20608 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17407) );
  AOI22_X1 U20609 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n9619), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20610 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n9596), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20611 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17404) );
  NAND4_X1 U20612 ( .A1(n17407), .A2(n17406), .A3(n17405), .A4(n17404), .ZN(
        n17413) );
  AOI22_X1 U20613 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n9586), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20614 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U20615 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U20616 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17408) );
  NAND4_X1 U20617 ( .A1(n17411), .A2(n17410), .A3(n17409), .A4(n17408), .ZN(
        n17412) );
  NOR2_X1 U20618 ( .A1(n17413), .A2(n17412), .ZN(n18231) );
  AOI22_X1 U20619 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U20620 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17416) );
  AOI22_X1 U20621 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17415) );
  AOI22_X1 U20622 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17414) );
  NAND4_X1 U20623 ( .A1(n17417), .A2(n17416), .A3(n17415), .A4(n17414), .ZN(
        n17424) );
  AOI22_X1 U20624 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9592), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20625 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U20626 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20627 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17419) );
  NAND4_X1 U20628 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17423) );
  NOR2_X1 U20629 ( .A1(n17424), .A2(n17423), .ZN(n18243) );
  AOI22_X1 U20630 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20631 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20632 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20633 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17425) );
  NAND4_X1 U20634 ( .A1(n17428), .A2(n17427), .A3(n17426), .A4(n17425), .ZN(
        n17434) );
  AOI22_X1 U20635 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20636 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20637 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20638 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20639 ( .A1(n17432), .A2(n17431), .A3(n17430), .A4(n17429), .ZN(
        n17433) );
  OR2_X1 U20640 ( .A1(n17434), .A2(n17433), .ZN(n18249) );
  INV_X1 U20641 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17435) );
  NOR2_X1 U20642 ( .A1(n17436), .A2(n17435), .ZN(n17441) );
  INV_X1 U20643 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17439) );
  INV_X1 U20644 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17437) );
  OAI22_X1 U20645 ( .A1(n9608), .A2(n17439), .B1(n17438), .B2(n17437), .ZN(
        n17440) );
  AOI211_X1 U20646 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n18428), .A(
        n17441), .B(n17440), .ZN(n17449) );
  AOI22_X1 U20647 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20648 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20649 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20650 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17442) );
  AND4_X1 U20651 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17448) );
  AOI22_X1 U20652 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20653 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17446) );
  NAND4_X1 U20654 ( .A1(n17449), .A2(n17448), .A3(n17447), .A4(n17446), .ZN(
        n18250) );
  NAND2_X1 U20655 ( .A1(n18249), .A2(n18250), .ZN(n18248) );
  NOR2_X1 U20656 ( .A1(n18243), .A2(n18248), .ZN(n18242) );
  AOI22_X1 U20657 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U20658 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20659 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U20660 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17450) );
  NAND4_X1 U20661 ( .A1(n17453), .A2(n17452), .A3(n17451), .A4(n17450), .ZN(
        n17459) );
  AOI22_X1 U20662 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20663 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20664 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20665 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17454) );
  NAND4_X1 U20666 ( .A1(n17457), .A2(n17456), .A3(n17455), .A4(n17454), .ZN(
        n17458) );
  OR2_X1 U20667 ( .A1(n17459), .A2(n17458), .ZN(n18237) );
  NAND2_X1 U20668 ( .A1(n18242), .A2(n18237), .ZN(n18236) );
  NOR2_X1 U20669 ( .A1(n18231), .A2(n18236), .ZN(n18230) );
  AOI22_X1 U20670 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U20671 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U20672 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20673 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17461) );
  NAND4_X1 U20674 ( .A1(n17464), .A2(n17463), .A3(n17462), .A4(n17461), .ZN(
        n17472) );
  AOI22_X1 U20675 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20676 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U20677 ( .A1(n18271), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20678 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17467) );
  NAND4_X1 U20679 ( .A1(n17470), .A2(n17469), .A3(n17468), .A4(n17467), .ZN(
        n17471) );
  OR2_X1 U20680 ( .A1(n17472), .A2(n17471), .ZN(n18227) );
  NAND2_X1 U20681 ( .A1(n18230), .A2(n18227), .ZN(n18226) );
  NOR2_X1 U20682 ( .A1(n17473), .A2(n18226), .ZN(n18221) );
  AOI21_X1 U20683 ( .B1(n17473), .B2(n18226), .A(n18221), .ZN(n18490) );
  AOI22_X1 U20684 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18224), .B1(n18490), 
        .B2(n18471), .ZN(n17474) );
  OAI21_X1 U20685 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17475), .A(n17474), .ZN(
        P3_U2675) );
  AOI22_X1 U20686 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20687 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20688 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20689 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17476) );
  NAND4_X1 U20690 ( .A1(n17479), .A2(n17478), .A3(n17477), .A4(n17476), .ZN(
        n17485) );
  AOI22_X1 U20691 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20692 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20693 ( .A1(n18410), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13057), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U20694 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17480) );
  NAND4_X1 U20695 ( .A1(n17483), .A2(n17482), .A3(n17481), .A4(n17480), .ZN(
        n17484) );
  NOR2_X1 U20696 ( .A1(n17485), .A2(n17484), .ZN(n18567) );
  OAI21_X1 U20697 ( .B1(n18389), .B2(n18377), .A(n18034), .ZN(n17486) );
  INV_X1 U20698 ( .A(n17486), .ZN(n17488) );
  NAND4_X1 U20699 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n18376), .A4(n18451), .ZN(n18375) );
  NAND2_X1 U20700 ( .A1(n18458), .A2(n18375), .ZN(n17487) );
  OAI22_X1 U20701 ( .A1(n18567), .A2(n18458), .B1(n17488), .B2(n17487), .ZN(
        P3_U2690) );
  INV_X1 U20702 ( .A(n19227), .ZN(n19145) );
  AOI21_X1 U20703 ( .B1(n19145), .B2(n18740), .A(n17489), .ZN(n17497) );
  AOI21_X1 U20704 ( .B1(n17491), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17490), .ZN(n17492) );
  XNOR2_X1 U20705 ( .A(n17492), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17700) );
  OAI22_X1 U20706 ( .A1(n19379), .A2(n17697), .B1(n19290), .B2(n17694), .ZN(
        n17493) );
  NOR2_X1 U20707 ( .A1(n17494), .A2(n17493), .ZN(n17539) );
  NOR2_X1 U20708 ( .A1(n17539), .A2(n19390), .ZN(n17496) );
  OAI22_X1 U20709 ( .A1(n17693), .A2(n19321), .B1(n17695), .B2(n19406), .ZN(
        n17495) );
  NOR2_X1 U20710 ( .A1(n19392), .A2(n17495), .ZN(n17541) );
  NAND2_X1 U20711 ( .A1(n19402), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17703) );
  INV_X1 U20712 ( .A(n17509), .ZN(n17512) );
  NOR2_X1 U20713 ( .A1(n17498), .A2(n21307), .ZN(n17499) );
  AND2_X1 U20714 ( .A1(n17500), .A2(n17499), .ZN(n17505) );
  AOI211_X1 U20715 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n17505), .A(
        n17502), .B(n17501), .ZN(n17503) );
  INV_X1 U20716 ( .A(n17503), .ZN(n17504) );
  OAI21_X1 U20717 ( .B1(n17505), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17504), .ZN(n17506) );
  AND2_X1 U20718 ( .A1(n21203), .A2(n17506), .ZN(n17507) );
  OAI222_X1 U20719 ( .A1(n17510), .A2(n17509), .B1(n17508), .B2(n17507), .C1(
        n21203), .C2(n17506), .ZN(n17511) );
  OAI21_X1 U20720 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17512), .A(
        n17511), .ZN(n17521) );
  INV_X1 U20721 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21154) );
  OAI21_X1 U20722 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17513), .ZN(n17516) );
  AND4_X1 U20723 ( .A1(n17516), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n17515), 
        .A4(n17514), .ZN(n17517) );
  NAND2_X1 U20724 ( .A1(n17518), .A2(n17517), .ZN(n17519) );
  AOI211_X1 U20725 ( .C1(n17521), .C2(n21154), .A(n17520), .B(n17519), .ZN(
        n17528) );
  NOR3_X1 U20726 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11775), .A3(n21389), 
        .ZN(n17524) );
  OAI22_X1 U20727 ( .A1(n17525), .A2(n17524), .B1(n17523), .B2(n17522), .ZN(
        n17631) );
  INV_X1 U20728 ( .A(n17631), .ZN(n17526) );
  OAI21_X1 U20729 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n17528), .A(n17526), 
        .ZN(n17531) );
  AOI22_X1 U20730 ( .A1(n17528), .A2(n17631), .B1(n17637), .B2(n17527), .ZN(
        n17530) );
  AOI211_X1 U20731 ( .C1(n21467), .C2(n11775), .A(n17530), .B(n17529), .ZN(
        n17535) );
  OAI21_X1 U20732 ( .B1(n17532), .B2(n17534), .A(n17531), .ZN(n17533) );
  AOI22_X1 U20733 ( .A1(n17535), .A2(n17534), .B1(n21369), .B2(n17533), .ZN(
        P1_U3161) );
  INV_X1 U20734 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17679) );
  NOR2_X1 U20735 ( .A1(n19400), .A2(n19995), .ZN(n17683) );
  NOR3_X1 U20736 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17539), .A3(
        n17538), .ZN(n17540) );
  NAND2_X1 U20737 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21379) );
  INV_X1 U20738 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21377) );
  NOR2_X1 U20739 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21377), .ZN(n21383) );
  NOR2_X1 U20740 ( .A1(n21377), .A2(n21389), .ZN(n21387) );
  AOI211_X1 U20741 ( .C1(HOLD), .C2(n21383), .A(n17543), .B(n21387), .ZN(
        n17544) );
  OAI221_X1 U20742 ( .B1(n21379), .B2(HOLD), .C1(n21379), .C2(
        P1_STATE_REG_2__SCAN_IN), .A(n17544), .ZN(P1_U3195) );
  AND2_X1 U20743 ( .A1(n21055), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U20744 ( .A1(n17545), .A2(n20892), .ZN(P2_U3047) );
  INV_X1 U20745 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18678) );
  NOR2_X1 U20746 ( .A1(n18475), .A2(n18678), .ZN(n18616) );
  NAND2_X1 U20747 ( .A1(n10457), .A2(n9967), .ZN(n18589) );
  AOI22_X1 U20748 ( .A1(n18613), .A2(BUF2_REG_0__SCAN_IN), .B1(n18612), .B2(
        n13905), .ZN(n17546) );
  OAI221_X1 U20749 ( .B1(n18616), .B2(n18678), .C1(n18616), .C2(n18589), .A(
        n17546), .ZN(P3_U2735) );
  INV_X1 U20750 ( .A(n17547), .ZN(n17548) );
  AOI22_X1 U20751 ( .A1(n21014), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n21018), 
        .B2(n17548), .ZN(n17559) );
  AOI22_X1 U20752 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21016), .B1(
        n21013), .B2(n17549), .ZN(n17558) );
  NAND3_X1 U20753 ( .A1(n17551), .A2(n17550), .A3(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n17554) );
  AOI21_X1 U20754 ( .B1(n17554), .B2(n17553), .A(n17552), .ZN(n17555) );
  AOI21_X1 U20755 ( .B1(n17556), .B2(n20989), .A(n17555), .ZN(n17557) );
  NAND4_X1 U20756 ( .A1(n17559), .A2(n17558), .A3(n17557), .A4(n20998), .ZN(
        P1_U2826) );
  AOI21_X1 U20757 ( .B1(n21016), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20952), .ZN(n17561) );
  NAND2_X1 U20758 ( .A1(n21014), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n17560) );
  OAI211_X1 U20759 ( .C1(n20983), .C2(n17562), .A(n17561), .B(n17560), .ZN(
        n17563) );
  AOI21_X1 U20760 ( .B1(n21013), .B2(n17564), .A(n17563), .ZN(n17568) );
  AOI22_X1 U20761 ( .A1(n17566), .A2(n20989), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n17565), .ZN(n17567) );
  OAI211_X1 U20762 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n17569), .A(n17568), 
        .B(n17567), .ZN(P1_U2829) );
  AOI22_X1 U20763 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n21133), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17576) );
  INV_X1 U20764 ( .A(n20973), .ZN(n17574) );
  NAND2_X1 U20765 ( .A1(n17571), .A2(n17570), .ZN(n17572) );
  XNOR2_X1 U20766 ( .A(n17573), .B(n17572), .ZN(n17606) );
  AOI22_X1 U20767 ( .A1(n21101), .A2(n17574), .B1(n17606), .B2(n21102), .ZN(
        n17575) );
  OAI211_X1 U20768 ( .C1(n21106), .C2(n20967), .A(n17576), .B(n17575), .ZN(
        P1_U2992) );
  AOI22_X1 U20769 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21133), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17581) );
  XNOR2_X1 U20770 ( .A(n17578), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17579) );
  XNOR2_X1 U20771 ( .A(n17577), .B(n17579), .ZN(n17616) );
  AOI22_X1 U20772 ( .A1(n21032), .A2(n21101), .B1(n17616), .B2(n21102), .ZN(
        n17580) );
  OAI211_X1 U20773 ( .C1(n21106), .C2(n20982), .A(n17581), .B(n17580), .ZN(
        P1_U2993) );
  AOI22_X1 U20774 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n21133), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17589) );
  INV_X1 U20775 ( .A(n17582), .ZN(n17587) );
  OAI21_X1 U20776 ( .B1(n17585), .B2(n17584), .A(n17583), .ZN(n17586) );
  INV_X1 U20777 ( .A(n17586), .ZN(n17624) );
  AOI22_X1 U20778 ( .A1(n17587), .A2(n21101), .B1(n17624), .B2(n21102), .ZN(
        n17588) );
  OAI211_X1 U20779 ( .C1(n21106), .C2(n17590), .A(n17589), .B(n17588), .ZN(
        P1_U2994) );
  NAND2_X1 U20780 ( .A1(n17593), .A2(n21113), .ZN(n17610) );
  INV_X1 U20781 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U20782 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17594), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15255), .ZN(n17605) );
  AOI21_X1 U20783 ( .B1(n21142), .B2(n17596), .A(n17595), .ZN(n17604) );
  INV_X1 U20784 ( .A(n17597), .ZN(n21122) );
  INV_X1 U20785 ( .A(n17598), .ZN(n17599) );
  OAI21_X1 U20786 ( .B1(n21122), .B2(n17600), .A(n17599), .ZN(n21117) );
  AOI21_X1 U20787 ( .B1(n21148), .B2(n17614), .A(n21117), .ZN(n17626) );
  OAI21_X1 U20788 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17601), .A(
        n17626), .ZN(n17607) );
  AOI22_X1 U20789 ( .A1(n17602), .A2(n21145), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17607), .ZN(n17603) );
  OAI211_X1 U20790 ( .C1(n17610), .C2(n17605), .A(n17604), .B(n17603), .ZN(
        P1_U3023) );
  AOI22_X1 U20791 ( .A1(n21142), .A2(n20977), .B1(n21133), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17609) );
  AOI22_X1 U20792 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17607), .B1(
        n17606), .B2(n21145), .ZN(n17608) );
  OAI211_X1 U20793 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17610), .A(
        n17609), .B(n17608), .ZN(P1_U3024) );
  OR2_X1 U20794 ( .A1(n17612), .A2(n17611), .ZN(n17613) );
  AND2_X1 U20795 ( .A1(n14494), .A2(n17613), .ZN(n21029) );
  AOI22_X1 U20796 ( .A1(n21142), .A2(n21029), .B1(n21133), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17618) );
  NOR2_X1 U20797 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17614), .ZN(
        n17615) );
  AOI22_X1 U20798 ( .A1(n17616), .A2(n21145), .B1(n21113), .B2(n17615), .ZN(
        n17617) );
  OAI211_X1 U20799 ( .C1(n17626), .C2(n17619), .A(n17618), .B(n17617), .ZN(
        P1_U3025) );
  NAND2_X1 U20800 ( .A1(n21112), .A2(n21113), .ZN(n17628) );
  OAI22_X1 U20801 ( .A1(n17622), .A2(n17621), .B1(n17620), .B2(n15176), .ZN(
        n17623) );
  AOI21_X1 U20802 ( .B1(n17624), .B2(n21145), .A(n17623), .ZN(n17625) );
  OAI221_X1 U20803 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17628), .C1(
        n17627), .C2(n17626), .A(n17625), .ZN(P1_U3026) );
  NAND4_X1 U20804 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n11775), .A4(n21389), .ZN(n17629) );
  NAND2_X1 U20805 ( .A1(n17630), .A2(n17629), .ZN(n21370) );
  OAI21_X1 U20806 ( .B1(n17632), .B2(n21370), .A(n17631), .ZN(n17633) );
  OAI21_X1 U20807 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n17637), .A(n17633), 
        .ZN(n17634) );
  AOI221_X1 U20808 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21468), .C1(n21467), 
        .C2(n21468), .A(n17634), .ZN(P1_U3162) );
  OAI21_X1 U20809 ( .B1(n17637), .B2(n17636), .A(n17635), .ZN(P1_U3466) );
  AOI22_X1 U20810 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n20179), .B1(n20209), 
        .B2(n17638), .ZN(n17643) );
  AOI222_X1 U20811 ( .A1(n17641), .A2(n20196), .B1(n20213), .B2(n17640), .C1(
        n20205), .C2(n17639), .ZN(n17642) );
  OAI211_X1 U20812 ( .C1(n17654), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        P2_U3009) );
  AOI22_X1 U20813 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n20179), .B1(n20209), 
        .B2(n17645), .ZN(n17653) );
  NAND3_X1 U20814 ( .A1(n17647), .A2(n17646), .A3(n20205), .ZN(n17648) );
  OAI21_X1 U20815 ( .B1(n20194), .B2(n17649), .A(n17648), .ZN(n17650) );
  AOI21_X1 U20816 ( .B1(n17651), .B2(n20196), .A(n17650), .ZN(n17652) );
  OAI211_X1 U20817 ( .C1(n17655), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P2_U3011) );
  OAI22_X1 U20818 ( .A1(n20242), .A2(n13666), .B1(n20227), .B2(n17656), .ZN(
        n17659) );
  INV_X1 U20819 ( .A(n17657), .ZN(n20246) );
  MUX2_X1 U20820 ( .A(n20236), .B(n20246), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n17658) );
  AOI211_X1 U20821 ( .C1(n17661), .C2(n17660), .A(n17659), .B(n17658), .ZN(
        n17663) );
  OAI211_X1 U20822 ( .C1(n20219), .C2(n17664), .A(n17663), .B(n17662), .ZN(
        P2_U3046) );
  OAI21_X1 U20823 ( .B1(n20917), .B2(n17666), .A(n17665), .ZN(n17674) );
  NOR2_X1 U20824 ( .A1(n20917), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17671) );
  INV_X1 U20825 ( .A(n20916), .ZN(n17670) );
  MUX2_X1 U20826 ( .A(n17668), .B(n17667), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17669) );
  AOI22_X1 U20827 ( .A1(n17672), .A2(n17671), .B1(n17670), .B2(n17669), .ZN(
        n17673) );
  AOI211_X1 U20828 ( .C1(n20898), .C2(n17675), .A(n17674), .B(n17673), .ZN(
        n17676) );
  OAI21_X1 U20829 ( .B1(n17678), .B2(n17677), .A(n17676), .ZN(P2_U3176) );
  NAND3_X1 U20830 ( .A1(n18744), .A2(n18902), .A3(n17679), .ZN(n17688) );
  AOI22_X1 U20831 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17681), .B1(
        n17680), .B2(n17836), .ZN(n17682) );
  AOI211_X1 U20832 ( .C1(n18935), .C2(n17835), .A(n17683), .B(n17682), .ZN(
        n17687) );
  OAI22_X1 U20833 ( .A1(n17695), .A2(n19100), .B1(n17693), .B2(n19009), .ZN(
        n17685) );
  AOI22_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17685), .B1(
        n19011), .B2(n17684), .ZN(n17686) );
  OAI211_X1 U20835 ( .C1(n17689), .C2(n17688), .A(n17687), .B(n17686), .ZN(
        P3_U2800) );
  INV_X1 U20836 ( .A(n17690), .ZN(n17692) );
  AOI22_X1 U20837 ( .A1(n9779), .A2(n17692), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17691), .ZN(n17705) );
  AOI211_X1 U20838 ( .C1(n17696), .C2(n17694), .A(n17693), .B(n19009), .ZN(
        n17699) );
  AOI211_X1 U20839 ( .C1(n17697), .C2(n17696), .A(n17695), .B(n19100), .ZN(
        n17698) );
  AOI211_X1 U20840 ( .C1(n19011), .C2(n17700), .A(n17699), .B(n17698), .ZN(
        n17704) );
  OAI21_X1 U20841 ( .B1(n17701), .B2(n18935), .A(n17844), .ZN(n17702) );
  NAND4_X1 U20842 ( .A1(n17705), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        P3_U2801) );
  NOR3_X1 U20843 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), .A3(
        P3_BE_N_REG_0__SCAN_IN), .ZN(n17707) );
  NOR4_X1 U20844 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_BE_N_REG_3__SCAN_IN), .A4(P3_D_C_N_REG_SCAN_IN), .ZN(n17706) );
  NAND4_X1 U20845 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17707), .A3(n17706), .A4(
        U215), .ZN(U213) );
  INV_X2 U20846 ( .A(U214), .ZN(n17764) );
  INV_X1 U20847 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17801) );
  OAI222_X1 U20848 ( .A1(U212), .A2(n20144), .B1(n17766), .B2(n20286), .C1(
        U214), .C2(n17801), .ZN(U216) );
  INV_X1 U20849 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20279) );
  AOI22_X1 U20850 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17753), .ZN(n17709) );
  OAI21_X1 U20851 ( .B1(n20279), .B2(n17766), .A(n17709), .ZN(U217) );
  INV_X1 U20852 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20272) );
  AOI22_X1 U20853 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17753), .ZN(n17710) );
  OAI21_X1 U20854 ( .B1(n20272), .B2(n17766), .A(n17710), .ZN(U218) );
  AOI22_X1 U20855 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17753), .ZN(n17711) );
  OAI21_X1 U20856 ( .B1(n17712), .B2(n17766), .A(n17711), .ZN(U219) );
  INV_X1 U20857 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n17713) );
  OAI222_X1 U20858 ( .A1(U212), .A2(n17795), .B1(n17766), .B2(n17714), .C1(
        U214), .C2(n17713), .ZN(U220) );
  AOI22_X1 U20859 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17753), .ZN(n17715) );
  OAI21_X1 U20860 ( .B1(n17716), .B2(n17766), .A(n17715), .ZN(U221) );
  AOI22_X1 U20861 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17753), .ZN(n17717) );
  OAI21_X1 U20862 ( .B1(n17718), .B2(n17766), .A(n17717), .ZN(U222) );
  AOI22_X1 U20863 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17753), .ZN(n17719) );
  OAI21_X1 U20864 ( .B1(n17720), .B2(n17766), .A(n17719), .ZN(U223) );
  AOI22_X1 U20865 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17753), .ZN(n17721) );
  OAI21_X1 U20866 ( .B1(n20291), .B2(n17766), .A(n17721), .ZN(U224) );
  INV_X1 U20867 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20281) );
  AOI22_X1 U20868 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17753), .ZN(n17722) );
  OAI21_X1 U20869 ( .B1(n20281), .B2(n17766), .A(n17722), .ZN(U225) );
  INV_X1 U20870 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n17723) );
  OAI222_X1 U20871 ( .A1(U214), .A2(n17723), .B1(U212), .B2(n17789), .C1(
        n20275), .C2(n17766), .ZN(U226) );
  AOI22_X1 U20872 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17753), .ZN(n17724) );
  OAI21_X1 U20873 ( .B1(n17725), .B2(n17766), .A(n17724), .ZN(U227) );
  AOI22_X1 U20874 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17753), .ZN(n17726) );
  OAI21_X1 U20875 ( .B1(n17727), .B2(n17766), .A(n17726), .ZN(U228) );
  AOI22_X1 U20876 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17753), .ZN(n17728) );
  OAI21_X1 U20877 ( .B1(n17729), .B2(n17766), .A(n17728), .ZN(U229) );
  AOI22_X1 U20878 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17753), .ZN(n17730) );
  OAI21_X1 U20879 ( .B1(n17731), .B2(n17766), .A(n17730), .ZN(U230) );
  AOI22_X1 U20880 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17753), .ZN(n17732) );
  OAI21_X1 U20881 ( .B1(n17733), .B2(n17766), .A(n17732), .ZN(U231) );
  AOI22_X1 U20882 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17753), .ZN(n17734) );
  OAI21_X1 U20883 ( .B1(n14438), .B2(n17766), .A(n17734), .ZN(U232) );
  INV_X1 U20884 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U20885 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17753), .ZN(n17735) );
  OAI21_X1 U20886 ( .B1(n17736), .B2(n17766), .A(n17735), .ZN(U233) );
  INV_X1 U20887 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n17738) );
  AOI22_X1 U20888 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17753), .ZN(n17737) );
  OAI21_X1 U20889 ( .B1(n17738), .B2(n17766), .A(n17737), .ZN(U234) );
  INV_X1 U20890 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U20891 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17753), .ZN(n17739) );
  OAI21_X1 U20892 ( .B1(n17740), .B2(n17766), .A(n17739), .ZN(U235) );
  INV_X1 U20893 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17742) );
  AOI22_X1 U20894 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17753), .ZN(n17741) );
  OAI21_X1 U20895 ( .B1(n17742), .B2(n17766), .A(n17741), .ZN(U236) );
  INV_X1 U20896 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17744) );
  AOI22_X1 U20897 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17753), .ZN(n17743) );
  OAI21_X1 U20898 ( .B1(n17744), .B2(n17766), .A(n17743), .ZN(U237) );
  INV_X1 U20899 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U20900 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17753), .ZN(n17745) );
  OAI21_X1 U20901 ( .B1(n17746), .B2(n17766), .A(n17745), .ZN(U238) );
  INV_X1 U20902 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17748) );
  AOI22_X1 U20903 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17753), .ZN(n17747) );
  OAI21_X1 U20904 ( .B1(n17748), .B2(n17766), .A(n17747), .ZN(U239) );
  INV_X1 U20905 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U20906 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17753), .ZN(n17749) );
  OAI21_X1 U20907 ( .B1(n17750), .B2(n17766), .A(n17749), .ZN(U240) );
  INV_X1 U20908 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17752) );
  AOI22_X1 U20909 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17753), .ZN(n17751) );
  OAI21_X1 U20910 ( .B1(n17752), .B2(n17766), .A(n17751), .ZN(U241) );
  AOI22_X1 U20911 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17753), .ZN(n17754) );
  OAI21_X1 U20912 ( .B1(n17755), .B2(n17766), .A(n17754), .ZN(U242) );
  INV_X1 U20913 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U20914 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17753), .ZN(n17756) );
  OAI21_X1 U20915 ( .B1(n17757), .B2(n17766), .A(n17756), .ZN(U243) );
  AOI22_X1 U20916 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17753), .ZN(n17758) );
  OAI21_X1 U20917 ( .B1(n17759), .B2(n17766), .A(n17758), .ZN(U244) );
  INV_X1 U20918 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U20919 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17753), .ZN(n17760) );
  OAI21_X1 U20920 ( .B1(n17761), .B2(n17766), .A(n17760), .ZN(U245) );
  INV_X1 U20921 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U20922 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17753), .ZN(n17762) );
  OAI21_X1 U20923 ( .B1(n17763), .B2(n17766), .A(n17762), .ZN(U246) );
  AOI22_X1 U20924 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17764), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17753), .ZN(n17765) );
  OAI21_X1 U20925 ( .B1(n12880), .B2(n17766), .A(n17765), .ZN(U247) );
  OAI22_X1 U20926 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17799), .ZN(n17767) );
  INV_X1 U20927 ( .A(n17767), .ZN(U251) );
  OAI22_X1 U20928 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17799), .ZN(n17768) );
  INV_X1 U20929 ( .A(n17768), .ZN(U252) );
  OAI22_X1 U20930 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17799), .ZN(n17769) );
  INV_X1 U20931 ( .A(n17769), .ZN(U253) );
  OAI22_X1 U20932 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17799), .ZN(n17770) );
  INV_X1 U20933 ( .A(n17770), .ZN(U254) );
  OAI22_X1 U20934 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17799), .ZN(n17771) );
  INV_X1 U20935 ( .A(n17771), .ZN(U255) );
  OAI22_X1 U20936 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17787), .ZN(n17772) );
  INV_X1 U20937 ( .A(n17772), .ZN(U256) );
  OAI22_X1 U20938 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n17799), .ZN(n17773) );
  INV_X1 U20939 ( .A(n17773), .ZN(U257) );
  OAI22_X1 U20940 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n17799), .ZN(n17774) );
  INV_X1 U20941 ( .A(n17774), .ZN(U258) );
  OAI22_X1 U20942 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17799), .ZN(n17775) );
  INV_X1 U20943 ( .A(n17775), .ZN(U259) );
  OAI22_X1 U20944 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17787), .ZN(n17776) );
  INV_X1 U20945 ( .A(n17776), .ZN(U260) );
  OAI22_X1 U20946 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17787), .ZN(n17777) );
  INV_X1 U20947 ( .A(n17777), .ZN(U261) );
  OAI22_X1 U20948 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17787), .ZN(n17778) );
  INV_X1 U20949 ( .A(n17778), .ZN(U262) );
  OAI22_X1 U20950 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17787), .ZN(n17779) );
  INV_X1 U20951 ( .A(n17779), .ZN(U263) );
  OAI22_X1 U20952 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17787), .ZN(n17780) );
  INV_X1 U20953 ( .A(n17780), .ZN(U264) );
  OAI22_X1 U20954 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17787), .ZN(n17781) );
  INV_X1 U20955 ( .A(n17781), .ZN(U265) );
  OAI22_X1 U20956 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17787), .ZN(n17782) );
  INV_X1 U20957 ( .A(n17782), .ZN(U266) );
  OAI22_X1 U20958 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17799), .ZN(n17783) );
  INV_X1 U20959 ( .A(n17783), .ZN(U267) );
  OAI22_X1 U20960 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17799), .ZN(n17784) );
  INV_X1 U20961 ( .A(n17784), .ZN(U268) );
  OAI22_X1 U20962 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17787), .ZN(n17785) );
  INV_X1 U20963 ( .A(n17785), .ZN(U269) );
  OAI22_X1 U20964 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17799), .ZN(n17786) );
  INV_X1 U20965 ( .A(n17786), .ZN(U270) );
  OAI22_X1 U20966 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17787), .ZN(n17788) );
  INV_X1 U20967 ( .A(n17788), .ZN(U271) );
  INV_X1 U20968 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20274) );
  AOI22_X1 U20969 ( .A1(n17799), .A2(n17789), .B1(n20274), .B2(U215), .ZN(U272) );
  OAI22_X1 U20970 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n17799), .ZN(n17790) );
  INV_X1 U20971 ( .A(n17790), .ZN(U273) );
  OAI22_X1 U20972 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17799), .ZN(n17791) );
  INV_X1 U20973 ( .A(n17791), .ZN(U274) );
  OAI22_X1 U20974 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17799), .ZN(n17792) );
  INV_X1 U20975 ( .A(n17792), .ZN(U275) );
  OAI22_X1 U20976 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17799), .ZN(n17793) );
  INV_X1 U20977 ( .A(n17793), .ZN(U276) );
  OAI22_X1 U20978 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17799), .ZN(n17794) );
  INV_X1 U20979 ( .A(n17794), .ZN(U277) );
  AOI22_X1 U20980 ( .A1(n17799), .A2(n17795), .B1(n16442), .B2(U215), .ZN(U278) );
  OAI22_X1 U20981 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17799), .ZN(n17796) );
  INV_X1 U20982 ( .A(n17796), .ZN(U279) );
  OAI22_X1 U20983 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17799), .ZN(n17797) );
  INV_X1 U20984 ( .A(n17797), .ZN(U280) );
  OAI22_X1 U20985 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17799), .ZN(n17798) );
  INV_X1 U20986 ( .A(n17798), .ZN(U281) );
  INV_X1 U20987 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20285) );
  AOI22_X1 U20988 ( .A1(n17799), .A2(n20144), .B1(n20285), .B2(U215), .ZN(U282) );
  INV_X1 U20989 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17800) );
  AOI222_X1 U20990 ( .A1(n17801), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20144), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17800), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17802) );
  INV_X2 U20991 ( .A(n17804), .ZN(n17803) );
  INV_X1 U20992 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19953) );
  INV_X1 U20993 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U20994 ( .A1(n17803), .A2(n19953), .B1(n20823), .B2(n17804), .ZN(
        U347) );
  INV_X1 U20995 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19951) );
  INV_X1 U20996 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U20997 ( .A1(n17802), .A2(n19951), .B1(n20822), .B2(n17804), .ZN(
        U348) );
  INV_X1 U20998 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19948) );
  INV_X1 U20999 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20820) );
  AOI22_X1 U21000 ( .A1(n17803), .A2(n19948), .B1(n20820), .B2(n17804), .ZN(
        U349) );
  INV_X1 U21001 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19947) );
  INV_X1 U21002 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20818) );
  AOI22_X1 U21003 ( .A1(n17803), .A2(n19947), .B1(n20818), .B2(n17804), .ZN(
        U350) );
  INV_X1 U21004 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19945) );
  INV_X1 U21005 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U21006 ( .A1(n17803), .A2(n19945), .B1(n20816), .B2(n17804), .ZN(
        U351) );
  INV_X1 U21007 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19942) );
  INV_X1 U21008 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20814) );
  AOI22_X1 U21009 ( .A1(n17803), .A2(n19942), .B1(n20814), .B2(n17804), .ZN(
        U352) );
  INV_X1 U21010 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19941) );
  INV_X1 U21011 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20813) );
  AOI22_X1 U21012 ( .A1(n17803), .A2(n19941), .B1(n20813), .B2(n17804), .ZN(
        U353) );
  INV_X1 U21013 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19939) );
  AOI22_X1 U21014 ( .A1(n17803), .A2(n19939), .B1(n20812), .B2(n17804), .ZN(
        U354) );
  INV_X1 U21015 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19994) );
  INV_X1 U21016 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U21017 ( .A1(n17803), .A2(n19994), .B1(n20857), .B2(n17804), .ZN(
        U355) );
  INV_X1 U21018 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19992) );
  INV_X1 U21019 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U21020 ( .A1(n17803), .A2(n19992), .B1(n20854), .B2(n17804), .ZN(
        U356) );
  INV_X1 U21021 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19989) );
  INV_X1 U21022 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20852) );
  AOI22_X1 U21023 ( .A1(n17803), .A2(n19989), .B1(n20852), .B2(n17804), .ZN(
        U357) );
  INV_X1 U21024 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19988) );
  INV_X1 U21025 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U21026 ( .A1(n17803), .A2(n19988), .B1(n20850), .B2(n17804), .ZN(
        U358) );
  INV_X1 U21027 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19986) );
  INV_X1 U21028 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20849) );
  AOI22_X1 U21029 ( .A1(n17803), .A2(n19986), .B1(n20849), .B2(n17804), .ZN(
        U359) );
  INV_X1 U21030 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U21031 ( .A1(n17803), .A2(n19983), .B1(n20847), .B2(n17804), .ZN(
        U360) );
  INV_X1 U21032 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19981) );
  INV_X1 U21033 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U21034 ( .A1(n17803), .A2(n19981), .B1(n20845), .B2(n17804), .ZN(
        U361) );
  INV_X1 U21035 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19978) );
  INV_X1 U21036 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20843) );
  AOI22_X1 U21037 ( .A1(n17803), .A2(n19978), .B1(n20843), .B2(n17804), .ZN(
        U362) );
  INV_X1 U21038 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19977) );
  INV_X1 U21039 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20841) );
  AOI22_X1 U21040 ( .A1(n17803), .A2(n19977), .B1(n20841), .B2(n17804), .ZN(
        U363) );
  INV_X1 U21041 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19975) );
  INV_X1 U21042 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U21043 ( .A1(n17803), .A2(n19975), .B1(n20840), .B2(n17804), .ZN(
        U364) );
  INV_X1 U21044 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19937) );
  INV_X1 U21045 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U21046 ( .A1(n17803), .A2(n19937), .B1(n20810), .B2(n17804), .ZN(
        U365) );
  INV_X1 U21047 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19973) );
  INV_X1 U21048 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U21049 ( .A1(n17803), .A2(n19973), .B1(n20838), .B2(n17804), .ZN(
        U366) );
  INV_X1 U21050 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19971) );
  INV_X1 U21051 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U21052 ( .A1(n17803), .A2(n19971), .B1(n20837), .B2(n17804), .ZN(
        U367) );
  INV_X1 U21053 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19969) );
  INV_X1 U21054 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20835) );
  AOI22_X1 U21055 ( .A1(n17803), .A2(n19969), .B1(n20835), .B2(n17804), .ZN(
        U368) );
  INV_X1 U21056 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19967) );
  INV_X1 U21057 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20833) );
  AOI22_X1 U21058 ( .A1(n17803), .A2(n19967), .B1(n20833), .B2(n17804), .ZN(
        U369) );
  INV_X1 U21059 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19964) );
  INV_X1 U21060 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U21061 ( .A1(n17803), .A2(n19964), .B1(n20831), .B2(n17804), .ZN(
        U370) );
  INV_X1 U21062 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19963) );
  INV_X1 U21063 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U21064 ( .A1(n17802), .A2(n19963), .B1(n20830), .B2(n17804), .ZN(
        U371) );
  INV_X1 U21065 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19960) );
  INV_X1 U21066 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20828) );
  AOI22_X1 U21067 ( .A1(n17803), .A2(n19960), .B1(n20828), .B2(n17804), .ZN(
        U372) );
  INV_X1 U21068 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19959) );
  INV_X1 U21069 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U21070 ( .A1(n17803), .A2(n19959), .B1(n20826), .B2(n17804), .ZN(
        U373) );
  INV_X1 U21071 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19957) );
  INV_X1 U21072 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U21073 ( .A1(n17803), .A2(n19957), .B1(n20825), .B2(n17804), .ZN(
        U374) );
  INV_X1 U21074 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19955) );
  INV_X1 U21075 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U21076 ( .A1(n17802), .A2(n19955), .B1(n20824), .B2(n17804), .ZN(
        U375) );
  INV_X1 U21077 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19935) );
  INV_X1 U21078 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20807) );
  AOI22_X1 U21079 ( .A1(n17802), .A2(n19935), .B1(n20807), .B2(n17804), .ZN(
        U376) );
  INV_X1 U21080 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19934) );
  NAND2_X1 U21081 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19934), .ZN(n19924) );
  AOI22_X1 U21082 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19924), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19932), .ZN(n20006) );
  OAI21_X1 U21083 ( .B1(n17805), .B2(n19932), .A(n20003), .ZN(P3_U2633) );
  NAND2_X1 U21084 ( .A1(n20039), .A2(n20009), .ZN(n17809) );
  INV_X1 U21085 ( .A(n17806), .ZN(n17815) );
  NOR2_X1 U21086 ( .A1(n17815), .A2(n17814), .ZN(n17807) );
  OAI21_X1 U21087 ( .B1(n17807), .B2(n18679), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17808) );
  OAI21_X1 U21088 ( .B1(n17809), .B2(n19910), .A(n17808), .ZN(P3_U2634) );
  AOI21_X1 U21089 ( .B1(n19932), .B2(n19934), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17810) );
  AOI22_X1 U21090 ( .A1(n20018), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17810), 
        .B2(n20037), .ZN(P3_U2635) );
  OAI21_X1 U21091 ( .B1(n17811), .B2(BS16), .A(n20006), .ZN(n20004) );
  OAI21_X1 U21092 ( .B1(n20006), .B2(n17812), .A(n20004), .ZN(P3_U2636) );
  OAI211_X1 U21093 ( .C1(n17815), .C2(n17814), .A(n19876), .B(n17813), .ZN(
        n19858) );
  NAND2_X1 U21094 ( .A1(n20026), .A2(n19858), .ZN(n20022) );
  AOI21_X1 U21095 ( .B1(n20022), .B2(P3_FLUSH_REG_SCAN_IN), .A(n17816), .ZN(
        n17817) );
  INV_X1 U21096 ( .A(n17817), .ZN(P3_U2637) );
  NOR4_X1 U21097 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17821) );
  NOR4_X1 U21098 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17820) );
  NOR4_X1 U21099 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17819) );
  NOR4_X1 U21100 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17818) );
  NAND4_X1 U21101 ( .A1(n17821), .A2(n17820), .A3(n17819), .A4(n17818), .ZN(
        n17827) );
  NOR4_X1 U21102 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n17825) );
  AOI211_X1 U21103 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n17824) );
  NOR4_X1 U21104 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17823) );
  NOR4_X1 U21105 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17822) );
  NAND4_X1 U21106 ( .A1(n17825), .A2(n17824), .A3(n17823), .A4(n17822), .ZN(
        n17826) );
  NOR2_X1 U21107 ( .A1(n17827), .A2(n17826), .ZN(n20017) );
  INV_X1 U21108 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17829) );
  NOR3_X1 U21109 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17830) );
  OAI21_X1 U21110 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17830), .A(n20017), .ZN(
        n17828) );
  OAI21_X1 U21111 ( .B1(n20017), .B2(n17829), .A(n17828), .ZN(P3_U2638) );
  INV_X1 U21112 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20010) );
  INV_X1 U21113 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20005) );
  AOI21_X1 U21114 ( .B1(n20010), .B2(n20005), .A(n17830), .ZN(n17832) );
  INV_X1 U21115 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17831) );
  INV_X1 U21116 ( .A(n20017), .ZN(n20012) );
  AOI22_X1 U21117 ( .A1(n20017), .A2(n17832), .B1(n17831), .B2(n20012), .ZN(
        P3_U2639) );
  OAI22_X1 U21118 ( .A1(n17849), .A2(n19995), .B1(n17836), .B2(n18157), .ZN(
        n17837) );
  OAI21_X1 U21119 ( .B1(n18132), .B2(n17839), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17840) );
  AOI22_X1 U21120 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n17848) );
  INV_X1 U21121 ( .A(n17841), .ZN(n17842) );
  AOI211_X1 U21122 ( .C1(n17844), .C2(n17843), .A(n17842), .B(n19913), .ZN(
        n17846) );
  NOR3_X1 U21123 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n19987), .A3(n17863), 
        .ZN(n17850) );
  AOI21_X1 U21124 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18132), .A(n17850), .ZN(
        n17858) );
  OAI21_X1 U21125 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17863), .A(n17880), 
        .ZN(n17856) );
  AOI211_X1 U21126 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17866), .A(n17851), .B(
        n18185), .ZN(n17855) );
  AOI211_X1 U21127 ( .C1(n18735), .C2(n17853), .A(n17852), .B(n19913), .ZN(
        n17854) );
  AOI211_X1 U21128 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17856), .A(n17855), 
        .B(n17854), .ZN(n17857) );
  OAI211_X1 U21129 ( .C1(n17859), .C2(n18157), .A(n17858), .B(n17857), .ZN(
        P3_U2643) );
  AOI211_X1 U21130 ( .C1(n17862), .C2(n17861), .A(n17860), .B(n19913), .ZN(
        n17865) );
  OAI22_X1 U21131 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17863), .B1(n18732), 
        .B2(n18157), .ZN(n17864) );
  AOI211_X1 U21132 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n18132), .A(n17865), .B(
        n17864), .ZN(n17869) );
  OAI211_X1 U21133 ( .C1(n17870), .C2(n17867), .A(n18170), .B(n17866), .ZN(
        n17868) );
  OAI211_X1 U21134 ( .C1(n17880), .C2(n19987), .A(n17869), .B(n17868), .ZN(
        P3_U2644) );
  AOI21_X1 U21135 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n17881), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n17879) );
  AOI22_X1 U21136 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17878) );
  AOI211_X1 U21137 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17871), .A(n17870), .B(
        n18185), .ZN(n17876) );
  INV_X1 U21138 ( .A(n17872), .ZN(n17873) );
  AOI211_X1 U21139 ( .C1(n18768), .C2(n17874), .A(n17873), .B(n19913), .ZN(
        n17875) );
  NOR2_X1 U21140 ( .A1(n17876), .A2(n17875), .ZN(n17877) );
  OAI211_X1 U21141 ( .C1(n17880), .C2(n17879), .A(n17878), .B(n17877), .ZN(
        P3_U2645) );
  INV_X1 U21142 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17896) );
  INV_X1 U21143 ( .A(n17881), .ZN(n17885) );
  NOR2_X1 U21144 ( .A1(n18189), .A2(n17996), .ZN(n18019) );
  INV_X1 U21145 ( .A(n18019), .ZN(n17882) );
  NOR2_X1 U21146 ( .A1(n18167), .A2(n18189), .ZN(n17995) );
  INV_X1 U21147 ( .A(n17995), .ZN(n18187) );
  OAI21_X1 U21148 ( .B1(n17883), .B2(n17882), .A(n18187), .ZN(n17919) );
  INV_X1 U21149 ( .A(n17919), .ZN(n17906) );
  NOR2_X1 U21150 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18179), .ZN(n17897) );
  NOR2_X1 U21151 ( .A1(n17906), .A2(n17897), .ZN(n17884) );
  MUX2_X1 U21152 ( .A(n17885), .B(n17884), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n17895) );
  INV_X1 U21153 ( .A(n17887), .ZN(n17886) );
  OAI21_X1 U21154 ( .B1(n18185), .B2(n17886), .A(n18186), .ZN(n17893) );
  NOR2_X1 U21155 ( .A1(n17887), .A2(n18185), .ZN(n17899) );
  AOI211_X1 U21156 ( .C1(n17890), .C2(n17889), .A(n17888), .B(n19913), .ZN(
        n17891) );
  AOI221_X1 U21157 ( .B1(n17893), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17899), 
        .C2(n17892), .A(n17891), .ZN(n17894) );
  OAI211_X1 U21158 ( .C1(n17896), .C2(n18157), .A(n17895), .B(n17894), .ZN(
        P3_U2646) );
  AOI22_X1 U21159 ( .A1(n18132), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17898), 
        .B2(n17897), .ZN(n17908) );
  INV_X1 U21160 ( .A(n17899), .ZN(n17900) );
  AOI21_X1 U21161 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17916), .A(n17900), .ZN(
        n17905) );
  AOI211_X1 U21162 ( .C1(n17903), .C2(n17902), .A(n17901), .B(n19913), .ZN(
        n17904) );
  AOI211_X1 U21163 ( .C1(n17906), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17905), 
        .B(n17904), .ZN(n17907) );
  OAI211_X1 U21164 ( .C1(n18790), .C2(n18157), .A(n17908), .B(n17907), .ZN(
        P3_U2647) );
  INV_X1 U21165 ( .A(n17924), .ZN(n17910) );
  NOR3_X1 U21166 ( .A1(n18179), .A2(n17996), .A3(n17909), .ZN(n17982) );
  NAND2_X1 U21167 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17982), .ZN(n17975) );
  NOR2_X1 U21168 ( .A1(n17910), .A2(n17975), .ZN(n17938) );
  AOI21_X1 U21169 ( .B1(n17926), .B2(n17938), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n17920) );
  AOI211_X1 U21170 ( .C1(n17913), .C2(n17912), .A(n17911), .B(n19913), .ZN(
        n17915) );
  NOR2_X1 U21171 ( .A1(n18186), .A2(n18241), .ZN(n17914) );
  AOI211_X1 U21172 ( .C1(n18176), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17915), .B(n17914), .ZN(n17918) );
  OAI211_X1 U21173 ( .C1(n17921), .C2(n18241), .A(n18170), .B(n17916), .ZN(
        n17917) );
  OAI211_X1 U21174 ( .C1(n17920), .C2(n17919), .A(n17918), .B(n17917), .ZN(
        P3_U2648) );
  AOI211_X1 U21175 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17939), .A(n17921), .B(
        n18185), .ZN(n17922) );
  AOI21_X1 U21176 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18132), .A(n17922), .ZN(
        n17932) );
  AOI21_X1 U21177 ( .B1(n17923), .B2(n18019), .A(n17995), .ZN(n17981) );
  INV_X1 U21178 ( .A(n17981), .ZN(n17974) );
  OAI21_X1 U21179 ( .B1(n17924), .B2(n17995), .A(n17974), .ZN(n17943) );
  INV_X1 U21180 ( .A(n17938), .ZN(n17925) );
  AOI211_X1 U21181 ( .C1(n19976), .C2(n19974), .A(n17926), .B(n17925), .ZN(
        n17930) );
  AOI211_X1 U21182 ( .C1(n18815), .C2(n17928), .A(n17927), .B(n19913), .ZN(
        n17929) );
  AOI211_X1 U21183 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17943), .A(n17930), 
        .B(n17929), .ZN(n17931) );
  OAI211_X1 U21184 ( .C1(n17933), .C2(n18157), .A(n17932), .B(n17931), .ZN(
        P3_U2649) );
  AOI22_X1 U21185 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17942) );
  AOI211_X1 U21186 ( .C1(n17936), .C2(n17935), .A(n17934), .B(n19913), .ZN(
        n17937) );
  AOI221_X1 U21187 ( .B1(n17938), .B2(n19974), .C1(n17943), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n17937), .ZN(n17941) );
  OAI211_X1 U21188 ( .C1(n17946), .C2(n18279), .A(n18170), .B(n17939), .ZN(
        n17940) );
  NAND3_X1 U21189 ( .A1(n17942), .A2(n17941), .A3(n17940), .ZN(P3_U2650) );
  NOR2_X1 U21190 ( .A1(n19968), .A2(n17975), .ZN(n17961) );
  NAND2_X1 U21191 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17961), .ZN(n17953) );
  INV_X1 U21192 ( .A(n17943), .ZN(n17952) );
  AOI211_X1 U21193 ( .C1(n18846), .C2(n17945), .A(n17944), .B(n19913), .ZN(
        n17950) );
  AOI211_X1 U21194 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17962), .A(n17946), .B(
        n18185), .ZN(n17949) );
  AOI22_X1 U21195 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n17947) );
  INV_X1 U21196 ( .A(n17947), .ZN(n17948) );
  NOR3_X1 U21197 ( .A1(n17950), .A2(n17949), .A3(n17948), .ZN(n17951) );
  OAI221_X1 U21198 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17953), .C1(n19972), 
        .C2(n17952), .A(n17951), .ZN(P3_U2651) );
  AOI22_X1 U21199 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17965) );
  OAI21_X1 U21200 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17975), .A(n17974), 
        .ZN(n17960) );
  INV_X1 U21201 ( .A(n17976), .ZN(n18853) );
  NAND2_X1 U21202 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18853), .ZN(
        n17966) );
  NAND3_X1 U21203 ( .A1(n17954), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18894) );
  NOR2_X1 U21204 ( .A1(n18912), .A2(n18894), .ZN(n18001) );
  AOI21_X1 U21205 ( .B1(n18001), .B2(n18190), .A(n9628), .ZN(n17991) );
  AOI21_X1 U21206 ( .B1(n10198), .B2(n17966), .A(n17991), .ZN(n17958) );
  INV_X1 U21207 ( .A(n17966), .ZN(n17956) );
  OAI21_X1 U21208 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17956), .A(
        n17955), .ZN(n18857) );
  OAI21_X1 U21209 ( .B1(n17958), .B2(n18857), .A(n18097), .ZN(n17957) );
  AOI21_X1 U21210 ( .B1(n17958), .B2(n18857), .A(n17957), .ZN(n17959) );
  AOI221_X1 U21211 ( .B1(n17961), .B2(n19970), .C1(n17960), .C2(
        P3_REIP_REG_19__SCAN_IN), .A(n17959), .ZN(n17964) );
  OAI211_X1 U21212 ( .C1(n17969), .C2(n18306), .A(n18170), .B(n17962), .ZN(
        n17963) );
  NAND4_X1 U21213 ( .A1(n17965), .A2(n17964), .A3(n19400), .A4(n17963), .ZN(
        P3_U2652) );
  OAI21_X1 U21214 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18853), .A(
        n17966), .ZN(n18866) );
  NOR2_X1 U21215 ( .A1(n10189), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18165) );
  INV_X1 U21216 ( .A(n18165), .ZN(n18137) );
  OAI21_X1 U21217 ( .B1(n18854), .B2(n18137), .A(n10198), .ZN(n17968) );
  OAI21_X1 U21218 ( .B1(n18866), .B2(n17968), .A(n18097), .ZN(n17967) );
  AOI21_X1 U21219 ( .B1(n18866), .B2(n17968), .A(n17967), .ZN(n17972) );
  AOI211_X1 U21220 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17983), .A(n17969), .B(
        n18185), .ZN(n17971) );
  OAI22_X1 U21221 ( .A1(n18869), .A2(n18157), .B1(n18186), .B2(n18320), .ZN(
        n17970) );
  NOR4_X1 U21222 ( .A1(n19402), .A2(n17972), .A3(n17971), .A4(n17970), .ZN(
        n17973) );
  OAI221_X1 U21223 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17975), .C1(n19968), 
        .C2(n17974), .A(n17973), .ZN(P3_U2653) );
  AOI22_X1 U21224 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18176), .B1(
        n18132), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n17987) );
  OAI21_X1 U21225 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17977), .A(
        n17976), .ZN(n18883) );
  OAI21_X1 U21226 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17989), .A(
        n10198), .ZN(n17979) );
  OAI21_X1 U21227 ( .B1(n18883), .B2(n17979), .A(n18097), .ZN(n17978) );
  AOI21_X1 U21228 ( .B1(n18883), .B2(n17979), .A(n17978), .ZN(n17980) );
  AOI221_X1 U21229 ( .B1(n17982), .B2(n19966), .C1(n17981), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n17980), .ZN(n17986) );
  OAI211_X1 U21230 ( .C1(n17992), .C2(n17984), .A(n18170), .B(n17983), .ZN(
        n17985) );
  NAND4_X1 U21231 ( .A1(n17987), .A2(n17986), .A3(n19400), .A4(n17985), .ZN(
        P3_U2654) );
  NOR3_X1 U21232 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n17996), .A3(n18179), 
        .ZN(n17988) );
  AOI22_X1 U21233 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18176), .B1(
        P3_REIP_REG_15__SCAN_IN), .B2(n17988), .ZN(n17999) );
  OAI21_X1 U21234 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18001), .A(
        n17989), .ZN(n17990) );
  INV_X1 U21235 ( .A(n17990), .ZN(n18895) );
  INV_X1 U21236 ( .A(n17991), .ZN(n18004) );
  AOI221_X1 U21237 ( .B1(n18895), .B2(n17991), .C1(n17990), .C2(n18004), .A(
        n19913), .ZN(n17994) );
  AOI211_X1 U21238 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18005), .A(n17992), .B(
        n18185), .ZN(n17993) );
  AOI211_X1 U21239 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18132), .A(n17994), .B(
        n17993), .ZN(n17998) );
  NOR2_X1 U21240 ( .A1(n17995), .A2(n18019), .ZN(n18021) );
  NOR3_X1 U21241 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n17996), .A3(n18179), 
        .ZN(n18003) );
  OAI21_X1 U21242 ( .B1(n18021), .B2(n18003), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n17997) );
  NAND4_X1 U21243 ( .A1(n17999), .A2(n17998), .A3(n19400), .A4(n17997), .ZN(
        P3_U2655) );
  NAND2_X1 U21244 ( .A1(n10198), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18000) );
  NAND2_X1 U21245 ( .A1(n18097), .A2(n18000), .ZN(n18184) );
  INV_X1 U21246 ( .A(n18894), .ZN(n18002) );
  AOI21_X1 U21247 ( .B1(n18912), .B2(n18894), .A(n18001), .ZN(n18910) );
  OAI21_X1 U21248 ( .B1(n18002), .B2(n9628), .A(n18910), .ZN(n18012) );
  AOI211_X1 U21249 ( .C1(n18132), .C2(P3_EBX_REG_15__SCAN_IN), .A(n19402), .B(
        n18003), .ZN(n18011) );
  NOR3_X1 U21250 ( .A1(n18910), .A2(n18004), .A3(n19913), .ZN(n18009) );
  OAI211_X1 U21251 ( .C1(n18014), .C2(n18006), .A(n18170), .B(n18005), .ZN(
        n18007) );
  OAI21_X1 U21252 ( .B1(n18157), .B2(n18912), .A(n18007), .ZN(n18008) );
  AOI211_X1 U21253 ( .C1(n18021), .C2(P3_REIP_REG_15__SCAN_IN), .A(n18009), 
        .B(n18008), .ZN(n18010) );
  OAI211_X1 U21254 ( .C1(n18184), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        P3_U2656) );
  NOR2_X1 U21255 ( .A1(n18013), .A2(n18137), .ZN(n18114) );
  AOI21_X1 U21256 ( .B1(n18026), .B2(n18114), .A(n9628), .ZN(n18045) );
  AOI21_X1 U21257 ( .B1(n10198), .B2(n18943), .A(n18045), .ZN(n18029) );
  AND2_X1 U21258 ( .A1(n17954), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18027) );
  OAI21_X1 U21259 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18027), .A(
        n18894), .ZN(n18922) );
  XNOR2_X1 U21260 ( .A(n18029), .B(n18922), .ZN(n18024) );
  AOI211_X1 U21261 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18030), .A(n18014), .B(
        n18185), .ZN(n18015) );
  AOI21_X1 U21262 ( .B1(n18176), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18015), .ZN(n18023) );
  NAND2_X1 U21263 ( .A1(n18167), .A2(n18016), .ZN(n18018) );
  OAI22_X1 U21264 ( .A1(n18019), .A2(n18018), .B1(n18186), .B2(n18017), .ZN(
        n18020) );
  AOI211_X1 U21265 ( .C1(P3_REIP_REG_14__SCAN_IN), .C2(n18021), .A(n19402), 
        .B(n18020), .ZN(n18022) );
  OAI211_X1 U21266 ( .C1(n19913), .C2(n18024), .A(n18023), .B(n18022), .ZN(
        P3_U2657) );
  INV_X1 U21267 ( .A(n18025), .ZN(n18047) );
  AOI21_X1 U21268 ( .B1(n18167), .B2(n18047), .A(n18189), .ZN(n18054) );
  INV_X1 U21269 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19956) );
  NAND2_X1 U21270 ( .A1(n18167), .A2(n19956), .ZN(n18046) );
  INV_X1 U21271 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U21272 ( .A1(n18963), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18121) );
  NOR2_X1 U21273 ( .A1(n19031), .A2(n18121), .ZN(n18108) );
  NAND2_X1 U21274 ( .A1(n18026), .A2(n18108), .ZN(n18931) );
  INV_X1 U21275 ( .A(n18931), .ZN(n18044) );
  NAND2_X1 U21276 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18044), .ZN(
        n18043) );
  INV_X1 U21277 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18035) );
  AOI21_X1 U21278 ( .B1(n18035), .B2(n18043), .A(n18027), .ZN(n18934) );
  INV_X1 U21279 ( .A(n18934), .ZN(n18028) );
  AOI211_X1 U21280 ( .C1(n10198), .C2(n18043), .A(n18028), .B(n18184), .ZN(
        n18039) );
  NOR3_X1 U21281 ( .A1(n18934), .A2(n18029), .A3(n19913), .ZN(n18038) );
  NAND2_X1 U21282 ( .A1(n18167), .A2(n19958), .ZN(n18032) );
  OAI211_X1 U21283 ( .C1(n18041), .C2(n18034), .A(n18170), .B(n18030), .ZN(
        n18031) );
  OAI211_X1 U21284 ( .C1(n18033), .C2(n18032), .A(n19400), .B(n18031), .ZN(
        n18037) );
  OAI22_X1 U21285 ( .A1(n18035), .A2(n18157), .B1(n18186), .B2(n18034), .ZN(
        n18036) );
  NOR4_X1 U21286 ( .A1(n18039), .A2(n18038), .A3(n18037), .A4(n18036), .ZN(
        n18040) );
  OAI221_X1 U21287 ( .B1(n19958), .B2(n18054), .C1(n19958), .C2(n18046), .A(
        n18040), .ZN(P3_U2658) );
  AOI211_X1 U21288 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18056), .A(n18041), .B(
        n18185), .ZN(n18042) );
  AOI21_X1 U21289 ( .B1(n18176), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n18042), .ZN(n18051) );
  OAI21_X1 U21290 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18044), .A(
        n18043), .ZN(n18961) );
  XNOR2_X1 U21291 ( .A(n18045), .B(n18961), .ZN(n18049) );
  OAI22_X1 U21292 ( .A1(n18389), .A2(n18186), .B1(n18047), .B2(n18046), .ZN(
        n18048) );
  AOI211_X1 U21293 ( .C1(n18097), .C2(n18049), .A(n19402), .B(n18048), .ZN(
        n18050) );
  OAI211_X1 U21294 ( .C1(n19956), .C2(n18054), .A(n18051), .B(n18050), .ZN(
        P3_U2659) );
  INV_X1 U21295 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18095) );
  NAND3_X1 U21296 ( .A1(n18052), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18096) );
  NOR2_X1 U21297 ( .A1(n18095), .A2(n18096), .ZN(n18087) );
  NAND2_X1 U21298 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18087), .ZN(
        n18074) );
  NOR2_X1 U21299 ( .A1(n18984), .A2(n18074), .ZN(n18067) );
  OAI21_X1 U21300 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18067), .A(
        n18931), .ZN(n18964) );
  AOI21_X1 U21301 ( .B1(n18067), .B2(n18190), .A(n9628), .ZN(n18053) );
  XNOR2_X1 U21302 ( .A(n18964), .B(n18053), .ZN(n18060) );
  NAND3_X1 U21303 ( .A1(n18167), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n18120), 
        .ZN(n18088) );
  AOI221_X1 U21304 ( .B1(n18055), .B2(n19954), .C1(n18088), .C2(n19954), .A(
        n18054), .ZN(n18059) );
  OAI211_X1 U21305 ( .C1(n18063), .C2(n18062), .A(n18170), .B(n18056), .ZN(
        n18057) );
  OAI21_X1 U21306 ( .B1(n18157), .B2(n18967), .A(n18057), .ZN(n18058) );
  AOI211_X1 U21307 ( .C1(n18060), .C2(n18097), .A(n18059), .B(n18058), .ZN(
        n18061) );
  OAI211_X1 U21308 ( .C1(n18186), .C2(n18062), .A(n18061), .B(n19400), .ZN(
        P3_U2660) );
  AOI211_X1 U21309 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18077), .A(n18063), .B(
        n18185), .ZN(n18064) );
  AOI211_X1 U21310 ( .C1(n18132), .C2(P3_EBX_REG_10__SCAN_IN), .A(n19402), .B(
        n18064), .ZN(n18073) );
  AOI21_X1 U21311 ( .B1(n18167), .B2(n18065), .A(n18189), .ZN(n18124) );
  OAI21_X1 U21312 ( .B1(n18066), .B2(n18179), .A(n18124), .ZN(n18089) );
  INV_X1 U21313 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19952) );
  INV_X1 U21314 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19950) );
  INV_X1 U21315 ( .A(n18088), .ZN(n18117) );
  NAND2_X1 U21316 ( .A1(n18066), .A2(n18117), .ZN(n18083) );
  AOI221_X1 U21317 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n19952), .C2(n19950), .A(n18083), .ZN(n18071) );
  AOI21_X1 U21318 ( .B1(n18984), .B2(n18074), .A(n18067), .ZN(n18982) );
  OAI21_X1 U21319 ( .B1(n18074), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10198), .ZN(n18076) );
  INV_X1 U21320 ( .A(n18076), .ZN(n18069) );
  OAI21_X1 U21321 ( .B1(n18982), .B2(n18069), .A(n18097), .ZN(n18068) );
  AOI21_X1 U21322 ( .B1(n18982), .B2(n18069), .A(n18068), .ZN(n18070) );
  AOI211_X1 U21323 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n18089), .A(n18071), 
        .B(n18070), .ZN(n18072) );
  OAI211_X1 U21324 ( .C1(n18984), .C2(n18157), .A(n18073), .B(n18072), .ZN(
        P3_U2661) );
  INV_X1 U21325 ( .A(n18089), .ZN(n18082) );
  OAI21_X1 U21326 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18087), .A(
        n18074), .ZN(n18996) );
  NOR2_X1 U21327 ( .A1(n19913), .A2(n10198), .ZN(n18142) );
  INV_X1 U21328 ( .A(n18142), .ZN(n18159) );
  AND2_X1 U21329 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18114), .ZN(
        n18086) );
  OAI221_X1 U21330 ( .B1(n18996), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n18996), .C2(n18086), .A(n18097), .ZN(n18075) );
  AOI22_X1 U21331 ( .A1(n18076), .A2(n18996), .B1(n18159), .B2(n18075), .ZN(
        n18080) );
  OAI211_X1 U21332 ( .C1(n18084), .C2(n18402), .A(n18170), .B(n18077), .ZN(
        n18078) );
  OAI211_X1 U21333 ( .C1(n18186), .C2(n18402), .A(n19400), .B(n18078), .ZN(
        n18079) );
  AOI211_X1 U21334 ( .C1(n18176), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n18080), .B(n18079), .ZN(n18081) );
  OAI221_X1 U21335 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n18083), .C1(n19950), 
        .C2(n18082), .A(n18081), .ZN(P3_U2662) );
  AOI211_X1 U21336 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18100), .A(n18084), .B(
        n18185), .ZN(n18085) );
  AOI211_X1 U21337 ( .C1(n18132), .C2(P3_EBX_REG_8__SCAN_IN), .A(n19402), .B(
        n18085), .ZN(n18094) );
  OR2_X1 U21338 ( .A1(n18086), .A2(n9628), .ZN(n18099) );
  AOI21_X1 U21339 ( .B1(n18095), .B2(n18096), .A(n18087), .ZN(n19005) );
  XNOR2_X1 U21340 ( .A(n18099), .B(n19005), .ZN(n18092) );
  NOR2_X1 U21341 ( .A1(n18105), .A2(n18088), .ZN(n18090) );
  MUX2_X1 U21342 ( .A(n18090), .B(n18089), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n18091) );
  AOI21_X1 U21343 ( .B1(n18092), .B2(n18097), .A(n18091), .ZN(n18093) );
  OAI211_X1 U21344 ( .C1(n18095), .C2(n18157), .A(n18094), .B(n18093), .ZN(
        P3_U2663) );
  INV_X1 U21345 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19946) );
  OAI21_X1 U21346 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18108), .A(
        n18096), .ZN(n19019) );
  OAI21_X1 U21347 ( .B1(n18114), .B2(n19019), .A(n18097), .ZN(n18098) );
  AOI22_X1 U21348 ( .A1(n19019), .A2(n18099), .B1(n18159), .B2(n18098), .ZN(
        n18104) );
  OAI211_X1 U21349 ( .C1(n18110), .C2(n18102), .A(n18170), .B(n18100), .ZN(
        n18101) );
  OAI211_X1 U21350 ( .C1(n18186), .C2(n18102), .A(n19400), .B(n18101), .ZN(
        n18103) );
  AOI211_X1 U21351 ( .C1(n18176), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n18104), .B(n18103), .ZN(n18107) );
  OAI211_X1 U21352 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n18117), .B(n18105), .ZN(n18106) );
  OAI211_X1 U21353 ( .C1(n18124), .C2(n19946), .A(n18107), .B(n18106), .ZN(
        P3_U2664) );
  INV_X1 U21354 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19944) );
  AOI21_X1 U21355 ( .B1(n19031), .B2(n18121), .A(n18108), .ZN(n19033) );
  INV_X1 U21356 ( .A(n19033), .ZN(n18109) );
  AOI211_X1 U21357 ( .C1(n10198), .C2(n18121), .A(n18109), .B(n18184), .ZN(
        n18112) );
  AOI211_X1 U21358 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18126), .A(n18110), .B(
        n18185), .ZN(n18111) );
  AOI211_X1 U21359 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18132), .A(n18112), .B(
        n18111), .ZN(n18119) );
  NOR3_X1 U21360 ( .A1(n19033), .A2(n18114), .A3(n18113), .ZN(n18116) );
  OAI21_X1 U21361 ( .B1(n19031), .B2(n18157), .A(n19400), .ZN(n18115) );
  AOI211_X1 U21362 ( .C1(n18117), .C2(n19944), .A(n18116), .B(n18115), .ZN(
        n18118) );
  OAI211_X1 U21363 ( .C1(n18124), .C2(n19944), .A(n18119), .B(n18118), .ZN(
        P3_U2665) );
  AOI21_X1 U21364 ( .B1(n18167), .B2(n18120), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n18123) );
  OAI21_X1 U21365 ( .B1(n19039), .B2(n18137), .A(n10198), .ZN(n18136) );
  NOR2_X1 U21366 ( .A1(n19039), .A2(n10189), .ZN(n18134) );
  OAI21_X1 U21367 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18134), .A(
        n18121), .ZN(n19043) );
  XNOR2_X1 U21368 ( .A(n18136), .B(n19043), .ZN(n18122) );
  OAI22_X1 U21369 ( .A1(n18124), .A2(n18123), .B1(n19913), .B2(n18122), .ZN(
        n18125) );
  AOI211_X1 U21370 ( .C1(n18132), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19402), .B(
        n18125), .ZN(n18128) );
  OAI211_X1 U21371 ( .C1(n18129), .C2(n18442), .A(n18170), .B(n18126), .ZN(
        n18127) );
  OAI211_X1 U21372 ( .C1(n18157), .C2(n19038), .A(n18128), .B(n18127), .ZN(
        P3_U2666) );
  INV_X1 U21373 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19058) );
  NOR3_X1 U21374 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18179), .A3(n18145), .ZN(
        n18131) );
  AOI211_X1 U21375 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18154), .A(n18129), .B(
        n18185), .ZN(n18130) );
  AOI211_X1 U21376 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18132), .A(n18131), .B(
        n18130), .ZN(n18144) );
  NAND2_X1 U21377 ( .A1(n18133), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18148) );
  AOI21_X1 U21378 ( .B1(n19058), .B2(n18148), .A(n18134), .ZN(n19060) );
  NAND2_X1 U21379 ( .A1(n19426), .A2(n20042), .ZN(n18193) );
  INV_X1 U21380 ( .A(n18193), .ZN(n20044) );
  OAI21_X1 U21381 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17465), .A(
        n20044), .ZN(n18135) );
  NAND2_X1 U21382 ( .A1(n18135), .A2(n19400), .ZN(n18141) );
  AOI21_X1 U21383 ( .B1(n18167), .B2(n18145), .A(n18189), .ZN(n18151) );
  NAND2_X1 U21384 ( .A1(n19058), .A2(n18133), .ZN(n19051) );
  OAI22_X1 U21385 ( .A1(n18137), .A2(n19051), .B1(n18136), .B2(n19060), .ZN(
        n18138) );
  INV_X1 U21386 ( .A(n18138), .ZN(n18139) );
  OAI22_X1 U21387 ( .A1(n18151), .A2(n19940), .B1(n18139), .B2(n19913), .ZN(
        n18140) );
  AOI211_X1 U21388 ( .C1(n19060), .C2(n18142), .A(n18141), .B(n18140), .ZN(
        n18143) );
  OAI211_X1 U21389 ( .C1(n19058), .C2(n18157), .A(n18144), .B(n18143), .ZN(
        P3_U2667) );
  NAND2_X1 U21390 ( .A1(n18167), .A2(n18145), .ZN(n18147) );
  NAND2_X1 U21391 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18166) );
  OAI22_X1 U21392 ( .A1(n18147), .A2(n18166), .B1(n18193), .B2(n18146), .ZN(
        n18153) );
  INV_X1 U21393 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19938) );
  NAND2_X1 U21394 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18158) );
  INV_X1 U21395 ( .A(n18158), .ZN(n18163) );
  OAI21_X1 U21396 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18163), .A(
        n18148), .ZN(n19068) );
  OAI21_X1 U21397 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18158), .A(
        n10198), .ZN(n18149) );
  XNOR2_X1 U21398 ( .A(n19068), .B(n18149), .ZN(n18150) );
  OAI22_X1 U21399 ( .A1(n18151), .A2(n19938), .B1(n19913), .B2(n18150), .ZN(
        n18152) );
  AOI211_X1 U21400 ( .C1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n18176), .A(
        n18153), .B(n18152), .ZN(n18156) );
  OAI211_X1 U21401 ( .C1(n18168), .C2(n18453), .A(n18170), .B(n18154), .ZN(
        n18155) );
  OAI211_X1 U21402 ( .C1(n18453), .C2(n18186), .A(n18156), .B(n18155), .ZN(
        P3_U2668) );
  OAI22_X1 U21403 ( .A1(n19082), .A2(n18157), .B1(n18186), .B2(n9829), .ZN(
        n18162) );
  OAI21_X1 U21404 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n18158), .ZN(n19079) );
  OAI22_X1 U21405 ( .A1(n18160), .A2(n18193), .B1(n19079), .B2(n18159), .ZN(
        n18161) );
  AOI211_X1 U21406 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(n18189), .A(n18162), .B(
        n18161), .ZN(n18175) );
  NAND2_X1 U21407 ( .A1(n18163), .A2(n18190), .ZN(n18164) );
  OAI211_X1 U21408 ( .C1(n18165), .C2(n19079), .A(n18177), .B(n18164), .ZN(
        n18174) );
  OAI211_X1 U21409 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18167), .B(n18166), .ZN(n18173) );
  NOR2_X1 U21410 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18171) );
  INV_X1 U21411 ( .A(n18168), .ZN(n18169) );
  OAI211_X1 U21412 ( .C1(n18171), .C2(n9829), .A(n18170), .B(n18169), .ZN(
        n18172) );
  NAND4_X1 U21413 ( .A1(n18175), .A2(n18174), .A3(n18173), .A4(n18172), .ZN(
        P3_U2669) );
  AOI21_X1 U21414 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18177), .A(
        n18176), .ZN(n18183) );
  OAI21_X1 U21415 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18462), .ZN(n18469) );
  OAI22_X1 U21416 ( .A1(n18186), .A2(n9830), .B1(n18185), .B2(n18469), .ZN(
        n18181) );
  OAI22_X1 U21417 ( .A1(n18179), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18193), 
        .B2(n18178), .ZN(n18180) );
  AOI211_X1 U21418 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n18189), .A(n18181), .B(
        n18180), .ZN(n18182) );
  OAI221_X1 U21419 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18184), .C1(
        n10189), .C2(n18183), .A(n18182), .ZN(P3_U2670) );
  NAND2_X1 U21420 ( .A1(n18186), .A2(n18185), .ZN(n18188) );
  AOI22_X1 U21421 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n18188), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n18187), .ZN(n18192) );
  OR3_X1 U21422 ( .A1(n18190), .A2(n20040), .A3(n18189), .ZN(n18191) );
  OAI211_X1 U21423 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18193), .A(
        n18192), .B(n18191), .ZN(P3_U2671) );
  AOI22_X1 U21424 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U21425 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18197) );
  AOI22_X1 U21426 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18196) );
  AOI22_X1 U21427 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18195) );
  NAND4_X1 U21428 ( .A1(n18198), .A2(n18197), .A3(n18196), .A4(n18195), .ZN(
        n18204) );
  AOI22_X1 U21429 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9593), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U21430 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U21431 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U21432 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18199) );
  NAND4_X1 U21433 ( .A1(n18202), .A2(n18201), .A3(n18200), .A4(n18199), .ZN(
        n18203) );
  NOR2_X1 U21434 ( .A1(n18204), .A2(n18203), .ZN(n18215) );
  AOI22_X1 U21435 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18208) );
  AOI22_X1 U21436 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U21437 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U21438 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18205) );
  NAND4_X1 U21439 ( .A1(n18208), .A2(n18207), .A3(n18206), .A4(n18205), .ZN(
        n18214) );
  AOI22_X1 U21440 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U21441 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U21442 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U21443 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18209) );
  NAND4_X1 U21444 ( .A1(n18212), .A2(n18211), .A3(n18210), .A4(n18209), .ZN(
        n18213) );
  OR2_X1 U21445 ( .A1(n18214), .A2(n18213), .ZN(n18220) );
  NAND2_X1 U21446 ( .A1(n18221), .A2(n18220), .ZN(n18219) );
  XNOR2_X1 U21447 ( .A(n18215), .B(n18219), .ZN(n18485) );
  NOR2_X1 U21448 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18216), .ZN(n18218) );
  OAI22_X1 U21449 ( .A1(n18485), .A2(n18458), .B1(n18218), .B2(n18217), .ZN(
        P3_U2673) );
  OAI21_X1 U21450 ( .B1(n18221), .B2(n18220), .A(n18219), .ZN(n18489) );
  NOR2_X1 U21451 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18222), .ZN(n18223) );
  AOI22_X1 U21452 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18224), .B1(n18246), 
        .B2(n18223), .ZN(n18225) );
  OAI21_X1 U21453 ( .B1(n18489), .B2(n18458), .A(n18225), .ZN(P3_U2674) );
  OAI21_X1 U21454 ( .B1(n18230), .B2(n18227), .A(n18226), .ZN(n18498) );
  NAND3_X1 U21455 ( .A1(n18229), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18458), 
        .ZN(n18228) );
  OAI221_X1 U21456 ( .B1(n18229), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18458), 
        .C2(n18498), .A(n18228), .ZN(P3_U2676) );
  INV_X1 U21457 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n18234) );
  AOI21_X1 U21458 ( .B1(n18231), .B2(n18236), .A(n18230), .ZN(n18499) );
  NAND2_X1 U21459 ( .A1(n18499), .A2(n18471), .ZN(n18232) );
  OAI221_X1 U21460 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18235), .C1(n18234), 
        .C2(n18233), .A(n18232), .ZN(P3_U2677) );
  AOI21_X1 U21461 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18458), .A(n18246), .ZN(
        n18238) );
  OAI21_X1 U21462 ( .B1(n18242), .B2(n18237), .A(n18236), .ZN(n18508) );
  OAI22_X1 U21463 ( .A1(n18239), .A2(n18238), .B1(n18508), .B2(n18458), .ZN(
        P3_U2678) );
  NOR2_X1 U21464 ( .A1(n18279), .A2(n18240), .ZN(n18253) );
  NAND2_X1 U21465 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18253), .ZN(n18247) );
  NOR2_X1 U21466 ( .A1(n18241), .A2(n18247), .ZN(n18252) );
  AOI21_X1 U21467 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18458), .A(n18252), .ZN(
        n18245) );
  AOI21_X1 U21468 ( .B1(n18243), .B2(n18248), .A(n18242), .ZN(n18509) );
  INV_X1 U21469 ( .A(n18509), .ZN(n18244) );
  OAI22_X1 U21470 ( .A1(n18246), .A2(n18245), .B1(n18458), .B2(n18244), .ZN(
        P3_U2679) );
  INV_X1 U21471 ( .A(n18247), .ZN(n18266) );
  AOI21_X1 U21472 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18458), .A(n18266), .ZN(
        n18251) );
  OAI21_X1 U21473 ( .B1(n18250), .B2(n18249), .A(n18248), .ZN(n18517) );
  OAI22_X1 U21474 ( .A1(n18252), .A2(n18251), .B1(n18458), .B2(n18517), .ZN(
        P3_U2680) );
  AOI21_X1 U21475 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18458), .A(n18253), .ZN(
        n18265) );
  AOI22_X1 U21476 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U21477 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U21478 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18255) );
  AOI22_X1 U21479 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18254) );
  NAND4_X1 U21480 ( .A1(n18257), .A2(n18256), .A3(n18255), .A4(n18254), .ZN(
        n18264) );
  AOI22_X1 U21481 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18262) );
  AOI22_X1 U21482 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18261) );
  AOI22_X1 U21483 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18260) );
  AOI22_X1 U21484 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18259) );
  NAND4_X1 U21485 ( .A1(n18262), .A2(n18261), .A3(n18260), .A4(n18259), .ZN(
        n18263) );
  NOR2_X1 U21486 ( .A1(n18264), .A2(n18263), .ZN(n18519) );
  OAI22_X1 U21487 ( .A1(n18266), .A2(n18265), .B1(n18519), .B2(n18458), .ZN(
        P3_U2681) );
  AOI22_X1 U21488 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U21489 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U21490 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18268) );
  AOI22_X1 U21491 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18267) );
  NAND4_X1 U21492 ( .A1(n18270), .A2(n18269), .A3(n18268), .A4(n18267), .ZN(
        n18277) );
  AOI22_X1 U21493 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U21494 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U21495 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18273) );
  AOI22_X1 U21496 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18272) );
  NAND4_X1 U21497 ( .A1(n18275), .A2(n18274), .A3(n18273), .A4(n18272), .ZN(
        n18276) );
  NOR2_X1 U21498 ( .A1(n18277), .A2(n18276), .ZN(n18527) );
  AND2_X1 U21499 ( .A1(n18458), .A2(n18278), .ZN(n18293) );
  AOI22_X1 U21500 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18293), .B1(n18280), 
        .B2(n18279), .ZN(n18281) );
  OAI21_X1 U21501 ( .B1(n18527), .B2(n18458), .A(n18281), .ZN(P3_U2682) );
  AOI22_X1 U21502 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18285) );
  AOI22_X1 U21503 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18258), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U21504 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U21505 ( .A1(n18426), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18282) );
  NAND4_X1 U21506 ( .A1(n18285), .A2(n18284), .A3(n18283), .A4(n18282), .ZN(
        n18292) );
  AOI22_X1 U21507 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U21508 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18428), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18289) );
  AOI22_X1 U21509 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18288) );
  AOI22_X1 U21510 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18287) );
  NAND4_X1 U21511 ( .A1(n18290), .A2(n18289), .A3(n18288), .A4(n18287), .ZN(
        n18291) );
  NOR2_X1 U21512 ( .A1(n18292), .A2(n18291), .ZN(n18532) );
  OAI21_X1 U21513 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18294), .A(n18293), .ZN(
        n18295) );
  OAI21_X1 U21514 ( .B1(n18532), .B2(n18458), .A(n18295), .ZN(P3_U2683) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n9620), .B1(n9597), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18299) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n9595), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U21517 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U21518 ( .A1(n18426), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18296) );
  NAND4_X1 U21519 ( .A1(n18299), .A2(n18298), .A3(n18297), .A4(n18296), .ZN(
        n18305) );
  AOI22_X1 U21520 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U21521 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18258), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18301) );
  AOI22_X1 U21523 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18300) );
  NAND4_X1 U21524 ( .A1(n18303), .A2(n18302), .A3(n18301), .A4(n18300), .ZN(
        n18304) );
  NOR2_X1 U21525 ( .A1(n18305), .A2(n18304), .ZN(n18539) );
  NOR2_X1 U21526 ( .A1(n18471), .A2(n18307), .ZN(n18321) );
  OAI222_X1 U21527 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n10457), .B1(
        P3_EBX_REG_19__SCAN_IN), .B2(n18307), .C1(n18321), .C2(n18306), .ZN(
        n18308) );
  OAI21_X1 U21528 ( .B1(n18539), .B2(n18458), .A(n18308), .ZN(P3_U2684) );
  AOI22_X1 U21529 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9620), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U21530 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U21531 ( .A1(n9593), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U21532 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18310) );
  NAND4_X1 U21533 ( .A1(n18313), .A2(n18312), .A3(n18311), .A4(n18310), .ZN(
        n18319) );
  AOI22_X1 U21534 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18317) );
  AOI22_X1 U21535 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18316) );
  AOI22_X1 U21536 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18315) );
  AOI22_X1 U21537 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18314) );
  NAND4_X1 U21538 ( .A1(n18317), .A2(n18316), .A3(n18315), .A4(n18314), .ZN(
        n18318) );
  NOR2_X1 U21539 ( .A1(n18319), .A2(n18318), .ZN(n18544) );
  NAND2_X1 U21540 ( .A1(n18320), .A2(n18335), .ZN(n18322) );
  NAND2_X1 U21541 ( .A1(n18322), .A2(n18321), .ZN(n18323) );
  OAI21_X1 U21542 ( .B1(n18544), .B2(n18458), .A(n18323), .ZN(P3_U2685) );
  AOI22_X1 U21543 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U21544 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18327) );
  AOI22_X1 U21545 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18326) );
  AOI22_X1 U21546 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18324), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18325) );
  NAND4_X1 U21547 ( .A1(n18328), .A2(n18327), .A3(n18326), .A4(n18325), .ZN(
        n18334) );
  AOI22_X1 U21548 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18332) );
  AOI22_X1 U21549 ( .A1(n18410), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18331) );
  AOI22_X1 U21550 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U21551 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18329) );
  NAND4_X1 U21552 ( .A1(n18332), .A2(n18331), .A3(n18330), .A4(n18329), .ZN(
        n18333) );
  NOR2_X1 U21553 ( .A1(n18334), .A2(n18333), .ZN(n18549) );
  OAI21_X1 U21554 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18350), .A(n18335), .ZN(
        n18336) );
  AOI22_X1 U21555 ( .A1(n18471), .A2(n18549), .B1(n18336), .B2(n18458), .ZN(
        P3_U2686) );
  OAI21_X1 U21556 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18337), .A(n18458), .ZN(
        n18349) );
  AOI22_X1 U21557 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18341) );
  AOI22_X1 U21558 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U21559 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U21560 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18338) );
  NAND4_X1 U21561 ( .A1(n18341), .A2(n18340), .A3(n18339), .A4(n18338), .ZN(
        n18348) );
  AOI22_X1 U21562 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18346) );
  AOI22_X1 U21563 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13081), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U21564 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U21565 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18342), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18343) );
  NAND4_X1 U21566 ( .A1(n18346), .A2(n18345), .A3(n18344), .A4(n18343), .ZN(
        n18347) );
  NOR2_X1 U21567 ( .A1(n18348), .A2(n18347), .ZN(n18555) );
  OAI22_X1 U21568 ( .A1(n18350), .A2(n18349), .B1(n18555), .B2(n18458), .ZN(
        P3_U2687) );
  AOI22_X1 U21569 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9593), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U21570 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U21571 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U21572 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18351) );
  NAND4_X1 U21573 ( .A1(n18354), .A2(n18353), .A3(n18352), .A4(n18351), .ZN(
        n18360) );
  AOI22_X1 U21574 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18358) );
  AOI22_X1 U21575 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18357) );
  AOI22_X1 U21576 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13081), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U21577 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18355) );
  NAND4_X1 U21578 ( .A1(n18358), .A2(n18357), .A3(n18356), .A4(n18355), .ZN(
        n18359) );
  NOR2_X1 U21579 ( .A1(n18360), .A2(n18359), .ZN(n18559) );
  OAI21_X1 U21580 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18362), .A(n18361), .ZN(
        n18363) );
  AOI22_X1 U21581 ( .A1(n18471), .A2(n18559), .B1(n18363), .B2(n18458), .ZN(
        P3_U2688) );
  AOI22_X1 U21582 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9591), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18367) );
  AOI22_X1 U21583 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18366) );
  AOI22_X1 U21584 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13081), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U21585 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18364) );
  NAND4_X1 U21586 ( .A1(n18367), .A2(n18366), .A3(n18365), .A4(n18364), .ZN(
        n18373) );
  AOI22_X1 U21587 ( .A1(n9599), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18371) );
  AOI22_X1 U21588 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18370) );
  AOI22_X1 U21589 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U21590 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18368) );
  NAND4_X1 U21591 ( .A1(n18371), .A2(n18370), .A3(n18369), .A4(n18368), .ZN(
        n18372) );
  NOR2_X1 U21592 ( .A1(n18373), .A2(n18372), .ZN(n18563) );
  NAND3_X1 U21593 ( .A1(n18375), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n18458), 
        .ZN(n18374) );
  OAI221_X1 U21594 ( .B1(n18375), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n18458), 
        .C2(n18563), .A(n18374), .ZN(P3_U2689) );
  NAND2_X1 U21595 ( .A1(n18376), .A2(n18451), .ZN(n18390) );
  NAND2_X1 U21596 ( .A1(n18458), .A2(n18377), .ZN(n18404) );
  AOI22_X1 U21597 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18381) );
  AOI22_X1 U21598 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18380) );
  AOI22_X1 U21599 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18271), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18379) );
  AOI22_X1 U21600 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18378) );
  NAND4_X1 U21601 ( .A1(n18381), .A2(n18380), .A3(n18379), .A4(n18378), .ZN(
        n18387) );
  AOI22_X1 U21602 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18385) );
  AOI22_X1 U21603 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18384) );
  AOI22_X1 U21604 ( .A1(n9591), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18383) );
  AOI22_X1 U21605 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18382) );
  NAND4_X1 U21606 ( .A1(n18385), .A2(n18384), .A3(n18383), .A4(n18382), .ZN(
        n18386) );
  NOR2_X1 U21607 ( .A1(n18387), .A2(n18386), .ZN(n18570) );
  OR2_X1 U21608 ( .A1(n18570), .A2(n18458), .ZN(n18388) );
  OAI221_X1 U21609 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18390), .C1(n18389), 
        .C2(n18404), .A(n18388), .ZN(P3_U2691) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n9620), .B1(
        n18258), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U21611 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18393) );
  AOI22_X1 U21612 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U21613 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18391) );
  NAND4_X1 U21614 ( .A1(n18394), .A2(n18393), .A3(n18392), .A4(n18391), .ZN(
        n18401) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n9595), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18399) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n9597), .B1(
        n18395), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18398) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18428), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18397) );
  AOI22_X1 U21618 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18396) );
  NAND4_X1 U21619 ( .A1(n18399), .A2(n18398), .A3(n18397), .A4(n18396), .ZN(
        n18400) );
  NOR2_X1 U21620 ( .A1(n18401), .A2(n18400), .ZN(n18573) );
  INV_X1 U21621 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n18417) );
  NOR2_X1 U21622 ( .A1(n18417), .A2(n18402), .ZN(n18403) );
  AOI21_X1 U21623 ( .B1(n18403), .B2(n18436), .A(P3_EBX_REG_11__SCAN_IN), .ZN(
        n18405) );
  OAI22_X1 U21624 ( .A1(n18573), .A2(n18458), .B1(n18405), .B2(n18404), .ZN(
        P3_U2692) );
  AOI22_X1 U21625 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18409) );
  AOI22_X1 U21626 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13081), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18408) );
  AOI22_X1 U21627 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18407) );
  AOI22_X1 U21628 ( .A1(n9620), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18406) );
  NAND4_X1 U21629 ( .A1(n18409), .A2(n18408), .A3(n18407), .A4(n18406), .ZN(
        n18416) );
  AOI22_X1 U21630 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18258), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18414) );
  AOI22_X1 U21631 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13868), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U21632 ( .A1(n17466), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U21633 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18411) );
  NAND4_X1 U21634 ( .A1(n18414), .A2(n18413), .A3(n18412), .A4(n18411), .ZN(
        n18415) );
  NOR2_X1 U21635 ( .A1(n18416), .A2(n18415), .ZN(n18580) );
  AOI21_X1 U21636 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18436), .A(n18471), .ZN(
        n18435) );
  NAND2_X1 U21637 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18435), .ZN(n18419) );
  NAND4_X1 U21638 ( .A1(n10457), .A2(P3_EBX_REG_9__SCAN_IN), .A3(n18436), .A4(
        n18417), .ZN(n18418) );
  OAI211_X1 U21639 ( .C1(n18580), .C2(n18458), .A(n18419), .B(n18418), .ZN(
        P3_U2693) );
  AOI22_X1 U21640 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U21641 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18424) );
  AOI22_X1 U21642 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13076), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18423) );
  AOI22_X1 U21643 ( .A1(n9619), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17466), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18422) );
  NAND4_X1 U21644 ( .A1(n18425), .A2(n18424), .A3(n18423), .A4(n18422), .ZN(
        n18434) );
  AOI22_X1 U21645 ( .A1(n9592), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18286), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18432) );
  AOI22_X1 U21646 ( .A1(n18258), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18426), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U21647 ( .A1(n13868), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U21648 ( .A1(n18428), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18427), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18429) );
  NAND4_X1 U21649 ( .A1(n18432), .A2(n18431), .A3(n18430), .A4(n18429), .ZN(
        n18433) );
  NOR2_X1 U21650 ( .A1(n18434), .A2(n18433), .ZN(n18582) );
  OAI21_X1 U21651 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18436), .A(n18435), .ZN(
        n18437) );
  OAI21_X1 U21652 ( .B1(n18582), .B2(n18458), .A(n18437), .ZN(P3_U2694) );
  NOR3_X1 U21653 ( .A1(n18470), .A2(n18450), .A3(n18438), .ZN(n18441) );
  AOI21_X1 U21654 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18458), .A(n18445), .ZN(
        n18440) );
  INV_X1 U21655 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18439) );
  OAI22_X1 U21656 ( .A1(n18441), .A2(n18440), .B1(n18439), .B2(n18458), .ZN(
        P3_U2696) );
  NOR3_X1 U21657 ( .A1(n18442), .A2(n18450), .A3(n18473), .ZN(n18449) );
  AOI21_X1 U21658 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18458), .A(n18449), .ZN(
        n18444) );
  INV_X1 U21659 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18443) );
  OAI22_X1 U21660 ( .A1(n18445), .A2(n18444), .B1(n18443), .B2(n18458), .ZN(
        P3_U2697) );
  NOR2_X1 U21661 ( .A1(n18470), .A2(n18450), .ZN(n18446) );
  OAI21_X1 U21662 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18446), .A(n18458), .ZN(
        n18448) );
  INV_X1 U21663 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18447) );
  OAI22_X1 U21664 ( .A1(n18449), .A2(n18448), .B1(n18447), .B2(n18458), .ZN(
        P3_U2698) );
  NOR2_X1 U21665 ( .A1(n18450), .A2(n18473), .ZN(n18456) );
  NAND2_X1 U21666 ( .A1(n18452), .A2(n18451), .ZN(n18457) );
  NOR2_X1 U21667 ( .A1(n18453), .A2(n18457), .ZN(n18461) );
  AOI21_X1 U21668 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18458), .A(n18461), .ZN(
        n18455) );
  INV_X1 U21669 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18454) );
  OAI22_X1 U21670 ( .A1(n18456), .A2(n18455), .B1(n18454), .B2(n18458), .ZN(
        P3_U2699) );
  INV_X1 U21671 ( .A(n18457), .ZN(n18464) );
  AOI21_X1 U21672 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18458), .A(n18464), .ZN(
        n18460) );
  INV_X1 U21673 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18459) );
  OAI22_X1 U21674 ( .A1(n18461), .A2(n18460), .B1(n18459), .B2(n18458), .ZN(
        P3_U2700) );
  OAI221_X1 U21675 ( .B1(n18462), .B2(n18470), .C1(n10457), .C2(n18470), .A(
        n9829), .ZN(n18463) );
  INV_X1 U21676 ( .A(n18463), .ZN(n18465) );
  AOI211_X1 U21677 ( .C1(n18471), .C2(n18466), .A(n18465), .B(n18464), .ZN(
        P3_U2701) );
  INV_X1 U21678 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18467) );
  OAI222_X1 U21679 ( .A1(n18469), .A2(n18473), .B1(n9830), .B2(n18468), .C1(
        n18467), .C2(n18458), .ZN(P3_U2702) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18471), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18470), .ZN(n18472) );
  OAI21_X1 U21681 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18473), .A(n18472), .ZN(
        P3_U2703) );
  INV_X1 U21682 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18624) );
  INV_X1 U21683 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18628) );
  INV_X1 U21684 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18660) );
  NAND2_X1 U21685 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n18597) );
  NAND4_X1 U21686 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n18474) );
  NAND4_X1 U21687 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n18564)
         );
  INV_X1 U21688 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18730) );
  INV_X1 U21689 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18638) );
  INV_X1 U21690 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18640) );
  NOR2_X1 U21691 ( .A1(n18638), .A2(n18640), .ZN(n18521) );
  NAND4_X1 U21692 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n18521), .ZN(n18526) );
  INV_X1 U21693 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18634) );
  NAND2_X1 U21694 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18510), .ZN(n18511) );
  NAND2_X1 U21695 ( .A1(n18482), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n18478) );
  NAND2_X1 U21696 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18550), .ZN(n18477) );
  OAI221_X1 U21697 ( .B1(n18482), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n18478), 
        .C2(n18576), .A(n18477), .ZN(P3_U2704) );
  NOR2_X2 U21698 ( .A1(n18479), .A2(n18615), .ZN(n18551) );
  AOI22_X1 U21699 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18550), .ZN(n18484) );
  NAND2_X1 U21700 ( .A1(n18482), .A2(n18481), .ZN(n18483) );
  OAI211_X1 U21701 ( .C1(n18485), .C2(n18607), .A(n18484), .B(n18483), .ZN(
        P3_U2705) );
  AOI22_X1 U21702 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18550), .ZN(n18488) );
  OAI211_X1 U21703 ( .C1(n9658), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18615), .B(
        n18486), .ZN(n18487) );
  OAI211_X1 U21704 ( .C1(n18489), .C2(n18607), .A(n18488), .B(n18487), .ZN(
        P3_U2706) );
  AOI22_X1 U21705 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18551), .B1(n18612), .B2(
        n18490), .ZN(n18493) );
  AOI211_X1 U21706 ( .C1(n18624), .C2(n18495), .A(n9658), .B(n18576), .ZN(
        n18491) );
  INV_X1 U21707 ( .A(n18491), .ZN(n18492) );
  OAI211_X1 U21708 ( .C1(n18531), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        P3_U2707) );
  AOI22_X1 U21709 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18550), .ZN(n18497) );
  OAI211_X1 U21710 ( .C1(n18500), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18615), .B(
        n18495), .ZN(n18496) );
  OAI211_X1 U21711 ( .C1(n18498), .C2(n18607), .A(n18497), .B(n18496), .ZN(
        P3_U2708) );
  AOI22_X1 U21712 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18551), .B1(n18612), .B2(
        n18499), .ZN(n18503) );
  AOI211_X1 U21713 ( .C1(n18628), .C2(n18504), .A(n18500), .B(n18576), .ZN(
        n18501) );
  INV_X1 U21714 ( .A(n18501), .ZN(n18502) );
  OAI211_X1 U21715 ( .C1(n18531), .C2(n16450), .A(n18503), .B(n18502), .ZN(
        P3_U2709) );
  AOI22_X1 U21716 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18550), .ZN(n18507) );
  OAI211_X1 U21717 ( .C1(n18505), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18615), .B(
        n18504), .ZN(n18506) );
  OAI211_X1 U21718 ( .C1(n18508), .C2(n18607), .A(n18507), .B(n18506), .ZN(
        P3_U2710) );
  AOI22_X1 U21719 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18551), .B1(n18612), .B2(
        n18509), .ZN(n18513) );
  OAI211_X1 U21720 ( .C1(n18510), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18615), .B(
        n18511), .ZN(n18512) );
  OAI211_X1 U21721 ( .C1(n18531), .C2(n16462), .A(n18513), .B(n18512), .ZN(
        P3_U2711) );
  AOI22_X1 U21722 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18550), .ZN(n18516) );
  OAI211_X1 U21723 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n9763), .A(n18615), .B(
        n18514), .ZN(n18515) );
  OAI211_X1 U21724 ( .C1(n18517), .C2(n18607), .A(n18516), .B(n18515), .ZN(
        P3_U2712) );
  NAND2_X1 U21725 ( .A1(n18546), .A2(n18634), .ZN(n18525) );
  INV_X1 U21726 ( .A(n18519), .ZN(n18520) );
  AOI22_X1 U21727 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18550), .B1(n18612), .B2(
        n18520), .ZN(n18524) );
  INV_X1 U21728 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18642) );
  NAND2_X1 U21729 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n18546), .ZN(n18545) );
  NAND2_X1 U21730 ( .A1(n18521), .A2(n18540), .ZN(n18530) );
  NAND2_X1 U21731 ( .A1(n18615), .A2(n18530), .ZN(n18535) );
  OAI21_X1 U21732 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18589), .A(n18535), .ZN(
        n18522) );
  AOI22_X1 U21733 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18551), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18522), .ZN(n18523) );
  OAI211_X1 U21734 ( .C1(n18526), .C2(n18525), .A(n18524), .B(n18523), .ZN(
        P3_U2713) );
  INV_X1 U21735 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18636) );
  OAI22_X1 U21736 ( .A1(n18527), .A2(n18607), .B1(n20274), .B2(n18531), .ZN(
        n18528) );
  AOI21_X1 U21737 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n18551), .A(n18528), .ZN(
        n18529) );
  OAI221_X1 U21738 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18530), .C1(n18636), 
        .C2(n18535), .A(n18529), .ZN(P3_U2714) );
  NAND2_X1 U21739 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18540), .ZN(n18536) );
  OAI22_X1 U21740 ( .A1(n18532), .A2(n18607), .B1(n16488), .B2(n18531), .ZN(
        n18533) );
  AOI21_X1 U21741 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n18551), .A(n18533), .ZN(
        n18534) );
  OAI221_X1 U21742 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n18536), .C1(n18638), 
        .C2(n18535), .A(n18534), .ZN(P3_U2715) );
  AOI22_X1 U21743 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18550), .ZN(n18538) );
  OAI211_X1 U21744 ( .C1(n18540), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18615), .B(
        n18536), .ZN(n18537) );
  OAI211_X1 U21745 ( .C1(n18539), .C2(n18607), .A(n18538), .B(n18537), .ZN(
        P3_U2716) );
  AOI22_X1 U21746 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18550), .ZN(n18543) );
  AOI211_X1 U21747 ( .C1(n18642), .C2(n18545), .A(n18540), .B(n18576), .ZN(
        n18541) );
  INV_X1 U21748 ( .A(n18541), .ZN(n18542) );
  OAI211_X1 U21749 ( .C1(n18544), .C2(n18607), .A(n18543), .B(n18542), .ZN(
        P3_U2717) );
  AOI22_X1 U21750 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18550), .ZN(n18548) );
  OAI211_X1 U21751 ( .C1(n18546), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18615), .B(
        n18545), .ZN(n18547) );
  OAI211_X1 U21752 ( .C1(n18549), .C2(n18607), .A(n18548), .B(n18547), .ZN(
        P3_U2718) );
  AOI22_X1 U21753 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18551), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18550), .ZN(n18554) );
  OAI211_X1 U21754 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18556), .A(n18615), .B(
        n18552), .ZN(n18553) );
  OAI211_X1 U21755 ( .C1(n18555), .C2(n18607), .A(n18554), .B(n18553), .ZN(
        P3_U2719) );
  AOI211_X1 U21756 ( .C1(n18730), .C2(n18560), .A(n18576), .B(n18556), .ZN(
        n18557) );
  AOI21_X1 U21757 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n18613), .A(n18557), .ZN(
        n18558) );
  OAI21_X1 U21758 ( .B1(n18559), .B2(n18607), .A(n18558), .ZN(P3_U2720) );
  OAI211_X1 U21759 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n9678), .A(n18615), .B(
        n18560), .ZN(n18562) );
  NAND2_X1 U21760 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18613), .ZN(n18561) );
  OAI211_X1 U21761 ( .C1(n18563), .C2(n18607), .A(n18562), .B(n18561), .ZN(
        P3_U2721) );
  NAND3_X1 U21762 ( .A1(n10457), .A2(P3_EAX_REG_8__SCAN_IN), .A3(n18593), .ZN(
        n18568) );
  NOR2_X1 U21763 ( .A1(n18564), .A2(n18568), .ZN(n18572) );
  AOI22_X1 U21764 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18613), .B1(n18572), .B2(
        n18723), .ZN(n18566) );
  OR3_X1 U21765 ( .A1(n18723), .A2(n18576), .A3(n18572), .ZN(n18565) );
  OAI211_X1 U21766 ( .C1(n18567), .C2(n18607), .A(n18566), .B(n18565), .ZN(
        P3_U2722) );
  NAND2_X1 U21767 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n18569) );
  INV_X1 U21768 ( .A(n18568), .ZN(n18581) );
  NAND2_X1 U21769 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18581), .ZN(n18577) );
  NOR2_X1 U21770 ( .A1(n18569), .A2(n18577), .ZN(n18575) );
  AOI21_X1 U21771 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18615), .A(n18575), .ZN(
        n18571) );
  OAI222_X1 U21772 ( .A1(n18610), .A2(n18721), .B1(n18572), .B2(n18571), .C1(
        n18607), .C2(n18570), .ZN(P3_U2723) );
  INV_X1 U21773 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18717) );
  INV_X1 U21774 ( .A(n18577), .ZN(n18584) );
  AOI22_X1 U21775 ( .A1(n18584), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n18615), .ZN(n18574) );
  OAI222_X1 U21776 ( .A1(n18610), .A2(n18717), .B1(n18575), .B2(n18574), .C1(
        n18607), .C2(n18573), .ZN(P3_U2724) );
  INV_X1 U21777 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18655) );
  AOI221_X1 U21778 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n18584), .C1(n18655), 
        .C2(n18577), .A(n18576), .ZN(n18578) );
  AOI21_X1 U21779 ( .B1(n18613), .B2(BUF2_REG_10__SCAN_IN), .A(n18578), .ZN(
        n18579) );
  OAI21_X1 U21780 ( .B1(n18580), .B2(n18607), .A(n18579), .ZN(P3_U2725) );
  INV_X1 U21781 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18713) );
  AOI21_X1 U21782 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18615), .A(n18581), .ZN(
        n18583) );
  OAI222_X1 U21783 ( .A1(n18610), .A2(n18713), .B1(n18584), .B2(n18583), .C1(
        n18607), .C2(n18582), .ZN(P3_U2726) );
  OAI211_X1 U21784 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n18593), .A(n18615), .B(
        n18585), .ZN(n18587) );
  NAND2_X1 U21785 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18613), .ZN(n18586) );
  OAI211_X1 U21786 ( .C1(n18588), .C2(n18607), .A(n18587), .B(n18586), .ZN(
        P3_U2727) );
  NOR2_X1 U21787 ( .A1(n18590), .A2(n18589), .ZN(n18600) );
  AOI22_X1 U21788 ( .A1(n18600), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n18615), .ZN(n18592) );
  OAI222_X1 U21789 ( .A1(n19452), .A2(n18610), .B1(n18593), .B2(n18592), .C1(
        n18607), .C2(n18591), .ZN(P3_U2728) );
  AND2_X1 U21790 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18600), .ZN(n18596) );
  AOI21_X1 U21791 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18615), .A(n18600), .ZN(
        n18595) );
  OAI222_X1 U21792 ( .A1(n13757), .A2(n18610), .B1(n18596), .B2(n18595), .C1(
        n18607), .C2(n18594), .ZN(P3_U2729) );
  INV_X1 U21793 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19445) );
  NOR2_X1 U21794 ( .A1(n18597), .A2(n18604), .ZN(n18603) );
  AOI21_X1 U21795 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18615), .A(n18603), .ZN(
        n18599) );
  OAI222_X1 U21796 ( .A1(n19445), .A2(n18610), .B1(n18600), .B2(n18599), .C1(
        n18607), .C2(n18598), .ZN(P3_U2730) );
  INV_X1 U21797 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19441) );
  AOI22_X1 U21798 ( .A1(n18605), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n18615), .ZN(n18602) );
  OAI222_X1 U21799 ( .A1(n19441), .A2(n18610), .B1(n18603), .B2(n18602), .C1(
        n18607), .C2(n18601), .ZN(P3_U2731) );
  INV_X1 U21800 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19437) );
  INV_X1 U21801 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18669) );
  NOR2_X1 U21802 ( .A1(n18669), .A2(n18604), .ZN(n18609) );
  AOI21_X1 U21803 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18615), .A(n18605), .ZN(
        n18608) );
  OAI222_X1 U21804 ( .A1(n19437), .A2(n18610), .B1(n18609), .B2(n18608), .C1(
        n18607), .C2(n18606), .ZN(P3_U2732) );
  AOI22_X1 U21805 ( .A1(n18613), .A2(BUF2_REG_1__SCAN_IN), .B1(n18612), .B2(
        n18611), .ZN(n18618) );
  OAI211_X1 U21806 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n18616), .A(n18615), .B(
        n18614), .ZN(n18617) );
  NAND2_X1 U21807 ( .A1(n18618), .A2(n18617), .ZN(P3_U2734) );
  NAND2_X1 U21808 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18932), .ZN(n18674) );
  INV_X2 U21809 ( .A(n18674), .ZN(n18675) );
  NOR2_X4 U21810 ( .A1(n18675), .A2(n18672), .ZN(n18661) );
  AND2_X1 U21811 ( .A1(n18661), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21812 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18699) );
  AOI22_X1 U21813 ( .A1(n18675), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18621) );
  OAI21_X1 U21814 ( .B1(n18699), .B2(n18645), .A(n18621), .ZN(P3_U2737) );
  INV_X1 U21815 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18697) );
  AOI22_X1 U21816 ( .A1(n18675), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18622) );
  OAI21_X1 U21817 ( .B1(n18697), .B2(n18645), .A(n18622), .ZN(P3_U2738) );
  AOI22_X1 U21818 ( .A1(n18675), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18623) );
  OAI21_X1 U21819 ( .B1(n18624), .B2(n18645), .A(n18623), .ZN(P3_U2739) );
  INV_X1 U21820 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18626) );
  AOI22_X1 U21821 ( .A1(n18675), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18625) );
  OAI21_X1 U21822 ( .B1(n18626), .B2(n18645), .A(n18625), .ZN(P3_U2740) );
  AOI22_X1 U21823 ( .A1(n18675), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18627) );
  OAI21_X1 U21824 ( .B1(n18628), .B2(n18645), .A(n18627), .ZN(P3_U2741) );
  AOI22_X1 U21825 ( .A1(n18675), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18629) );
  OAI21_X1 U21826 ( .B1(n18630), .B2(n18645), .A(n18629), .ZN(P3_U2742) );
  INV_X1 U21827 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18691) );
  AOI22_X1 U21828 ( .A1(n18675), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18631) );
  OAI21_X1 U21829 ( .B1(n18691), .B2(n18645), .A(n18631), .ZN(P3_U2743) );
  AOI22_X1 U21830 ( .A1(n18675), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18632) );
  OAI21_X1 U21831 ( .B1(n9971), .B2(n18645), .A(n18632), .ZN(P3_U2744) );
  AOI22_X1 U21832 ( .A1(n18675), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18633) );
  OAI21_X1 U21833 ( .B1(n18634), .B2(n18645), .A(n18633), .ZN(P3_U2745) );
  AOI22_X1 U21834 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(n18661), .B1(n18675), 
        .B2(P3_UWORD_REG_5__SCAN_IN), .ZN(n18635) );
  OAI21_X1 U21835 ( .B1(n18636), .B2(n18645), .A(n18635), .ZN(P3_U2746) );
  AOI22_X1 U21836 ( .A1(n18675), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18637) );
  OAI21_X1 U21837 ( .B1(n18638), .B2(n18645), .A(n18637), .ZN(P3_U2747) );
  AOI22_X1 U21838 ( .A1(n18675), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18639) );
  OAI21_X1 U21839 ( .B1(n18640), .B2(n18645), .A(n18639), .ZN(P3_U2748) );
  AOI22_X1 U21840 ( .A1(n18675), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18641) );
  OAI21_X1 U21841 ( .B1(n18642), .B2(n18645), .A(n18641), .ZN(P3_U2749) );
  INV_X1 U21842 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18683) );
  AOI22_X1 U21843 ( .A1(n18675), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18643) );
  OAI21_X1 U21844 ( .B1(n18683), .B2(n18645), .A(n18643), .ZN(P3_U2750) );
  INV_X1 U21845 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18646) );
  AOI22_X1 U21846 ( .A1(n18675), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18644) );
  OAI21_X1 U21847 ( .B1(n18646), .B2(n18645), .A(n18644), .ZN(P3_U2751) );
  AOI22_X1 U21848 ( .A1(n18675), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18647) );
  OAI21_X1 U21849 ( .B1(n18730), .B2(n18677), .A(n18647), .ZN(P3_U2752) );
  INV_X1 U21850 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18725) );
  AOI22_X1 U21851 ( .A1(n18675), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18648) );
  OAI21_X1 U21852 ( .B1(n18725), .B2(n18677), .A(n18648), .ZN(P3_U2753) );
  AOI22_X1 U21853 ( .A1(n18675), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18649) );
  OAI21_X1 U21854 ( .B1(n18723), .B2(n18677), .A(n18649), .ZN(P3_U2754) );
  INV_X1 U21855 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18651) );
  AOI22_X1 U21856 ( .A1(n18675), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18650) );
  OAI21_X1 U21857 ( .B1(n18651), .B2(n18677), .A(n18650), .ZN(P3_U2755) );
  INV_X1 U21858 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18653) );
  AOI22_X1 U21859 ( .A1(n18675), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18652) );
  OAI21_X1 U21860 ( .B1(n18653), .B2(n18677), .A(n18652), .ZN(P3_U2756) );
  AOI22_X1 U21861 ( .A1(n18675), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18654) );
  OAI21_X1 U21862 ( .B1(n18655), .B2(n18677), .A(n18654), .ZN(P3_U2757) );
  INV_X1 U21863 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18657) );
  AOI22_X1 U21864 ( .A1(n18675), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18656) );
  OAI21_X1 U21865 ( .B1(n18657), .B2(n18677), .A(n18656), .ZN(P3_U2758) );
  INV_X1 U21866 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18711) );
  AOI22_X1 U21867 ( .A1(n18675), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18658) );
  OAI21_X1 U21868 ( .B1(n18711), .B2(n18677), .A(n18658), .ZN(P3_U2759) );
  AOI22_X1 U21869 ( .A1(n18675), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18659) );
  OAI21_X1 U21870 ( .B1(n18660), .B2(n18677), .A(n18659), .ZN(P3_U2760) );
  AOI22_X1 U21871 ( .A1(n18675), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18662) );
  OAI21_X1 U21872 ( .B1(n18663), .B2(n18677), .A(n18662), .ZN(P3_U2761) );
  INV_X1 U21873 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18665) );
  AOI22_X1 U21874 ( .A1(n18675), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18664) );
  OAI21_X1 U21875 ( .B1(n18665), .B2(n18677), .A(n18664), .ZN(P3_U2762) );
  INV_X1 U21876 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18667) );
  AOI22_X1 U21877 ( .A1(n18675), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18666) );
  OAI21_X1 U21878 ( .B1(n18667), .B2(n18677), .A(n18666), .ZN(P3_U2763) );
  AOI22_X1 U21879 ( .A1(n18675), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18668) );
  OAI21_X1 U21880 ( .B1(n18669), .B2(n18677), .A(n18668), .ZN(P3_U2764) );
  INV_X1 U21881 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18671) );
  AOI22_X1 U21882 ( .A1(n18675), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18670) );
  OAI21_X1 U21883 ( .B1(n18671), .B2(n18677), .A(n18670), .ZN(P3_U2765) );
  AOI22_X1 U21884 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n18672), .B1(n18661), .B2(
        P3_DATAO_REG_1__SCAN_IN), .ZN(n18673) );
  OAI21_X1 U21885 ( .B1(n18702), .B2(n18674), .A(n18673), .ZN(P3_U2766) );
  AOI22_X1 U21886 ( .A1(n18675), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18661), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18676) );
  OAI21_X1 U21887 ( .B1(n18678), .B2(n18677), .A(n18676), .ZN(P3_U2767) );
  INV_X1 U21888 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19422) );
  AOI22_X1 U21889 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18726), .ZN(n18681) );
  OAI21_X1 U21890 ( .B1(n19422), .B2(n18720), .A(n18681), .ZN(P3_U2768) );
  AOI22_X1 U21891 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18727), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18726), .ZN(n18682) );
  OAI21_X1 U21892 ( .B1(n18683), .B2(n18729), .A(n18682), .ZN(P3_U2769) );
  AOI22_X1 U21893 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18726), .ZN(n18684) );
  OAI21_X1 U21894 ( .B1(n19433), .B2(n18720), .A(n18684), .ZN(P3_U2770) );
  AOI22_X1 U21895 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18726), .ZN(n18685) );
  OAI21_X1 U21896 ( .B1(n19437), .B2(n18720), .A(n18685), .ZN(P3_U2771) );
  AOI22_X1 U21897 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18726), .ZN(n18686) );
  OAI21_X1 U21898 ( .B1(n19441), .B2(n18720), .A(n18686), .ZN(P3_U2772) );
  AOI22_X1 U21899 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18726), .ZN(n18687) );
  OAI21_X1 U21900 ( .B1(n19445), .B2(n18720), .A(n18687), .ZN(P3_U2773) );
  AOI22_X1 U21901 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18726), .ZN(n18688) );
  OAI21_X1 U21902 ( .B1(n13757), .B2(n18720), .A(n18688), .ZN(P3_U2774) );
  AOI22_X1 U21903 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18726), .ZN(n18689) );
  OAI21_X1 U21904 ( .B1(n19452), .B2(n18720), .A(n18689), .ZN(P3_U2775) );
  AOI22_X1 U21905 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18727), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18726), .ZN(n18690) );
  OAI21_X1 U21906 ( .B1(n18691), .B2(n18729), .A(n18690), .ZN(P3_U2776) );
  AOI22_X1 U21907 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18726), .ZN(n18692) );
  OAI21_X1 U21908 ( .B1(n18713), .B2(n18720), .A(n18692), .ZN(P3_U2777) );
  INV_X1 U21909 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18715) );
  AOI22_X1 U21910 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18726), .ZN(n18693) );
  OAI21_X1 U21911 ( .B1(n18715), .B2(n18720), .A(n18693), .ZN(P3_U2778) );
  AOI22_X1 U21912 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18726), .ZN(n18694) );
  OAI21_X1 U21913 ( .B1(n18717), .B2(n18720), .A(n18694), .ZN(P3_U2779) );
  AOI22_X1 U21914 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18718), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18726), .ZN(n18695) );
  OAI21_X1 U21915 ( .B1(n18721), .B2(n18720), .A(n18695), .ZN(P3_U2780) );
  AOI22_X1 U21916 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18727), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18726), .ZN(n18696) );
  OAI21_X1 U21917 ( .B1(n18697), .B2(n18729), .A(n18696), .ZN(P3_U2781) );
  AOI22_X1 U21918 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18727), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18726), .ZN(n18698) );
  OAI21_X1 U21919 ( .B1(n18699), .B2(n18729), .A(n18698), .ZN(P3_U2782) );
  AOI22_X1 U21920 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18726), .ZN(n18700) );
  OAI21_X1 U21921 ( .B1(n19422), .B2(n18720), .A(n18700), .ZN(P3_U2783) );
  AOI22_X1 U21922 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18727), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n18718), .ZN(n18701) );
  OAI21_X1 U21923 ( .B1(n18703), .B2(n18702), .A(n18701), .ZN(P3_U2784) );
  AOI22_X1 U21924 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18726), .ZN(n18704) );
  OAI21_X1 U21925 ( .B1(n19433), .B2(n18720), .A(n18704), .ZN(P3_U2785) );
  AOI22_X1 U21926 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18726), .ZN(n18705) );
  OAI21_X1 U21927 ( .B1(n19437), .B2(n18720), .A(n18705), .ZN(P3_U2786) );
  AOI22_X1 U21928 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18726), .ZN(n18706) );
  OAI21_X1 U21929 ( .B1(n19441), .B2(n18720), .A(n18706), .ZN(P3_U2787) );
  AOI22_X1 U21930 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18726), .ZN(n18707) );
  OAI21_X1 U21931 ( .B1(n19445), .B2(n18720), .A(n18707), .ZN(P3_U2788) );
  AOI22_X1 U21932 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18726), .ZN(n18708) );
  OAI21_X1 U21933 ( .B1(n13757), .B2(n18720), .A(n18708), .ZN(P3_U2789) );
  AOI22_X1 U21934 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18726), .ZN(n18709) );
  OAI21_X1 U21935 ( .B1(n19452), .B2(n18720), .A(n18709), .ZN(P3_U2790) );
  AOI22_X1 U21936 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18727), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18726), .ZN(n18710) );
  OAI21_X1 U21937 ( .B1(n18711), .B2(n18729), .A(n18710), .ZN(P3_U2791) );
  AOI22_X1 U21938 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18726), .ZN(n18712) );
  OAI21_X1 U21939 ( .B1(n18713), .B2(n18720), .A(n18712), .ZN(P3_U2792) );
  AOI22_X1 U21940 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18726), .ZN(n18714) );
  OAI21_X1 U21941 ( .B1(n18715), .B2(n18720), .A(n18714), .ZN(P3_U2793) );
  AOI22_X1 U21942 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18726), .ZN(n18716) );
  OAI21_X1 U21943 ( .B1(n18717), .B2(n18720), .A(n18716), .ZN(P3_U2794) );
  AOI22_X1 U21944 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18718), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18726), .ZN(n18719) );
  OAI21_X1 U21945 ( .B1(n18721), .B2(n18720), .A(n18719), .ZN(P3_U2795) );
  AOI22_X1 U21946 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18727), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18726), .ZN(n18722) );
  OAI21_X1 U21947 ( .B1(n18723), .B2(n18729), .A(n18722), .ZN(P3_U2796) );
  AOI22_X1 U21948 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18727), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18726), .ZN(n18724) );
  OAI21_X1 U21949 ( .B1(n18725), .B2(n18729), .A(n18724), .ZN(P3_U2797) );
  AOI22_X1 U21950 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18727), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18726), .ZN(n18728) );
  OAI21_X1 U21951 ( .B1(n18730), .B2(n18729), .A(n18728), .ZN(P3_U2798) );
  NOR4_X1 U21952 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18942), .A3(
        n18732), .A4(n18731), .ZN(n18734) );
  AOI211_X1 U21953 ( .C1(n18935), .C2(n18735), .A(n18734), .B(n18733), .ZN(
        n18750) );
  OAI211_X1 U21954 ( .C1(n18738), .C2(n18737), .A(n18736), .B(n19011), .ZN(
        n18743) );
  INV_X1 U21955 ( .A(n18739), .ZN(n18741) );
  NAND3_X1 U21956 ( .A1(n18902), .A2(n18741), .A3(n18740), .ZN(n18742) );
  AND2_X1 U21957 ( .A1(n18743), .A2(n18742), .ZN(n18749) );
  NAND2_X1 U21958 ( .A1(n19100), .A2(n19009), .ZN(n18841) );
  AOI22_X1 U21959 ( .A1(n19088), .A2(n19105), .B1(n18970), .B2(n19104), .ZN(
        n18773) );
  NAND2_X1 U21960 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18773), .ZN(
        n18760) );
  NAND3_X1 U21961 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18841), .A3(
        n18760), .ZN(n18748) );
  NOR3_X1 U21962 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18942), .A3(
        n18731), .ZN(n18758) );
  OAI21_X1 U21963 ( .B1(n18745), .B2(n19095), .A(n19096), .ZN(n18746) );
  AOI21_X1 U21964 ( .B1(n19004), .B2(n18731), .A(n18746), .ZN(n18766) );
  OAI21_X1 U21965 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18880), .A(
        n18766), .ZN(n18759) );
  OAI21_X1 U21966 ( .B1(n18758), .B2(n18759), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18747) );
  NAND4_X1 U21967 ( .A1(n18750), .A2(n18749), .A3(n18748), .A4(n18747), .ZN(
        P3_U2802) );
  NAND2_X1 U21968 ( .A1(n18751), .A2(n18752), .ZN(n18753) );
  MUX2_X1 U21969 ( .A(n18753), .B(n18752), .S(n18890), .Z(n18755) );
  NAND2_X1 U21970 ( .A1(n18755), .A2(n18754), .ZN(n19113) );
  OAI22_X1 U21971 ( .A1(n19400), .A2(n19987), .B1(n18962), .B2(n18756), .ZN(
        n18757) );
  AOI211_X1 U21972 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n18759), .A(
        n18758), .B(n18757), .ZN(n18763) );
  INV_X1 U21973 ( .A(n18902), .ZN(n18836) );
  NOR2_X1 U21974 ( .A1(n19101), .A2(n18836), .ZN(n18761) );
  OAI21_X1 U21975 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18761), .A(
        n18760), .ZN(n18762) );
  OAI211_X1 U21976 ( .C1(n19113), .C2(n18991), .A(n18763), .B(n18762), .ZN(
        P3_U2803) );
  AOI21_X1 U21977 ( .B1(n19801), .B2(n18764), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18765) );
  INV_X1 U21978 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19985) );
  OAI22_X1 U21979 ( .A1(n18766), .A2(n18765), .B1(n19400), .B2(n19985), .ZN(
        n18767) );
  AOI221_X1 U21980 ( .B1(n18935), .B2(n18768), .C1(n9612), .C2(n18768), .A(
        n18767), .ZN(n18772) );
  XNOR2_X1 U21981 ( .A(n18769), .B(n19110), .ZN(n19114) );
  NOR2_X1 U21982 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18770), .ZN(
        n19115) );
  AOI22_X1 U21983 ( .A1(n19114), .A2(n19011), .B1(n18902), .B2(n19115), .ZN(
        n18771) );
  OAI211_X1 U21984 ( .C1(n18773), .C2(n19110), .A(n18772), .B(n18771), .ZN(
        P3_U2804) );
  NAND2_X1 U21985 ( .A1(n19157), .A2(n19125), .ZN(n18774) );
  XOR2_X1 U21986 ( .A(n18774), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n19128) );
  OAI21_X1 U21987 ( .B1(n18802), .B2(n19095), .A(n19096), .ZN(n18775) );
  AOI21_X1 U21988 ( .B1(n19801), .B2(n13007), .A(n18775), .ZN(n18800) );
  OAI21_X1 U21989 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18880), .A(
        n18800), .ZN(n18789) );
  NOR2_X1 U21990 ( .A1(n18942), .A2(n13007), .ZN(n18791) );
  OAI211_X1 U21991 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18791), .B(n18776), .ZN(n18777) );
  NAND2_X1 U21992 ( .A1(n19402), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n19133) );
  OAI211_X1 U21993 ( .C1(n18962), .C2(n18778), .A(n18777), .B(n19133), .ZN(
        n18785) );
  NAND2_X1 U21994 ( .A1(n19125), .A2(n19158), .ZN(n18779) );
  XOR2_X1 U21995 ( .A(n18779), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n19130) );
  INV_X1 U21996 ( .A(n18780), .ZN(n18782) );
  NOR2_X1 U21997 ( .A1(n18782), .A2(n18781), .ZN(n18783) );
  XNOR2_X1 U21998 ( .A(n18783), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19129) );
  OAI22_X1 U21999 ( .A1(n19100), .A2(n19130), .B1(n18991), .B2(n19129), .ZN(
        n18784) );
  AOI211_X1 U22000 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18789), .A(
        n18785), .B(n18784), .ZN(n18786) );
  OAI21_X1 U22001 ( .B1(n19009), .B2(n19128), .A(n18786), .ZN(P3_U2805) );
  OR2_X1 U22002 ( .A1(n18792), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n19149) );
  INV_X1 U22003 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19980) );
  OAI22_X1 U22004 ( .A1(n19400), .A2(n19980), .B1(n18962), .B2(n18787), .ZN(
        n18788) );
  AOI221_X1 U22005 ( .B1(n18791), .B2(n18790), .C1(n18789), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18788), .ZN(n18796) );
  INV_X1 U22006 ( .A(n19158), .ZN(n19235) );
  NOR2_X1 U22007 ( .A1(n19235), .A2(n18792), .ZN(n19140) );
  INV_X1 U22008 ( .A(n19157), .ZN(n19234) );
  NOR2_X1 U22009 ( .A1(n18792), .A2(n19234), .ZN(n19136) );
  OAI22_X1 U22010 ( .A1(n19140), .A2(n19100), .B1(n19136), .B2(n19009), .ZN(
        n18808) );
  OAI21_X1 U22011 ( .B1(n9754), .B2(n18794), .A(n18793), .ZN(n19135) );
  AOI22_X1 U22012 ( .A1(n18808), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19011), .B2(n19135), .ZN(n18795) );
  OAI211_X1 U22013 ( .C1(n18836), .C2(n19149), .A(n18796), .B(n18795), .ZN(
        P3_U2806) );
  NOR2_X1 U22014 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18880), .ZN(
        n18803) );
  AOI21_X1 U22015 ( .B1(n18797), .B2(n19801), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18799) );
  OAI22_X1 U22016 ( .A1(n18800), .A2(n18799), .B1(n18962), .B2(n18798), .ZN(
        n18801) );
  AOI21_X1 U22017 ( .B1(n18803), .B2(n18802), .A(n18801), .ZN(n18811) );
  NAND2_X1 U22018 ( .A1(n19006), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18805) );
  OAI211_X1 U22019 ( .C1(n18806), .C2(n18816), .A(n18848), .B(n18805), .ZN(
        n18807) );
  XNOR2_X1 U22020 ( .A(n18807), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19150) );
  AOI22_X1 U22021 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18808), .B1(
        n19011), .B2(n19150), .ZN(n18810) );
  NAND3_X1 U22022 ( .A1(n19121), .A2(n18902), .A3(n19141), .ZN(n18809) );
  NAND2_X1 U22023 ( .A1(n19402), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n19155) );
  NAND4_X1 U22024 ( .A1(n18811), .A2(n18810), .A3(n18809), .A4(n19155), .ZN(
        P3_U2807) );
  OAI21_X1 U22025 ( .B1(n18813), .B2(n19095), .A(n19096), .ZN(n18814) );
  AOI21_X1 U22026 ( .B1(n19004), .B2(n18812), .A(n18814), .ZN(n18844) );
  OAI21_X1 U22027 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18880), .A(
        n18844), .ZN(n18828) );
  AOI22_X1 U22028 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18828), .B1(
        n18935), .B2(n18815), .ZN(n18825) );
  AND3_X1 U22029 ( .A1(n18873), .A2(n19165), .A3(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18817) );
  OAI21_X1 U22030 ( .B1(n18817), .B2(n18816), .A(n18848), .ZN(n18818) );
  XNOR2_X1 U22031 ( .A(n18818), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19170) );
  NOR2_X1 U22032 ( .A1(n19168), .A2(n18836), .ZN(n18820) );
  OAI22_X1 U22033 ( .A1(n19158), .A2(n19100), .B1(n19157), .B2(n19009), .ZN(
        n18901) );
  AOI21_X1 U22034 ( .B1(n19168), .B2(n18841), .A(n18901), .ZN(n18840) );
  INV_X1 U22035 ( .A(n18840), .ZN(n18819) );
  MUX2_X1 U22036 ( .A(n18820), .B(n18819), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18821) );
  AOI21_X1 U22037 ( .B1(n19011), .B2(n19170), .A(n18821), .ZN(n18824) );
  NAND2_X1 U22038 ( .A1(n19402), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19172) );
  NOR2_X1 U22039 ( .A1(n18942), .A2(n18812), .ZN(n18830) );
  OAI211_X1 U22040 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18830), .B(n18822), .ZN(n18823) );
  NAND4_X1 U22041 ( .A1(n18825), .A2(n18824), .A3(n19172), .A4(n18823), .ZN(
        P3_U2808) );
  INV_X1 U22042 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18829) );
  OAI22_X1 U22043 ( .A1(n19400), .A2(n19974), .B1(n18962), .B2(n18826), .ZN(
        n18827) );
  AOI221_X1 U22044 ( .B1(n18830), .B2(n18829), .C1(n18828), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18827), .ZN(n18838) );
  INV_X1 U22045 ( .A(n18891), .ZN(n18832) );
  INV_X1 U22046 ( .A(n18831), .ZN(n19202) );
  NAND2_X1 U22047 ( .A1(n18890), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18872) );
  NOR3_X1 U22048 ( .A1(n18832), .A2(n19202), .A3(n18872), .ZN(n18849) );
  INV_X1 U22049 ( .A(n18849), .ZN(n18859) );
  OAI22_X1 U22050 ( .A1(n18859), .A2(n18835), .B1(n18833), .B2(n18873), .ZN(
        n18834) );
  XOR2_X1 U22051 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18834), .Z(
        n19182) );
  NOR2_X1 U22052 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18835), .ZN(
        n19181) );
  NOR2_X1 U22053 ( .A1(n19164), .A2(n18836), .ZN(n18861) );
  AOI22_X1 U22054 ( .A1(n19011), .A2(n19182), .B1(n19181), .B2(n18861), .ZN(
        n18837) );
  OAI211_X1 U22055 ( .C1(n18840), .C2(n18839), .A(n18838), .B(n18837), .ZN(
        P3_U2809) );
  NAND2_X1 U22056 ( .A1(n19179), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n19190) );
  AOI21_X1 U22057 ( .B1(n18841), .B2(n19190), .A(n18901), .ZN(n18865) );
  AOI21_X1 U22058 ( .B1(n19801), .B2(n18842), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18843) );
  OAI22_X1 U22059 ( .A1(n18844), .A2(n18843), .B1(n19400), .B2(n19972), .ZN(
        n18845) );
  AOI221_X1 U22060 ( .B1(n18935), .B2(n18846), .C1(n9612), .C2(n18846), .A(
        n18845), .ZN(n18852) );
  NAND2_X1 U22061 ( .A1(n18871), .A2(n18864), .ZN(n18847) );
  OAI211_X1 U22062 ( .C1(n18849), .C2(n18864), .A(n18848), .B(n18847), .ZN(
        n18850) );
  XNOR2_X1 U22063 ( .A(n18850), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n19187) );
  NOR2_X1 U22064 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19190), .ZN(
        n19185) );
  AOI22_X1 U22065 ( .A1(n19011), .A2(n19187), .B1(n18902), .B2(n19185), .ZN(
        n18851) );
  OAI211_X1 U22066 ( .C1(n18865), .C2(n19162), .A(n18852), .B(n18851), .ZN(
        P3_U2810) );
  AOI21_X1 U22067 ( .B1(n19004), .B2(n18854), .A(n19083), .ZN(n18887) );
  OAI21_X1 U22068 ( .B1(n18853), .B2(n19095), .A(n18887), .ZN(n18868) );
  NOR2_X1 U22069 ( .A1(n18942), .A2(n18854), .ZN(n18870) );
  OAI211_X1 U22070 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18870), .B(n18855), .ZN(n18856) );
  NAND2_X1 U22071 ( .A1(n19402), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19198) );
  OAI211_X1 U22072 ( .C1(n18962), .C2(n18857), .A(n18856), .B(n19198), .ZN(
        n18858) );
  AOI21_X1 U22073 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18868), .A(
        n18858), .ZN(n18863) );
  OAI21_X1 U22074 ( .B1(n18873), .B2(n18871), .A(n18859), .ZN(n18860) );
  XOR2_X1 U22075 ( .A(n18860), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n19196) );
  AOI22_X1 U22076 ( .A1(n19011), .A2(n19196), .B1(n18861), .B2(n18864), .ZN(
        n18862) );
  OAI211_X1 U22077 ( .C1(n18865), .C2(n18864), .A(n18863), .B(n18862), .ZN(
        P3_U2811) );
  AOI21_X1 U22078 ( .B1(n18902), .B2(n19202), .A(n18901), .ZN(n18882) );
  OAI22_X1 U22079 ( .A1(n19400), .A2(n19968), .B1(n18962), .B2(n18866), .ZN(
        n18867) );
  AOI221_X1 U22080 ( .B1(n18870), .B2(n18869), .C1(n18868), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18867), .ZN(n18876) );
  NAND2_X1 U22081 ( .A1(n18872), .A2(n18871), .ZN(n18874) );
  XOR2_X1 U22082 ( .A(n18874), .B(n18873), .Z(n19212) );
  NOR2_X1 U22083 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n19202), .ZN(
        n19211) );
  AOI22_X1 U22084 ( .A1(n19011), .A2(n19212), .B1(n18902), .B2(n19211), .ZN(
        n18875) );
  OAI211_X1 U22085 ( .C1(n18882), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P3_U2812) );
  AOI21_X1 U22086 ( .B1(n18878), .B2(n19801), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18888) );
  XNOR2_X1 U22087 ( .A(n18879), .B(n19217), .ZN(n19215) );
  OR2_X2 U22088 ( .A1(n18935), .A2(n9612), .ZN(n19089) );
  AOI21_X1 U22089 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18902), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18881) );
  OAI22_X1 U22090 ( .A1(n19080), .A2(n18883), .B1(n18882), .B2(n18881), .ZN(
        n18884) );
  AOI21_X1 U22091 ( .B1(n19011), .B2(n19215), .A(n18884), .ZN(n18886) );
  NAND2_X1 U22092 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n19402), .ZN(n18885) );
  OAI211_X1 U22093 ( .C1(n18888), .C2(n18887), .A(n18886), .B(n18885), .ZN(
        P3_U2813) );
  NOR2_X1 U22094 ( .A1(n19006), .A2(n10273), .ZN(n18889) );
  NAND2_X1 U22095 ( .A1(n18905), .A2(n18889), .ZN(n18993) );
  OAI22_X1 U22096 ( .A1(n18891), .A2(n18890), .B1(n18993), .B2(n19210), .ZN(
        n18892) );
  XOR2_X1 U22097 ( .A(n19228), .B(n18892), .Z(n19233) );
  AOI21_X1 U22098 ( .B1(n18896), .B2(n19004), .A(n19083), .ZN(n18893) );
  INV_X1 U22099 ( .A(n18893), .ZN(n18920) );
  AOI21_X1 U22100 ( .B1(n18932), .B2(n18894), .A(n18920), .ZN(n18913) );
  AOI22_X1 U22101 ( .A1(n19402), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18935), 
        .B2(n18895), .ZN(n18898) );
  NOR2_X1 U22102 ( .A1(n18942), .A2(n18896), .ZN(n18909) );
  OAI221_X1 U22103 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C1(n18899), .C2(n18912), .A(
        n18909), .ZN(n18897) );
  OAI211_X1 U22104 ( .C1(n18913), .C2(n18899), .A(n18898), .B(n18897), .ZN(
        n18900) );
  AOI221_X1 U22105 ( .B1(n18902), .B2(n19228), .C1(n18901), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n18900), .ZN(n18903) );
  OAI21_X1 U22106 ( .B1(n19233), .B2(n18991), .A(n18903), .ZN(P3_U2814) );
  AND2_X1 U22107 ( .A1(n18918), .A2(n17304), .ZN(n19240) );
  NAND2_X1 U22108 ( .A1(n19088), .A2(n19235), .ZN(n18917) );
  NOR3_X1 U22109 ( .A1(n19280), .A2(n18927), .A3(n10273), .ZN(n18904) );
  AOI21_X1 U22110 ( .B1(n18905), .B2(n18904), .A(n18939), .ZN(n18907) );
  MUX2_X1 U22111 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n19006), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18906) );
  AOI211_X1 U22112 ( .C1(n18973), .C2(n18939), .A(n18907), .B(n18906), .ZN(
        n18908) );
  XNOR2_X1 U22113 ( .A(n18908), .B(n17304), .ZN(n19244) );
  NOR2_X1 U22114 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18924), .ZN(
        n19242) );
  NOR3_X1 U22115 ( .A1(n19157), .A2(n19242), .A3(n19009), .ZN(n18915) );
  AOI22_X1 U22116 ( .A1(n18910), .A2(n18935), .B1(n18909), .B2(n18912), .ZN(
        n18911) );
  NAND2_X1 U22117 ( .A1(n19402), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n19246) );
  OAI211_X1 U22118 ( .C1(n18913), .C2(n18912), .A(n18911), .B(n19246), .ZN(
        n18914) );
  AOI211_X1 U22119 ( .C1(n19244), .C2(n19011), .A(n18915), .B(n18914), .ZN(
        n18916) );
  OAI21_X1 U22120 ( .B1(n19240), .B2(n18917), .A(n18916), .ZN(P3_U2815) );
  OAI21_X1 U22121 ( .B1(n18919), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18918), .ZN(n19262) );
  OAI221_X1 U22122 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17954), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19801), .A(n18920), .ZN(
        n18921) );
  OAI21_X1 U22123 ( .B1(n19080), .B2(n18922), .A(n18921), .ZN(n18923) );
  AOI21_X1 U22124 ( .B1(n19402), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18923), 
        .ZN(n18930) );
  AOI221_X1 U22125 ( .B1(n18969), .B2(n18927), .C1(n19249), .C2(n18927), .A(
        n18924), .ZN(n19258) );
  NOR2_X1 U22126 ( .A1(n18993), .A2(n17301), .ZN(n18978) );
  AND2_X1 U22127 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18925) );
  AND2_X1 U22128 ( .A1(n18978), .A2(n18925), .ZN(n18951) );
  NAND2_X1 U22129 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18951), .ZN(
        n18938) );
  INV_X1 U22130 ( .A(n18952), .ZN(n18926) );
  NAND2_X1 U22131 ( .A1(n18926), .A2(n18939), .ZN(n18937) );
  OAI21_X1 U22132 ( .B1(n18938), .B2(n18939), .A(n18937), .ZN(n18928) );
  XNOR2_X1 U22133 ( .A(n18928), .B(n18927), .ZN(n19257) );
  AOI22_X1 U22134 ( .A1(n18970), .A2(n19258), .B1(n19011), .B2(n19257), .ZN(
        n18929) );
  OAI211_X1 U22135 ( .C1(n19100), .C2(n19262), .A(n18930), .B(n18929), .ZN(
        P3_U2816) );
  AOI22_X1 U22136 ( .A1(n18932), .A2(n18931), .B1(n19004), .B2(n18941), .ZN(
        n18933) );
  NAND2_X1 U22137 ( .A1(n18933), .A2(n19096), .ZN(n18948) );
  AOI22_X1 U22138 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18948), .B1(
        n18935), .B2(n18934), .ZN(n18947) );
  NAND3_X1 U22139 ( .A1(n18952), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n18938), .ZN(n18936) );
  OAI211_X1 U22140 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18938), .A(
        n18937), .B(n18936), .ZN(n19263) );
  NAND2_X1 U22141 ( .A1(n19251), .A2(n18939), .ZN(n19273) );
  NAND2_X1 U22142 ( .A1(n19251), .A2(n19291), .ZN(n19264) );
  AOI22_X1 U22143 ( .A1(n19088), .A2(n19266), .B1(n18970), .B2(n19264), .ZN(
        n18955) );
  OAI22_X1 U22144 ( .A1(n19003), .A2(n19273), .B1(n18955), .B2(n18939), .ZN(
        n18940) );
  AOI21_X1 U22145 ( .B1(n19011), .B2(n19263), .A(n18940), .ZN(n18946) );
  NAND2_X1 U22146 ( .A1(n19402), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18945) );
  NOR2_X1 U22147 ( .A1(n18942), .A2(n18941), .ZN(n18950) );
  OAI211_X1 U22148 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18950), .B(n18943), .ZN(n18944) );
  NAND4_X1 U22149 ( .A1(n18947), .A2(n18946), .A3(n18945), .A4(n18944), .ZN(
        P3_U2817) );
  INV_X1 U22150 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18949) );
  NOR2_X1 U22151 ( .A1(n19400), .A2(n19956), .ZN(n19284) );
  AOI221_X1 U22152 ( .B1(n18950), .B2(n18949), .C1(n18948), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n19284), .ZN(n18960) );
  INV_X1 U22153 ( .A(n18951), .ZN(n18954) );
  NAND3_X1 U22154 ( .A1(n18954), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n18973), .ZN(n18953) );
  OAI211_X1 U22155 ( .C1(n18954), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18953), .B(n18952), .ZN(n19282) );
  NOR2_X1 U22156 ( .A1(n19003), .A2(n19280), .ZN(n18957) );
  INV_X1 U22157 ( .A(n18955), .ZN(n18956) );
  MUX2_X1 U22158 ( .A(n18957), .B(n18956), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n18958) );
  AOI21_X1 U22159 ( .B1(n19011), .B2(n19282), .A(n18958), .ZN(n18959) );
  OAI211_X1 U22160 ( .C1(n18962), .C2(n18961), .A(n18960), .B(n18959), .ZN(
        P3_U2818) );
  NAND2_X1 U22161 ( .A1(n18972), .A2(n17303), .ZN(n19302) );
  INV_X1 U22162 ( .A(n19027), .ZN(n19090) );
  AND2_X1 U22163 ( .A1(n19801), .A2(n18963), .ZN(n19032) );
  NAND2_X1 U22164 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19032), .ZN(
        n19024) );
  NOR2_X1 U22165 ( .A1(n19012), .A2(n19024), .ZN(n18995) );
  NAND2_X1 U22166 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18995), .ZN(
        n18983) );
  INV_X1 U22167 ( .A(n18983), .ZN(n18998) );
  NAND2_X1 U22168 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18998), .ZN(
        n18986) );
  INV_X1 U22169 ( .A(n18986), .ZN(n18966) );
  NOR2_X1 U22170 ( .A1(n18967), .A2(n18966), .ZN(n18968) );
  OAI22_X1 U22171 ( .A1(n19080), .A2(n18964), .B1(n19400), .B2(n19954), .ZN(
        n18965) );
  AOI221_X1 U22172 ( .B1(n19090), .B2(n18968), .C1(n18967), .C2(n18966), .A(
        n18965), .ZN(n18977) );
  AOI22_X1 U22173 ( .A1(n19088), .A2(n18971), .B1(n18970), .B2(n18969), .ZN(
        n19002) );
  OAI21_X1 U22174 ( .B1(n18972), .B2(n19003), .A(n19002), .ZN(n18988) );
  NAND2_X1 U22175 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18978), .ZN(
        n18975) );
  NAND3_X1 U22176 ( .A1(n9768), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18975), .ZN(n18974) );
  OAI211_X1 U22177 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n18975), .A(
        n18974), .B(n18973), .ZN(n19288) );
  AOI22_X1 U22178 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18988), .B1(
        n19011), .B2(n19288), .ZN(n18976) );
  OAI211_X1 U22179 ( .C1(n19003), .C2(n19302), .A(n18977), .B(n18976), .ZN(
        P3_U2819) );
  INV_X1 U22180 ( .A(n18978), .ZN(n18980) );
  NAND2_X1 U22181 ( .A1(n18980), .A2(n18979), .ZN(n18981) );
  XNOR2_X1 U22182 ( .A(n18981), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19311) );
  AOI22_X1 U22183 ( .A1(n19402), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18982), 
        .B2(n19089), .ZN(n18990) );
  OAI21_X1 U22184 ( .B1(n19003), .B2(n17301), .A(n10282), .ZN(n18987) );
  OAI21_X1 U22185 ( .B1(n19027), .B2(n18984), .A(n18983), .ZN(n18985) );
  AOI22_X1 U22186 ( .A1(n18988), .A2(n18987), .B1(n18986), .B2(n18985), .ZN(
        n18989) );
  OAI211_X1 U22187 ( .C1(n19311), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P3_U2820) );
  NAND2_X1 U22188 ( .A1(n18993), .A2(n18992), .ZN(n18994) );
  XOR2_X1 U22189 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18994), .Z(
        n19317) );
  NOR2_X1 U22190 ( .A1(n19400), .A2(n19950), .ZN(n19000) );
  AOI21_X1 U22191 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19090), .A(
        n18995), .ZN(n18997) );
  OAI22_X1 U22192 ( .A1(n18998), .A2(n18997), .B1(n19080), .B2(n18996), .ZN(
        n18999) );
  AOI211_X1 U22193 ( .C1(n19011), .C2(n19317), .A(n19000), .B(n18999), .ZN(
        n19001) );
  OAI221_X1 U22194 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19003), .C1(
        n17301), .C2(n19002), .A(n19001), .ZN(P3_U2821) );
  INV_X1 U22195 ( .A(n19004), .ZN(n19056) );
  OAI21_X1 U22196 ( .B1(n18052), .B2(n19056), .A(n19096), .ZN(n19017) );
  AOI22_X1 U22197 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19017), .B1(
        n19005), .B2(n19089), .ZN(n19016) );
  XNOR2_X1 U22198 ( .A(n19322), .B(n19006), .ZN(n19325) );
  OAI21_X1 U22199 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n19008), .A(
        n19007), .ZN(n19323) );
  OAI22_X1 U22200 ( .A1(n19323), .A2(n19100), .B1(n19322), .B2(n19009), .ZN(
        n19010) );
  AOI21_X1 U22201 ( .B1(n19011), .B2(n19325), .A(n19010), .ZN(n19015) );
  NAND2_X1 U22202 ( .A1(n19402), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19331) );
  AND2_X1 U22203 ( .A1(n18052), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19013) );
  OAI211_X1 U22204 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n19013), .A(
        n19801), .B(n19012), .ZN(n19014) );
  NAND4_X1 U22205 ( .A1(n19016), .A2(n19015), .A3(n19331), .A4(n19014), .ZN(
        P3_U2822) );
  AOI22_X1 U22206 ( .A1(n19402), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19017), .ZN(n19023) );
  OAI22_X1 U22207 ( .A1(n19080), .A2(n19019), .B1(n19018), .B2(n19099), .ZN(
        n19020) );
  AOI21_X1 U22208 ( .B1(n19088), .B2(n19021), .A(n19020), .ZN(n19022) );
  OAI211_X1 U22209 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19024), .A(
        n19023), .B(n19022), .ZN(P3_U2823) );
  OAI21_X1 U22210 ( .B1(n19026), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n19025), .ZN(n19335) );
  NOR2_X1 U22211 ( .A1(n19027), .A2(n19032), .ZN(n19046) );
  XNOR2_X1 U22212 ( .A(n19029), .B(n19028), .ZN(n19334) );
  OAI22_X1 U22213 ( .A1(n19099), .A2(n19334), .B1(n19944), .B2(n19400), .ZN(
        n19030) );
  AOI221_X1 U22214 ( .B1(n19046), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C1(
        n19032), .C2(n19031), .A(n19030), .ZN(n19035) );
  NAND2_X1 U22215 ( .A1(n19033), .A2(n19089), .ZN(n19034) );
  OAI211_X1 U22216 ( .C1(n19335), .C2(n19100), .A(n19035), .B(n19034), .ZN(
        P3_U2824) );
  OAI21_X1 U22217 ( .B1(n19083), .B2(n19039), .A(n19038), .ZN(n19045) );
  XNOR2_X1 U22218 ( .A(n19040), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19041) );
  XNOR2_X1 U22219 ( .A(n19042), .B(n19041), .ZN(n19341) );
  OAI22_X1 U22220 ( .A1(n19080), .A2(n19043), .B1(n19099), .B2(n19341), .ZN(
        n19044) );
  AOI21_X1 U22221 ( .B1(n19046), .B2(n19045), .A(n19044), .ZN(n19048) );
  INV_X1 U22222 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19943) );
  NOR2_X1 U22223 ( .A1(n19400), .A2(n19943), .ZN(n19344) );
  INV_X1 U22224 ( .A(n19344), .ZN(n19047) );
  OAI211_X1 U22225 ( .C1(n19100), .C2(n19342), .A(n19048), .B(n19047), .ZN(
        P3_U2825) );
  OAI21_X1 U22226 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19050), .A(
        n19049), .ZN(n19358) );
  OAI22_X1 U22227 ( .A1(n19400), .A2(n19940), .B1(n19479), .B2(n19051), .ZN(
        n19052) );
  INV_X1 U22228 ( .A(n19052), .ZN(n19062) );
  XNOR2_X1 U22229 ( .A(n19053), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19054) );
  XNOR2_X1 U22230 ( .A(n19055), .B(n19054), .ZN(n19351) );
  OAI21_X1 U22231 ( .B1(n19056), .B2(n18133), .A(n19096), .ZN(n19071) );
  INV_X1 U22232 ( .A(n19071), .ZN(n19057) );
  OAI22_X1 U22233 ( .A1(n19099), .A2(n19351), .B1(n19058), .B2(n19057), .ZN(
        n19059) );
  AOI21_X1 U22234 ( .B1(n19060), .B2(n19089), .A(n19059), .ZN(n19061) );
  OAI211_X1 U22235 ( .C1(n19100), .C2(n19358), .A(n19062), .B(n19061), .ZN(
        P3_U2826) );
  OAI21_X1 U22236 ( .B1(n19065), .B2(n19064), .A(n19063), .ZN(n19361) );
  NOR2_X1 U22237 ( .A1(n19083), .A2(n19082), .ZN(n19070) );
  XNOR2_X1 U22238 ( .A(n19067), .B(n19066), .ZN(n19360) );
  OAI22_X1 U22239 ( .A1(n19080), .A2(n19068), .B1(n19099), .B2(n19360), .ZN(
        n19069) );
  AOI221_X1 U22240 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19071), .C1(
        n19070), .C2(n19071), .A(n19069), .ZN(n19072) );
  NAND2_X1 U22241 ( .A1(n19402), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19365) );
  OAI211_X1 U22242 ( .C1(n19100), .C2(n19361), .A(n19072), .B(n19365), .ZN(
        P3_U2827) );
  OR2_X1 U22243 ( .A1(n19074), .A2(n19073), .ZN(n19076) );
  NAND2_X1 U22244 ( .A1(n19076), .A2(n19075), .ZN(n19378) );
  XNOR2_X1 U22245 ( .A(n19078), .B(n19077), .ZN(n19377) );
  OAI22_X1 U22246 ( .A1(n19080), .A2(n19079), .B1(n19377), .B2(n19099), .ZN(
        n19081) );
  AOI221_X1 U22247 ( .B1(n19083), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19801), .C2(n19082), .A(n19081), .ZN(n19084) );
  NAND2_X1 U22248 ( .A1(n19402), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19383) );
  OAI211_X1 U22249 ( .C1(n19100), .C2(n19378), .A(n19084), .B(n19383), .ZN(
        P3_U2828) );
  OAI21_X1 U22250 ( .B1(n19086), .B2(n19093), .A(n19085), .ZN(n19395) );
  NAND2_X1 U22251 ( .A1(n19396), .A2(n19094), .ZN(n19087) );
  XNOR2_X1 U22252 ( .A(n19087), .B(n19086), .ZN(n19388) );
  AOI22_X1 U22253 ( .A1(n19088), .A2(n19388), .B1(n19402), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n19092) );
  AOI22_X1 U22254 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n10189), .ZN(n19091) );
  OAI211_X1 U22255 ( .C1(n19099), .C2(n19395), .A(n19092), .B(n19091), .ZN(
        P3_U2829) );
  AOI21_X1 U22256 ( .B1(n19094), .B2(n19396), .A(n19093), .ZN(n19407) );
  INV_X1 U22257 ( .A(n19407), .ZN(n19405) );
  NAND3_X1 U22258 ( .A1(n19895), .A2(n19096), .A3(n19095), .ZN(n19097) );
  AOI22_X1 U22259 ( .A1(n19402), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19097), .ZN(n19098) );
  OAI221_X1 U22260 ( .B1(n19407), .B2(n19100), .C1(n19405), .C2(n19099), .A(
        n19098), .ZN(P3_U2830) );
  NOR2_X1 U22261 ( .A1(n19169), .A2(n19101), .ZN(n19111) );
  OAI22_X1 U22262 ( .A1(n19398), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n19314), .B2(n19102), .ZN(n19103) );
  INV_X1 U22263 ( .A(n19103), .ZN(n19109) );
  INV_X1 U22264 ( .A(n19290), .ZN(n19265) );
  NOR2_X1 U22265 ( .A1(n19371), .A2(n19161), .ZN(n19204) );
  NAND2_X1 U22266 ( .A1(n19121), .A2(n19204), .ZN(n19120) );
  NAND2_X1 U22267 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19123) );
  INV_X1 U22268 ( .A(n19369), .ZN(n19208) );
  OAI21_X1 U22269 ( .B1(n19120), .B2(n19123), .A(n19208), .ZN(n19106) );
  NAND4_X1 U22270 ( .A1(n19109), .A2(n19108), .A3(n19107), .A4(n19106), .ZN(
        n19116) );
  NAND2_X1 U22271 ( .A1(n19402), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n19112) );
  OAI211_X1 U22272 ( .C1(n19113), .C2(n19310), .A(n9728), .B(n19112), .ZN(
        P3_U2835) );
  AOI22_X1 U22273 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19392), .B1(
        n19402), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n19119) );
  AOI22_X1 U22274 ( .A1(n19186), .A2(n19115), .B1(n19326), .B2(n19114), .ZN(
        n19118) );
  NAND3_X1 U22275 ( .A1(n19397), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n19116), .ZN(n19117) );
  NAND3_X1 U22276 ( .A1(n19119), .A2(n19118), .A3(n19117), .ZN(P3_U2836) );
  NAND2_X1 U22277 ( .A1(n19208), .A2(n19120), .ZN(n19138) );
  INV_X1 U22278 ( .A(n19121), .ZN(n19151) );
  OAI21_X1 U22279 ( .B1(n19151), .B2(n19159), .A(n19880), .ZN(n19142) );
  NAND2_X1 U22280 ( .A1(n19138), .A2(n19142), .ZN(n19122) );
  OAI211_X1 U22281 ( .C1(n19123), .C2(n19122), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n19145), .ZN(n19127) );
  NAND3_X1 U22282 ( .A1(n19125), .A2(n10268), .A3(n19124), .ZN(n19126) );
  OAI211_X1 U22283 ( .C1(n19128), .C2(n19290), .A(n19127), .B(n19126), .ZN(
        n19132) );
  OAI22_X1 U22284 ( .A1(n19406), .A2(n19130), .B1(n19310), .B2(n19129), .ZN(
        n19131) );
  AOI21_X1 U22285 ( .B1(n19397), .B2(n19132), .A(n19131), .ZN(n19134) );
  OAI211_X1 U22286 ( .C1(n19384), .C2(n10268), .A(n19134), .B(n19133), .ZN(
        P3_U2837) );
  AOI22_X1 U22287 ( .A1(n19135), .A2(n19326), .B1(n19402), .B2(
        P3_REIP_REG_24__SCAN_IN), .ZN(n19147) );
  INV_X1 U22288 ( .A(n19136), .ZN(n19137) );
  AOI21_X1 U22289 ( .B1(n19265), .B2(n19137), .A(n19392), .ZN(n19139) );
  OAI211_X1 U22290 ( .C1(n19140), .C2(n19379), .A(n19139), .B(n19138), .ZN(
        n19144) );
  NOR2_X1 U22291 ( .A1(n19141), .A2(n19144), .ZN(n19143) );
  AOI21_X1 U22292 ( .B1(n19143), .B2(n19142), .A(n19402), .ZN(n19152) );
  OAI211_X1 U22293 ( .C1(n19145), .C2(n19144), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n19152), .ZN(n19146) );
  OAI211_X1 U22294 ( .C1(n19149), .C2(n19148), .A(n19147), .B(n19146), .ZN(
        P3_U2838) );
  INV_X1 U22295 ( .A(n19150), .ZN(n19156) );
  NOR3_X1 U22296 ( .A1(n19392), .A2(n19169), .A3(n19151), .ZN(n19153) );
  OAI21_X1 U22297 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n19153), .A(
        n19152), .ZN(n19154) );
  OAI211_X1 U22298 ( .C1(n19156), .C2(n19310), .A(n19155), .B(n19154), .ZN(
        P3_U2839) );
  OAI22_X1 U22299 ( .A1(n19158), .A2(n19379), .B1(n19157), .B2(n19290), .ZN(
        n19175) );
  INV_X1 U22300 ( .A(n19159), .ZN(n19201) );
  AOI21_X1 U22301 ( .B1(n19179), .B2(n19201), .A(n19375), .ZN(n19160) );
  AOI221_X1 U22302 ( .B1(n19161), .B2(n19224), .C1(n19190), .C2(n19224), .A(
        n19160), .ZN(n19192) );
  NAND2_X1 U22303 ( .A1(n19379), .A2(n19290), .ZN(n19296) );
  AOI22_X1 U22304 ( .A1(n19224), .A2(n19162), .B1(n19168), .B2(n19296), .ZN(
        n19163) );
  NAND2_X1 U22305 ( .A1(n19192), .A2(n19163), .ZN(n19178) );
  OAI21_X1 U22306 ( .B1(n19164), .B2(n19221), .A(n19277), .ZN(n19188) );
  OAI211_X1 U22307 ( .C1(n19227), .C2(n19165), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n19188), .ZN(n19166) );
  NOR3_X1 U22308 ( .A1(n19175), .A2(n19178), .A3(n19166), .ZN(n19167) );
  AOI221_X1 U22309 ( .B1(n19169), .B2(n19174), .C1(n19168), .C2(n19174), .A(
        n19167), .ZN(n19171) );
  AOI22_X1 U22310 ( .A1(n19397), .A2(n19171), .B1(n19326), .B2(n19170), .ZN(
        n19173) );
  OAI211_X1 U22311 ( .C1(n19384), .C2(n19174), .A(n19173), .B(n19172), .ZN(
        P3_U2840) );
  NOR2_X1 U22312 ( .A1(n19880), .A2(n19277), .ZN(n19391) );
  OAI211_X1 U22313 ( .C1(n19176), .C2(n19391), .A(n19226), .B(n19188), .ZN(
        n19177) );
  OAI21_X1 U22314 ( .B1(n19178), .B2(n19177), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19184) );
  NAND2_X1 U22315 ( .A1(n19179), .A2(n19186), .ZN(n19200) );
  INV_X1 U22316 ( .A(n19200), .ZN(n19180) );
  AOI22_X1 U22317 ( .A1(n19326), .A2(n19182), .B1(n19181), .B2(n19180), .ZN(
        n19183) );
  OAI221_X1 U22318 ( .B1(n19402), .B2(n19184), .C1(n19400), .C2(n19974), .A(
        n19183), .ZN(P3_U2841) );
  AOI22_X1 U22319 ( .A1(n19326), .A2(n19187), .B1(n19186), .B2(n19185), .ZN(
        n19195) );
  NAND2_X1 U22320 ( .A1(n19226), .A2(n19188), .ZN(n19189) );
  AOI21_X1 U22321 ( .B1(n19190), .B2(n19296), .A(n19189), .ZN(n19191) );
  AOI21_X1 U22322 ( .B1(n19192), .B2(n19191), .A(n19402), .ZN(n19197) );
  NOR3_X1 U22323 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19391), .A3(
        n20039), .ZN(n19193) );
  OAI21_X1 U22324 ( .B1(n19197), .B2(n19193), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19194) );
  OAI211_X1 U22325 ( .C1(n19972), .C2(n19400), .A(n19195), .B(n19194), .ZN(
        P3_U2842) );
  AOI22_X1 U22326 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19197), .B1(
        n19326), .B2(n19196), .ZN(n19199) );
  OAI211_X1 U22327 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19200), .A(
        n19199), .B(n19198), .ZN(P3_U2843) );
  NOR2_X1 U22328 ( .A1(n19201), .A2(n19375), .ZN(n19203) );
  OAI22_X1 U22329 ( .A1(n19880), .A2(n19296), .B1(n19203), .B2(n19202), .ZN(
        n19207) );
  AOI21_X1 U22330 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19204), .A(
        n19369), .ZN(n19205) );
  INV_X1 U22331 ( .A(n19205), .ZN(n19206) );
  NAND3_X1 U22332 ( .A1(n19226), .A2(n19207), .A3(n19206), .ZN(n19216) );
  OAI221_X1 U22333 ( .B1(n19216), .B2(n19217), .C1(n19216), .C2(n19208), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19214) );
  NOR2_X1 U22334 ( .A1(n19359), .A2(n19209), .ZN(n19275) );
  OAI21_X1 U22335 ( .B1(n19275), .B2(n19274), .A(n19397), .ZN(n19320) );
  NOR2_X1 U22336 ( .A1(n19210), .A2(n19320), .ZN(n19229) );
  AOI22_X1 U22337 ( .A1(n19326), .A2(n19212), .B1(n19211), .B2(n19229), .ZN(
        n19213) );
  OAI221_X1 U22338 ( .B1(n19402), .B2(n19214), .C1(n19400), .C2(n19968), .A(
        n19213), .ZN(P3_U2844) );
  AOI22_X1 U22339 ( .A1(n19215), .A2(n19326), .B1(n19402), .B2(
        P3_REIP_REG_17__SCAN_IN), .ZN(n19220) );
  NAND3_X1 U22340 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19400), .A3(
        n19216), .ZN(n19219) );
  NAND3_X1 U22341 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19229), .A3(
        n19217), .ZN(n19218) );
  NAND3_X1 U22342 ( .A1(n19220), .A2(n19219), .A3(n19218), .ZN(P3_U2845) );
  INV_X1 U22343 ( .A(n19221), .ZN(n19222) );
  AOI21_X1 U22344 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19314), .A(
        n19222), .ZN(n19225) );
  OR2_X1 U22345 ( .A1(n19223), .A2(n19375), .ZN(n19293) );
  NAND2_X1 U22346 ( .A1(n19224), .A2(n19250), .ZN(n19313) );
  NAND2_X1 U22347 ( .A1(n19293), .A2(n19313), .ZN(n19248) );
  AOI211_X1 U22348 ( .C1(n19304), .C2(n19236), .A(n19225), .B(n19248), .ZN(
        n19238) );
  AOI221_X1 U22349 ( .B1(n19227), .B2(n19226), .C1(n19238), .C2(n19226), .A(
        n19402), .ZN(n19230) );
  AOI22_X1 U22350 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19228), .ZN(n19232) );
  NAND2_X1 U22351 ( .A1(n19402), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n19231) );
  OAI211_X1 U22352 ( .C1(n19233), .C2(n19310), .A(n19232), .B(n19231), .ZN(
        P3_U2846) );
  NAND2_X1 U22353 ( .A1(n19265), .A2(n19234), .ZN(n19243) );
  NAND2_X1 U22354 ( .A1(n19878), .A2(n19235), .ZN(n19241) );
  INV_X1 U22355 ( .A(n19236), .ZN(n19237) );
  AOI21_X1 U22356 ( .B1(n19237), .B2(n19275), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19239) );
  OAI222_X1 U22357 ( .A1(n19243), .A2(n19242), .B1(n19241), .B2(n19240), .C1(
        n19239), .C2(n19238), .ZN(n19245) );
  AOI22_X1 U22358 ( .A1(n19397), .A2(n19245), .B1(n19326), .B2(n19244), .ZN(
        n19247) );
  OAI211_X1 U22359 ( .C1(n19384), .C2(n17304), .A(n19247), .B(n19246), .ZN(
        P3_U2847) );
  AOI211_X1 U22360 ( .C1(n19304), .C2(n19249), .A(n18927), .B(n19248), .ZN(
        n19252) );
  NOR2_X1 U22361 ( .A1(n19396), .A2(n19250), .ZN(n19312) );
  NAND2_X1 U22362 ( .A1(n19251), .A2(n19312), .ZN(n19278) );
  NAND2_X1 U22363 ( .A1(n19277), .A2(n19278), .ZN(n19268) );
  OAI211_X1 U22364 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n19391), .A(
        n19252), .B(n19268), .ZN(n19253) );
  OAI221_X1 U22365 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19254), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n19275), .A(n19253), .ZN(
        n19255) );
  OAI22_X1 U22366 ( .A1(n18927), .A2(n19384), .B1(n19390), .B2(n19255), .ZN(
        n19256) );
  AOI21_X1 U22367 ( .B1(n19402), .B2(P3_REIP_REG_14__SCAN_IN), .A(n19256), 
        .ZN(n19261) );
  AOI22_X1 U22368 ( .A1(n19259), .A2(n19258), .B1(n19326), .B2(n19257), .ZN(
        n19260) );
  OAI211_X1 U22369 ( .C1(n19406), .C2(n19262), .A(n19261), .B(n19260), .ZN(
        P3_U2848) );
  AOI22_X1 U22370 ( .A1(n19402), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19326), 
        .B2(n19263), .ZN(n19272) );
  INV_X1 U22371 ( .A(n19313), .ZN(n19303) );
  AOI21_X1 U22372 ( .B1(n19304), .B2(n19280), .A(n19303), .ZN(n19298) );
  AOI22_X1 U22373 ( .A1(n19878), .A2(n19266), .B1(n19265), .B2(n19264), .ZN(
        n19267) );
  NAND3_X1 U22374 ( .A1(n19298), .A2(n19267), .A3(n19293), .ZN(n19276) );
  OAI211_X1 U22375 ( .C1(n19269), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19397), .B(n19268), .ZN(n19270) );
  OAI211_X1 U22376 ( .C1(n19276), .C2(n19270), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19400), .ZN(n19271) );
  OAI211_X1 U22377 ( .C1(n19320), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P3_U2849) );
  NOR2_X1 U22378 ( .A1(n19275), .A2(n19274), .ZN(n19281) );
  AOI211_X1 U22379 ( .C1(n19278), .C2(n19277), .A(n19276), .B(n19287), .ZN(
        n19279) );
  AOI221_X1 U22380 ( .B1(n19281), .B2(n19287), .C1(n19280), .C2(n19287), .A(
        n19279), .ZN(n19283) );
  AOI22_X1 U22381 ( .A1(n19397), .A2(n19283), .B1(n19326), .B2(n19282), .ZN(
        n19286) );
  INV_X1 U22382 ( .A(n19284), .ZN(n19285) );
  OAI211_X1 U22383 ( .C1(n19384), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P3_U2850) );
  AOI22_X1 U22384 ( .A1(n19402), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19326), 
        .B2(n19288), .ZN(n19301) );
  AOI21_X1 U22385 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19312), .A(
        n19314), .ZN(n19295) );
  OAI22_X1 U22386 ( .A1(n19291), .A2(n19290), .B1(n19379), .B2(n19289), .ZN(
        n19292) );
  NOR2_X1 U22387 ( .A1(n19390), .A2(n19292), .ZN(n19294) );
  NAND2_X1 U22388 ( .A1(n19294), .A2(n19293), .ZN(n19315) );
  AOI211_X1 U22389 ( .C1(n19297), .C2(n19296), .A(n19295), .B(n19315), .ZN(
        n19306) );
  OAI211_X1 U22390 ( .C1(n19314), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n19298), .B(n19306), .ZN(n19299) );
  NAND3_X1 U22391 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19400), .A3(
        n19299), .ZN(n19300) );
  OAI211_X1 U22392 ( .C1(n19320), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P3_U2851) );
  AOI21_X1 U22393 ( .B1(n19304), .B2(n17301), .A(n19303), .ZN(n19305) );
  AOI21_X1 U22394 ( .B1(n19306), .B2(n19305), .A(n10282), .ZN(n19308) );
  NOR3_X1 U22395 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17301), .A3(
        n19320), .ZN(n19307) );
  AOI221_X1 U22396 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n19402), .C1(n19308), 
        .C2(n19400), .A(n19307), .ZN(n19309) );
  OAI21_X1 U22397 ( .B1(n19311), .B2(n19310), .A(n19309), .ZN(P3_U2852) );
  AOI21_X1 U22398 ( .B1(n19314), .B2(n19313), .A(n19312), .ZN(n19316) );
  OAI21_X1 U22399 ( .B1(n19316), .B2(n19315), .A(n19400), .ZN(n19319) );
  AOI22_X1 U22400 ( .A1(n19402), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19326), 
        .B2(n19317), .ZN(n19318) );
  OAI221_X1 U22401 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19320), .C1(
        n17301), .C2(n19319), .A(n19318), .ZN(P3_U2853) );
  OAI22_X1 U22402 ( .A1(n19323), .A2(n19406), .B1(n19322), .B2(n19321), .ZN(
        n19324) );
  AOI21_X1 U22403 ( .B1(n19326), .B2(n19325), .A(n19324), .ZN(n19332) );
  OAI21_X1 U22404 ( .B1(n19392), .B2(n19327), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19330) );
  NOR2_X1 U22405 ( .A1(n19359), .A2(n19390), .ZN(n19349) );
  NAND3_X1 U22406 ( .A1(n19328), .A2(n19349), .A3(n10273), .ZN(n19329) );
  NAND4_X1 U22407 ( .A1(n19332), .A2(n19331), .A3(n19330), .A4(n19329), .ZN(
        P3_U2854) );
  OAI21_X1 U22408 ( .B1(n19333), .B2(n19385), .A(n19384), .ZN(n19345) );
  OAI22_X1 U22409 ( .A1(n19406), .A2(n19335), .B1(n19404), .B2(n19334), .ZN(
        n19336) );
  AOI21_X1 U22410 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19345), .A(
        n19336), .ZN(n19340) );
  NAND3_X1 U22411 ( .A1(n19338), .A2(n19349), .A3(n19337), .ZN(n19339) );
  OAI211_X1 U22412 ( .C1(n19944), .C2(n19400), .A(n19340), .B(n19339), .ZN(
        P3_U2856) );
  OAI22_X1 U22413 ( .A1(n19406), .A2(n19342), .B1(n19404), .B2(n19341), .ZN(
        n19343) );
  AOI211_X1 U22414 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n19345), .A(
        n19344), .B(n19343), .ZN(n19348) );
  NAND4_X1 U22415 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n19349), .A4(n19346), .ZN(
        n19347) );
  NAND2_X1 U22416 ( .A1(n19348), .A2(n19347), .ZN(P3_U2857) );
  AND2_X1 U22417 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19349), .ZN(
        n19355) );
  AOI21_X1 U22418 ( .B1(n19350), .B2(n19364), .A(n19392), .ZN(n19352) );
  OAI22_X1 U22419 ( .A1(n19352), .A2(n19354), .B1(n19404), .B2(n19351), .ZN(
        n19353) );
  AOI21_X1 U22420 ( .B1(n19355), .B2(n19354), .A(n19353), .ZN(n19357) );
  NAND2_X1 U22421 ( .A1(n19402), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n19356) );
  OAI211_X1 U22422 ( .C1(n19406), .C2(n19358), .A(n19357), .B(n19356), .ZN(
        P3_U2858) );
  AOI21_X1 U22423 ( .B1(n19359), .B2(n19367), .A(n19390), .ZN(n19363) );
  OAI22_X1 U22424 ( .A1(n19406), .A2(n19361), .B1(n19404), .B2(n19360), .ZN(
        n19362) );
  AOI21_X1 U22425 ( .B1(n19364), .B2(n19363), .A(n19362), .ZN(n19366) );
  OAI211_X1 U22426 ( .C1(n19384), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P3_U2859) );
  NAND2_X1 U22427 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19368) );
  OAI22_X1 U22428 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19369), .B1(
        n19375), .B2(n19368), .ZN(n19370) );
  OAI21_X1 U22429 ( .B1(n19371), .B2(n19370), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19374) );
  NAND3_X1 U22430 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19372), .A3(
        n13945), .ZN(n19373) );
  OAI211_X1 U22431 ( .C1(n19376), .C2(n19375), .A(n19374), .B(n19373), .ZN(
        n19381) );
  OAI22_X1 U22432 ( .A1(n19379), .A2(n19378), .B1(n19377), .B2(n19875), .ZN(
        n19380) );
  OAI21_X1 U22433 ( .B1(n19381), .B2(n19380), .A(n19397), .ZN(n19382) );
  OAI211_X1 U22434 ( .C1(n19384), .C2(n13945), .A(n19383), .B(n19382), .ZN(
        P3_U2860) );
  NOR2_X1 U22435 ( .A1(n19400), .A2(n20010), .ZN(n19387) );
  AOI211_X1 U22436 ( .C1(n19398), .C2(n19396), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n19385), .ZN(n19386) );
  AOI211_X1 U22437 ( .C1(n19389), .C2(n19388), .A(n19387), .B(n19386), .ZN(
        n19394) );
  NOR3_X1 U22438 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19391), .A3(
        n19390), .ZN(n19399) );
  OAI21_X1 U22439 ( .B1(n19392), .B2(n19399), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19393) );
  OAI211_X1 U22440 ( .C1(n19395), .C2(n19404), .A(n19394), .B(n19393), .ZN(
        P3_U2861) );
  AOI21_X1 U22441 ( .B1(n19398), .B2(n19397), .A(n19396), .ZN(n19401) );
  AOI221_X1 U22442 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n19402), .C1(n19401), 
        .C2(n19400), .A(n19399), .ZN(n19403) );
  OAI221_X1 U22443 ( .B1(n19407), .B2(n19406), .C1(n19405), .C2(n19404), .A(
        n19403), .ZN(P3_U2862) );
  AOI211_X1 U22444 ( .C1(n19409), .C2(n19408), .A(n20039), .B(n19895), .ZN(
        n19900) );
  OAI21_X1 U22445 ( .B1(n19900), .B2(n19458), .A(n19419), .ZN(n19410) );
  OAI221_X1 U22446 ( .B1(n13148), .B2(n20025), .C1(n13148), .C2(n19419), .A(
        n19410), .ZN(P3_U2863) );
  AOI221_X1 U22447 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19866), .C1(n19412), 
        .C2(n19866), .A(n19411), .ZN(n19418) );
  NOR2_X1 U22448 ( .A1(n19413), .A2(n19866), .ZN(n19415) );
  OAI21_X1 U22449 ( .B1(n19415), .B2(n19414), .A(n19419), .ZN(n19416) );
  AOI22_X1 U22450 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19418), .B1(
        n19416), .B2(n19882), .ZN(P3_U2865) );
  NAND2_X1 U22451 ( .A1(n19860), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19566) );
  INV_X1 U22452 ( .A(n19566), .ZN(n19590) );
  NOR2_X1 U22453 ( .A1(n19860), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19635) );
  NOR2_X1 U22454 ( .A1(n19590), .A2(n19635), .ZN(n19417) );
  OAI22_X1 U22455 ( .A1(n19418), .A2(n19860), .B1(n19417), .B2(n19416), .ZN(
        P3_U2866) );
  NOR2_X1 U22456 ( .A1(n19861), .A2(n19419), .ZN(P3_U2867) );
  NOR2_X1 U22457 ( .A1(n19882), .A2(n19860), .ZN(n19731) );
  INV_X1 U22458 ( .A(n19731), .ZN(n19420) );
  NOR2_X1 U22459 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19420), .ZN(
        n19800) );
  NAND2_X1 U22460 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19800), .ZN(
        n19838) );
  NOR2_X1 U22461 ( .A1(n16462), .A2(n19479), .ZN(n19797) );
  NOR2_X1 U22462 ( .A1(n19866), .A2(n19420), .ZN(n19799) );
  NAND2_X1 U22463 ( .A1(n13148), .A2(n19799), .ZN(n19477) );
  NOR2_X2 U22464 ( .A1(n19479), .A2(n19421), .ZN(n19802) );
  NOR2_X2 U22465 ( .A1(n19523), .A2(n19422), .ZN(n19796) );
  INV_X1 U22466 ( .A(n19729), .ZN(n19908) );
  NOR2_X1 U22467 ( .A1(n19866), .A2(n13148), .ZN(n19864) );
  NAND2_X1 U22468 ( .A1(n19864), .A2(n19731), .ZN(n19806) );
  INV_X1 U22469 ( .A(n19806), .ZN(n19850) );
  NOR2_X1 U22470 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19611) );
  NOR2_X1 U22471 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19501) );
  NAND2_X1 U22472 ( .A1(n19611), .A2(n19501), .ZN(n19516) );
  NOR2_X1 U22473 ( .A1(n19850), .A2(n19518), .ZN(n19480) );
  NOR2_X1 U22474 ( .A1(n19908), .A2(n19480), .ZN(n19453) );
  AOI22_X1 U22475 ( .A1(n19790), .A2(n19802), .B1(n19796), .B2(n19453), .ZN(
        n19428) );
  INV_X1 U22476 ( .A(n19838), .ZN(n19848) );
  NOR2_X1 U22477 ( .A1(n19848), .A2(n19790), .ZN(n19755) );
  INV_X1 U22478 ( .A(n19523), .ZN(n19759) );
  OAI21_X1 U22479 ( .B1(n13148), .B2(n20009), .A(n19759), .ZN(n19612) );
  OAI22_X1 U22480 ( .A1(n19479), .A2(n19755), .B1(n19612), .B2(n19480), .ZN(
        n19423) );
  NAND2_X1 U22481 ( .A1(n19425), .A2(n19424), .ZN(n19454) );
  NOR2_X1 U22482 ( .A1(n19426), .A2(n19454), .ZN(n19760) );
  AOI22_X1 U22483 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19760), .ZN(n19427) );
  OAI211_X1 U22484 ( .C1(n19838), .C2(n19763), .A(n19428), .B(n19427), .ZN(
        P3_U2868) );
  NOR2_X1 U22485 ( .A1(n19429), .A2(n19479), .ZN(n19764) );
  NAND2_X1 U22486 ( .A1(n19801), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19767) );
  INV_X1 U22487 ( .A(n19767), .ZN(n19808) );
  AOI22_X1 U22488 ( .A1(n19790), .A2(n19808), .B1(n19453), .B2(n19807), .ZN(
        n19432) );
  NOR2_X2 U22489 ( .A1(n19430), .A2(n19454), .ZN(n19809) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19809), .ZN(n19431) );
  OAI211_X1 U22491 ( .C1(n19838), .C2(n19812), .A(n19432), .B(n19431), .ZN(
        P3_U2869) );
  NOR2_X1 U22492 ( .A1(n19479), .A2(n16505), .ZN(n19768) );
  INV_X1 U22493 ( .A(n19768), .ZN(n19818) );
  NAND2_X1 U22494 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19801), .ZN(n19771) );
  INV_X1 U22495 ( .A(n19771), .ZN(n19814) );
  NOR2_X2 U22496 ( .A1(n19523), .A2(n19433), .ZN(n19813) );
  AOI22_X1 U22497 ( .A1(n19848), .A2(n19814), .B1(n19453), .B2(n19813), .ZN(
        n19436) );
  NOR2_X2 U22498 ( .A1(n19434), .A2(n19454), .ZN(n19815) );
  AOI22_X1 U22499 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19815), .ZN(n19435) );
  OAI211_X1 U22500 ( .C1(n19477), .C2(n19818), .A(n19436), .B(n19435), .ZN(
        P3_U2870) );
  NOR2_X1 U22501 ( .A1(n16442), .A2(n19479), .ZN(n19820) );
  INV_X1 U22502 ( .A(n19820), .ZN(n19775) );
  NAND2_X1 U22503 ( .A1(n19801), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19824) );
  INV_X1 U22504 ( .A(n19824), .ZN(n19772) );
  NOR2_X2 U22505 ( .A1(n19523), .A2(n19437), .ZN(n19819) );
  AOI22_X1 U22506 ( .A1(n19790), .A2(n19772), .B1(n19453), .B2(n19819), .ZN(
        n19440) );
  NOR2_X2 U22507 ( .A1(n19438), .A2(n19454), .ZN(n19821) );
  AOI22_X1 U22508 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19821), .ZN(n19439) );
  OAI211_X1 U22509 ( .C1(n19838), .C2(n19775), .A(n19440), .B(n19439), .ZN(
        P3_U2871) );
  NOR2_X1 U22510 ( .A1(n19479), .A2(n16488), .ZN(n19826) );
  NAND2_X1 U22511 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19801), .ZN(n19830) );
  NOR2_X2 U22512 ( .A1(n19523), .A2(n19441), .ZN(n19825) );
  AOI22_X1 U22513 ( .A1(n19848), .A2(n19742), .B1(n19453), .B2(n19825), .ZN(
        n19444) );
  NOR2_X2 U22514 ( .A1(n19442), .A2(n19454), .ZN(n19827) );
  AOI22_X1 U22515 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19827), .ZN(n19443) );
  OAI211_X1 U22516 ( .C1(n19477), .C2(n19745), .A(n19444), .B(n19443), .ZN(
        P3_U2872) );
  NOR2_X1 U22517 ( .A1(n19479), .A2(n20274), .ZN(n19778) );
  INV_X1 U22518 ( .A(n19778), .ZN(n19837) );
  NAND2_X1 U22519 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19801), .ZN(n19782) );
  INV_X1 U22520 ( .A(n19782), .ZN(n19833) );
  NOR2_X2 U22521 ( .A1(n19523), .A2(n19445), .ZN(n19831) );
  AOI22_X1 U22522 ( .A1(n19848), .A2(n19833), .B1(n19453), .B2(n19831), .ZN(
        n19448) );
  NOR2_X2 U22523 ( .A1(n19446), .A2(n19454), .ZN(n19834) );
  AOI22_X1 U22524 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19834), .ZN(n19447) );
  OAI211_X1 U22525 ( .C1(n19477), .C2(n19837), .A(n19448), .B(n19447), .ZN(
        P3_U2873) );
  NOR2_X1 U22526 ( .A1(n19479), .A2(n16475), .ZN(n19840) );
  INV_X1 U22527 ( .A(n19840), .ZN(n19786) );
  NAND2_X1 U22528 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19801), .ZN(n19844) );
  INV_X1 U22529 ( .A(n19844), .ZN(n19783) );
  NOR2_X2 U22530 ( .A1(n19523), .A2(n13757), .ZN(n19839) );
  AOI22_X1 U22531 ( .A1(n19848), .A2(n19783), .B1(n19453), .B2(n19839), .ZN(
        n19451) );
  NOR2_X2 U22532 ( .A1(n19449), .A2(n19454), .ZN(n19841) );
  AOI22_X1 U22533 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19841), .ZN(n19450) );
  OAI211_X1 U22534 ( .C1(n19477), .C2(n19786), .A(n19451), .B(n19450), .ZN(
        P3_U2874) );
  NOR2_X1 U22535 ( .A1(n19479), .A2(n16469), .ZN(n19847) );
  INV_X1 U22536 ( .A(n19847), .ZN(n19794) );
  NAND2_X1 U22537 ( .A1(n19801), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19855) );
  INV_X1 U22538 ( .A(n19855), .ZN(n19789) );
  NOR2_X2 U22539 ( .A1(n19523), .A2(n19452), .ZN(n19846) );
  AOI22_X1 U22540 ( .A1(n19848), .A2(n19789), .B1(n19453), .B2(n19846), .ZN(
        n19457) );
  NOR2_X2 U22541 ( .A1(n10457), .A2(n19454), .ZN(n19849) );
  AOI22_X1 U22542 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19455), .B1(
        n19518), .B2(n19849), .ZN(n19456) );
  OAI211_X1 U22543 ( .C1(n19477), .C2(n19794), .A(n19457), .B(n19456), .ZN(
        P3_U2875) );
  INV_X1 U22544 ( .A(n19501), .ZN(n19478) );
  NAND2_X1 U22545 ( .A1(n19866), .A2(n19729), .ZN(n19636) );
  NOR2_X1 U22546 ( .A1(n19478), .A2(n19636), .ZN(n19473) );
  AOI22_X1 U22547 ( .A1(n19850), .A2(n19802), .B1(n19796), .B2(n19473), .ZN(
        n19460) );
  NOR2_X1 U22548 ( .A1(n19523), .A2(n19458), .ZN(n19798) );
  INV_X1 U22549 ( .A(n19798), .ZN(n19500) );
  NOR2_X1 U22550 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19500), .ZN(
        n19730) );
  AOI22_X1 U22551 ( .A1(n19801), .A2(n19799), .B1(n19501), .B2(n19730), .ZN(
        n19474) );
  NAND2_X1 U22552 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19866), .ZN(
        n19638) );
  NOR2_X2 U22553 ( .A1(n19478), .A2(n19638), .ZN(n19535) );
  AOI22_X1 U22554 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19474), .B1(
        n19760), .B2(n19535), .ZN(n19459) );
  OAI211_X1 U22555 ( .C1(n19477), .C2(n19763), .A(n19460), .B(n19459), .ZN(
        P3_U2876) );
  AOI22_X1 U22556 ( .A1(n19850), .A2(n19808), .B1(n19807), .B2(n19473), .ZN(
        n19462) );
  AOI22_X1 U22557 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19474), .B1(
        n19809), .B2(n19535), .ZN(n19461) );
  OAI211_X1 U22558 ( .C1(n19477), .C2(n19812), .A(n19462), .B(n19461), .ZN(
        P3_U2877) );
  AOI22_X1 U22559 ( .A1(n19850), .A2(n19768), .B1(n19813), .B2(n19473), .ZN(
        n19464) );
  AOI22_X1 U22560 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19474), .B1(
        n19815), .B2(n19535), .ZN(n19463) );
  OAI211_X1 U22561 ( .C1(n19477), .C2(n19771), .A(n19464), .B(n19463), .ZN(
        P3_U2878) );
  AOI22_X1 U22562 ( .A1(n19850), .A2(n19772), .B1(n19819), .B2(n19473), .ZN(
        n19466) );
  AOI22_X1 U22563 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19474), .B1(
        n19821), .B2(n19535), .ZN(n19465) );
  OAI211_X1 U22564 ( .C1(n19477), .C2(n19775), .A(n19466), .B(n19465), .ZN(
        P3_U2879) );
  AOI22_X1 U22565 ( .A1(n19850), .A2(n19826), .B1(n19825), .B2(n19473), .ZN(
        n19468) );
  AOI22_X1 U22566 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19474), .B1(
        n19827), .B2(n19535), .ZN(n19467) );
  OAI211_X1 U22567 ( .C1(n19477), .C2(n19830), .A(n19468), .B(n19467), .ZN(
        P3_U2880) );
  AOI22_X1 U22568 ( .A1(n19790), .A2(n19833), .B1(n19831), .B2(n19473), .ZN(
        n19470) );
  AOI22_X1 U22569 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19474), .B1(
        n19834), .B2(n19535), .ZN(n19469) );
  OAI211_X1 U22570 ( .C1(n19806), .C2(n19837), .A(n19470), .B(n19469), .ZN(
        P3_U2881) );
  AOI22_X1 U22571 ( .A1(n19790), .A2(n19783), .B1(n19839), .B2(n19473), .ZN(
        n19472) );
  AOI22_X1 U22572 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19474), .B1(
        n19841), .B2(n19535), .ZN(n19471) );
  OAI211_X1 U22573 ( .C1(n19806), .C2(n19786), .A(n19472), .B(n19471), .ZN(
        P3_U2882) );
  AOI22_X1 U22574 ( .A1(n19850), .A2(n19847), .B1(n19846), .B2(n19473), .ZN(
        n19476) );
  AOI22_X1 U22575 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19474), .B1(
        n19849), .B2(n19535), .ZN(n19475) );
  OAI211_X1 U22576 ( .C1(n19477), .C2(n19855), .A(n19476), .B(n19475), .ZN(
        P3_U2883) );
  INV_X1 U22577 ( .A(n19760), .ZN(n19805) );
  NOR2_X1 U22578 ( .A1(n19866), .A2(n19478), .ZN(n19545) );
  NAND2_X1 U22579 ( .A1(n19545), .A2(n13148), .ZN(n19565) );
  AOI21_X1 U22580 ( .B1(n19544), .B2(n19565), .A(n19908), .ZN(n19496) );
  AOI22_X1 U22581 ( .A1(n19850), .A2(n19797), .B1(n19796), .B2(n19496), .ZN(
        n19483) );
  INV_X1 U22582 ( .A(n19565), .ZN(n19554) );
  OAI21_X1 U22583 ( .B1(n19535), .B2(n19554), .A(n19759), .ZN(n19522) );
  OAI21_X1 U22584 ( .B1(n19480), .B2(n19479), .A(n19522), .ZN(n19481) );
  OAI21_X1 U22585 ( .B1(n19554), .B2(n20009), .A(n19481), .ZN(n19497) );
  AOI22_X1 U22586 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19497), .B1(
        n19518), .B2(n19802), .ZN(n19482) );
  OAI211_X1 U22587 ( .C1(n19805), .C2(n19565), .A(n19483), .B(n19482), .ZN(
        P3_U2884) );
  AOI22_X1 U22588 ( .A1(n19518), .A2(n19808), .B1(n19807), .B2(n19496), .ZN(
        n19485) );
  AOI22_X1 U22589 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19497), .B1(
        n19809), .B2(n19554), .ZN(n19484) );
  OAI211_X1 U22590 ( .C1(n19806), .C2(n19812), .A(n19485), .B(n19484), .ZN(
        P3_U2885) );
  AOI22_X1 U22591 ( .A1(n19850), .A2(n19814), .B1(n19813), .B2(n19496), .ZN(
        n19487) );
  AOI22_X1 U22592 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19497), .B1(
        n19815), .B2(n19554), .ZN(n19486) );
  OAI211_X1 U22593 ( .C1(n19516), .C2(n19818), .A(n19487), .B(n19486), .ZN(
        P3_U2886) );
  AOI22_X1 U22594 ( .A1(n19850), .A2(n19820), .B1(n19819), .B2(n19496), .ZN(
        n19489) );
  AOI22_X1 U22595 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19497), .B1(
        n19821), .B2(n19554), .ZN(n19488) );
  OAI211_X1 U22596 ( .C1(n19516), .C2(n19824), .A(n19489), .B(n19488), .ZN(
        P3_U2887) );
  AOI22_X1 U22597 ( .A1(n19850), .A2(n19742), .B1(n19825), .B2(n19496), .ZN(
        n19491) );
  AOI22_X1 U22598 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19497), .B1(
        n19827), .B2(n19554), .ZN(n19490) );
  OAI211_X1 U22599 ( .C1(n19516), .C2(n19745), .A(n19491), .B(n19490), .ZN(
        P3_U2888) );
  AOI22_X1 U22600 ( .A1(n19518), .A2(n19778), .B1(n19831), .B2(n19496), .ZN(
        n19493) );
  AOI22_X1 U22601 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19497), .B1(
        n19834), .B2(n19554), .ZN(n19492) );
  OAI211_X1 U22602 ( .C1(n19806), .C2(n19782), .A(n19493), .B(n19492), .ZN(
        P3_U2889) );
  AOI22_X1 U22603 ( .A1(n19850), .A2(n19783), .B1(n19839), .B2(n19496), .ZN(
        n19495) );
  AOI22_X1 U22604 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19497), .B1(
        n19841), .B2(n19554), .ZN(n19494) );
  OAI211_X1 U22605 ( .C1(n19516), .C2(n19786), .A(n19495), .B(n19494), .ZN(
        P3_U2890) );
  AOI22_X1 U22606 ( .A1(n19518), .A2(n19847), .B1(n19846), .B2(n19496), .ZN(
        n19499) );
  AOI22_X1 U22607 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19497), .B1(
        n19849), .B2(n19554), .ZN(n19498) );
  OAI211_X1 U22608 ( .C1(n19806), .C2(n19855), .A(n19499), .B(n19498), .ZN(
        P3_U2891) );
  AND2_X1 U22609 ( .A1(n19729), .A2(n19545), .ZN(n19517) );
  AOI22_X1 U22610 ( .A1(n19802), .A2(n19535), .B1(n19796), .B2(n19517), .ZN(
        n19503) );
  AOI21_X1 U22611 ( .B1(n19866), .B2(n19756), .A(n19500), .ZN(n19589) );
  NAND2_X1 U22612 ( .A1(n19501), .A2(n19589), .ZN(n19519) );
  NAND2_X1 U22613 ( .A1(n19864), .A2(n19501), .ZN(n19588) );
  AOI22_X1 U22614 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19519), .B1(
        n19760), .B2(n19575), .ZN(n19502) );
  OAI211_X1 U22615 ( .C1(n19516), .C2(n19763), .A(n19503), .B(n19502), .ZN(
        P3_U2892) );
  AOI22_X1 U22616 ( .A1(n19808), .A2(n19535), .B1(n19807), .B2(n19517), .ZN(
        n19505) );
  AOI22_X1 U22617 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19519), .B1(
        n19809), .B2(n19575), .ZN(n19504) );
  OAI211_X1 U22618 ( .C1(n19516), .C2(n19812), .A(n19505), .B(n19504), .ZN(
        P3_U2893) );
  AOI22_X1 U22619 ( .A1(n19518), .A2(n19814), .B1(n19813), .B2(n19517), .ZN(
        n19507) );
  AOI22_X1 U22620 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19519), .B1(
        n19815), .B2(n19575), .ZN(n19506) );
  OAI211_X1 U22621 ( .C1(n19818), .C2(n19544), .A(n19507), .B(n19506), .ZN(
        P3_U2894) );
  AOI22_X1 U22622 ( .A1(n19772), .A2(n19535), .B1(n19819), .B2(n19517), .ZN(
        n19509) );
  AOI22_X1 U22623 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19519), .B1(
        n19821), .B2(n19575), .ZN(n19508) );
  OAI211_X1 U22624 ( .C1(n19516), .C2(n19775), .A(n19509), .B(n19508), .ZN(
        P3_U2895) );
  AOI22_X1 U22625 ( .A1(n19518), .A2(n19742), .B1(n19825), .B2(n19517), .ZN(
        n19511) );
  AOI22_X1 U22626 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19519), .B1(
        n19827), .B2(n19575), .ZN(n19510) );
  OAI211_X1 U22627 ( .C1(n19745), .C2(n19544), .A(n19511), .B(n19510), .ZN(
        P3_U2896) );
  AOI22_X1 U22628 ( .A1(n19518), .A2(n19833), .B1(n19831), .B2(n19517), .ZN(
        n19513) );
  AOI22_X1 U22629 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19519), .B1(
        n19834), .B2(n19575), .ZN(n19512) );
  OAI211_X1 U22630 ( .C1(n19837), .C2(n19544), .A(n19513), .B(n19512), .ZN(
        P3_U2897) );
  AOI22_X1 U22631 ( .A1(n19840), .A2(n19535), .B1(n19839), .B2(n19517), .ZN(
        n19515) );
  AOI22_X1 U22632 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19519), .B1(
        n19841), .B2(n19575), .ZN(n19514) );
  OAI211_X1 U22633 ( .C1(n19516), .C2(n19844), .A(n19515), .B(n19514), .ZN(
        P3_U2898) );
  AOI22_X1 U22634 ( .A1(n19518), .A2(n19789), .B1(n19846), .B2(n19517), .ZN(
        n19521) );
  AOI22_X1 U22635 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19519), .B1(
        n19849), .B2(n19575), .ZN(n19520) );
  OAI211_X1 U22636 ( .C1(n19794), .C2(n19544), .A(n19521), .B(n19520), .ZN(
        P3_U2899) );
  INV_X1 U22637 ( .A(n19611), .ZN(n19870) );
  NOR2_X2 U22638 ( .A1(n19870), .A2(n19566), .ZN(n19603) );
  INV_X1 U22639 ( .A(n19603), .ZN(n19610) );
  NOR2_X1 U22640 ( .A1(n19575), .A2(n19603), .ZN(n19567) );
  NOR2_X1 U22641 ( .A1(n19908), .A2(n19567), .ZN(n19540) );
  AOI22_X1 U22642 ( .A1(n19797), .A2(n19535), .B1(n19796), .B2(n19540), .ZN(
        n19526) );
  OAI22_X1 U22643 ( .A1(n19567), .A2(n19523), .B1(n19756), .B2(n19522), .ZN(
        n19524) );
  OAI21_X1 U22644 ( .B1(n19603), .B2(n20009), .A(n19524), .ZN(n19541) );
  AOI22_X1 U22645 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19541), .B1(
        n19802), .B2(n19554), .ZN(n19525) );
  OAI211_X1 U22646 ( .C1(n19805), .C2(n19610), .A(n19526), .B(n19525), .ZN(
        P3_U2900) );
  AOI22_X1 U22647 ( .A1(n19764), .A2(n19535), .B1(n19807), .B2(n19540), .ZN(
        n19528) );
  AOI22_X1 U22648 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19541), .B1(
        n19809), .B2(n19603), .ZN(n19527) );
  OAI211_X1 U22649 ( .C1(n19767), .C2(n19565), .A(n19528), .B(n19527), .ZN(
        P3_U2901) );
  AOI22_X1 U22650 ( .A1(n19768), .A2(n19554), .B1(n19813), .B2(n19540), .ZN(
        n19530) );
  AOI22_X1 U22651 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19541), .B1(
        n19815), .B2(n19603), .ZN(n19529) );
  OAI211_X1 U22652 ( .C1(n19771), .C2(n19544), .A(n19530), .B(n19529), .ZN(
        P3_U2902) );
  AOI22_X1 U22653 ( .A1(n19820), .A2(n19535), .B1(n19819), .B2(n19540), .ZN(
        n19532) );
  AOI22_X1 U22654 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19541), .B1(
        n19821), .B2(n19603), .ZN(n19531) );
  OAI211_X1 U22655 ( .C1(n19824), .C2(n19565), .A(n19532), .B(n19531), .ZN(
        P3_U2903) );
  AOI22_X1 U22656 ( .A1(n19826), .A2(n19554), .B1(n19825), .B2(n19540), .ZN(
        n19534) );
  AOI22_X1 U22657 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19541), .B1(
        n19827), .B2(n19603), .ZN(n19533) );
  OAI211_X1 U22658 ( .C1(n19830), .C2(n19544), .A(n19534), .B(n19533), .ZN(
        P3_U2904) );
  AOI22_X1 U22659 ( .A1(n19833), .A2(n19535), .B1(n19831), .B2(n19540), .ZN(
        n19537) );
  AOI22_X1 U22660 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19541), .B1(
        n19834), .B2(n19603), .ZN(n19536) );
  OAI211_X1 U22661 ( .C1(n19837), .C2(n19565), .A(n19537), .B(n19536), .ZN(
        P3_U2905) );
  AOI22_X1 U22662 ( .A1(n19840), .A2(n19554), .B1(n19839), .B2(n19540), .ZN(
        n19539) );
  AOI22_X1 U22663 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19541), .B1(
        n19841), .B2(n19603), .ZN(n19538) );
  OAI211_X1 U22664 ( .C1(n19844), .C2(n19544), .A(n19539), .B(n19538), .ZN(
        P3_U2906) );
  AOI22_X1 U22665 ( .A1(n19847), .A2(n19554), .B1(n19846), .B2(n19540), .ZN(
        n19543) );
  AOI22_X1 U22666 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19541), .B1(
        n19849), .B2(n19603), .ZN(n19542) );
  OAI211_X1 U22667 ( .C1(n19855), .C2(n19544), .A(n19543), .B(n19542), .ZN(
        P3_U2907) );
  NOR2_X1 U22668 ( .A1(n19636), .A2(n19566), .ZN(n19561) );
  AOI22_X1 U22669 ( .A1(n19802), .A2(n19575), .B1(n19796), .B2(n19561), .ZN(
        n19547) );
  AOI22_X1 U22670 ( .A1(n19801), .A2(n19545), .B1(n19730), .B2(n19590), .ZN(
        n19562) );
  NOR2_X2 U22671 ( .A1(n19638), .A2(n19566), .ZN(n19621) );
  AOI22_X1 U22672 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19562), .B1(
        n19760), .B2(n19621), .ZN(n19546) );
  OAI211_X1 U22673 ( .C1(n19763), .C2(n19565), .A(n19547), .B(n19546), .ZN(
        P3_U2908) );
  AOI22_X1 U22674 ( .A1(n19808), .A2(n19575), .B1(n19807), .B2(n19561), .ZN(
        n19549) );
  AOI22_X1 U22675 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19562), .B1(
        n19809), .B2(n19621), .ZN(n19548) );
  OAI211_X1 U22676 ( .C1(n19812), .C2(n19565), .A(n19549), .B(n19548), .ZN(
        P3_U2909) );
  AOI22_X1 U22677 ( .A1(n19768), .A2(n19575), .B1(n19813), .B2(n19561), .ZN(
        n19551) );
  AOI22_X1 U22678 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19562), .B1(
        n19815), .B2(n19621), .ZN(n19550) );
  OAI211_X1 U22679 ( .C1(n19771), .C2(n19565), .A(n19551), .B(n19550), .ZN(
        P3_U2910) );
  AOI22_X1 U22680 ( .A1(n19820), .A2(n19554), .B1(n19819), .B2(n19561), .ZN(
        n19553) );
  AOI22_X1 U22681 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19562), .B1(
        n19821), .B2(n19621), .ZN(n19552) );
  OAI211_X1 U22682 ( .C1(n19824), .C2(n19588), .A(n19553), .B(n19552), .ZN(
        P3_U2911) );
  AOI22_X1 U22683 ( .A1(n19742), .A2(n19554), .B1(n19825), .B2(n19561), .ZN(
        n19556) );
  AOI22_X1 U22684 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19562), .B1(
        n19827), .B2(n19621), .ZN(n19555) );
  OAI211_X1 U22685 ( .C1(n19745), .C2(n19588), .A(n19556), .B(n19555), .ZN(
        P3_U2912) );
  AOI22_X1 U22686 ( .A1(n19778), .A2(n19575), .B1(n19831), .B2(n19561), .ZN(
        n19558) );
  AOI22_X1 U22687 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19562), .B1(
        n19834), .B2(n19621), .ZN(n19557) );
  OAI211_X1 U22688 ( .C1(n19782), .C2(n19565), .A(n19558), .B(n19557), .ZN(
        P3_U2913) );
  AOI22_X1 U22689 ( .A1(n19840), .A2(n19575), .B1(n19839), .B2(n19561), .ZN(
        n19560) );
  AOI22_X1 U22690 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19562), .B1(
        n19841), .B2(n19621), .ZN(n19559) );
  OAI211_X1 U22691 ( .C1(n19844), .C2(n19565), .A(n19560), .B(n19559), .ZN(
        P3_U2914) );
  AOI22_X1 U22692 ( .A1(n19847), .A2(n19575), .B1(n19846), .B2(n19561), .ZN(
        n19564) );
  AOI22_X1 U22693 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19562), .B1(
        n19849), .B2(n19621), .ZN(n19563) );
  OAI211_X1 U22694 ( .C1(n19855), .C2(n19565), .A(n19564), .B(n19563), .ZN(
        P3_U2915) );
  NOR2_X1 U22695 ( .A1(n19866), .A2(n19566), .ZN(n19637) );
  NAND2_X1 U22696 ( .A1(n13148), .A2(n19637), .ZN(n19653) );
  NOR2_X1 U22697 ( .A1(n19621), .A2(n19655), .ZN(n19613) );
  NOR2_X1 U22698 ( .A1(n19908), .A2(n19613), .ZN(n19584) );
  AOI22_X1 U22699 ( .A1(n19802), .A2(n19603), .B1(n19796), .B2(n19584), .ZN(
        n19570) );
  OAI21_X1 U22700 ( .B1(n19567), .B2(n19756), .A(n19613), .ZN(n19568) );
  OAI211_X1 U22701 ( .C1(n19655), .C2(n20009), .A(n19759), .B(n19568), .ZN(
        n19585) );
  AOI22_X1 U22702 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19585), .B1(
        n19760), .B2(n19655), .ZN(n19569) );
  OAI211_X1 U22703 ( .C1(n19763), .C2(n19588), .A(n19570), .B(n19569), .ZN(
        P3_U2916) );
  AOI22_X1 U22704 ( .A1(n19764), .A2(n19575), .B1(n19807), .B2(n19584), .ZN(
        n19572) );
  AOI22_X1 U22705 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19585), .B1(
        n19809), .B2(n19655), .ZN(n19571) );
  OAI211_X1 U22706 ( .C1(n19767), .C2(n19610), .A(n19572), .B(n19571), .ZN(
        P3_U2917) );
  AOI22_X1 U22707 ( .A1(n19814), .A2(n19575), .B1(n19813), .B2(n19584), .ZN(
        n19574) );
  AOI22_X1 U22708 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19585), .B1(
        n19815), .B2(n19655), .ZN(n19573) );
  OAI211_X1 U22709 ( .C1(n19818), .C2(n19610), .A(n19574), .B(n19573), .ZN(
        P3_U2918) );
  AOI22_X1 U22710 ( .A1(n19820), .A2(n19575), .B1(n19819), .B2(n19584), .ZN(
        n19577) );
  AOI22_X1 U22711 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19585), .B1(
        n19821), .B2(n19655), .ZN(n19576) );
  OAI211_X1 U22712 ( .C1(n19824), .C2(n19610), .A(n19577), .B(n19576), .ZN(
        P3_U2919) );
  AOI22_X1 U22713 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19585), .B1(
        n19825), .B2(n19584), .ZN(n19579) );
  AOI22_X1 U22714 ( .A1(n19826), .A2(n19603), .B1(n19827), .B2(n19655), .ZN(
        n19578) );
  OAI211_X1 U22715 ( .C1(n19830), .C2(n19588), .A(n19579), .B(n19578), .ZN(
        P3_U2920) );
  AOI22_X1 U22716 ( .A1(n19778), .A2(n19603), .B1(n19831), .B2(n19584), .ZN(
        n19581) );
  AOI22_X1 U22717 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19585), .B1(
        n19834), .B2(n19655), .ZN(n19580) );
  OAI211_X1 U22718 ( .C1(n19782), .C2(n19588), .A(n19581), .B(n19580), .ZN(
        P3_U2921) );
  AOI22_X1 U22719 ( .A1(n19840), .A2(n19603), .B1(n19839), .B2(n19584), .ZN(
        n19583) );
  AOI22_X1 U22720 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19585), .B1(
        n19841), .B2(n19655), .ZN(n19582) );
  OAI211_X1 U22721 ( .C1(n19844), .C2(n19588), .A(n19583), .B(n19582), .ZN(
        P3_U2922) );
  AOI22_X1 U22722 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19585), .B1(
        n19846), .B2(n19584), .ZN(n19587) );
  AOI22_X1 U22723 ( .A1(n19847), .A2(n19603), .B1(n19849), .B2(n19655), .ZN(
        n19586) );
  OAI211_X1 U22724 ( .C1(n19855), .C2(n19588), .A(n19587), .B(n19586), .ZN(
        P3_U2923) );
  AND2_X1 U22725 ( .A1(n19729), .A2(n19637), .ZN(n19606) );
  AOI22_X1 U22726 ( .A1(n19802), .A2(n19621), .B1(n19796), .B2(n19606), .ZN(
        n19592) );
  NAND2_X1 U22727 ( .A1(n19589), .A2(n19590), .ZN(n19607) );
  NAND2_X1 U22728 ( .A1(n19864), .A2(n19590), .ZN(n19680) );
  INV_X1 U22729 ( .A(n19680), .ZN(n19671) );
  AOI22_X1 U22730 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19607), .B1(
        n19760), .B2(n19671), .ZN(n19591) );
  OAI211_X1 U22731 ( .C1(n19763), .C2(n19610), .A(n19592), .B(n19591), .ZN(
        P3_U2924) );
  AOI22_X1 U22732 ( .A1(n19764), .A2(n19603), .B1(n19807), .B2(n19606), .ZN(
        n19594) );
  AOI22_X1 U22733 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19607), .B1(
        n19809), .B2(n19671), .ZN(n19593) );
  OAI211_X1 U22734 ( .C1(n19767), .C2(n19634), .A(n19594), .B(n19593), .ZN(
        P3_U2925) );
  AOI22_X1 U22735 ( .A1(n19768), .A2(n19621), .B1(n19813), .B2(n19606), .ZN(
        n19596) );
  AOI22_X1 U22736 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19607), .B1(
        n19815), .B2(n19671), .ZN(n19595) );
  OAI211_X1 U22737 ( .C1(n19771), .C2(n19610), .A(n19596), .B(n19595), .ZN(
        P3_U2926) );
  AOI22_X1 U22738 ( .A1(n19820), .A2(n19603), .B1(n19819), .B2(n19606), .ZN(
        n19598) );
  AOI22_X1 U22739 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19607), .B1(
        n19821), .B2(n19671), .ZN(n19597) );
  OAI211_X1 U22740 ( .C1(n19824), .C2(n19634), .A(n19598), .B(n19597), .ZN(
        P3_U2927) );
  AOI22_X1 U22741 ( .A1(n19742), .A2(n19603), .B1(n19825), .B2(n19606), .ZN(
        n19600) );
  AOI22_X1 U22742 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19607), .B1(
        n19827), .B2(n19671), .ZN(n19599) );
  OAI211_X1 U22743 ( .C1(n19745), .C2(n19634), .A(n19600), .B(n19599), .ZN(
        P3_U2928) );
  AOI22_X1 U22744 ( .A1(n19833), .A2(n19603), .B1(n19831), .B2(n19606), .ZN(
        n19602) );
  AOI22_X1 U22745 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19607), .B1(
        n19834), .B2(n19671), .ZN(n19601) );
  OAI211_X1 U22746 ( .C1(n19837), .C2(n19634), .A(n19602), .B(n19601), .ZN(
        P3_U2929) );
  AOI22_X1 U22747 ( .A1(n19783), .A2(n19603), .B1(n19839), .B2(n19606), .ZN(
        n19605) );
  AOI22_X1 U22748 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19607), .B1(
        n19841), .B2(n19671), .ZN(n19604) );
  OAI211_X1 U22749 ( .C1(n19786), .C2(n19634), .A(n19605), .B(n19604), .ZN(
        P3_U2930) );
  AOI22_X1 U22750 ( .A1(n19847), .A2(n19621), .B1(n19846), .B2(n19606), .ZN(
        n19609) );
  AOI22_X1 U22751 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19607), .B1(
        n19849), .B2(n19671), .ZN(n19608) );
  OAI211_X1 U22752 ( .C1(n19855), .C2(n19610), .A(n19609), .B(n19608), .ZN(
        P3_U2931) );
  NAND2_X1 U22753 ( .A1(n19611), .A2(n19635), .ZN(n19696) );
  NOR2_X1 U22754 ( .A1(n19671), .A2(n19702), .ZN(n19659) );
  NOR2_X1 U22755 ( .A1(n19908), .A2(n19659), .ZN(n19630) );
  AOI22_X1 U22756 ( .A1(n19802), .A2(n19655), .B1(n19796), .B2(n19630), .ZN(
        n19616) );
  AOI221_X1 U22757 ( .B1(n19659), .B2(n19756), .C1(n19659), .C2(n19613), .A(
        n19612), .ZN(n19614) );
  INV_X1 U22758 ( .A(n19614), .ZN(n19631) );
  AOI22_X1 U22759 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19631), .B1(
        n19760), .B2(n19702), .ZN(n19615) );
  OAI211_X1 U22760 ( .C1(n19763), .C2(n19634), .A(n19616), .B(n19615), .ZN(
        P3_U2932) );
  AOI22_X1 U22761 ( .A1(n19808), .A2(n19655), .B1(n19807), .B2(n19630), .ZN(
        n19618) );
  AOI22_X1 U22762 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19631), .B1(
        n19809), .B2(n19702), .ZN(n19617) );
  OAI211_X1 U22763 ( .C1(n19812), .C2(n19634), .A(n19618), .B(n19617), .ZN(
        P3_U2933) );
  AOI22_X1 U22764 ( .A1(n19768), .A2(n19655), .B1(n19813), .B2(n19630), .ZN(
        n19620) );
  AOI22_X1 U22765 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19631), .B1(
        n19815), .B2(n19702), .ZN(n19619) );
  OAI211_X1 U22766 ( .C1(n19771), .C2(n19634), .A(n19620), .B(n19619), .ZN(
        P3_U2934) );
  AOI22_X1 U22767 ( .A1(n19820), .A2(n19621), .B1(n19819), .B2(n19630), .ZN(
        n19623) );
  AOI22_X1 U22768 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19631), .B1(
        n19821), .B2(n19702), .ZN(n19622) );
  OAI211_X1 U22769 ( .C1(n19824), .C2(n19653), .A(n19623), .B(n19622), .ZN(
        P3_U2935) );
  AOI22_X1 U22770 ( .A1(n19826), .A2(n19655), .B1(n19825), .B2(n19630), .ZN(
        n19625) );
  AOI22_X1 U22771 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19631), .B1(
        n19827), .B2(n19702), .ZN(n19624) );
  OAI211_X1 U22772 ( .C1(n19830), .C2(n19634), .A(n19625), .B(n19624), .ZN(
        P3_U2936) );
  AOI22_X1 U22773 ( .A1(n19778), .A2(n19655), .B1(n19831), .B2(n19630), .ZN(
        n19627) );
  AOI22_X1 U22774 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19631), .B1(
        n19834), .B2(n19702), .ZN(n19626) );
  OAI211_X1 U22775 ( .C1(n19782), .C2(n19634), .A(n19627), .B(n19626), .ZN(
        P3_U2937) );
  AOI22_X1 U22776 ( .A1(n19840), .A2(n19655), .B1(n19839), .B2(n19630), .ZN(
        n19629) );
  AOI22_X1 U22777 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19631), .B1(
        n19841), .B2(n19702), .ZN(n19628) );
  OAI211_X1 U22778 ( .C1(n19844), .C2(n19634), .A(n19629), .B(n19628), .ZN(
        P3_U2938) );
  AOI22_X1 U22779 ( .A1(n19847), .A2(n19655), .B1(n19846), .B2(n19630), .ZN(
        n19633) );
  AOI22_X1 U22780 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19631), .B1(
        n19849), .B2(n19702), .ZN(n19632) );
  OAI211_X1 U22781 ( .C1(n19855), .C2(n19634), .A(n19633), .B(n19632), .ZN(
        P3_U2939) );
  NOR2_X1 U22782 ( .A1(n19636), .A2(n19681), .ZN(n19654) );
  AOI22_X1 U22783 ( .A1(n19802), .A2(n19671), .B1(n19796), .B2(n19654), .ZN(
        n19640) );
  NOR2_X1 U22784 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19681), .ZN(
        n19683) );
  AOI22_X1 U22785 ( .A1(n19801), .A2(n19637), .B1(n19798), .B2(n19683), .ZN(
        n19656) );
  NOR2_X2 U22786 ( .A1(n19638), .A2(n19681), .ZN(n19717) );
  AOI22_X1 U22787 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19656), .B1(
        n19760), .B2(n19717), .ZN(n19639) );
  OAI211_X1 U22788 ( .C1(n19763), .C2(n19653), .A(n19640), .B(n19639), .ZN(
        P3_U2940) );
  AOI22_X1 U22789 ( .A1(n19808), .A2(n19671), .B1(n19807), .B2(n19654), .ZN(
        n19642) );
  AOI22_X1 U22790 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19656), .B1(
        n19809), .B2(n19717), .ZN(n19641) );
  OAI211_X1 U22791 ( .C1(n19812), .C2(n19653), .A(n19642), .B(n19641), .ZN(
        P3_U2941) );
  AOI22_X1 U22792 ( .A1(n19814), .A2(n19655), .B1(n19813), .B2(n19654), .ZN(
        n19644) );
  AOI22_X1 U22793 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19656), .B1(
        n19815), .B2(n19717), .ZN(n19643) );
  OAI211_X1 U22794 ( .C1(n19818), .C2(n19680), .A(n19644), .B(n19643), .ZN(
        P3_U2942) );
  AOI22_X1 U22795 ( .A1(n19772), .A2(n19671), .B1(n19819), .B2(n19654), .ZN(
        n19646) );
  AOI22_X1 U22796 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19656), .B1(
        n19821), .B2(n19717), .ZN(n19645) );
  OAI211_X1 U22797 ( .C1(n19775), .C2(n19653), .A(n19646), .B(n19645), .ZN(
        P3_U2943) );
  AOI22_X1 U22798 ( .A1(n19742), .A2(n19655), .B1(n19825), .B2(n19654), .ZN(
        n19648) );
  AOI22_X1 U22799 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19656), .B1(
        n19827), .B2(n19717), .ZN(n19647) );
  OAI211_X1 U22800 ( .C1(n19745), .C2(n19680), .A(n19648), .B(n19647), .ZN(
        P3_U2944) );
  AOI22_X1 U22801 ( .A1(n19778), .A2(n19671), .B1(n19831), .B2(n19654), .ZN(
        n19650) );
  AOI22_X1 U22802 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19656), .B1(
        n19834), .B2(n19717), .ZN(n19649) );
  OAI211_X1 U22803 ( .C1(n19782), .C2(n19653), .A(n19650), .B(n19649), .ZN(
        P3_U2945) );
  AOI22_X1 U22804 ( .A1(n19840), .A2(n19671), .B1(n19839), .B2(n19654), .ZN(
        n19652) );
  AOI22_X1 U22805 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19656), .B1(
        n19841), .B2(n19717), .ZN(n19651) );
  OAI211_X1 U22806 ( .C1(n19844), .C2(n19653), .A(n19652), .B(n19651), .ZN(
        P3_U2946) );
  AOI22_X1 U22807 ( .A1(n19789), .A2(n19655), .B1(n19846), .B2(n19654), .ZN(
        n19658) );
  AOI22_X1 U22808 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19656), .B1(
        n19849), .B2(n19717), .ZN(n19657) );
  OAI211_X1 U22809 ( .C1(n19794), .C2(n19680), .A(n19658), .B(n19657), .ZN(
        P3_U2947) );
  NOR2_X1 U22810 ( .A1(n19866), .A2(n19681), .ZN(n19732) );
  NAND2_X1 U22811 ( .A1(n13148), .A2(n19732), .ZN(n19754) );
  INV_X1 U22812 ( .A(n19754), .ZN(n19741) );
  NOR2_X1 U22813 ( .A1(n19717), .A2(n19741), .ZN(n19706) );
  OAI21_X1 U22814 ( .B1(n19659), .B2(n19756), .A(n19706), .ZN(n19660) );
  OAI211_X1 U22815 ( .C1(n19741), .C2(n20009), .A(n19759), .B(n19660), .ZN(
        n19677) );
  NOR2_X1 U22816 ( .A1(n19908), .A2(n19706), .ZN(n19676) );
  AOI22_X1 U22817 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19677), .B1(
        n19796), .B2(n19676), .ZN(n19662) );
  AOI22_X1 U22818 ( .A1(n19760), .A2(n19741), .B1(n19802), .B2(n19702), .ZN(
        n19661) );
  OAI211_X1 U22819 ( .C1(n19763), .C2(n19680), .A(n19662), .B(n19661), .ZN(
        P3_U2948) );
  AOI22_X1 U22820 ( .A1(n19808), .A2(n19702), .B1(n19807), .B2(n19676), .ZN(
        n19664) );
  AOI22_X1 U22821 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19677), .B1(
        n19809), .B2(n19741), .ZN(n19663) );
  OAI211_X1 U22822 ( .C1(n19812), .C2(n19680), .A(n19664), .B(n19663), .ZN(
        P3_U2949) );
  AOI22_X1 U22823 ( .A1(n19814), .A2(n19671), .B1(n19813), .B2(n19676), .ZN(
        n19666) );
  AOI22_X1 U22824 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19677), .B1(
        n19815), .B2(n19741), .ZN(n19665) );
  OAI211_X1 U22825 ( .C1(n19818), .C2(n19696), .A(n19666), .B(n19665), .ZN(
        P3_U2950) );
  AOI22_X1 U22826 ( .A1(n19820), .A2(n19671), .B1(n19819), .B2(n19676), .ZN(
        n19668) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19677), .B1(
        n19821), .B2(n19741), .ZN(n19667) );
  OAI211_X1 U22828 ( .C1(n19824), .C2(n19696), .A(n19668), .B(n19667), .ZN(
        P3_U2951) );
  AOI22_X1 U22829 ( .A1(n19826), .A2(n19702), .B1(n19825), .B2(n19676), .ZN(
        n19670) );
  AOI22_X1 U22830 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19677), .B1(
        n19827), .B2(n19741), .ZN(n19669) );
  OAI211_X1 U22831 ( .C1(n19830), .C2(n19680), .A(n19670), .B(n19669), .ZN(
        P3_U2952) );
  AOI22_X1 U22832 ( .A1(n19833), .A2(n19671), .B1(n19831), .B2(n19676), .ZN(
        n19673) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19677), .B1(
        n19834), .B2(n19741), .ZN(n19672) );
  OAI211_X1 U22834 ( .C1(n19837), .C2(n19696), .A(n19673), .B(n19672), .ZN(
        P3_U2953) );
  AOI22_X1 U22835 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19677), .B1(
        n19839), .B2(n19676), .ZN(n19675) );
  AOI22_X1 U22836 ( .A1(n19840), .A2(n19702), .B1(n19841), .B2(n19741), .ZN(
        n19674) );
  OAI211_X1 U22837 ( .C1(n19844), .C2(n19680), .A(n19675), .B(n19674), .ZN(
        P3_U2954) );
  AOI22_X1 U22838 ( .A1(n19847), .A2(n19702), .B1(n19846), .B2(n19676), .ZN(
        n19679) );
  AOI22_X1 U22839 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19677), .B1(
        n19849), .B2(n19741), .ZN(n19678) );
  OAI211_X1 U22840 ( .C1(n19855), .C2(n19680), .A(n19679), .B(n19678), .ZN(
        P3_U2955) );
  INV_X1 U22841 ( .A(n19864), .ZN(n19682) );
  NOR2_X2 U22842 ( .A1(n19682), .A2(n19681), .ZN(n19788) );
  AND2_X1 U22843 ( .A1(n19729), .A2(n19732), .ZN(n19701) );
  AOI22_X1 U22844 ( .A1(n19797), .A2(n19702), .B1(n19796), .B2(n19701), .ZN(
        n19685) );
  AOI22_X1 U22845 ( .A1(n19801), .A2(n19683), .B1(n19798), .B2(n19732), .ZN(
        n19703) );
  AOI22_X1 U22846 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19703), .B1(
        n19802), .B2(n19717), .ZN(n19684) );
  OAI211_X1 U22847 ( .C1(n19805), .C2(n19781), .A(n19685), .B(n19684), .ZN(
        P3_U2956) );
  INV_X1 U22848 ( .A(n19809), .ZN(n19688) );
  AOI22_X1 U22849 ( .A1(n19764), .A2(n19702), .B1(n19807), .B2(n19701), .ZN(
        n19687) );
  AOI22_X1 U22850 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19703), .B1(
        n19808), .B2(n19717), .ZN(n19686) );
  OAI211_X1 U22851 ( .C1(n19688), .C2(n19781), .A(n19687), .B(n19686), .ZN(
        P3_U2957) );
  INV_X1 U22852 ( .A(n19815), .ZN(n19714) );
  AOI22_X1 U22853 ( .A1(n19814), .A2(n19702), .B1(n19813), .B2(n19701), .ZN(
        n19690) );
  AOI22_X1 U22854 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19703), .B1(
        n19768), .B2(n19717), .ZN(n19689) );
  OAI211_X1 U22855 ( .C1(n19714), .C2(n19781), .A(n19690), .B(n19689), .ZN(
        P3_U2958) );
  INV_X1 U22856 ( .A(n19821), .ZN(n19693) );
  AOI22_X1 U22857 ( .A1(n19820), .A2(n19702), .B1(n19819), .B2(n19701), .ZN(
        n19692) );
  AOI22_X1 U22858 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19703), .B1(
        n19772), .B2(n19717), .ZN(n19691) );
  OAI211_X1 U22859 ( .C1(n19693), .C2(n19781), .A(n19692), .B(n19691), .ZN(
        P3_U2959) );
  AOI22_X1 U22860 ( .A1(n19826), .A2(n19717), .B1(n19825), .B2(n19701), .ZN(
        n19695) );
  AOI22_X1 U22861 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19703), .B1(
        n19827), .B2(n19788), .ZN(n19694) );
  OAI211_X1 U22862 ( .C1(n19830), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P3_U2960) );
  INV_X1 U22863 ( .A(n19717), .ZN(n19728) );
  AOI22_X1 U22864 ( .A1(n19833), .A2(n19702), .B1(n19831), .B2(n19701), .ZN(
        n19698) );
  AOI22_X1 U22865 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19703), .B1(
        n19834), .B2(n19788), .ZN(n19697) );
  OAI211_X1 U22866 ( .C1(n19837), .C2(n19728), .A(n19698), .B(n19697), .ZN(
        P3_U2961) );
  AOI22_X1 U22867 ( .A1(n19783), .A2(n19702), .B1(n19839), .B2(n19701), .ZN(
        n19700) );
  AOI22_X1 U22868 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19703), .B1(
        n19841), .B2(n19788), .ZN(n19699) );
  OAI211_X1 U22869 ( .C1(n19786), .C2(n19728), .A(n19700), .B(n19699), .ZN(
        P3_U2962) );
  AOI22_X1 U22870 ( .A1(n19789), .A2(n19702), .B1(n19846), .B2(n19701), .ZN(
        n19705) );
  AOI22_X1 U22871 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19703), .B1(
        n19849), .B2(n19788), .ZN(n19704) );
  OAI211_X1 U22872 ( .C1(n19794), .C2(n19728), .A(n19705), .B(n19704), .ZN(
        P3_U2963) );
  NAND2_X1 U22873 ( .A1(n19800), .A2(n13148), .ZN(n19854) );
  INV_X1 U22874 ( .A(n19854), .ZN(n19832) );
  NOR2_X1 U22875 ( .A1(n19788), .A2(n19832), .ZN(n19757) );
  NOR2_X1 U22876 ( .A1(n19908), .A2(n19757), .ZN(n19724) );
  AOI22_X1 U22877 ( .A1(n19797), .A2(n19717), .B1(n19796), .B2(n19724), .ZN(
        n19709) );
  OAI21_X1 U22878 ( .B1(n19706), .B2(n19756), .A(n19757), .ZN(n19707) );
  OAI211_X1 U22879 ( .C1(n19832), .C2(n20009), .A(n19759), .B(n19707), .ZN(
        n19725) );
  AOI22_X1 U22880 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19725), .B1(
        n19802), .B2(n19741), .ZN(n19708) );
  OAI211_X1 U22881 ( .C1(n19805), .C2(n19854), .A(n19709), .B(n19708), .ZN(
        P3_U2964) );
  AOI22_X1 U22882 ( .A1(n19808), .A2(n19741), .B1(n19807), .B2(n19724), .ZN(
        n19711) );
  AOI22_X1 U22883 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19725), .B1(
        n19809), .B2(n19832), .ZN(n19710) );
  OAI211_X1 U22884 ( .C1(n19812), .C2(n19728), .A(n19711), .B(n19710), .ZN(
        P3_U2965) );
  AOI22_X1 U22885 ( .A1(n19814), .A2(n19717), .B1(n19813), .B2(n19724), .ZN(
        n19713) );
  AOI22_X1 U22886 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19725), .B1(
        n19768), .B2(n19741), .ZN(n19712) );
  OAI211_X1 U22887 ( .C1(n19714), .C2(n19854), .A(n19713), .B(n19712), .ZN(
        P3_U2966) );
  AOI22_X1 U22888 ( .A1(n19772), .A2(n19741), .B1(n19819), .B2(n19724), .ZN(
        n19716) );
  AOI22_X1 U22889 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19725), .B1(
        n19821), .B2(n19832), .ZN(n19715) );
  OAI211_X1 U22890 ( .C1(n19775), .C2(n19728), .A(n19716), .B(n19715), .ZN(
        P3_U2967) );
  AOI22_X1 U22891 ( .A1(n19742), .A2(n19717), .B1(n19825), .B2(n19724), .ZN(
        n19719) );
  AOI22_X1 U22892 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19725), .B1(
        n19827), .B2(n19832), .ZN(n19718) );
  OAI211_X1 U22893 ( .C1(n19745), .C2(n19754), .A(n19719), .B(n19718), .ZN(
        P3_U2968) );
  AOI22_X1 U22894 ( .A1(n19778), .A2(n19741), .B1(n19831), .B2(n19724), .ZN(
        n19721) );
  AOI22_X1 U22895 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19725), .B1(
        n19834), .B2(n19832), .ZN(n19720) );
  OAI211_X1 U22896 ( .C1(n19782), .C2(n19728), .A(n19721), .B(n19720), .ZN(
        P3_U2969) );
  AOI22_X1 U22897 ( .A1(n19840), .A2(n19741), .B1(n19839), .B2(n19724), .ZN(
        n19723) );
  AOI22_X1 U22898 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19725), .B1(
        n19841), .B2(n19832), .ZN(n19722) );
  OAI211_X1 U22899 ( .C1(n19844), .C2(n19728), .A(n19723), .B(n19722), .ZN(
        P3_U2970) );
  AOI22_X1 U22900 ( .A1(n19847), .A2(n19741), .B1(n19846), .B2(n19724), .ZN(
        n19727) );
  AOI22_X1 U22901 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19725), .B1(
        n19849), .B2(n19832), .ZN(n19726) );
  OAI211_X1 U22902 ( .C1(n19855), .C2(n19728), .A(n19727), .B(n19726), .ZN(
        P3_U2971) );
  AND2_X1 U22903 ( .A1(n19729), .A2(n19800), .ZN(n19750) );
  AOI22_X1 U22904 ( .A1(n19797), .A2(n19741), .B1(n19796), .B2(n19750), .ZN(
        n19734) );
  AOI22_X1 U22905 ( .A1(n19801), .A2(n19732), .B1(n19731), .B2(n19730), .ZN(
        n19751) );
  AOI22_X1 U22906 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19751), .B1(
        n19802), .B2(n19788), .ZN(n19733) );
  OAI211_X1 U22907 ( .C1(n19838), .C2(n19805), .A(n19734), .B(n19733), .ZN(
        P3_U2972) );
  AOI22_X1 U22908 ( .A1(n19808), .A2(n19788), .B1(n19807), .B2(n19750), .ZN(
        n19736) );
  AOI22_X1 U22909 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19809), .ZN(n19735) );
  OAI211_X1 U22910 ( .C1(n19812), .C2(n19754), .A(n19736), .B(n19735), .ZN(
        P3_U2973) );
  AOI22_X1 U22911 ( .A1(n19768), .A2(n19788), .B1(n19813), .B2(n19750), .ZN(
        n19738) );
  AOI22_X1 U22912 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19815), .ZN(n19737) );
  OAI211_X1 U22913 ( .C1(n19771), .C2(n19754), .A(n19738), .B(n19737), .ZN(
        P3_U2974) );
  AOI22_X1 U22914 ( .A1(n19820), .A2(n19741), .B1(n19819), .B2(n19750), .ZN(
        n19740) );
  AOI22_X1 U22915 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19821), .ZN(n19739) );
  OAI211_X1 U22916 ( .C1(n19824), .C2(n19781), .A(n19740), .B(n19739), .ZN(
        P3_U2975) );
  AOI22_X1 U22917 ( .A1(n19742), .A2(n19741), .B1(n19825), .B2(n19750), .ZN(
        n19744) );
  AOI22_X1 U22918 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19827), .ZN(n19743) );
  OAI211_X1 U22919 ( .C1(n19745), .C2(n19781), .A(n19744), .B(n19743), .ZN(
        P3_U2976) );
  AOI22_X1 U22920 ( .A1(n19778), .A2(n19788), .B1(n19831), .B2(n19750), .ZN(
        n19747) );
  AOI22_X1 U22921 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19834), .ZN(n19746) );
  OAI211_X1 U22922 ( .C1(n19782), .C2(n19754), .A(n19747), .B(n19746), .ZN(
        P3_U2977) );
  AOI22_X1 U22923 ( .A1(n19840), .A2(n19788), .B1(n19839), .B2(n19750), .ZN(
        n19749) );
  AOI22_X1 U22924 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19841), .ZN(n19748) );
  OAI211_X1 U22925 ( .C1(n19844), .C2(n19754), .A(n19749), .B(n19748), .ZN(
        P3_U2978) );
  AOI22_X1 U22926 ( .A1(n19847), .A2(n19788), .B1(n19846), .B2(n19750), .ZN(
        n19753) );
  AOI22_X1 U22927 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19751), .B1(
        n19848), .B2(n19849), .ZN(n19752) );
  OAI211_X1 U22928 ( .C1(n19855), .C2(n19754), .A(n19753), .B(n19752), .ZN(
        P3_U2979) );
  NOR2_X1 U22929 ( .A1(n19908), .A2(n19755), .ZN(n19787) );
  AOI22_X1 U22930 ( .A1(n19802), .A2(n19832), .B1(n19796), .B2(n19787), .ZN(
        n19762) );
  OAI21_X1 U22931 ( .B1(n19757), .B2(n19756), .A(n19755), .ZN(n19758) );
  OAI211_X1 U22932 ( .C1(n19790), .C2(n20009), .A(n19759), .B(n19758), .ZN(
        n19791) );
  AOI22_X1 U22933 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19760), .ZN(n19761) );
  OAI211_X1 U22934 ( .C1(n19763), .C2(n19781), .A(n19762), .B(n19761), .ZN(
        P3_U2980) );
  AOI22_X1 U22935 ( .A1(n19764), .A2(n19788), .B1(n19807), .B2(n19787), .ZN(
        n19766) );
  AOI22_X1 U22936 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19809), .ZN(n19765) );
  OAI211_X1 U22937 ( .C1(n19767), .C2(n19854), .A(n19766), .B(n19765), .ZN(
        P3_U2981) );
  AOI22_X1 U22938 ( .A1(n19768), .A2(n19832), .B1(n19813), .B2(n19787), .ZN(
        n19770) );
  AOI22_X1 U22939 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19815), .ZN(n19769) );
  OAI211_X1 U22940 ( .C1(n19771), .C2(n19781), .A(n19770), .B(n19769), .ZN(
        P3_U2982) );
  AOI22_X1 U22941 ( .A1(n19772), .A2(n19832), .B1(n19819), .B2(n19787), .ZN(
        n19774) );
  AOI22_X1 U22942 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19821), .ZN(n19773) );
  OAI211_X1 U22943 ( .C1(n19775), .C2(n19781), .A(n19774), .B(n19773), .ZN(
        P3_U2983) );
  AOI22_X1 U22944 ( .A1(n19826), .A2(n19832), .B1(n19825), .B2(n19787), .ZN(
        n19777) );
  AOI22_X1 U22945 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19827), .ZN(n19776) );
  OAI211_X1 U22946 ( .C1(n19830), .C2(n19781), .A(n19777), .B(n19776), .ZN(
        P3_U2984) );
  AOI22_X1 U22947 ( .A1(n19778), .A2(n19832), .B1(n19831), .B2(n19787), .ZN(
        n19780) );
  AOI22_X1 U22948 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19834), .ZN(n19779) );
  OAI211_X1 U22949 ( .C1(n19782), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        P3_U2985) );
  AOI22_X1 U22950 ( .A1(n19783), .A2(n19788), .B1(n19839), .B2(n19787), .ZN(
        n19785) );
  AOI22_X1 U22951 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19841), .ZN(n19784) );
  OAI211_X1 U22952 ( .C1(n19786), .C2(n19854), .A(n19785), .B(n19784), .ZN(
        P3_U2986) );
  AOI22_X1 U22953 ( .A1(n19789), .A2(n19788), .B1(n19846), .B2(n19787), .ZN(
        n19793) );
  AOI22_X1 U22954 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19791), .B1(
        n19790), .B2(n19849), .ZN(n19792) );
  OAI211_X1 U22955 ( .C1(n19794), .C2(n19854), .A(n19793), .B(n19792), .ZN(
        P3_U2987) );
  INV_X1 U22956 ( .A(n19799), .ZN(n19795) );
  NOR2_X1 U22957 ( .A1(n19908), .A2(n19795), .ZN(n19845) );
  AOI22_X1 U22958 ( .A1(n19797), .A2(n19832), .B1(n19796), .B2(n19845), .ZN(
        n19804) );
  AOI22_X1 U22959 ( .A1(n19801), .A2(n19800), .B1(n19799), .B2(n19798), .ZN(
        n19851) );
  AOI22_X1 U22960 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19851), .B1(
        n19848), .B2(n19802), .ZN(n19803) );
  OAI211_X1 U22961 ( .C1(n19806), .C2(n19805), .A(n19804), .B(n19803), .ZN(
        P3_U2988) );
  AOI22_X1 U22962 ( .A1(n19848), .A2(n19808), .B1(n19807), .B2(n19845), .ZN(
        n19811) );
  AOI22_X1 U22963 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19809), .ZN(n19810) );
  OAI211_X1 U22964 ( .C1(n19812), .C2(n19854), .A(n19811), .B(n19810), .ZN(
        P3_U2989) );
  AOI22_X1 U22965 ( .A1(n19814), .A2(n19832), .B1(n19813), .B2(n19845), .ZN(
        n19817) );
  AOI22_X1 U22966 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19815), .ZN(n19816) );
  OAI211_X1 U22967 ( .C1(n19838), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P3_U2990) );
  AOI22_X1 U22968 ( .A1(n19820), .A2(n19832), .B1(n19819), .B2(n19845), .ZN(
        n19823) );
  AOI22_X1 U22969 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19821), .ZN(n19822) );
  OAI211_X1 U22970 ( .C1(n19838), .C2(n19824), .A(n19823), .B(n19822), .ZN(
        P3_U2991) );
  AOI22_X1 U22971 ( .A1(n19848), .A2(n19826), .B1(n19825), .B2(n19845), .ZN(
        n19829) );
  AOI22_X1 U22972 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19827), .ZN(n19828) );
  OAI211_X1 U22973 ( .C1(n19830), .C2(n19854), .A(n19829), .B(n19828), .ZN(
        P3_U2992) );
  AOI22_X1 U22974 ( .A1(n19833), .A2(n19832), .B1(n19831), .B2(n19845), .ZN(
        n19836) );
  AOI22_X1 U22975 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19834), .ZN(n19835) );
  OAI211_X1 U22976 ( .C1(n19838), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        P3_U2993) );
  AOI22_X1 U22977 ( .A1(n19848), .A2(n19840), .B1(n19839), .B2(n19845), .ZN(
        n19843) );
  AOI22_X1 U22978 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19841), .ZN(n19842) );
  OAI211_X1 U22979 ( .C1(n19844), .C2(n19854), .A(n19843), .B(n19842), .ZN(
        P3_U2994) );
  AOI22_X1 U22980 ( .A1(n19848), .A2(n19847), .B1(n19846), .B2(n19845), .ZN(
        n19853) );
  AOI22_X1 U22981 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19849), .ZN(n19852) );
  OAI211_X1 U22982 ( .C1(n19855), .C2(n19854), .A(n19853), .B(n19852), .ZN(
        P3_U2995) );
  NOR2_X1 U22983 ( .A1(P3_MORE_REG_SCAN_IN), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(
        n19859) );
  OAI211_X1 U22984 ( .C1(n19859), .C2(n19858), .A(n19857), .B(n19856), .ZN(
        n19893) );
  NAND2_X1 U22985 ( .A1(n19861), .A2(n19860), .ZN(n19891) );
  NOR2_X1 U22986 ( .A1(n19884), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n19862) );
  AOI21_X1 U22987 ( .B1(n19863), .B2(n19884), .A(n19862), .ZN(n19888) );
  NAND2_X1 U22988 ( .A1(n19865), .A2(n19864), .ZN(n19868) );
  INV_X1 U22989 ( .A(n19865), .ZN(n19867) );
  AOI22_X1 U22990 ( .A1(n19869), .A2(n19868), .B1(n19867), .B2(n19866), .ZN(
        n19871) );
  OAI21_X1 U22991 ( .B1(n19871), .B2(n19894), .A(n19870), .ZN(n19881) );
  AND2_X1 U22992 ( .A1(n19881), .A2(n19882), .ZN(n19872) );
  OAI22_X1 U22993 ( .A1(n19888), .A2(n19872), .B1(n19882), .B2(n19881), .ZN(
        n19890) );
  AOI221_X1 U22994 ( .B1(n19876), .B2(n19875), .C1(n19874), .C2(n19875), .A(
        n19873), .ZN(n19877) );
  AOI221_X1 U22995 ( .B1(n19880), .B2(n19879), .C1(n19878), .C2(n19879), .A(
        n19877), .ZN(n20021) );
  NAND2_X1 U22996 ( .A1(n19882), .A2(n19881), .ZN(n19883) );
  AOI21_X1 U22997 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n19883), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19887) );
  MUX2_X1 U22998 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n19885), .S(
        n19884), .Z(n19886) );
  OAI21_X1 U22999 ( .B1(n19888), .B2(n19887), .A(n19886), .ZN(n19889) );
  OAI211_X1 U23000 ( .C1(n19891), .C2(n19890), .A(n20021), .B(n19889), .ZN(
        n19892) );
  AOI211_X1 U23001 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19894), .A(
        n19893), .B(n19892), .ZN(n19907) );
  NAND2_X1 U23002 ( .A1(n20039), .A2(n19895), .ZN(n19916) );
  INV_X1 U23003 ( .A(n19916), .ZN(n20033) );
  AOI22_X1 U23004 ( .A1(n19896), .A2(n20033), .B1(n20028), .B2(n18675), .ZN(
        n19897) );
  INV_X1 U23005 ( .A(n19897), .ZN(n19902) );
  OAI211_X1 U23006 ( .C1(n19899), .C2(n19898), .A(n20026), .B(n19907), .ZN(
        n20008) );
  OAI21_X1 U23007 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n20023), .A(n20008), 
        .ZN(n19909) );
  NOR2_X1 U23008 ( .A1(n19900), .A2(n19909), .ZN(n19901) );
  MUX2_X1 U23009 ( .A(n19902), .B(n19901), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19905) );
  INV_X1 U23010 ( .A(n19903), .ZN(n19904) );
  OAI211_X1 U23011 ( .C1(n19907), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P3_U2996) );
  NAND2_X1 U23012 ( .A1(n20028), .A2(n18675), .ZN(n19912) );
  NAND4_X1 U23013 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n20028), .A4(n20039), .ZN(n19914) );
  OR3_X1 U23014 ( .A1(n19910), .A2(n19909), .A3(n19908), .ZN(n19911) );
  NAND4_X1 U23015 ( .A1(n19913), .A2(n19912), .A3(n19914), .A4(n19911), .ZN(
        P3_U2997) );
  AND4_X1 U23016 ( .A1(n19916), .A2(n19915), .A3(n19914), .A4(n20007), .ZN(
        P3_U2998) );
  AND2_X1 U23017 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20003), .ZN(
        P3_U2999) );
  AND2_X1 U23018 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20003), .ZN(
        P3_U3000) );
  AND2_X1 U23019 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20003), .ZN(
        P3_U3001) );
  AND2_X1 U23020 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20003), .ZN(
        P3_U3002) );
  AND2_X1 U23021 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20003), .ZN(
        P3_U3003) );
  AND2_X1 U23022 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20003), .ZN(
        P3_U3004) );
  AND2_X1 U23023 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n20003), .ZN(
        P3_U3005) );
  AND2_X1 U23024 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n20003), .ZN(
        P3_U3006) );
  AND2_X1 U23025 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20003), .ZN(
        P3_U3007) );
  AND2_X1 U23026 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20003), .ZN(
        P3_U3008) );
  AND2_X1 U23027 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n20003), .ZN(
        P3_U3009) );
  AND2_X1 U23028 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20003), .ZN(
        P3_U3010) );
  AND2_X1 U23029 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20003), .ZN(
        P3_U3011) );
  AND2_X1 U23030 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20003), .ZN(
        P3_U3012) );
  AND2_X1 U23031 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20003), .ZN(
        P3_U3013) );
  AND2_X1 U23032 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20003), .ZN(
        P3_U3014) );
  AND2_X1 U23033 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20003), .ZN(
        P3_U3015) );
  AND2_X1 U23034 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20003), .ZN(
        P3_U3016) );
  AND2_X1 U23035 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20003), .ZN(
        P3_U3017) );
  AND2_X1 U23036 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20003), .ZN(
        P3_U3018) );
  AND2_X1 U23037 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20003), .ZN(
        P3_U3019) );
  AND2_X1 U23038 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n20003), .ZN(
        P3_U3020) );
  AND2_X1 U23039 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20003), .ZN(P3_U3021) );
  AND2_X1 U23040 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20003), .ZN(P3_U3022) );
  AND2_X1 U23041 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20003), .ZN(P3_U3023) );
  AND2_X1 U23042 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20003), .ZN(P3_U3024) );
  AND2_X1 U23043 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n20003), .ZN(P3_U3025) );
  AND2_X1 U23044 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20003), .ZN(P3_U3026) );
  AND2_X1 U23045 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20003), .ZN(P3_U3027) );
  AND2_X1 U23046 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20003), .ZN(P3_U3028) );
  AOI21_X1 U23047 ( .B1(HOLD), .B2(n19917), .A(n20035), .ZN(n19920) );
  NOR2_X1 U23048 ( .A1(n19918), .A2(n20023), .ZN(n19927) );
  OAI21_X1 U23049 ( .B1(n19927), .B2(n19932), .A(n19934), .ZN(n19919) );
  NAND3_X1 U23050 ( .A1(NA), .A2(n19918), .A3(n19932), .ZN(n19926) );
  OAI211_X1 U23051 ( .C1(n20018), .C2(n19920), .A(n19919), .B(n19926), .ZN(
        P3_U3029) );
  INV_X1 U23052 ( .A(HOLD), .ZN(n19925) );
  NOR2_X1 U23053 ( .A1(n19934), .A2(n19925), .ZN(n19930) );
  NOR3_X1 U23054 ( .A1(n19930), .A2(n19932), .A3(n20035), .ZN(n19921) );
  NOR2_X1 U23055 ( .A1(n19921), .A2(n19927), .ZN(n19923) );
  OAI211_X1 U23056 ( .C1(n19925), .C2(n19924), .A(n19923), .B(n19922), .ZN(
        P3_U3030) );
  AOI21_X1 U23057 ( .B1(n19932), .B2(n19926), .A(n19927), .ZN(n19933) );
  INV_X1 U23058 ( .A(n19927), .ZN(n19928) );
  OAI22_X1 U23059 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19928), .ZN(n19929) );
  OAI22_X1 U23060 ( .A1(n19930), .A2(n19929), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19931) );
  OAI22_X1 U23061 ( .A1(n19933), .A2(n19934), .B1(n19932), .B2(n19931), .ZN(
        P3_U3031) );
  INV_X1 U23062 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19936) );
  OAI222_X1 U23063 ( .A1(n20010), .A2(n19996), .B1(n19935), .B2(n20018), .C1(
        n19936), .C2(n19982), .ZN(P3_U3032) );
  OAI222_X1 U23064 ( .A1(n19982), .A2(n19938), .B1(n19937), .B2(n20018), .C1(
        n19936), .C2(n19996), .ZN(P3_U3033) );
  OAI222_X1 U23065 ( .A1(n19982), .A2(n19940), .B1(n19939), .B2(n20018), .C1(
        n19938), .C2(n19996), .ZN(P3_U3034) );
  OAI222_X1 U23066 ( .A1(n19982), .A2(n19943), .B1(n19941), .B2(n20018), .C1(
        n19940), .C2(n19996), .ZN(P3_U3035) );
  OAI222_X1 U23067 ( .A1(n19943), .A2(n19996), .B1(n19942), .B2(n20018), .C1(
        n19944), .C2(n19982), .ZN(P3_U3036) );
  OAI222_X1 U23068 ( .A1(n19982), .A2(n19946), .B1(n19945), .B2(n20018), .C1(
        n19944), .C2(n19996), .ZN(P3_U3037) );
  OAI222_X1 U23069 ( .A1(n19982), .A2(n19949), .B1(n19947), .B2(n20018), .C1(
        n19946), .C2(n19996), .ZN(P3_U3038) );
  OAI222_X1 U23070 ( .A1(n19949), .A2(n19996), .B1(n19948), .B2(n20018), .C1(
        n19950), .C2(n19982), .ZN(P3_U3039) );
  OAI222_X1 U23071 ( .A1(n19982), .A2(n19952), .B1(n19951), .B2(n20018), .C1(
        n19950), .C2(n19996), .ZN(P3_U3040) );
  OAI222_X1 U23072 ( .A1(n19982), .A2(n19954), .B1(n19953), .B2(n20018), .C1(
        n19952), .C2(n19996), .ZN(P3_U3041) );
  OAI222_X1 U23073 ( .A1(n19982), .A2(n19956), .B1(n19955), .B2(n20018), .C1(
        n19954), .C2(n19996), .ZN(P3_U3042) );
  OAI222_X1 U23074 ( .A1(n19982), .A2(n19958), .B1(n19957), .B2(n20018), .C1(
        n19956), .C2(n19996), .ZN(P3_U3043) );
  INV_X1 U23075 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19961) );
  OAI222_X1 U23076 ( .A1(n19982), .A2(n19961), .B1(n19959), .B2(n20018), .C1(
        n19958), .C2(n19996), .ZN(P3_U3044) );
  INV_X1 U23077 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19962) );
  OAI222_X1 U23078 ( .A1(n19961), .A2(n19996), .B1(n19960), .B2(n20018), .C1(
        n19962), .C2(n19982), .ZN(P3_U3045) );
  INV_X1 U23079 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19965) );
  OAI222_X1 U23080 ( .A1(n19982), .A2(n19965), .B1(n19963), .B2(n20018), .C1(
        n19962), .C2(n19996), .ZN(P3_U3046) );
  OAI222_X1 U23081 ( .A1(n19996), .A2(n19965), .B1(n19964), .B2(n20018), .C1(
        n19966), .C2(n19982), .ZN(P3_U3047) );
  OAI222_X1 U23082 ( .A1(n19982), .A2(n19968), .B1(n19967), .B2(n20018), .C1(
        n19966), .C2(n19996), .ZN(P3_U3048) );
  OAI222_X1 U23083 ( .A1(n19982), .A2(n19970), .B1(n19969), .B2(n20018), .C1(
        n19968), .C2(n19996), .ZN(P3_U3049) );
  OAI222_X1 U23084 ( .A1(n19982), .A2(n19972), .B1(n19971), .B2(n20018), .C1(
        n19970), .C2(n19996), .ZN(P3_U3050) );
  OAI222_X1 U23085 ( .A1(n19982), .A2(n19974), .B1(n19973), .B2(n20018), .C1(
        n19972), .C2(n19996), .ZN(P3_U3051) );
  OAI222_X1 U23086 ( .A1(n19982), .A2(n19976), .B1(n19975), .B2(n20018), .C1(
        n19974), .C2(n19996), .ZN(P3_U3052) );
  INV_X1 U23087 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19979) );
  OAI222_X1 U23088 ( .A1(n19982), .A2(n19979), .B1(n19977), .B2(n20018), .C1(
        n19976), .C2(n19996), .ZN(P3_U3053) );
  OAI222_X1 U23089 ( .A1(n19979), .A2(n19996), .B1(n19978), .B2(n20018), .C1(
        n19980), .C2(n19982), .ZN(P3_U3054) );
  INV_X1 U23090 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19984) );
  OAI222_X1 U23091 ( .A1(n19982), .A2(n19984), .B1(n19981), .B2(n20018), .C1(
        n19980), .C2(n19996), .ZN(P3_U3055) );
  OAI222_X1 U23092 ( .A1(n19984), .A2(n19996), .B1(n19983), .B2(n20018), .C1(
        n19985), .C2(n19982), .ZN(P3_U3056) );
  OAI222_X1 U23093 ( .A1(n19982), .A2(n19987), .B1(n19986), .B2(n20018), .C1(
        n19985), .C2(n19996), .ZN(P3_U3057) );
  OAI222_X1 U23094 ( .A1(n19982), .A2(n19990), .B1(n19988), .B2(n20018), .C1(
        n19987), .C2(n19996), .ZN(P3_U3058) );
  OAI222_X1 U23095 ( .A1(n19990), .A2(n19996), .B1(n19989), .B2(n20018), .C1(
        n19991), .C2(n19982), .ZN(P3_U3059) );
  OAI222_X1 U23096 ( .A1(n19982), .A2(n19995), .B1(n19992), .B2(n20018), .C1(
        n19991), .C2(n19996), .ZN(P3_U3060) );
  OAI222_X1 U23097 ( .A1(n19996), .A2(n19995), .B1(n19994), .B2(n20018), .C1(
        n19993), .C2(n19982), .ZN(P3_U3061) );
  OAI22_X1 U23098 ( .A1(n20037), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n20018), .ZN(n19997) );
  INV_X1 U23099 ( .A(n19997), .ZN(P3_U3274) );
  OAI22_X1 U23100 ( .A1(n20037), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n20018), .ZN(n19998) );
  INV_X1 U23101 ( .A(n19998), .ZN(P3_U3275) );
  OAI22_X1 U23102 ( .A1(n20037), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n20018), .ZN(n19999) );
  INV_X1 U23103 ( .A(n19999), .ZN(P3_U3276) );
  OAI22_X1 U23104 ( .A1(n20037), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n20018), .ZN(n20000) );
  INV_X1 U23105 ( .A(n20000), .ZN(P3_U3277) );
  INV_X1 U23106 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20002) );
  INV_X1 U23107 ( .A(n20004), .ZN(n20001) );
  AOI21_X1 U23108 ( .B1(n20003), .B2(n20002), .A(n20001), .ZN(P3_U3280) );
  OAI21_X1 U23109 ( .B1(n20006), .B2(n20005), .A(n20004), .ZN(P3_U3281) );
  OAI221_X1 U23110 ( .B1(n20009), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n20009), 
        .C2(n20008), .A(n20007), .ZN(P3_U3282) );
  AOI21_X1 U23111 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20011) );
  AOI22_X1 U23112 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n20011), .B2(n20010), .ZN(n20014) );
  INV_X1 U23113 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U23114 ( .A1(n20017), .A2(n20014), .B1(n20013), .B2(n20012), .ZN(
        P3_U3292) );
  INV_X1 U23115 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20016) );
  OAI21_X1 U23116 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n20017), .ZN(n20015) );
  OAI21_X1 U23117 ( .B1(n20017), .B2(n20016), .A(n20015), .ZN(P3_U3293) );
  INV_X1 U23118 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20043) );
  OAI22_X1 U23119 ( .A1(n20037), .A2(n20043), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n20018), .ZN(n20019) );
  INV_X1 U23120 ( .A(n20019), .ZN(P3_U3294) );
  NAND2_X1 U23121 ( .A1(n20022), .A2(P3_MORE_REG_SCAN_IN), .ZN(n20020) );
  OAI21_X1 U23122 ( .B1(n20022), .B2(n20021), .A(n20020), .ZN(P3_U3295) );
  AOI21_X1 U23123 ( .B1(n18675), .B2(n20023), .A(n20042), .ZN(n20024) );
  OAI21_X1 U23124 ( .B1(n20026), .B2(n20025), .A(n20024), .ZN(n20036) );
  OAI21_X1 U23125 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n14057), .A(n20027), 
        .ZN(n20029) );
  AOI211_X1 U23126 ( .C1(n20041), .C2(n20029), .A(n20028), .B(n20039), .ZN(
        n20031) );
  NOR2_X1 U23127 ( .A1(n20031), .A2(n20030), .ZN(n20032) );
  OAI21_X1 U23128 ( .B1(n20033), .B2(n20032), .A(n20036), .ZN(n20034) );
  OAI21_X1 U23129 ( .B1(n20036), .B2(n20035), .A(n20034), .ZN(P3_U3296) );
  OAI22_X1 U23130 ( .A1(n20037), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n20018), .ZN(n20038) );
  INV_X1 U23131 ( .A(n20038), .ZN(P3_U3297) );
  AOI21_X1 U23132 ( .B1(n20040), .B2(n20039), .A(n20042), .ZN(n20046) );
  AOI22_X1 U23133 ( .A1(n20046), .A2(n20043), .B1(n20042), .B2(n20041), .ZN(
        P3_U3298) );
  INV_X1 U23134 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20045) );
  AOI21_X1 U23135 ( .B1(n20046), .B2(n20045), .A(n20044), .ZN(P3_U3299) );
  NAND2_X1 U23136 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20806), .ZN(n20796) );
  AOI22_X1 U23137 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20796), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20789), .ZN(n20867) );
  AOI21_X1 U23138 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20867), .ZN(n20047) );
  INV_X1 U23139 ( .A(n20047), .ZN(P2_U2815) );
  NAND2_X1 U23140 ( .A1(n20789), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20924) );
  NAND2_X1 U23141 ( .A1(n20049), .A2(n20924), .ZN(n20792) );
  AOI21_X1 U23142 ( .B1(n20789), .B2(n20792), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n20048) );
  AOI21_X1 U23143 ( .B1(n20856), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n20048), 
        .ZN(P2_U2817) );
  INV_X1 U23144 ( .A(n20049), .ZN(n20798) );
  OAI21_X1 U23145 ( .B1(n20798), .B2(BS16), .A(n20867), .ZN(n20865) );
  OAI21_X1 U23146 ( .B1(n20867), .B2(n20050), .A(n20865), .ZN(P2_U2818) );
  NOR4_X1 U23147 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20054) );
  NOR4_X1 U23148 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20053) );
  NOR4_X1 U23149 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20052) );
  NOR4_X1 U23150 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20051) );
  NAND4_X1 U23151 ( .A1(n20054), .A2(n20053), .A3(n20052), .A4(n20051), .ZN(
        n20060) );
  NOR4_X1 U23152 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20058) );
  AOI211_X1 U23153 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20057) );
  NOR4_X1 U23154 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20056) );
  NOR4_X1 U23155 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20055) );
  NAND4_X1 U23156 ( .A1(n20058), .A2(n20057), .A3(n20056), .A4(n20055), .ZN(
        n20059) );
  NOR2_X1 U23157 ( .A1(n20060), .A2(n20059), .ZN(n20070) );
  INV_X1 U23158 ( .A(n20070), .ZN(n20068) );
  NOR2_X1 U23159 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n20068), .ZN(n20062) );
  AOI22_X1 U23160 ( .A1(n20062), .A2(n20063), .B1(n20061), .B2(n20068), .ZN(
        P2_U2820) );
  OR3_X1 U23161 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20067) );
  INV_X1 U23162 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U23163 ( .A1(n20062), .A2(n20067), .B1(n20068), .B2(n20862), .ZN(
        P2_U2821) );
  INV_X1 U23164 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U23165 ( .A1(n20062), .A2(n20866), .ZN(n20066) );
  OAI21_X1 U23166 ( .B1(n20063), .B2(n20808), .A(n20070), .ZN(n20064) );
  OAI21_X1 U23167 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20070), .A(n20064), 
        .ZN(n20065) );
  OAI221_X1 U23168 ( .B1(n20066), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20066), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20065), .ZN(P2_U2822) );
  INV_X1 U23169 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20069) );
  OAI221_X1 U23170 ( .B1(n20070), .B2(n20069), .C1(n20068), .C2(n20067), .A(
        n20066), .ZN(P2_U2823) );
  OAI22_X1 U23171 ( .A1(n20074), .A2(n20073), .B1(n20072), .B2(n20071), .ZN(
        n20075) );
  AOI211_X1 U23172 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n20076), .A(n20179), .B(
        n20075), .ZN(n20091) );
  OR2_X1 U23173 ( .A1(n20078), .A2(n20077), .ZN(n20086) );
  NOR2_X1 U23174 ( .A1(n20080), .A2(n20079), .ZN(n20082) );
  XNOR2_X1 U23175 ( .A(n20082), .B(n20081), .ZN(n20084) );
  NAND2_X1 U23176 ( .A1(n20084), .A2(n20083), .ZN(n20085) );
  OAI211_X1 U23177 ( .C1(n20088), .C2(n20087), .A(n20086), .B(n20085), .ZN(
        n20089) );
  INV_X1 U23178 ( .A(n20089), .ZN(n20090) );
  OAI211_X1 U23179 ( .C1(n10301), .C2(n20092), .A(n20091), .B(n20090), .ZN(
        P2_U2849) );
  XNOR2_X1 U23180 ( .A(n20094), .B(n20093), .ZN(n20096) );
  AOI22_X1 U23181 ( .A1(n20096), .A2(n20108), .B1(n20112), .B2(n20095), .ZN(
        n20097) );
  OAI21_X1 U23182 ( .B1(n20112), .B2(n20098), .A(n20097), .ZN(P2_U2875) );
  INV_X1 U23183 ( .A(n20099), .ZN(n20102) );
  AOI211_X1 U23184 ( .C1(n20103), .C2(n20102), .A(n20101), .B(n20100), .ZN(
        n20104) );
  AOI21_X1 U23185 ( .B1(n20105), .B2(n20112), .A(n20104), .ZN(n20106) );
  OAI21_X1 U23186 ( .B1(n20112), .B2(n20107), .A(n20106), .ZN(P2_U2877) );
  INV_X1 U23187 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U23188 ( .A1(n20109), .A2(n20108), .B1(n20112), .B2(n20181), .ZN(
        n20110) );
  OAI21_X1 U23189 ( .B1(n20112), .B2(n20111), .A(n20110), .ZN(P2_U2883) );
  AOI22_X1 U23190 ( .A1(n20114), .A2(n20113), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n20133), .ZN(n20123) );
  AOI22_X1 U23191 ( .A1(n20116), .A2(BUF1_REG_16__SCAN_IN), .B1(n20115), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n20122) );
  INV_X1 U23192 ( .A(n20117), .ZN(n20120) );
  INV_X1 U23193 ( .A(n20118), .ZN(n20119) );
  AOI22_X1 U23194 ( .A1(n20120), .A2(n20134), .B1(n20128), .B2(n20119), .ZN(
        n20121) );
  NAND3_X1 U23195 ( .A1(n20123), .A2(n20122), .A3(n20121), .ZN(P2_U2903) );
  INV_X1 U23196 ( .A(n20124), .ZN(n20125) );
  AOI22_X1 U23197 ( .A1(n20125), .A2(n20134), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20133), .ZN(n20131) );
  XNOR2_X1 U23198 ( .A(n20127), .B(n20126), .ZN(n20129) );
  NAND2_X1 U23199 ( .A1(n20129), .A2(n20128), .ZN(n20130) );
  OAI211_X1 U23200 ( .C1(n20132), .C2(n20142), .A(n20131), .B(n20130), .ZN(
        P2_U2915) );
  AOI22_X1 U23201 ( .A1(n20134), .A2(n20878), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20133), .ZN(n20141) );
  AOI21_X1 U23202 ( .B1(n20137), .B2(n20136), .A(n20135), .ZN(n20139) );
  OR2_X1 U23203 ( .A1(n20139), .A2(n20138), .ZN(n20140) );
  OAI211_X1 U23204 ( .C1(n20143), .C2(n20142), .A(n20141), .B(n20140), .ZN(
        P2_U2916) );
  NOR2_X1 U23205 ( .A1(n20145), .A2(n20144), .ZN(P2_U2920) );
  AOI22_X1 U23206 ( .A1(n20176), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n20146) );
  OAI21_X1 U23207 ( .B1(n13672), .B2(n20178), .A(n20146), .ZN(P2_U2936) );
  AOI22_X1 U23208 ( .A1(n20176), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n20147) );
  OAI21_X1 U23209 ( .B1(n20148), .B2(n20178), .A(n20147), .ZN(P2_U2937) );
  AOI22_X1 U23210 ( .A1(n20176), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n20149) );
  OAI21_X1 U23211 ( .B1(n20150), .B2(n20178), .A(n20149), .ZN(P2_U2938) );
  AOI22_X1 U23212 ( .A1(n20176), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n20151) );
  OAI21_X1 U23213 ( .B1(n20152), .B2(n20178), .A(n20151), .ZN(P2_U2939) );
  AOI22_X1 U23214 ( .A1(n20176), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n20153) );
  OAI21_X1 U23215 ( .B1(n20154), .B2(n20178), .A(n20153), .ZN(P2_U2940) );
  AOI22_X1 U23216 ( .A1(n20176), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n20155) );
  OAI21_X1 U23217 ( .B1(n20156), .B2(n20178), .A(n20155), .ZN(P2_U2941) );
  AOI22_X1 U23218 ( .A1(n20176), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U23219 ( .B1(n20158), .B2(n20178), .A(n20157), .ZN(P2_U2942) );
  AOI22_X1 U23220 ( .A1(n20176), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n20159) );
  OAI21_X1 U23221 ( .B1(n20160), .B2(n20178), .A(n20159), .ZN(P2_U2943) );
  AOI22_X1 U23222 ( .A1(n20176), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n20161) );
  OAI21_X1 U23223 ( .B1(n20162), .B2(n20178), .A(n20161), .ZN(P2_U2944) );
  AOI22_X1 U23224 ( .A1(n20176), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n20163) );
  OAI21_X1 U23225 ( .B1(n20164), .B2(n20178), .A(n20163), .ZN(P2_U2945) );
  INV_X1 U23226 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U23227 ( .A1(n20176), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n20165) );
  OAI21_X1 U23228 ( .B1(n20166), .B2(n20178), .A(n20165), .ZN(P2_U2946) );
  INV_X1 U23229 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20168) );
  AOI22_X1 U23230 ( .A1(n20176), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n20167) );
  OAI21_X1 U23231 ( .B1(n20168), .B2(n20178), .A(n20167), .ZN(P2_U2947) );
  INV_X1 U23232 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20170) );
  AOI22_X1 U23233 ( .A1(n20176), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n20169) );
  OAI21_X1 U23234 ( .B1(n20170), .B2(n20178), .A(n20169), .ZN(P2_U2948) );
  AOI22_X1 U23235 ( .A1(n20176), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n20171) );
  OAI21_X1 U23236 ( .B1(n20172), .B2(n20178), .A(n20171), .ZN(P2_U2949) );
  AOI22_X1 U23237 ( .A1(n20176), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n20173) );
  OAI21_X1 U23238 ( .B1(n20174), .B2(n20178), .A(n20173), .ZN(P2_U2950) );
  AOI22_X1 U23239 ( .A1(n20176), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n20175), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n20177) );
  OAI21_X1 U23240 ( .B1(n11299), .B2(n20178), .A(n20177), .ZN(P2_U2951) );
  AOI22_X1 U23241 ( .A1(n20204), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n20179), .ZN(n20184) );
  AOI222_X1 U23242 ( .A1(n20182), .A2(n20196), .B1(n20213), .B2(n20181), .C1(
        n20180), .C2(n20205), .ZN(n20183) );
  OAI211_X1 U23243 ( .C1(n20199), .C2(n20185), .A(n20184), .B(n20183), .ZN(
        P2_U3010) );
  XNOR2_X1 U23244 ( .A(n20186), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20188) );
  XNOR2_X1 U23245 ( .A(n20188), .B(n20187), .ZN(n20226) );
  OAI21_X1 U23246 ( .B1(n20191), .B2(n20190), .A(n20189), .ZN(n20220) );
  INV_X1 U23247 ( .A(n20220), .ZN(n20192) );
  NOR2_X1 U23248 ( .A1(n20207), .A2(n20809), .ZN(n20223) );
  AOI21_X1 U23249 ( .B1(n20192), .B2(n20205), .A(n20223), .ZN(n20193) );
  OAI21_X1 U23250 ( .B1(n20221), .B2(n20194), .A(n20193), .ZN(n20195) );
  AOI21_X1 U23251 ( .B1(n20196), .B2(n20226), .A(n20195), .ZN(n20198) );
  NAND2_X1 U23252 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20204), .ZN(
        n20197) );
  OAI211_X1 U23253 ( .C1(n20200), .C2(n20199), .A(n20198), .B(n20197), .ZN(
        P2_U3012) );
  AOI21_X1 U23254 ( .B1(n20203), .B2(n20202), .A(n20201), .ZN(n20239) );
  AOI22_X1 U23255 ( .A1(n20239), .A2(n20205), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20204), .ZN(n20216) );
  XNOR2_X1 U23256 ( .A(n20206), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20240) );
  NOR2_X1 U23257 ( .A1(n20207), .A2(n20808), .ZN(n20245) );
  AOI21_X1 U23258 ( .B1(n20209), .B2(n20208), .A(n20245), .ZN(n20210) );
  OAI21_X1 U23259 ( .B1(n20240), .B2(n20211), .A(n20210), .ZN(n20212) );
  AOI21_X1 U23260 ( .B1(n20214), .B2(n20213), .A(n20212), .ZN(n20215) );
  NAND2_X1 U23261 ( .A1(n20216), .A2(n20215), .ZN(P2_U3013) );
  INV_X1 U23262 ( .A(n20217), .ZN(n20225) );
  INV_X1 U23263 ( .A(n20218), .ZN(n20224) );
  OAI22_X1 U23264 ( .A1(n20242), .A2(n20221), .B1(n20220), .B2(n20219), .ZN(
        n20222) );
  AOI211_X1 U23265 ( .C1(n20225), .C2(n20224), .A(n20223), .B(n20222), .ZN(
        n20233) );
  INV_X1 U23266 ( .A(n20226), .ZN(n20228) );
  OAI22_X1 U23267 ( .A1(n20241), .A2(n20228), .B1(n20887), .B2(n20227), .ZN(
        n20229) );
  AOI211_X1 U23268 ( .C1(n20250), .C2(n20231), .A(n20230), .B(n20229), .ZN(
        n20232) );
  OAI211_X1 U23269 ( .C1(n20235), .C2(n20234), .A(n20233), .B(n20232), .ZN(
        P2_U3044) );
  OAI21_X1 U23270 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n20236), .ZN(n20249) );
  AOI22_X1 U23271 ( .A1(n12495), .A2(n20239), .B1(n20238), .B2(n20237), .ZN(
        n20248) );
  OAI22_X1 U23272 ( .A1(n20243), .A2(n20242), .B1(n20241), .B2(n20240), .ZN(
        n20244) );
  AOI211_X1 U23273 ( .C1(n20246), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20245), .B(n20244), .ZN(n20247) );
  OAI211_X1 U23274 ( .C1(n20250), .C2(n20249), .A(n20248), .B(n20247), .ZN(
        P2_U3045) );
  NOR2_X1 U23275 ( .A1(n20881), .A2(n20310), .ZN(n20252) );
  OR2_X1 U23276 ( .A1(n20881), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20873) );
  INV_X1 U23277 ( .A(n20873), .ZN(n20493) );
  AOI21_X1 U23278 ( .B1(n20256), .B2(n20252), .A(n20493), .ZN(n20254) );
  AOI22_X1 U23279 ( .A1(n20254), .A2(n20257), .B1(n20559), .B2(n20728), .ZN(
        n20255) );
  AND2_X1 U23280 ( .A1(n20253), .A2(n20679), .ZN(n20288) );
  INV_X1 U23281 ( .A(n20254), .ZN(n20259) );
  AOI22_X1 U23282 ( .A1(n20738), .A2(n20724), .B1(n20288), .B2(n20729), .ZN(
        n20262) );
  AOI21_X1 U23283 ( .B1(n9601), .B2(n11308), .A(n20906), .ZN(n20258) );
  AOI21_X1 U23284 ( .B1(n20259), .B2(n20728), .A(n20258), .ZN(n20260) );
  OAI21_X1 U23285 ( .B1(n20260), .B2(n20288), .A(n20731), .ZN(n20292) );
  AOI22_X1 U23286 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20683), .ZN(n20261) );
  OAI211_X1 U23287 ( .C1(n20295), .C2(n20691), .A(n20262), .B(n20261), .ZN(
        P2_U3048) );
  INV_X1 U23288 ( .A(n20743), .ZN(n20695) );
  AOI22_X1 U23289 ( .A1(n20744), .A2(n20724), .B1(n20288), .B2(n20742), .ZN(
        n20264) );
  AOI22_X1 U23290 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20692), .ZN(n20263) );
  OAI211_X1 U23291 ( .C1(n20295), .C2(n20695), .A(n20264), .B(n20263), .ZN(
        P2_U3049) );
  AOI22_X1 U23292 ( .A1(n20750), .A2(n20724), .B1(n20748), .B2(n20288), .ZN(
        n20266) );
  AOI22_X1 U23293 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20696), .ZN(n20265) );
  OAI211_X1 U23294 ( .C1(n20295), .C2(n20699), .A(n20266), .B(n20265), .ZN(
        P2_U3050) );
  INV_X1 U23295 ( .A(n20755), .ZN(n20703) );
  AOI22_X1 U23296 ( .A1(n20756), .A2(n20724), .B1(n20754), .B2(n20288), .ZN(
        n20268) );
  AOI22_X1 U23297 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20700), .ZN(n20267) );
  OAI211_X1 U23298 ( .C1(n20295), .C2(n20703), .A(n20268), .B(n20267), .ZN(
        P2_U3051) );
  INV_X1 U23299 ( .A(n20761), .ZN(n20707) );
  AOI22_X1 U23300 ( .A1(n20762), .A2(n20724), .B1(n20288), .B2(n20760), .ZN(
        n20270) );
  AOI22_X1 U23301 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20704), .ZN(n20269) );
  OAI211_X1 U23302 ( .C1(n20295), .C2(n20707), .A(n20270), .B(n20269), .ZN(
        P2_U3052) );
  INV_X1 U23303 ( .A(n20767), .ZN(n20711) );
  OAI22_X2 U23304 ( .A1(n20272), .A2(n20290), .B1(n16428), .B2(n20289), .ZN(
        n20768) );
  AOI22_X1 U23305 ( .A1(n20768), .A2(n20724), .B1(n20288), .B2(n9787), .ZN(
        n20277) );
  AOI22_X1 U23306 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20708), .ZN(n20276) );
  OAI211_X1 U23307 ( .C1(n20295), .C2(n20711), .A(n20277), .B(n20276), .ZN(
        P2_U3053) );
  OAI22_X2 U23308 ( .A1(n20279), .A2(n20290), .B1(n13596), .B2(n20289), .ZN(
        n20774) );
  NOR2_X2 U23309 ( .A1(n13230), .A2(n20280), .ZN(n20772) );
  AOI22_X1 U23310 ( .A1(n20774), .A2(n20724), .B1(n20288), .B2(n20772), .ZN(
        n20283) );
  OAI22_X2 U23311 ( .A1(n20281), .A2(n20290), .B1(n16475), .B2(n20289), .ZN(
        n20712) );
  AOI22_X1 U23312 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20712), .ZN(n20282) );
  OAI211_X1 U23313 ( .C1(n20295), .C2(n20715), .A(n20283), .B(n20282), .ZN(
        P2_U3054) );
  INV_X1 U23314 ( .A(n20780), .ZN(n20722) );
  OAI22_X2 U23315 ( .A1(n20286), .A2(n20290), .B1(n20285), .B2(n20289), .ZN(
        n20782) );
  AOI22_X1 U23316 ( .A1(n20782), .A2(n20724), .B1(n20288), .B2(n20778), .ZN(
        n20294) );
  AOI22_X1 U23317 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20292), .B1(
        n20310), .B2(n20717), .ZN(n20293) );
  OAI211_X1 U23318 ( .C1(n20295), .C2(n20722), .A(n20294), .B(n20293), .ZN(
        P2_U3055) );
  INV_X1 U23319 ( .A(n20342), .ZN(n20314) );
  AOI22_X1 U23320 ( .A1(n20309), .A2(n20749), .B1(n20748), .B2(n20308), .ZN(
        n20297) );
  AOI22_X1 U23321 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20750), .ZN(n20296) );
  OAI211_X1 U23322 ( .C1(n20753), .C2(n20314), .A(n20297), .B(n20296), .ZN(
        P2_U3058) );
  AOI22_X1 U23323 ( .A1(n20309), .A2(n20755), .B1(n20754), .B2(n20308), .ZN(
        n20299) );
  AOI22_X1 U23324 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20756), .ZN(n20298) );
  OAI211_X1 U23325 ( .C1(n20759), .C2(n20314), .A(n20299), .B(n20298), .ZN(
        P2_U3059) );
  AOI22_X1 U23326 ( .A1(n20309), .A2(n20761), .B1(n20760), .B2(n20308), .ZN(
        n20301) );
  AOI22_X1 U23327 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20762), .ZN(n20300) );
  OAI211_X1 U23328 ( .C1(n20765), .C2(n20314), .A(n20301), .B(n20300), .ZN(
        P2_U3060) );
  AOI22_X1 U23329 ( .A1(n20309), .A2(n20767), .B1(n20308), .B2(n20766), .ZN(
        n20303) );
  AOI22_X1 U23330 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20768), .ZN(n20302) );
  OAI211_X1 U23331 ( .C1(n20771), .C2(n20314), .A(n20303), .B(n20302), .ZN(
        P2_U3061) );
  AOI22_X1 U23332 ( .A1(n20309), .A2(n20773), .B1(n20308), .B2(n20772), .ZN(
        n20305) );
  AOI22_X1 U23333 ( .A1(n20342), .A2(n20712), .B1(n20310), .B2(n20774), .ZN(
        n20304) );
  OAI211_X1 U23334 ( .C1(n20307), .C2(n20306), .A(n20305), .B(n20304), .ZN(
        P2_U3062) );
  AOI22_X1 U23335 ( .A1(n20309), .A2(n20780), .B1(n20308), .B2(n20778), .ZN(
        n20313) );
  AOI22_X1 U23336 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20311), .B1(
        n20310), .B2(n20782), .ZN(n20312) );
  OAI211_X1 U23337 ( .C1(n20787), .C2(n20314), .A(n20313), .B(n20312), .ZN(
        P2_U3063) );
  NOR2_X1 U23338 ( .A1(n20555), .A2(n20322), .ZN(n20340) );
  OAI21_X1 U23339 ( .B1(n20316), .B2(n20340), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20317) );
  OAI21_X1 U23340 ( .B1(n20322), .B2(n20557), .A(n20317), .ZN(n20341) );
  AOI22_X1 U23341 ( .A1(n20341), .A2(n20730), .B1(n20340), .B2(n20729), .ZN(
        n20327) );
  INV_X1 U23342 ( .A(n20340), .ZN(n20318) );
  OAI211_X1 U23343 ( .C1(n20319), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20318), 
        .B(n20881), .ZN(n20325) );
  INV_X1 U23344 ( .A(n20377), .ZN(n20320) );
  OAI21_X1 U23345 ( .B1(n20342), .B2(n20320), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20321) );
  OAI21_X1 U23346 ( .B1(n20323), .B2(n20322), .A(n20321), .ZN(n20324) );
  NAND3_X1 U23347 ( .A1(n20325), .A2(n20731), .A3(n20324), .ZN(n20343) );
  AOI22_X1 U23348 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20738), .ZN(n20326) );
  OAI211_X1 U23349 ( .C1(n20741), .C2(n20377), .A(n20327), .B(n20326), .ZN(
        P2_U3064) );
  AOI22_X1 U23350 ( .A1(n20341), .A2(n20743), .B1(n20742), .B2(n20340), .ZN(
        n20329) );
  AOI22_X1 U23351 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20744), .ZN(n20328) );
  OAI211_X1 U23352 ( .C1(n20747), .C2(n20377), .A(n20329), .B(n20328), .ZN(
        P2_U3065) );
  AOI22_X1 U23353 ( .A1(n20341), .A2(n20749), .B1(n20748), .B2(n20340), .ZN(
        n20331) );
  AOI22_X1 U23354 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20750), .ZN(n20330) );
  OAI211_X1 U23355 ( .C1(n20753), .C2(n20377), .A(n20331), .B(n20330), .ZN(
        P2_U3066) );
  AOI22_X1 U23356 ( .A1(n20341), .A2(n20755), .B1(n20754), .B2(n20340), .ZN(
        n20333) );
  AOI22_X1 U23357 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20756), .ZN(n20332) );
  OAI211_X1 U23358 ( .C1(n20759), .C2(n20377), .A(n20333), .B(n20332), .ZN(
        P2_U3067) );
  AOI22_X1 U23359 ( .A1(n20341), .A2(n20761), .B1(n20760), .B2(n20340), .ZN(
        n20335) );
  AOI22_X1 U23360 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20762), .ZN(n20334) );
  OAI211_X1 U23361 ( .C1(n20765), .C2(n20377), .A(n20335), .B(n20334), .ZN(
        P2_U3068) );
  AOI22_X1 U23362 ( .A1(n20341), .A2(n20767), .B1(n9787), .B2(n20340), .ZN(
        n20337) );
  AOI22_X1 U23363 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20768), .ZN(n20336) );
  OAI211_X1 U23364 ( .C1(n20771), .C2(n20377), .A(n20337), .B(n20336), .ZN(
        P2_U3069) );
  AOI22_X1 U23365 ( .A1(n20341), .A2(n20773), .B1(n20772), .B2(n20340), .ZN(
        n20339) );
  AOI22_X1 U23366 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20774), .ZN(n20338) );
  OAI211_X1 U23367 ( .C1(n20777), .C2(n20377), .A(n20339), .B(n20338), .ZN(
        P2_U3070) );
  AOI22_X1 U23368 ( .A1(n20341), .A2(n20780), .B1(n20778), .B2(n20340), .ZN(
        n20345) );
  AOI22_X1 U23369 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20343), .B1(
        n20342), .B2(n20782), .ZN(n20344) );
  OAI211_X1 U23370 ( .C1(n20787), .C2(n20377), .A(n20345), .B(n20344), .ZN(
        P2_U3071) );
  INV_X1 U23371 ( .A(n20738), .ZN(n20471) );
  AND2_X1 U23372 ( .A1(n20462), .A2(n20349), .ZN(n20372) );
  AOI22_X1 U23373 ( .A1(n20683), .A2(n9650), .B1(n20372), .B2(n20729), .ZN(
        n20359) );
  INV_X1 U23374 ( .A(n20372), .ZN(n20347) );
  OAI21_X1 U23375 ( .B1(n20348), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20347), 
        .ZN(n20351) );
  NAND2_X1 U23376 ( .A1(n20464), .A2(n20870), .ZN(n20355) );
  NAND2_X1 U23377 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20349), .ZN(
        n20353) );
  NAND2_X1 U23378 ( .A1(n20355), .A2(n20353), .ZN(n20350) );
  MUX2_X1 U23379 ( .A(n20351), .B(n20350), .S(n20906), .Z(n20352) );
  NAND2_X1 U23380 ( .A1(n20352), .A2(n20731), .ZN(n20374) );
  INV_X1 U23381 ( .A(n20353), .ZN(n20354) );
  NAND3_X1 U23382 ( .A1(n20355), .A2(n20906), .A3(n20354), .ZN(n20357) );
  NAND2_X1 U23383 ( .A1(n20357), .A2(n20356), .ZN(n20373) );
  AOI22_X1 U23384 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20374), .B1(
        n20730), .B2(n20373), .ZN(n20358) );
  OAI211_X1 U23385 ( .C1(n20471), .C2(n20377), .A(n20359), .B(n20358), .ZN(
        P2_U3072) );
  INV_X1 U23386 ( .A(n20744), .ZN(n20474) );
  AOI22_X1 U23387 ( .A1(n20692), .A2(n9650), .B1(n20372), .B2(n20742), .ZN(
        n20361) );
  AOI22_X1 U23388 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20374), .B1(
        n20743), .B2(n20373), .ZN(n20360) );
  OAI211_X1 U23389 ( .C1(n20474), .C2(n20377), .A(n20361), .B(n20360), .ZN(
        P2_U3073) );
  INV_X1 U23390 ( .A(n20750), .ZN(n20591) );
  AOI22_X1 U23391 ( .A1(n20696), .A2(n9650), .B1(n20748), .B2(n20372), .ZN(
        n20363) );
  AOI22_X1 U23392 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20374), .B1(
        n20749), .B2(n20373), .ZN(n20362) );
  OAI211_X1 U23393 ( .C1(n20591), .C2(n20377), .A(n20363), .B(n20362), .ZN(
        P2_U3074) );
  INV_X1 U23394 ( .A(n20756), .ZN(n20479) );
  AOI22_X1 U23395 ( .A1(n20700), .A2(n9650), .B1(n20754), .B2(n20372), .ZN(
        n20365) );
  AOI22_X1 U23396 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20374), .B1(
        n20755), .B2(n20373), .ZN(n20364) );
  OAI211_X1 U23397 ( .C1(n20479), .C2(n20377), .A(n20365), .B(n20364), .ZN(
        P2_U3075) );
  INV_X1 U23398 ( .A(n20762), .ZN(n20482) );
  AOI22_X1 U23399 ( .A1(n20704), .A2(n9650), .B1(n20372), .B2(n20760), .ZN(
        n20367) );
  AOI22_X1 U23400 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20374), .B1(
        n20761), .B2(n20373), .ZN(n20366) );
  OAI211_X1 U23401 ( .C1(n20482), .C2(n20377), .A(n20367), .B(n20366), .ZN(
        P2_U3076) );
  INV_X1 U23402 ( .A(n20768), .ZN(n20598) );
  AOI22_X1 U23403 ( .A1(n20708), .A2(n9650), .B1(n20372), .B2(n9787), .ZN(
        n20369) );
  AOI22_X1 U23404 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20374), .B1(
        n20767), .B2(n20373), .ZN(n20368) );
  OAI211_X1 U23405 ( .C1(n20598), .C2(n20377), .A(n20369), .B(n20368), .ZN(
        P2_U3077) );
  INV_X1 U23406 ( .A(n20774), .ZN(n20601) );
  AOI22_X1 U23407 ( .A1(n20712), .A2(n9650), .B1(n20372), .B2(n20772), .ZN(
        n20371) );
  AOI22_X1 U23408 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20374), .B1(
        n20773), .B2(n20373), .ZN(n20370) );
  OAI211_X1 U23409 ( .C1(n20601), .C2(n20377), .A(n20371), .B(n20370), .ZN(
        P2_U3078) );
  INV_X1 U23410 ( .A(n20782), .ZN(n20608) );
  AOI22_X1 U23411 ( .A1(n20717), .A2(n9650), .B1(n20372), .B2(n20778), .ZN(
        n20376) );
  AOI22_X1 U23412 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20374), .B1(
        n20780), .B2(n20373), .ZN(n20375) );
  OAI211_X1 U23413 ( .C1(n20608), .C2(n20377), .A(n20376), .B(n20375), .ZN(
        P2_U3079) );
  INV_X1 U23414 ( .A(n20378), .ZN(n20380) );
  AND2_X1 U23415 ( .A1(n20379), .A2(n20679), .ZN(n20404) );
  NOR3_X1 U23416 ( .A1(n20380), .A2(n20404), .A3(n20559), .ZN(n20383) );
  NOR3_X1 U23417 ( .A1(n20381), .A2(n20434), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20384) );
  AOI21_X1 U23418 ( .B1(n20384), .B2(n11308), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20382) );
  AOI22_X1 U23419 ( .A1(n20405), .A2(n20730), .B1(n20404), .B2(n20729), .ZN(
        n20391) );
  INV_X1 U23420 ( .A(n20383), .ZN(n20389) );
  INV_X1 U23421 ( .A(n20384), .ZN(n20387) );
  OAI21_X1 U23422 ( .B1(n9650), .B2(n20427), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20386) );
  INV_X1 U23423 ( .A(n20404), .ZN(n20385) );
  AOI22_X1 U23424 ( .A1(n20387), .A2(n20386), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20385), .ZN(n20388) );
  NAND3_X1 U23425 ( .A1(n20389), .A2(n20388), .A3(n20731), .ZN(n20406) );
  AOI22_X1 U23426 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20738), .ZN(n20390) );
  OAI211_X1 U23427 ( .C1(n20741), .C2(n20425), .A(n20391), .B(n20390), .ZN(
        P2_U3080) );
  AOI22_X1 U23428 ( .A1(n20405), .A2(n20743), .B1(n20742), .B2(n20404), .ZN(
        n20393) );
  AOI22_X1 U23429 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20744), .ZN(n20392) );
  OAI211_X1 U23430 ( .C1(n20747), .C2(n20425), .A(n20393), .B(n20392), .ZN(
        P2_U3081) );
  AOI22_X1 U23431 ( .A1(n20405), .A2(n20749), .B1(n20748), .B2(n20404), .ZN(
        n20395) );
  AOI22_X1 U23432 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20750), .ZN(n20394) );
  OAI211_X1 U23433 ( .C1(n20753), .C2(n20425), .A(n20395), .B(n20394), .ZN(
        P2_U3082) );
  AOI22_X1 U23434 ( .A1(n20405), .A2(n20755), .B1(n20754), .B2(n20404), .ZN(
        n20397) );
  AOI22_X1 U23435 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20756), .ZN(n20396) );
  OAI211_X1 U23436 ( .C1(n20759), .C2(n20425), .A(n20397), .B(n20396), .ZN(
        P2_U3083) );
  AOI22_X1 U23437 ( .A1(n20405), .A2(n20761), .B1(n20760), .B2(n20404), .ZN(
        n20399) );
  AOI22_X1 U23438 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20762), .ZN(n20398) );
  OAI211_X1 U23439 ( .C1(n20765), .C2(n20425), .A(n20399), .B(n20398), .ZN(
        P2_U3084) );
  AOI22_X1 U23440 ( .A1(n20405), .A2(n20767), .B1(n9787), .B2(n20404), .ZN(
        n20401) );
  AOI22_X1 U23441 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20768), .ZN(n20400) );
  OAI211_X1 U23442 ( .C1(n20771), .C2(n20425), .A(n20401), .B(n20400), .ZN(
        P2_U3085) );
  AOI22_X1 U23443 ( .A1(n20405), .A2(n20773), .B1(n20772), .B2(n20404), .ZN(
        n20403) );
  AOI22_X1 U23444 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20774), .ZN(n20402) );
  OAI211_X1 U23445 ( .C1(n20777), .C2(n20425), .A(n20403), .B(n20402), .ZN(
        P2_U3086) );
  AOI22_X1 U23446 ( .A1(n20405), .A2(n20780), .B1(n20778), .B2(n20404), .ZN(
        n20408) );
  AOI22_X1 U23447 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20406), .B1(
        n9650), .B2(n20782), .ZN(n20407) );
  OAI211_X1 U23448 ( .C1(n20787), .C2(n20425), .A(n20408), .B(n20407), .ZN(
        P2_U3087) );
  AOI22_X1 U23449 ( .A1(n20738), .A2(n20427), .B1(n20426), .B2(n20729), .ZN(
        n20411) );
  AOI22_X1 U23450 ( .A1(n20730), .A2(n20428), .B1(n20457), .B2(n20683), .ZN(
        n20410) );
  OAI211_X1 U23451 ( .C1(n20432), .C2(n20412), .A(n20411), .B(n20410), .ZN(
        P2_U3088) );
  INV_X1 U23452 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U23453 ( .A1(n20744), .A2(n20427), .B1(n20426), .B2(n20742), .ZN(
        n20414) );
  AOI22_X1 U23454 ( .A1(n20743), .A2(n20428), .B1(n20457), .B2(n20692), .ZN(
        n20413) );
  OAI211_X1 U23455 ( .C1(n20432), .C2(n20415), .A(n20414), .B(n20413), .ZN(
        P2_U3089) );
  AOI22_X1 U23456 ( .A1(n20696), .A2(n20457), .B1(n20748), .B2(n20426), .ZN(
        n20417) );
  AOI22_X1 U23457 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20422), .B1(
        n20749), .B2(n20428), .ZN(n20416) );
  OAI211_X1 U23458 ( .C1(n20591), .C2(n20425), .A(n20417), .B(n20416), .ZN(
        P2_U3090) );
  AOI22_X1 U23459 ( .A1(n20700), .A2(n20457), .B1(n20754), .B2(n20426), .ZN(
        n20419) );
  AOI22_X1 U23460 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20422), .B1(
        n20755), .B2(n20428), .ZN(n20418) );
  OAI211_X1 U23461 ( .C1(n20479), .C2(n20425), .A(n20419), .B(n20418), .ZN(
        P2_U3091) );
  AOI22_X1 U23462 ( .A1(n20708), .A2(n20457), .B1(n20426), .B2(n20766), .ZN(
        n20421) );
  AOI22_X1 U23463 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20422), .B1(
        n20767), .B2(n20428), .ZN(n20420) );
  OAI211_X1 U23464 ( .C1(n20598), .C2(n20425), .A(n20421), .B(n20420), .ZN(
        P2_U3093) );
  AOI22_X1 U23465 ( .A1(n20712), .A2(n20457), .B1(n20426), .B2(n20772), .ZN(
        n20424) );
  AOI22_X1 U23466 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20422), .B1(
        n20773), .B2(n20428), .ZN(n20423) );
  OAI211_X1 U23467 ( .C1(n20601), .C2(n20425), .A(n20424), .B(n20423), .ZN(
        P2_U3094) );
  INV_X1 U23468 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n20431) );
  AOI22_X1 U23469 ( .A1(n20782), .A2(n20427), .B1(n20426), .B2(n20778), .ZN(
        n20430) );
  AOI22_X1 U23470 ( .A1(n20780), .A2(n20428), .B1(n20457), .B2(n20717), .ZN(
        n20429) );
  OAI211_X1 U23471 ( .C1(n20432), .C2(n20431), .A(n20430), .B(n20429), .ZN(
        P2_U3095) );
  NAND2_X1 U23472 ( .A1(n20434), .A2(n20461), .ZN(n20439) );
  NOR3_X1 U23473 ( .A1(n20436), .A2(n10465), .A3(n20559), .ZN(n20438) );
  AOI211_X2 U23474 ( .C1(n20559), .C2(n20439), .A(n20463), .B(n20438), .ZN(
        n20456) );
  AOI22_X1 U23475 ( .A1(n20456), .A2(n20730), .B1(n10465), .B2(n20729), .ZN(
        n20443) );
  OAI21_X1 U23476 ( .B1(n20457), .B2(n20437), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20440) );
  AOI211_X1 U23477 ( .C1(n20440), .C2(n20439), .A(n20636), .B(n20438), .ZN(
        n20441) );
  AOI22_X1 U23478 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20738), .ZN(n20442) );
  OAI211_X1 U23479 ( .C1(n20741), .C2(n20491), .A(n20443), .B(n20442), .ZN(
        P2_U3096) );
  AOI22_X1 U23480 ( .A1(n20456), .A2(n20743), .B1(n10465), .B2(n20742), .ZN(
        n20445) );
  AOI22_X1 U23481 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20744), .ZN(n20444) );
  OAI211_X1 U23482 ( .C1(n20747), .C2(n20491), .A(n20445), .B(n20444), .ZN(
        P2_U3097) );
  AOI22_X1 U23483 ( .A1(n20456), .A2(n20749), .B1(n20748), .B2(n10465), .ZN(
        n20447) );
  AOI22_X1 U23484 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20750), .ZN(n20446) );
  OAI211_X1 U23485 ( .C1(n20753), .C2(n20491), .A(n20447), .B(n20446), .ZN(
        P2_U3098) );
  AOI22_X1 U23486 ( .A1(n20456), .A2(n20755), .B1(n20754), .B2(n10465), .ZN(
        n20449) );
  AOI22_X1 U23487 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20756), .ZN(n20448) );
  OAI211_X1 U23488 ( .C1(n20759), .C2(n20491), .A(n20449), .B(n20448), .ZN(
        P2_U3099) );
  AOI22_X1 U23489 ( .A1(n20456), .A2(n20761), .B1(n10465), .B2(n20760), .ZN(
        n20451) );
  AOI22_X1 U23490 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20762), .ZN(n20450) );
  OAI211_X1 U23491 ( .C1(n20765), .C2(n20491), .A(n20451), .B(n20450), .ZN(
        P2_U3100) );
  AOI22_X1 U23492 ( .A1(n20456), .A2(n20767), .B1(n10465), .B2(n20766), .ZN(
        n20453) );
  AOI22_X1 U23493 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20768), .ZN(n20452) );
  OAI211_X1 U23494 ( .C1(n20771), .C2(n20491), .A(n20453), .B(n20452), .ZN(
        P2_U3101) );
  AOI22_X1 U23495 ( .A1(n20456), .A2(n20773), .B1(n10465), .B2(n20772), .ZN(
        n20455) );
  AOI22_X1 U23496 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20774), .ZN(n20454) );
  OAI211_X1 U23497 ( .C1(n20777), .C2(n20491), .A(n20455), .B(n20454), .ZN(
        P2_U3102) );
  AOI22_X1 U23498 ( .A1(n20456), .A2(n20780), .B1(n10465), .B2(n20778), .ZN(
        n20460) );
  AOI22_X1 U23499 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20458), .B1(
        n20457), .B2(n20782), .ZN(n20459) );
  OAI211_X1 U23500 ( .C1(n20787), .C2(n20491), .A(n20460), .B(n20459), .ZN(
        P2_U3103) );
  NAND3_X1 U23501 ( .A1(n20885), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20466) );
  NOR3_X1 U23502 ( .A1(n10817), .A2(n20501), .A3(n20559), .ZN(n20465) );
  AOI211_X2 U23503 ( .C1(n20559), .C2(n20466), .A(n20463), .B(n20465), .ZN(
        n20487) );
  AOI22_X1 U23504 ( .A1(n20487), .A2(n20730), .B1(n20501), .B2(n20729), .ZN(
        n20470) );
  INV_X1 U23505 ( .A(n20673), .ZN(n20736) );
  NAND2_X1 U23506 ( .A1(n20464), .A2(n20736), .ZN(n20882) );
  AOI211_X1 U23507 ( .C1(n20882), .C2(n20466), .A(n20636), .B(n20465), .ZN(
        n20467) );
  AOI22_X1 U23508 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20683), .ZN(n20469) );
  OAI211_X1 U23509 ( .C1(n20471), .C2(n20491), .A(n20470), .B(n20469), .ZN(
        P2_U3104) );
  AOI22_X1 U23510 ( .A1(n20487), .A2(n20743), .B1(n20501), .B2(n20742), .ZN(
        n20473) );
  AOI22_X1 U23511 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20692), .ZN(n20472) );
  OAI211_X1 U23512 ( .C1(n20474), .C2(n20491), .A(n20473), .B(n20472), .ZN(
        P2_U3105) );
  AOI22_X1 U23513 ( .A1(n20487), .A2(n20749), .B1(n20748), .B2(n20501), .ZN(
        n20476) );
  AOI22_X1 U23514 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20696), .ZN(n20475) );
  OAI211_X1 U23515 ( .C1(n20591), .C2(n20491), .A(n20476), .B(n20475), .ZN(
        P2_U3106) );
  AOI22_X1 U23516 ( .A1(n20487), .A2(n20755), .B1(n20754), .B2(n20501), .ZN(
        n20478) );
  AOI22_X1 U23517 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20700), .ZN(n20477) );
  OAI211_X1 U23518 ( .C1(n20479), .C2(n20491), .A(n20478), .B(n20477), .ZN(
        P2_U3107) );
  AOI22_X1 U23519 ( .A1(n20487), .A2(n20761), .B1(n20501), .B2(n20760), .ZN(
        n20481) );
  AOI22_X1 U23520 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20704), .ZN(n20480) );
  OAI211_X1 U23521 ( .C1(n20482), .C2(n20491), .A(n20481), .B(n20480), .ZN(
        P2_U3108) );
  AOI22_X1 U23522 ( .A1(n20487), .A2(n20767), .B1(n20501), .B2(n20766), .ZN(
        n20484) );
  AOI22_X1 U23523 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20708), .ZN(n20483) );
  OAI211_X1 U23524 ( .C1(n20598), .C2(n20491), .A(n20484), .B(n20483), .ZN(
        P2_U3109) );
  AOI22_X1 U23525 ( .A1(n20487), .A2(n20773), .B1(n20501), .B2(n20772), .ZN(
        n20486) );
  AOI22_X1 U23526 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20712), .ZN(n20485) );
  OAI211_X1 U23527 ( .C1(n20601), .C2(n20491), .A(n20486), .B(n20485), .ZN(
        P2_U3110) );
  AOI22_X1 U23528 ( .A1(n20487), .A2(n20780), .B1(n20501), .B2(n20778), .ZN(
        n20490) );
  AOI22_X1 U23529 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20488), .B1(
        n20520), .B2(n20717), .ZN(n20489) );
  OAI211_X1 U23530 ( .C1(n20608), .C2(n20491), .A(n20490), .B(n20489), .ZN(
        P2_U3111) );
  INV_X1 U23531 ( .A(n20501), .ZN(n20494) );
  NOR2_X1 U23532 ( .A1(n20500), .A2(n20494), .ZN(n20499) );
  INV_X1 U23533 ( .A(n20495), .ZN(n20558) );
  OR2_X1 U23534 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20558), .ZN(
        n20531) );
  NOR2_X1 U23535 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20531), .ZN(
        n20519) );
  INV_X1 U23536 ( .A(n20519), .ZN(n20496) );
  OAI21_X1 U23537 ( .B1(n20503), .B2(n20559), .A(n20496), .ZN(n20498) );
  INV_X1 U23538 ( .A(n20500), .ZN(n20497) );
  AOI22_X1 U23539 ( .A1(n20683), .A2(n20550), .B1(n20519), .B2(n20729), .ZN(
        n20506) );
  AOI22_X1 U23540 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20738), .ZN(n20505) );
  OAI211_X1 U23541 ( .C1(n20524), .C2(n20691), .A(n20506), .B(n20505), .ZN(
        P2_U3112) );
  AOI22_X1 U23542 ( .A1(n20692), .A2(n20550), .B1(n20519), .B2(n20742), .ZN(
        n20508) );
  AOI22_X1 U23543 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20744), .ZN(n20507) );
  OAI211_X1 U23544 ( .C1(n20524), .C2(n20695), .A(n20508), .B(n20507), .ZN(
        P2_U3113) );
  AOI22_X1 U23545 ( .A1(n20696), .A2(n20550), .B1(n20748), .B2(n20519), .ZN(
        n20510) );
  AOI22_X1 U23546 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20750), .ZN(n20509) );
  OAI211_X1 U23547 ( .C1(n20524), .C2(n20699), .A(n20510), .B(n20509), .ZN(
        P2_U3114) );
  AOI22_X1 U23548 ( .A1(n20700), .A2(n20550), .B1(n20754), .B2(n20519), .ZN(
        n20512) );
  AOI22_X1 U23549 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20756), .ZN(n20511) );
  OAI211_X1 U23550 ( .C1(n20524), .C2(n20703), .A(n20512), .B(n20511), .ZN(
        P2_U3115) );
  AOI22_X1 U23551 ( .A1(n20704), .A2(n20550), .B1(n20519), .B2(n20760), .ZN(
        n20514) );
  AOI22_X1 U23552 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20762), .ZN(n20513) );
  OAI211_X1 U23553 ( .C1(n20524), .C2(n20707), .A(n20514), .B(n20513), .ZN(
        P2_U3116) );
  AOI22_X1 U23554 ( .A1(n20708), .A2(n20550), .B1(n20519), .B2(n20766), .ZN(
        n20516) );
  AOI22_X1 U23555 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20768), .ZN(n20515) );
  OAI211_X1 U23556 ( .C1(n20524), .C2(n20711), .A(n20516), .B(n20515), .ZN(
        P2_U3117) );
  AOI22_X1 U23557 ( .A1(n20712), .A2(n20550), .B1(n20519), .B2(n20772), .ZN(
        n20518) );
  AOI22_X1 U23558 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20774), .ZN(n20517) );
  OAI211_X1 U23559 ( .C1(n20524), .C2(n20715), .A(n20518), .B(n20517), .ZN(
        P2_U3118) );
  AOI22_X1 U23560 ( .A1(n20717), .A2(n20550), .B1(n20519), .B2(n20778), .ZN(
        n20523) );
  AOI22_X1 U23561 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20782), .ZN(n20522) );
  OAI211_X1 U23562 ( .C1(n20524), .C2(n20722), .A(n20523), .B(n20522), .ZN(
        P2_U3119) );
  NOR2_X1 U23563 ( .A1(n20881), .A2(n20531), .ZN(n20527) );
  NOR2_X1 U23564 ( .A1(n20525), .A2(n20558), .ZN(n20549) );
  INV_X1 U23565 ( .A(n20549), .ZN(n20562) );
  AOI21_X1 U23566 ( .B1(n20528), .B2(n20562), .A(n20559), .ZN(n20526) );
  NOR2_X1 U23567 ( .A1(n20527), .A2(n20526), .ZN(n20554) );
  AOI22_X1 U23568 ( .A1(n20738), .A2(n20550), .B1(n20549), .B2(n20729), .ZN(
        n20536) );
  AOI21_X1 U23569 ( .B1(n20528), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20533) );
  NAND2_X1 U23570 ( .A1(n20735), .A2(n20529), .ZN(n20530) );
  NAND2_X1 U23571 ( .A1(n20531), .A2(n20530), .ZN(n20532) );
  OAI211_X1 U23572 ( .C1(n20549), .C2(n20533), .A(n20532), .B(n20731), .ZN(
        n20551) );
  AOI22_X1 U23573 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20551), .B1(
        n10477), .B2(n20683), .ZN(n20535) );
  OAI211_X1 U23574 ( .C1(n20554), .C2(n20691), .A(n20536), .B(n20535), .ZN(
        P2_U3120) );
  AOI22_X1 U23575 ( .A1(n20692), .A2(n10477), .B1(n20549), .B2(n20742), .ZN(
        n20538) );
  AOI22_X1 U23576 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20551), .B1(
        n20550), .B2(n20744), .ZN(n20537) );
  OAI211_X1 U23577 ( .C1(n20554), .C2(n20695), .A(n20538), .B(n20537), .ZN(
        P2_U3121) );
  AOI22_X1 U23578 ( .A1(n20696), .A2(n10477), .B1(n20748), .B2(n20549), .ZN(
        n20540) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20551), .B1(
        n20550), .B2(n20750), .ZN(n20539) );
  OAI211_X1 U23580 ( .C1(n20554), .C2(n20699), .A(n20540), .B(n20539), .ZN(
        P2_U3122) );
  AOI22_X1 U23581 ( .A1(n20756), .A2(n20550), .B1(n20754), .B2(n20549), .ZN(
        n20542) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20551), .B1(
        n10477), .B2(n20700), .ZN(n20541) );
  OAI211_X1 U23583 ( .C1(n20554), .C2(n20703), .A(n20542), .B(n20541), .ZN(
        P2_U3123) );
  AOI22_X1 U23584 ( .A1(n20704), .A2(n10477), .B1(n20549), .B2(n20760), .ZN(
        n20544) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20551), .B1(
        n20550), .B2(n20762), .ZN(n20543) );
  OAI211_X1 U23586 ( .C1(n20554), .C2(n20707), .A(n20544), .B(n20543), .ZN(
        P2_U3124) );
  AOI22_X1 U23587 ( .A1(n20708), .A2(n10477), .B1(n20549), .B2(n20766), .ZN(
        n20546) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20551), .B1(
        n20550), .B2(n20768), .ZN(n20545) );
  OAI211_X1 U23589 ( .C1(n20554), .C2(n20711), .A(n20546), .B(n20545), .ZN(
        P2_U3125) );
  AOI22_X1 U23590 ( .A1(n20712), .A2(n10477), .B1(n20549), .B2(n20772), .ZN(
        n20548) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20551), .B1(
        n20550), .B2(n20774), .ZN(n20547) );
  OAI211_X1 U23592 ( .C1(n20554), .C2(n20715), .A(n20548), .B(n20547), .ZN(
        P2_U3126) );
  AOI22_X1 U23593 ( .A1(n20782), .A2(n20550), .B1(n20549), .B2(n20778), .ZN(
        n20553) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20551), .B1(
        n10477), .B2(n20717), .ZN(n20552) );
  OAI211_X1 U23595 ( .C1(n20554), .C2(n20722), .A(n20553), .B(n20552), .ZN(
        P2_U3127) );
  NOR2_X1 U23596 ( .A1(n20555), .A2(n20558), .ZN(n20579) );
  OAI21_X1 U23597 ( .B1(n20560), .B2(n20579), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20556) );
  AOI22_X1 U23598 ( .A1(n20580), .A2(n20730), .B1(n20579), .B2(n20729), .ZN(
        n20566) );
  OAI21_X1 U23599 ( .B1(n10477), .B2(n20592), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20563) );
  OAI21_X1 U23600 ( .B1(n20560), .B2(n20559), .A(n11308), .ZN(n20561) );
  AOI21_X1 U23601 ( .B1(n20563), .B2(n20562), .A(n20561), .ZN(n20564) );
  OAI21_X1 U23602 ( .B1(n20564), .B2(n20579), .A(n20731), .ZN(n20581) );
  AOI22_X1 U23603 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20738), .ZN(n20565) );
  OAI211_X1 U23604 ( .C1(n20741), .C2(n20607), .A(n20566), .B(n20565), .ZN(
        P2_U3128) );
  AOI22_X1 U23605 ( .A1(n20580), .A2(n20743), .B1(n20579), .B2(n20742), .ZN(
        n20568) );
  AOI22_X1 U23606 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20744), .ZN(n20567) );
  OAI211_X1 U23607 ( .C1(n20747), .C2(n20607), .A(n20568), .B(n20567), .ZN(
        P2_U3129) );
  AOI22_X1 U23608 ( .A1(n20580), .A2(n20749), .B1(n20748), .B2(n20579), .ZN(
        n20570) );
  AOI22_X1 U23609 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20750), .ZN(n20569) );
  OAI211_X1 U23610 ( .C1(n20753), .C2(n20607), .A(n20570), .B(n20569), .ZN(
        P2_U3130) );
  AOI22_X1 U23611 ( .A1(n20580), .A2(n20755), .B1(n20754), .B2(n20579), .ZN(
        n20572) );
  AOI22_X1 U23612 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20756), .ZN(n20571) );
  OAI211_X1 U23613 ( .C1(n20759), .C2(n20607), .A(n20572), .B(n20571), .ZN(
        P2_U3131) );
  AOI22_X1 U23614 ( .A1(n20580), .A2(n20761), .B1(n20579), .B2(n20760), .ZN(
        n20574) );
  AOI22_X1 U23615 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20762), .ZN(n20573) );
  OAI211_X1 U23616 ( .C1(n20765), .C2(n20607), .A(n20574), .B(n20573), .ZN(
        P2_U3132) );
  AOI22_X1 U23617 ( .A1(n20580), .A2(n20767), .B1(n20579), .B2(n9787), .ZN(
        n20576) );
  AOI22_X1 U23618 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20768), .ZN(n20575) );
  OAI211_X1 U23619 ( .C1(n20771), .C2(n20607), .A(n20576), .B(n20575), .ZN(
        P2_U3133) );
  AOI22_X1 U23620 ( .A1(n20580), .A2(n20773), .B1(n20579), .B2(n20772), .ZN(
        n20578) );
  AOI22_X1 U23621 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20774), .ZN(n20577) );
  OAI211_X1 U23622 ( .C1(n20777), .C2(n20607), .A(n20578), .B(n20577), .ZN(
        P2_U3134) );
  AOI22_X1 U23623 ( .A1(n20580), .A2(n20780), .B1(n20579), .B2(n20778), .ZN(
        n20583) );
  AOI22_X1 U23624 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20581), .B1(
        n10477), .B2(n20782), .ZN(n20582) );
  OAI211_X1 U23625 ( .C1(n20787), .C2(n20607), .A(n20583), .B(n20582), .ZN(
        P2_U3135) );
  INV_X1 U23626 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20586) );
  AOI22_X1 U23627 ( .A1(n20603), .A2(n20730), .B1(n20602), .B2(n20729), .ZN(
        n20585) );
  AOI22_X1 U23628 ( .A1(n20622), .A2(n20683), .B1(n20592), .B2(n20738), .ZN(
        n20584) );
  OAI211_X1 U23629 ( .C1(n20595), .C2(n20586), .A(n20585), .B(n20584), .ZN(
        P2_U3136) );
  AOI22_X1 U23630 ( .A1(n20603), .A2(n20743), .B1(n20602), .B2(n20742), .ZN(
        n20588) );
  AOI22_X1 U23631 ( .A1(n20622), .A2(n20692), .B1(n20592), .B2(n20744), .ZN(
        n20587) );
  OAI211_X1 U23632 ( .C1(n20595), .C2(n10719), .A(n20588), .B(n20587), .ZN(
        P2_U3137) );
  AOI22_X1 U23633 ( .A1(n20603), .A2(n20749), .B1(n20748), .B2(n20602), .ZN(
        n20590) );
  AOI22_X1 U23634 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20604), .B1(
        n20622), .B2(n20696), .ZN(n20589) );
  OAI211_X1 U23635 ( .C1(n20591), .C2(n20607), .A(n20590), .B(n20589), .ZN(
        P2_U3138) );
  AOI22_X1 U23636 ( .A1(n20603), .A2(n20761), .B1(n20602), .B2(n20760), .ZN(
        n20594) );
  AOI22_X1 U23637 ( .A1(n20622), .A2(n20704), .B1(n20592), .B2(n20762), .ZN(
        n20593) );
  OAI211_X1 U23638 ( .C1(n20595), .C2(n11436), .A(n20594), .B(n20593), .ZN(
        P2_U3140) );
  AOI22_X1 U23639 ( .A1(n20603), .A2(n20767), .B1(n20602), .B2(n9787), .ZN(
        n20597) );
  AOI22_X1 U23640 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20604), .B1(
        n20622), .B2(n20708), .ZN(n20596) );
  OAI211_X1 U23641 ( .C1(n20598), .C2(n20607), .A(n20597), .B(n20596), .ZN(
        P2_U3141) );
  AOI22_X1 U23642 ( .A1(n20603), .A2(n20773), .B1(n20602), .B2(n20772), .ZN(
        n20600) );
  AOI22_X1 U23643 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20604), .B1(
        n20622), .B2(n20712), .ZN(n20599) );
  OAI211_X1 U23644 ( .C1(n20601), .C2(n20607), .A(n20600), .B(n20599), .ZN(
        P2_U3142) );
  AOI22_X1 U23645 ( .A1(n20603), .A2(n20780), .B1(n20602), .B2(n20778), .ZN(
        n20606) );
  AOI22_X1 U23646 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20604), .B1(
        n20622), .B2(n20717), .ZN(n20605) );
  OAI211_X1 U23647 ( .C1(n20608), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        P2_U3143) );
  INV_X1 U23648 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n20611) );
  AOI22_X1 U23649 ( .A1(n20621), .A2(n20730), .B1(n20620), .B2(n20729), .ZN(
        n20610) );
  AOI22_X1 U23650 ( .A1(n20669), .A2(n20683), .B1(n20622), .B2(n20738), .ZN(
        n20609) );
  OAI211_X1 U23651 ( .C1(n20626), .C2(n20611), .A(n20610), .B(n20609), .ZN(
        P2_U3144) );
  AOI22_X1 U23652 ( .A1(n20621), .A2(n20743), .B1(n20620), .B2(n20742), .ZN(
        n20613) );
  AOI22_X1 U23653 ( .A1(n20669), .A2(n20692), .B1(n20622), .B2(n20744), .ZN(
        n20612) );
  OAI211_X1 U23654 ( .C1(n20626), .C2(n13418), .A(n20613), .B(n20612), .ZN(
        P2_U3145) );
  AOI22_X1 U23655 ( .A1(n20621), .A2(n20761), .B1(n20620), .B2(n20760), .ZN(
        n20615) );
  AOI22_X1 U23656 ( .A1(n20669), .A2(n20704), .B1(n20622), .B2(n20762), .ZN(
        n20614) );
  OAI211_X1 U23657 ( .C1(n20626), .C2(n13491), .A(n20615), .B(n20614), .ZN(
        P2_U3148) );
  AOI22_X1 U23658 ( .A1(n20621), .A2(n20767), .B1(n20620), .B2(n9787), .ZN(
        n20617) );
  AOI22_X1 U23659 ( .A1(n20669), .A2(n20708), .B1(n20622), .B2(n20768), .ZN(
        n20616) );
  OAI211_X1 U23660 ( .C1(n20626), .C2(n13515), .A(n20617), .B(n20616), .ZN(
        P2_U3149) );
  AOI22_X1 U23661 ( .A1(n20621), .A2(n20773), .B1(n20620), .B2(n20772), .ZN(
        n20619) );
  AOI22_X1 U23662 ( .A1(n20669), .A2(n20712), .B1(n20622), .B2(n20774), .ZN(
        n20618) );
  OAI211_X1 U23663 ( .C1(n20626), .C2(n13533), .A(n20619), .B(n20618), .ZN(
        P2_U3150) );
  INV_X1 U23664 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20625) );
  AOI22_X1 U23665 ( .A1(n20621), .A2(n20780), .B1(n20620), .B2(n20778), .ZN(
        n20624) );
  AOI22_X1 U23666 ( .A1(n20669), .A2(n20717), .B1(n20622), .B2(n20782), .ZN(
        n20623) );
  OAI211_X1 U23667 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P2_U3151) );
  NAND2_X1 U23668 ( .A1(n20638), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20686) );
  NAND2_X1 U23669 ( .A1(n20686), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20628) );
  NOR2_X1 U23670 ( .A1(n20629), .A2(n20628), .ZN(n20635) );
  AOI21_X1 U23671 ( .B1(n20638), .B2(n11308), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20630) );
  OR2_X1 U23672 ( .A1(n20635), .A2(n20630), .ZN(n20667) );
  OAI22_X1 U23673 ( .A1(n20667), .A2(n20691), .B1(n20686), .B2(n20631), .ZN(
        n20632) );
  INV_X1 U23674 ( .A(n20632), .ZN(n20641) );
  INV_X1 U23675 ( .A(n20735), .ZN(n20634) );
  NOR2_X1 U23676 ( .A1(n20634), .A2(n20633), .ZN(n20639) );
  AOI211_X1 U23677 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20686), .A(n20636), 
        .B(n20635), .ZN(n20637) );
  AOI22_X1 U23678 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20738), .ZN(n20640) );
  OAI211_X1 U23679 ( .C1(n20741), .C2(n20675), .A(n20641), .B(n20640), .ZN(
        P2_U3152) );
  OAI22_X1 U23680 ( .A1(n20667), .A2(n20695), .B1(n20686), .B2(n20642), .ZN(
        n20643) );
  INV_X1 U23681 ( .A(n20643), .ZN(n20645) );
  AOI22_X1 U23682 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20744), .ZN(n20644) );
  OAI211_X1 U23683 ( .C1(n20747), .C2(n20675), .A(n20645), .B(n20644), .ZN(
        P2_U3153) );
  INV_X1 U23684 ( .A(n20748), .ZN(n20646) );
  OAI22_X1 U23685 ( .A1(n20667), .A2(n20699), .B1(n20646), .B2(n20686), .ZN(
        n20647) );
  INV_X1 U23686 ( .A(n20647), .ZN(n20649) );
  AOI22_X1 U23687 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20750), .ZN(n20648) );
  OAI211_X1 U23688 ( .C1(n20753), .C2(n20675), .A(n20649), .B(n20648), .ZN(
        P2_U3154) );
  INV_X1 U23689 ( .A(n20754), .ZN(n20650) );
  OAI22_X1 U23690 ( .A1(n20667), .A2(n20703), .B1(n20650), .B2(n20686), .ZN(
        n20651) );
  INV_X1 U23691 ( .A(n20651), .ZN(n20653) );
  AOI22_X1 U23692 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20756), .ZN(n20652) );
  OAI211_X1 U23693 ( .C1(n20759), .C2(n20675), .A(n20653), .B(n20652), .ZN(
        P2_U3155) );
  OAI22_X1 U23694 ( .A1(n20667), .A2(n20707), .B1(n20686), .B2(n20654), .ZN(
        n20655) );
  INV_X1 U23695 ( .A(n20655), .ZN(n20657) );
  AOI22_X1 U23696 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20762), .ZN(n20656) );
  OAI211_X1 U23697 ( .C1(n20765), .C2(n20675), .A(n20657), .B(n20656), .ZN(
        P2_U3156) );
  INV_X1 U23698 ( .A(n20766), .ZN(n20658) );
  OAI22_X1 U23699 ( .A1(n20667), .A2(n20711), .B1(n20686), .B2(n20658), .ZN(
        n20659) );
  INV_X1 U23700 ( .A(n20659), .ZN(n20661) );
  AOI22_X1 U23701 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20768), .ZN(n20660) );
  OAI211_X1 U23702 ( .C1(n20771), .C2(n20675), .A(n20661), .B(n20660), .ZN(
        P2_U3157) );
  INV_X1 U23703 ( .A(n20772), .ZN(n20662) );
  OAI22_X1 U23704 ( .A1(n20667), .A2(n20715), .B1(n20686), .B2(n20662), .ZN(
        n20663) );
  INV_X1 U23705 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23706 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20774), .ZN(n20664) );
  OAI211_X1 U23707 ( .C1(n20777), .C2(n20675), .A(n20665), .B(n20664), .ZN(
        P2_U3158) );
  INV_X1 U23708 ( .A(n20778), .ZN(n20666) );
  OAI22_X1 U23709 ( .A1(n20667), .A2(n20722), .B1(n20686), .B2(n20666), .ZN(
        n20668) );
  INV_X1 U23710 ( .A(n20668), .ZN(n20672) );
  AOI22_X1 U23711 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20782), .ZN(n20671) );
  OAI211_X1 U23712 ( .C1(n20787), .C2(n20675), .A(n20672), .B(n20671), .ZN(
        P2_U3159) );
  NAND3_X1 U23713 ( .A1(n20682), .A2(n20675), .A3(n20906), .ZN(n20676) );
  AOI22_X1 U23714 ( .A1(n20680), .A2(n20677), .B1(n20559), .B2(n20686), .ZN(
        n20681) );
  AND2_X1 U23715 ( .A1(n20678), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20737) );
  AND2_X1 U23716 ( .A1(n20737), .A2(n20679), .ZN(n20716) );
  AOI22_X1 U23717 ( .A1(n20683), .A2(n20783), .B1(n20716), .B2(n20729), .ZN(
        n20690) );
  AOI21_X1 U23718 ( .B1(n20684), .B2(n11308), .A(n20906), .ZN(n20685) );
  AOI21_X1 U23719 ( .B1(n20687), .B2(n20686), .A(n20685), .ZN(n20688) );
  OAI21_X1 U23720 ( .B1(n20688), .B2(n20716), .A(n20731), .ZN(n20719) );
  AOI22_X1 U23721 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20719), .B1(
        n20718), .B2(n20738), .ZN(n20689) );
  OAI211_X1 U23722 ( .C1(n20723), .C2(n20691), .A(n20690), .B(n20689), .ZN(
        P2_U3160) );
  AOI22_X1 U23723 ( .A1(n20744), .A2(n20718), .B1(n20716), .B2(n20742), .ZN(
        n20694) );
  AOI22_X1 U23724 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20719), .B1(
        n20783), .B2(n20692), .ZN(n20693) );
  OAI211_X1 U23725 ( .C1(n20723), .C2(n20695), .A(n20694), .B(n20693), .ZN(
        P2_U3161) );
  AOI22_X1 U23726 ( .A1(n20696), .A2(n20783), .B1(n20748), .B2(n20716), .ZN(
        n20698) );
  AOI22_X1 U23727 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20719), .B1(
        n20718), .B2(n20750), .ZN(n20697) );
  OAI211_X1 U23728 ( .C1(n20723), .C2(n20699), .A(n20698), .B(n20697), .ZN(
        P2_U3162) );
  AOI22_X1 U23729 ( .A1(n20756), .A2(n20718), .B1(n20754), .B2(n20716), .ZN(
        n20702) );
  AOI22_X1 U23730 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20719), .B1(
        n20783), .B2(n20700), .ZN(n20701) );
  OAI211_X1 U23731 ( .C1(n20723), .C2(n20703), .A(n20702), .B(n20701), .ZN(
        P2_U3163) );
  AOI22_X1 U23732 ( .A1(n20704), .A2(n20783), .B1(n20716), .B2(n20760), .ZN(
        n20706) );
  AOI22_X1 U23733 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20719), .B1(
        n20718), .B2(n20762), .ZN(n20705) );
  OAI211_X1 U23734 ( .C1(n20723), .C2(n20707), .A(n20706), .B(n20705), .ZN(
        P2_U3164) );
  AOI22_X1 U23735 ( .A1(n20768), .A2(n20718), .B1(n20716), .B2(n9787), .ZN(
        n20710) );
  AOI22_X1 U23736 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20719), .B1(
        n20783), .B2(n20708), .ZN(n20709) );
  OAI211_X1 U23737 ( .C1(n20723), .C2(n20711), .A(n20710), .B(n20709), .ZN(
        P2_U3165) );
  AOI22_X1 U23738 ( .A1(n20774), .A2(n20718), .B1(n20716), .B2(n20772), .ZN(
        n20714) );
  AOI22_X1 U23739 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20719), .B1(
        n20783), .B2(n20712), .ZN(n20713) );
  OAI211_X1 U23740 ( .C1(n20723), .C2(n20715), .A(n20714), .B(n20713), .ZN(
        P2_U3166) );
  AOI22_X1 U23741 ( .A1(n20717), .A2(n20783), .B1(n20716), .B2(n20778), .ZN(
        n20721) );
  AOI22_X1 U23742 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20719), .B1(
        n20718), .B2(n20782), .ZN(n20720) );
  OAI211_X1 U23743 ( .C1(n20723), .C2(n20722), .A(n20721), .B(n20720), .ZN(
        P2_U3167) );
  NAND2_X1 U23744 ( .A1(n20728), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20725) );
  NOR2_X1 U23745 ( .A1(n20726), .A2(n20725), .ZN(n20733) );
  AOI21_X1 U23746 ( .B1(n20737), .B2(n11308), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20727) );
  INV_X1 U23747 ( .A(n20728), .ZN(n20779) );
  AOI22_X1 U23748 ( .A1(n20781), .A2(n20730), .B1(n20779), .B2(n20729), .ZN(
        n20740) );
  OAI21_X1 U23749 ( .B1(n20779), .B2(n11308), .A(n20731), .ZN(n20732) );
  NOR2_X1 U23750 ( .A1(n20733), .A2(n20732), .ZN(n20734) );
  OAI221_X1 U23751 ( .B1(n20737), .B2(n20736), .C1(n20737), .C2(n20735), .A(
        n20734), .ZN(n20784) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20738), .ZN(n20739) );
  OAI211_X1 U23753 ( .C1(n20741), .C2(n20256), .A(n20740), .B(n20739), .ZN(
        P2_U3168) );
  AOI22_X1 U23754 ( .A1(n20781), .A2(n20743), .B1(n20779), .B2(n20742), .ZN(
        n20746) );
  AOI22_X1 U23755 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20744), .ZN(n20745) );
  OAI211_X1 U23756 ( .C1(n20747), .C2(n20256), .A(n20746), .B(n20745), .ZN(
        P2_U3169) );
  AOI22_X1 U23757 ( .A1(n20781), .A2(n20749), .B1(n20779), .B2(n20748), .ZN(
        n20752) );
  AOI22_X1 U23758 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20750), .ZN(n20751) );
  OAI211_X1 U23759 ( .C1(n20753), .C2(n20256), .A(n20752), .B(n20751), .ZN(
        P2_U3170) );
  AOI22_X1 U23760 ( .A1(n20781), .A2(n20755), .B1(n20779), .B2(n20754), .ZN(
        n20758) );
  AOI22_X1 U23761 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20756), .ZN(n20757) );
  OAI211_X1 U23762 ( .C1(n20759), .C2(n20256), .A(n20758), .B(n20757), .ZN(
        P2_U3171) );
  AOI22_X1 U23763 ( .A1(n20781), .A2(n20761), .B1(n20779), .B2(n20760), .ZN(
        n20764) );
  AOI22_X1 U23764 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20762), .ZN(n20763) );
  OAI211_X1 U23765 ( .C1(n20765), .C2(n20256), .A(n20764), .B(n20763), .ZN(
        P2_U3172) );
  AOI22_X1 U23766 ( .A1(n20781), .A2(n20767), .B1(n20779), .B2(n9787), .ZN(
        n20770) );
  AOI22_X1 U23767 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20768), .ZN(n20769) );
  OAI211_X1 U23768 ( .C1(n20771), .C2(n20256), .A(n20770), .B(n20769), .ZN(
        P2_U3173) );
  AOI22_X1 U23769 ( .A1(n20781), .A2(n20773), .B1(n20779), .B2(n20772), .ZN(
        n20776) );
  AOI22_X1 U23770 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20774), .ZN(n20775) );
  OAI211_X1 U23771 ( .C1(n20777), .C2(n20256), .A(n20776), .B(n20775), .ZN(
        P2_U3174) );
  AOI22_X1 U23772 ( .A1(n20781), .A2(n20780), .B1(n20779), .B2(n20778), .ZN(
        n20786) );
  AOI22_X1 U23773 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20784), .B1(
        n20783), .B2(n20782), .ZN(n20785) );
  OAI211_X1 U23774 ( .C1(n20787), .C2(n20256), .A(n20786), .B(n20785), .ZN(
        P2_U3175) );
  AND2_X1 U23775 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20788), .ZN(
        P2_U3179) );
  AND2_X1 U23776 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20788), .ZN(
        P2_U3180) );
  AND2_X1 U23777 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20788), .ZN(
        P2_U3181) );
  AND2_X1 U23778 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20788), .ZN(
        P2_U3182) );
  AND2_X1 U23779 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20788), .ZN(
        P2_U3183) );
  AND2_X1 U23780 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20788), .ZN(
        P2_U3184) );
  AND2_X1 U23781 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20788), .ZN(
        P2_U3185) );
  AND2_X1 U23782 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20788), .ZN(
        P2_U3186) );
  AND2_X1 U23783 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20788), .ZN(
        P2_U3187) );
  AND2_X1 U23784 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20788), .ZN(
        P2_U3188) );
  AND2_X1 U23785 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20788), .ZN(
        P2_U3189) );
  AND2_X1 U23786 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20788), .ZN(
        P2_U3190) );
  AND2_X1 U23787 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20788), .ZN(
        P2_U3191) );
  AND2_X1 U23788 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20788), .ZN(
        P2_U3192) );
  AND2_X1 U23789 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20788), .ZN(
        P2_U3193) );
  AND2_X1 U23790 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20788), .ZN(
        P2_U3194) );
  AND2_X1 U23791 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20788), .ZN(
        P2_U3195) );
  AND2_X1 U23792 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20788), .ZN(
        P2_U3196) );
  AND2_X1 U23793 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20788), .ZN(
        P2_U3197) );
  AND2_X1 U23794 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20788), .ZN(
        P2_U3198) );
  AND2_X1 U23795 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20788), .ZN(
        P2_U3199) );
  AND2_X1 U23796 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20788), .ZN(
        P2_U3200) );
  AND2_X1 U23797 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20788), .ZN(P2_U3201) );
  AND2_X1 U23798 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20788), .ZN(P2_U3202) );
  AND2_X1 U23799 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20788), .ZN(P2_U3203) );
  AND2_X1 U23800 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20788), .ZN(P2_U3204) );
  AND2_X1 U23801 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20788), .ZN(P2_U3205) );
  AND2_X1 U23802 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20788), .ZN(P2_U3206) );
  AND2_X1 U23803 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20788), .ZN(P2_U3207) );
  AND2_X1 U23804 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20788), .ZN(P2_U3208) );
  INV_X1 U23805 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20921) );
  NOR2_X1 U23806 ( .A1(n20917), .A2(n20799), .ZN(n20797) );
  OR3_X1 U23807 ( .A1(n20921), .A2(n20789), .A3(n20797), .ZN(n20790) );
  INV_X1 U23808 ( .A(NA), .ZN(n21388) );
  NOR3_X1 U23809 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21388), .ZN(n20803) );
  AOI21_X1 U23810 ( .B1(n20806), .B2(n20790), .A(n20803), .ZN(n20791) );
  OAI221_X1 U23811 ( .B1(n20792), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20792), .C2(n19925), .A(n20791), .ZN(P2_U3209) );
  AOI21_X1 U23812 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19925), .A(n20806), 
        .ZN(n20800) );
  NOR3_X1 U23813 ( .A1(n20800), .A2(n20921), .A3(n20789), .ZN(n20793) );
  NOR2_X1 U23814 ( .A1(n20793), .A2(n20797), .ZN(n20795) );
  OAI211_X1 U23815 ( .C1(n19925), .C2(n20796), .A(n20795), .B(n20794), .ZN(
        P2_U3210) );
  AOI22_X1 U23816 ( .A1(n20798), .A2(n20921), .B1(n20797), .B2(n21388), .ZN(
        n20805) );
  OAI21_X1 U23817 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20804) );
  NOR2_X1 U23818 ( .A1(n20799), .A2(n20806), .ZN(n20801) );
  AOI21_X1 U23819 ( .B1(n20801), .B2(n20910), .A(n20800), .ZN(n20802) );
  OAI22_X1 U23820 ( .A1(n20805), .A2(n20804), .B1(n20803), .B2(n20802), .ZN(
        P2_U3211) );
  NAND2_X2 U23821 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20856), .ZN(n20855) );
  NAND2_X2 U23822 ( .A1(n20856), .A2(n20806), .ZN(n20859) );
  OAI222_X1 U23823 ( .A1(n20855), .A2(n20808), .B1(n20807), .B2(n20856), .C1(
        n20809), .C2(n20859), .ZN(P2_U3212) );
  OAI222_X1 U23824 ( .A1(n20859), .A2(n20811), .B1(n20810), .B2(n20856), .C1(
        n20809), .C2(n20855), .ZN(P2_U3213) );
  OAI222_X1 U23825 ( .A1(n20859), .A2(n11104), .B1(n20812), .B2(n20856), .C1(
        n20811), .C2(n20855), .ZN(P2_U3214) );
  OAI222_X1 U23826 ( .A1(n20859), .A2(n11346), .B1(n20813), .B2(n20856), .C1(
        n11104), .C2(n20855), .ZN(P2_U3215) );
  OAI222_X1 U23827 ( .A1(n20859), .A2(n20815), .B1(n20814), .B2(n20856), .C1(
        n11346), .C2(n20855), .ZN(P2_U3216) );
  OAI222_X1 U23828 ( .A1(n20859), .A2(n20817), .B1(n20816), .B2(n20856), .C1(
        n20815), .C2(n20855), .ZN(P2_U3217) );
  OAI222_X1 U23829 ( .A1(n20859), .A2(n20819), .B1(n20818), .B2(n20856), .C1(
        n20817), .C2(n20855), .ZN(P2_U3218) );
  OAI222_X1 U23830 ( .A1(n20859), .A2(n20821), .B1(n20820), .B2(n20856), .C1(
        n20819), .C2(n20855), .ZN(P2_U3219) );
  OAI222_X1 U23831 ( .A1(n20859), .A2(n16721), .B1(n20822), .B2(n20856), .C1(
        n20821), .C2(n20855), .ZN(P2_U3220) );
  OAI222_X1 U23832 ( .A1(n20859), .A2(n16706), .B1(n20823), .B2(n20856), .C1(
        n16721), .C2(n20855), .ZN(P2_U3221) );
  OAI222_X1 U23833 ( .A1(n20859), .A2(n16685), .B1(n20824), .B2(n20856), .C1(
        n16706), .C2(n20855), .ZN(P2_U3222) );
  OAI222_X1 U23834 ( .A1(n20859), .A2(n16675), .B1(n20825), .B2(n20856), .C1(
        n16685), .C2(n20855), .ZN(P2_U3223) );
  OAI222_X1 U23835 ( .A1(n20859), .A2(n20827), .B1(n20826), .B2(n20856), .C1(
        n16675), .C2(n20855), .ZN(P2_U3224) );
  OAI222_X1 U23836 ( .A1(n20859), .A2(n20829), .B1(n20828), .B2(n20856), .C1(
        n20827), .C2(n20855), .ZN(P2_U3225) );
  OAI222_X1 U23837 ( .A1(n20859), .A2(n16643), .B1(n20830), .B2(n20856), .C1(
        n20829), .C2(n20855), .ZN(P2_U3226) );
  OAI222_X1 U23838 ( .A1(n20859), .A2(n20832), .B1(n20831), .B2(n20856), .C1(
        n16643), .C2(n20855), .ZN(P2_U3227) );
  OAI222_X1 U23839 ( .A1(n20859), .A2(n20834), .B1(n20833), .B2(n20856), .C1(
        n20832), .C2(n20855), .ZN(P2_U3228) );
  OAI222_X1 U23840 ( .A1(n20859), .A2(n20836), .B1(n20835), .B2(n20856), .C1(
        n20834), .C2(n20855), .ZN(P2_U3229) );
  OAI222_X1 U23841 ( .A1(n20859), .A2(n16000), .B1(n20837), .B2(n20856), .C1(
        n20836), .C2(n20855), .ZN(P2_U3230) );
  OAI222_X1 U23842 ( .A1(n20859), .A2(n20839), .B1(n20838), .B2(n20856), .C1(
        n16000), .C2(n20855), .ZN(P2_U3231) );
  OAI222_X1 U23843 ( .A1(n20859), .A2(n16589), .B1(n20840), .B2(n20856), .C1(
        n20839), .C2(n20855), .ZN(P2_U3232) );
  OAI222_X1 U23844 ( .A1(n20859), .A2(n20842), .B1(n20841), .B2(n20856), .C1(
        n16589), .C2(n20855), .ZN(P2_U3233) );
  OAI222_X1 U23845 ( .A1(n20859), .A2(n20844), .B1(n20843), .B2(n20856), .C1(
        n20842), .C2(n20855), .ZN(P2_U3234) );
  OAI222_X1 U23846 ( .A1(n20859), .A2(n20846), .B1(n20845), .B2(n20856), .C1(
        n20844), .C2(n20855), .ZN(P2_U3235) );
  OAI222_X1 U23847 ( .A1(n20859), .A2(n20848), .B1(n20847), .B2(n20856), .C1(
        n20846), .C2(n20855), .ZN(P2_U3236) );
  OAI222_X1 U23848 ( .A1(n20859), .A2(n20851), .B1(n20849), .B2(n20856), .C1(
        n20848), .C2(n20855), .ZN(P2_U3237) );
  OAI222_X1 U23849 ( .A1(n20855), .A2(n20851), .B1(n20850), .B2(n20856), .C1(
        n15868), .C2(n20859), .ZN(P2_U3238) );
  OAI222_X1 U23850 ( .A1(n20859), .A2(n20853), .B1(n20852), .B2(n20856), .C1(
        n15868), .C2(n20855), .ZN(P2_U3239) );
  OAI222_X1 U23851 ( .A1(n20859), .A2(n12844), .B1(n20854), .B2(n20856), .C1(
        n20853), .C2(n20855), .ZN(P2_U3240) );
  OAI222_X1 U23852 ( .A1(n20859), .A2(n20858), .B1(n20857), .B2(n20856), .C1(
        n12844), .C2(n20855), .ZN(P2_U3241) );
  OAI22_X1 U23853 ( .A1(n20924), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20856), .ZN(n20860) );
  INV_X1 U23854 ( .A(n20860), .ZN(P2_U3585) );
  MUX2_X1 U23855 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20924), .Z(P2_U3586) );
  AOI22_X1 U23856 ( .A1(n20856), .A2(n20862), .B1(n20861), .B2(n20924), .ZN(
        P2_U3587) );
  OAI22_X1 U23857 ( .A1(n20924), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20856), .ZN(n20863) );
  INV_X1 U23858 ( .A(n20863), .ZN(P2_U3588) );
  OAI21_X1 U23859 ( .B1(n20867), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20865), 
        .ZN(n20864) );
  INV_X1 U23860 ( .A(n20864), .ZN(P2_U3591) );
  OAI21_X1 U23861 ( .B1(n20867), .B2(n20866), .A(n20865), .ZN(P2_U3592) );
  INV_X1 U23862 ( .A(n20892), .ZN(n20895) );
  INV_X1 U23863 ( .A(n20868), .ZN(n20869) );
  NAND2_X1 U23864 ( .A1(n20870), .A2(n20869), .ZN(n20886) );
  OR2_X1 U23865 ( .A1(n20871), .A2(n20881), .ZN(n20875) );
  AND2_X1 U23866 ( .A1(n20873), .A2(n20872), .ZN(n20874) );
  AND2_X1 U23867 ( .A1(n20875), .A2(n20874), .ZN(n20888) );
  NAND2_X1 U23868 ( .A1(n20886), .A2(n20888), .ZN(n20877) );
  NAND2_X1 U23869 ( .A1(n20877), .A2(n20876), .ZN(n20880) );
  NAND2_X1 U23870 ( .A1(n20878), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20879) );
  OAI211_X1 U23871 ( .C1(n20882), .C2(n20881), .A(n20880), .B(n20879), .ZN(
        n20883) );
  INV_X1 U23872 ( .A(n20883), .ZN(n20884) );
  AOI22_X1 U23873 ( .A1(n20895), .A2(n20885), .B1(n20884), .B2(n20892), .ZN(
        P2_U3602) );
  INV_X1 U23874 ( .A(n20886), .ZN(n20891) );
  OAI22_X1 U23875 ( .A1(n20889), .A2(n20888), .B1(n20887), .B2(n11308), .ZN(
        n20890) );
  NOR2_X1 U23876 ( .A1(n20891), .A2(n20890), .ZN(n20893) );
  AOI22_X1 U23877 ( .A1(n20895), .A2(n20894), .B1(n20893), .B2(n20892), .ZN(
        P2_U3603) );
  AOI22_X1 U23878 ( .A1(n20856), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20896), 
        .B2(n20924), .ZN(P2_U3608) );
  INV_X1 U23879 ( .A(n20897), .ZN(n20905) );
  INV_X1 U23880 ( .A(n20898), .ZN(n20901) );
  INV_X1 U23881 ( .A(n20899), .ZN(n20900) );
  AOI21_X1 U23882 ( .B1(n20902), .B2(n20901), .A(n20900), .ZN(n20904) );
  NAND2_X1 U23883 ( .A1(n20905), .A2(P2_MORE_REG_SCAN_IN), .ZN(n20903) );
  OAI21_X1 U23884 ( .B1(n20905), .B2(n20904), .A(n20903), .ZN(P2_U3609) );
  AOI21_X1 U23885 ( .B1(n10130), .B2(n11308), .A(n20906), .ZN(n20907) );
  OAI211_X1 U23886 ( .C1(n20910), .C2(n20909), .A(n20908), .B(n20907), .ZN(
        n20922) );
  OAI22_X1 U23887 ( .A1(n20913), .A2(P2_STATEBS16_REG_SCAN_IN), .B1(n20912), 
        .B2(n20911), .ZN(n20914) );
  AND2_X1 U23888 ( .A1(n20915), .A2(n20914), .ZN(n20919) );
  AOI21_X1 U23889 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20917), .A(n20916), 
        .ZN(n20918) );
  OAI21_X1 U23890 ( .B1(n20919), .B2(n20918), .A(n20922), .ZN(n20920) );
  OAI21_X1 U23891 ( .B1(n20922), .B2(n20921), .A(n20920), .ZN(P2_U3610) );
  OAI22_X1 U23892 ( .A1(n20924), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20856), .ZN(n20925) );
  INV_X1 U23893 ( .A(n20925), .ZN(P2_U3611) );
  NOR2_X1 U23894 ( .A1(n21383), .A2(n21390), .ZN(n21392) );
  INV_X1 U23895 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20926) );
  AOI21_X1 U23896 ( .B1(n21392), .B2(n20926), .A(n21461), .ZN(P1_U2802) );
  OAI21_X1 U23897 ( .B1(n20928), .B2(n20927), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20929) );
  OAI21_X1 U23898 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20930), .A(n20929), 
        .ZN(P1_U2803) );
  INV_X2 U23899 ( .A(n21461), .ZN(n21476) );
  NOR2_X1 U23900 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21382) );
  OAI21_X1 U23901 ( .B1(n21382), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21476), .ZN(
        n20931) );
  OAI21_X1 U23902 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21476), .A(n20931), 
        .ZN(P1_U2804) );
  OAI21_X1 U23903 ( .B1(BS16), .B2(n21382), .A(n21450), .ZN(n21448) );
  OAI21_X1 U23904 ( .B1(n21450), .B2(n21204), .A(n21448), .ZN(P1_U2805) );
  OAI21_X1 U23905 ( .B1(n20934), .B2(n20933), .A(n20932), .ZN(P1_U2806) );
  AOI211_X1 U23906 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20935) );
  NAND4_X1 U23907 ( .A1(n20936), .A2(n20935), .A3(n21374), .A4(n21376), .ZN(
        n20944) );
  OR4_X1 U23908 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20943) );
  OR4_X1 U23909 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20942) );
  NOR4_X1 U23910 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20940) );
  NOR4_X1 U23911 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20939) );
  NOR4_X1 U23912 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20938) );
  NOR4_X1 U23913 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20937) );
  NAND4_X1 U23914 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20941) );
  NOR4_X2 U23915 ( .A1(n20944), .A2(n20943), .A3(n20942), .A4(n20941), .ZN(
        n21459) );
  INV_X1 U23916 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20946) );
  NOR3_X1 U23917 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20947) );
  OAI21_X1 U23918 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20947), .A(n21459), .ZN(
        n20945) );
  OAI21_X1 U23919 ( .B1(n21459), .B2(n20946), .A(n20945), .ZN(P1_U2807) );
  INV_X1 U23920 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20949) );
  NOR2_X1 U23921 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21453) );
  OAI21_X1 U23922 ( .B1(n20947), .B2(n21453), .A(n21459), .ZN(n20948) );
  OAI21_X1 U23923 ( .B1(n21459), .B2(n20949), .A(n20948), .ZN(P1_U2808) );
  AOI22_X1 U23924 ( .A1(n20951), .A2(n21018), .B1(n21013), .B2(n20950), .ZN(
        n20962) );
  AOI21_X1 U23925 ( .B1(n21016), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20952), .ZN(n20953) );
  OAI21_X1 U23926 ( .B1(n21006), .B2(n20954), .A(n20953), .ZN(n20955) );
  AOI21_X1 U23927 ( .B1(n20957), .B2(n20956), .A(n20955), .ZN(n20961) );
  AOI22_X1 U23928 ( .A1(n20959), .A2(n20989), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20958), .ZN(n20960) );
  NAND3_X1 U23929 ( .A1(n20962), .A2(n20961), .A3(n20960), .ZN(P1_U2831) );
  NOR3_X1 U23930 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20968), .A3(n20963), .ZN(
        n20966) );
  OAI21_X1 U23931 ( .B1(n21006), .B2(n20964), .A(n20998), .ZN(n20965) );
  NOR2_X1 U23932 ( .A1(n20966), .A2(n20965), .ZN(n20979) );
  NOR2_X1 U23933 ( .A1(n20967), .A2(n20983), .ZN(n20976) );
  INV_X1 U23934 ( .A(n20968), .ZN(n20969) );
  NOR2_X1 U23935 ( .A1(n20970), .A2(n20969), .ZN(n20971) );
  NOR2_X1 U23936 ( .A1(n20972), .A2(n20971), .ZN(n20984) );
  OAI22_X1 U23937 ( .A1(n20974), .A2(n20973), .B1(n20984), .B2(n21406), .ZN(
        n20975) );
  AOI211_X1 U23938 ( .C1(n20977), .C2(n21013), .A(n20976), .B(n20975), .ZN(
        n20978) );
  OAI211_X1 U23939 ( .C1(n20981), .C2(n20980), .A(n20979), .B(n20978), .ZN(
        P1_U2833) );
  AOI22_X1 U23940 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n21016), .B1(
        n21013), .B2(n21029), .ZN(n20991) );
  OAI22_X1 U23941 ( .A1(n20983), .A2(n20982), .B1(n21034), .B2(n21006), .ZN(
        n20988) );
  INV_X1 U23942 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20986) );
  AOI21_X1 U23943 ( .B1(n20986), .B2(n20985), .A(n20984), .ZN(n20987) );
  AOI211_X1 U23944 ( .C1(n20989), .C2(n21032), .A(n20988), .B(n20987), .ZN(
        n20990) );
  NAND3_X1 U23945 ( .A1(n20991), .A2(n20990), .A3(n20998), .ZN(P1_U2834) );
  INV_X1 U23946 ( .A(n21105), .ZN(n20992) );
  NAND2_X1 U23947 ( .A1(n21018), .A2(n20992), .ZN(n20999) );
  INV_X1 U23948 ( .A(n21020), .ZN(n20993) );
  NAND2_X1 U23949 ( .A1(n20994), .A2(n20993), .ZN(n20997) );
  NAND2_X1 U23950 ( .A1(n21016), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20996) );
  AND4_X1 U23951 ( .A1(n20999), .A2(n20998), .A3(n20997), .A4(n20996), .ZN(
        n21010) );
  NOR2_X1 U23952 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21000), .ZN(n21001) );
  NAND2_X1 U23953 ( .A1(n21002), .A2(n21001), .ZN(n21005) );
  INV_X1 U23954 ( .A(n21003), .ZN(n21107) );
  NAND2_X1 U23955 ( .A1(n21013), .A2(n21107), .ZN(n21004) );
  OAI211_X1 U23956 ( .C1(n21007), .C2(n21006), .A(n21005), .B(n21004), .ZN(
        n21008) );
  AOI21_X1 U23957 ( .B1(n21100), .B2(n21024), .A(n21008), .ZN(n21009) );
  OAI211_X1 U23958 ( .C1(n21011), .C2(n21399), .A(n21010), .B(n21009), .ZN(
        P1_U2836) );
  INV_X1 U23959 ( .A(n21012), .ZN(n21125) );
  AOI22_X1 U23960 ( .A1(n21014), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n21013), .B2(
        n21125), .ZN(n21027) );
  INV_X1 U23961 ( .A(n21015), .ZN(n21017) );
  AOI22_X1 U23962 ( .A1(n21018), .A2(n21017), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n21016), .ZN(n21019) );
  OAI21_X1 U23963 ( .B1(n14232), .B2(n21020), .A(n21019), .ZN(n21023) );
  INV_X1 U23964 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21397) );
  NOR2_X1 U23965 ( .A1(n21021), .A2(n21397), .ZN(n21022) );
  AOI211_X1 U23966 ( .C1(n21025), .C2(n21024), .A(n21023), .B(n21022), .ZN(
        n21026) );
  OAI211_X1 U23967 ( .C1(n14111), .C2(n21028), .A(n21027), .B(n21026), .ZN(
        P1_U2838) );
  AOI22_X1 U23968 ( .A1(n21032), .A2(n21031), .B1(n21030), .B2(n21029), .ZN(
        n21033) );
  OAI21_X1 U23969 ( .B1(n21035), .B2(n21034), .A(n21033), .ZN(P1_U2866) );
  AOI22_X1 U23970 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21036) );
  OAI21_X1 U23971 ( .B1(n21037), .B2(n21069), .A(n21036), .ZN(P1_U2921) );
  INV_X1 U23972 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21039) );
  AOI22_X1 U23973 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21038) );
  OAI21_X1 U23974 ( .B1(n21039), .B2(n21069), .A(n21038), .ZN(P1_U2922) );
  INV_X1 U23975 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U23976 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21040) );
  OAI21_X1 U23977 ( .B1(n21041), .B2(n21069), .A(n21040), .ZN(P1_U2923) );
  AOI22_X1 U23978 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21042) );
  OAI21_X1 U23979 ( .B1(n21043), .B2(n21069), .A(n21042), .ZN(P1_U2924) );
  AOI22_X1 U23980 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n21044), .B1(n21055), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21045) );
  OAI21_X1 U23981 ( .B1(n21046), .B2(n21466), .A(n21045), .ZN(P1_U2925) );
  INV_X1 U23982 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21048) );
  AOI22_X1 U23983 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21047) );
  OAI21_X1 U23984 ( .B1(n21048), .B2(n21069), .A(n21047), .ZN(P1_U2926) );
  INV_X1 U23985 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U23986 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n21049) );
  OAI21_X1 U23987 ( .B1(n21050), .B2(n21069), .A(n21049), .ZN(P1_U2927) );
  AOI22_X1 U23988 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21051) );
  OAI21_X1 U23989 ( .B1(n21052), .B2(n21069), .A(n21051), .ZN(P1_U2928) );
  AOI22_X1 U23990 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n21053) );
  OAI21_X1 U23991 ( .B1(n21054), .B2(n21069), .A(n21053), .ZN(P1_U2929) );
  AOI22_X1 U23992 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21056) );
  OAI21_X1 U23993 ( .B1(n21057), .B2(n21069), .A(n21056), .ZN(P1_U2930) );
  AOI22_X1 U23994 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21058) );
  OAI21_X1 U23995 ( .B1(n11875), .B2(n21069), .A(n21058), .ZN(P1_U2931) );
  AOI22_X1 U23996 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21059) );
  OAI21_X1 U23997 ( .B1(n21060), .B2(n21069), .A(n21059), .ZN(P1_U2932) );
  AOI22_X1 U23998 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21061) );
  OAI21_X1 U23999 ( .B1(n21062), .B2(n21069), .A(n21061), .ZN(P1_U2933) );
  AOI22_X1 U24000 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21063) );
  OAI21_X1 U24001 ( .B1(n21064), .B2(n21069), .A(n21063), .ZN(P1_U2934) );
  AOI22_X1 U24002 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n21065) );
  OAI21_X1 U24003 ( .B1(n21066), .B2(n21069), .A(n21065), .ZN(P1_U2935) );
  AOI22_X1 U24004 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21067), .B1(n21055), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n21068) );
  OAI21_X1 U24005 ( .B1(n21070), .B2(n21069), .A(n21068), .ZN(P1_U2936) );
  AOI22_X1 U24006 ( .A1(n21091), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n21090), .ZN(n21072) );
  NAND2_X1 U24007 ( .A1(n21080), .A2(n21071), .ZN(n21082) );
  NAND2_X1 U24008 ( .A1(n21072), .A2(n21082), .ZN(P1_U2946) );
  AOI22_X1 U24009 ( .A1(n21091), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n21090), .ZN(n21074) );
  NAND2_X1 U24010 ( .A1(n21080), .A2(n21073), .ZN(n21084) );
  NAND2_X1 U24011 ( .A1(n21074), .A2(n21084), .ZN(P1_U2947) );
  AOI22_X1 U24012 ( .A1(n21091), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n21090), .ZN(n21076) );
  NAND2_X1 U24013 ( .A1(n21080), .A2(n21075), .ZN(n21086) );
  NAND2_X1 U24014 ( .A1(n21076), .A2(n21086), .ZN(P1_U2948) );
  AOI22_X1 U24015 ( .A1(n21091), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n21090), .ZN(n21078) );
  NAND2_X1 U24016 ( .A1(n21080), .A2(n21077), .ZN(n21088) );
  NAND2_X1 U24017 ( .A1(n21078), .A2(n21088), .ZN(P1_U2950) );
  AOI22_X1 U24018 ( .A1(n21091), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n21090), .ZN(n21081) );
  NAND2_X1 U24019 ( .A1(n21080), .A2(n21079), .ZN(n21092) );
  NAND2_X1 U24020 ( .A1(n21081), .A2(n21092), .ZN(P1_U2951) );
  AOI22_X1 U24021 ( .A1(n21091), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21090), .ZN(n21083) );
  NAND2_X1 U24022 ( .A1(n21083), .A2(n21082), .ZN(P1_U2961) );
  AOI22_X1 U24023 ( .A1(n21091), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n21090), .ZN(n21085) );
  NAND2_X1 U24024 ( .A1(n21085), .A2(n21084), .ZN(P1_U2962) );
  AOI22_X1 U24025 ( .A1(n21091), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n21090), .ZN(n21087) );
  NAND2_X1 U24026 ( .A1(n21087), .A2(n21086), .ZN(P1_U2963) );
  AOI22_X1 U24027 ( .A1(n21091), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n21090), .ZN(n21089) );
  NAND2_X1 U24028 ( .A1(n21089), .A2(n21088), .ZN(P1_U2965) );
  AOI22_X1 U24029 ( .A1(n21091), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n21090), .ZN(n21093) );
  NAND2_X1 U24030 ( .A1(n21093), .A2(n21092), .ZN(P1_U2966) );
  AOI22_X1 U24031 ( .A1(n21094), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n21133), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n21104) );
  AOI21_X1 U24032 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21096), .A(
        n21095), .ZN(n21099) );
  XNOR2_X1 U24033 ( .A(n21097), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n21098) );
  XNOR2_X1 U24034 ( .A(n21099), .B(n21098), .ZN(n21108) );
  AOI22_X1 U24035 ( .A1(n21108), .A2(n21102), .B1(n21101), .B2(n21100), .ZN(
        n21103) );
  OAI211_X1 U24036 ( .C1(n21106), .C2(n21105), .A(n21104), .B(n21103), .ZN(
        P1_U2995) );
  OAI21_X1 U24037 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21113), .ZN(n21111) );
  AOI22_X1 U24038 ( .A1(n21142), .A2(n21107), .B1(n21133), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n21110) );
  AOI22_X1 U24039 ( .A1(n21108), .A2(n21145), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21117), .ZN(n21109) );
  OAI211_X1 U24040 ( .C1(n21112), .C2(n21111), .A(n21110), .B(n21109), .ZN(
        P1_U3027) );
  INV_X1 U24041 ( .A(n21113), .ZN(n21121) );
  INV_X1 U24042 ( .A(n21114), .ZN(n21116) );
  AOI21_X1 U24043 ( .B1(n21142), .B2(n21116), .A(n21115), .ZN(n21120) );
  AOI22_X1 U24044 ( .A1(n21118), .A2(n21145), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21117), .ZN(n21119) );
  OAI211_X1 U24045 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n21121), .A(
        n21120), .B(n21119), .ZN(P1_U3028) );
  NAND2_X1 U24046 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21124) );
  OAI21_X1 U24047 ( .B1(n21124), .B2(n21123), .A(n21122), .ZN(n21126) );
  AOI22_X1 U24048 ( .A1(n21127), .A2(n21126), .B1(n21142), .B2(n21125), .ZN(
        n21138) );
  INV_X1 U24049 ( .A(n21128), .ZN(n21132) );
  OAI21_X1 U24050 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21130), .A(
        n21129), .ZN(n21131) );
  AOI22_X1 U24051 ( .A1(n21132), .A2(n21145), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21131), .ZN(n21137) );
  NAND2_X1 U24052 ( .A1(n21133), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n21136) );
  OR3_X1 U24053 ( .A1(n21149), .A2(n21134), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21135) );
  NAND4_X1 U24054 ( .A1(n21138), .A2(n21137), .A3(n21136), .A4(n21135), .ZN(
        P1_U3029) );
  INV_X1 U24055 ( .A(n21139), .ZN(n21141) );
  AOI21_X1 U24056 ( .B1(n21142), .B2(n21141), .A(n21140), .ZN(n21152) );
  INV_X1 U24057 ( .A(n21143), .ZN(n21146) );
  AOI22_X1 U24058 ( .A1(n21146), .A2(n21145), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21144), .ZN(n21151) );
  NAND3_X1 U24059 ( .A1(n21149), .A2(n21148), .A3(n21147), .ZN(n21150) );
  NAND3_X1 U24060 ( .A1(n21152), .A2(n21151), .A3(n21150), .ZN(P1_U3030) );
  NOR2_X1 U24061 ( .A1(n21154), .A2(n21153), .ZN(P1_U3032) );
  AOI22_X1 U24062 ( .A1(n21164), .A2(n21215), .B1(n21163), .B2(n21322), .ZN(
        n21157) );
  AOI22_X1 U24063 ( .A1(n21323), .A2(n21165), .B1(n21155), .B2(n21324), .ZN(
        n21156) );
  OAI211_X1 U24064 ( .C1(n21158), .C2(n11771), .A(n21157), .B(n21156), .ZN(
        P1_U3034) );
  AOI22_X1 U24065 ( .A1(n21164), .A2(n21231), .B1(n21163), .B2(n21346), .ZN(
        n21160) );
  INV_X1 U24066 ( .A(n21158), .ZN(n21166) );
  AOI22_X1 U24067 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21166), .B1(
        n21347), .B2(n21165), .ZN(n21159) );
  OAI211_X1 U24068 ( .C1(n21234), .C2(n21198), .A(n21160), .B(n21159), .ZN(
        P1_U3038) );
  AOI22_X1 U24069 ( .A1(n21164), .A2(n21235), .B1(n21163), .B2(n21352), .ZN(
        n21162) );
  AOI22_X1 U24070 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21166), .B1(
        n21353), .B2(n21165), .ZN(n21161) );
  OAI211_X1 U24071 ( .C1(n21238), .C2(n21198), .A(n21162), .B(n21161), .ZN(
        P1_U3039) );
  AOI22_X1 U24072 ( .A1(n21164), .A2(n21241), .B1(n21163), .B2(n21359), .ZN(
        n21168) );
  AOI22_X1 U24073 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21166), .B1(
        n21361), .B2(n21165), .ZN(n21167) );
  OAI211_X1 U24074 ( .C1(n21246), .C2(n21198), .A(n21168), .B(n21167), .ZN(
        P1_U3040) );
  OR2_X1 U24075 ( .A1(n21170), .A2(n21309), .ZN(n21172) );
  NOR2_X1 U24076 ( .A1(n21307), .A2(n21173), .ZN(n21192) );
  INV_X1 U24077 ( .A(n21192), .ZN(n21171) );
  OAI22_X1 U24078 ( .A1(n21174), .A2(n21311), .B1(n21173), .B2(n11775), .ZN(
        n21193) );
  AOI22_X1 U24079 ( .A1(n21314), .A2(n21193), .B1(n21313), .B2(n21192), .ZN(
        n21179) );
  OAI21_X1 U24080 ( .B1(n21175), .B2(n21281), .A(n21174), .ZN(n21176) );
  OAI221_X1 U24081 ( .B1(n21285), .B2(n21177), .C1(n21311), .C2(n21176), .A(
        n21315), .ZN(n21195) );
  AOI22_X1 U24082 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21318), .ZN(n21178) );
  OAI211_X1 U24083 ( .C1(n21321), .C2(n21198), .A(n21179), .B(n21178), .ZN(
        P1_U3041) );
  AOI22_X1 U24084 ( .A1(n21323), .A2(n21193), .B1(n21322), .B2(n21192), .ZN(
        n21181) );
  AOI22_X1 U24085 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21324), .ZN(n21180) );
  OAI211_X1 U24086 ( .C1(n21327), .C2(n21198), .A(n21181), .B(n21180), .ZN(
        P1_U3042) );
  AOI22_X1 U24087 ( .A1(n21329), .A2(n21193), .B1(n21328), .B2(n21192), .ZN(
        n21183) );
  AOI22_X1 U24088 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21330), .ZN(n21182) );
  OAI211_X1 U24089 ( .C1(n21333), .C2(n21198), .A(n21183), .B(n21182), .ZN(
        P1_U3043) );
  AOI22_X1 U24090 ( .A1(n21335), .A2(n21193), .B1(n21334), .B2(n21192), .ZN(
        n21185) );
  AOI22_X1 U24091 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21336), .ZN(n21184) );
  OAI211_X1 U24092 ( .C1(n21339), .C2(n21198), .A(n21185), .B(n21184), .ZN(
        P1_U3044) );
  AOI22_X1 U24093 ( .A1(n21341), .A2(n21193), .B1(n21340), .B2(n21192), .ZN(
        n21187) );
  AOI22_X1 U24094 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21342), .ZN(n21186) );
  OAI211_X1 U24095 ( .C1(n21345), .C2(n21198), .A(n21187), .B(n21186), .ZN(
        P1_U3045) );
  AOI22_X1 U24096 ( .A1(n21347), .A2(n21193), .B1(n21346), .B2(n21192), .ZN(
        n21189) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21348), .ZN(n21188) );
  OAI211_X1 U24098 ( .C1(n21351), .C2(n21198), .A(n21189), .B(n21188), .ZN(
        P1_U3046) );
  AOI22_X1 U24099 ( .A1(n21353), .A2(n21193), .B1(n21352), .B2(n21192), .ZN(
        n21191) );
  AOI22_X1 U24100 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21354), .ZN(n21190) );
  OAI211_X1 U24101 ( .C1(n21357), .C2(n21198), .A(n21191), .B(n21190), .ZN(
        P1_U3047) );
  AOI22_X1 U24102 ( .A1(n21361), .A2(n21193), .B1(n21359), .B2(n21192), .ZN(
        n21197) );
  AOI22_X1 U24103 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21195), .B1(
        n21194), .B2(n21362), .ZN(n21196) );
  OAI211_X1 U24104 ( .C1(n21368), .C2(n21198), .A(n21197), .B(n21196), .ZN(
        P1_U3048) );
  NAND3_X1 U24105 ( .A1(n21248), .A2(n21285), .A3(n21206), .ZN(n21200) );
  NOR3_X1 U24106 ( .A1(n21203), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21254) );
  INV_X1 U24107 ( .A(n21254), .ZN(n21249) );
  NOR2_X1 U24108 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21249), .ZN(
        n21239) );
  AOI22_X1 U24109 ( .A1(n21314), .A2(n21240), .B1(n21313), .B2(n21239), .ZN(
        n21213) );
  AOI21_X1 U24110 ( .B1(n21210), .B2(n21275), .A(n21204), .ZN(n21205) );
  AOI21_X1 U24111 ( .B1(n21248), .B2(n21206), .A(n21205), .ZN(n21207) );
  NOR2_X1 U24112 ( .A1(n21207), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21209) );
  AOI22_X1 U24113 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n21242), .B2(n21211), .ZN(n21212) );
  OAI211_X1 U24114 ( .C1(n21214), .C2(n21275), .A(n21213), .B(n21212), .ZN(
        P1_U3065) );
  AOI22_X1 U24115 ( .A1(n21323), .A2(n21240), .B1(n21322), .B2(n21239), .ZN(
        n21217) );
  AOI22_X1 U24116 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n21242), .B2(n21215), .ZN(n21216) );
  OAI211_X1 U24117 ( .C1(n21218), .C2(n21275), .A(n21217), .B(n21216), .ZN(
        P1_U3066) );
  AOI22_X1 U24118 ( .A1(n21329), .A2(n21240), .B1(n21328), .B2(n21239), .ZN(
        n21221) );
  AOI22_X1 U24119 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n21242), .B2(n21219), .ZN(n21220) );
  OAI211_X1 U24120 ( .C1(n21222), .C2(n21275), .A(n21221), .B(n21220), .ZN(
        P1_U3067) );
  AOI22_X1 U24121 ( .A1(n21335), .A2(n21240), .B1(n21334), .B2(n21239), .ZN(
        n21225) );
  AOI22_X1 U24122 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n21242), .B2(n21223), .ZN(n21224) );
  OAI211_X1 U24123 ( .C1(n21226), .C2(n21275), .A(n21225), .B(n21224), .ZN(
        P1_U3068) );
  AOI22_X1 U24124 ( .A1(n21341), .A2(n21240), .B1(n21340), .B2(n21239), .ZN(
        n21229) );
  AOI22_X1 U24125 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n21242), .B2(n21227), .ZN(n21228) );
  OAI211_X1 U24126 ( .C1(n21230), .C2(n21275), .A(n21229), .B(n21228), .ZN(
        P1_U3069) );
  AOI22_X1 U24127 ( .A1(n21347), .A2(n21240), .B1(n21346), .B2(n21239), .ZN(
        n21233) );
  AOI22_X1 U24128 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n21242), .B2(n21231), .ZN(n21232) );
  OAI211_X1 U24129 ( .C1(n21234), .C2(n21275), .A(n21233), .B(n21232), .ZN(
        P1_U3070) );
  AOI22_X1 U24130 ( .A1(n21353), .A2(n21240), .B1(n21352), .B2(n21239), .ZN(
        n21237) );
  AOI22_X1 U24131 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n21242), .B2(n21235), .ZN(n21236) );
  OAI211_X1 U24132 ( .C1(n21238), .C2(n21275), .A(n21237), .B(n21236), .ZN(
        P1_U3071) );
  AOI22_X1 U24133 ( .A1(n21361), .A2(n21240), .B1(n21359), .B2(n21239), .ZN(
        n21245) );
  AOI22_X1 U24134 ( .A1(n21243), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n21242), .B2(n21241), .ZN(n21244) );
  OAI211_X1 U24135 ( .C1(n21246), .C2(n21275), .A(n21245), .B(n21244), .ZN(
        P1_U3072) );
  INV_X1 U24136 ( .A(n21309), .ZN(n21247) );
  NOR2_X1 U24137 ( .A1(n21307), .A2(n21249), .ZN(n21269) );
  AOI21_X1 U24138 ( .B1(n21248), .B2(n21247), .A(n21269), .ZN(n21251) );
  OAI22_X1 U24139 ( .A1(n21251), .A2(n21311), .B1(n21249), .B2(n11775), .ZN(
        n21270) );
  AOI22_X1 U24140 ( .A1(n21314), .A2(n21270), .B1(n21313), .B2(n21269), .ZN(
        n21256) );
  INV_X1 U24141 ( .A(n21250), .ZN(n21252) );
  OAI21_X1 U24142 ( .B1(n21252), .B2(n21281), .A(n21251), .ZN(n21253) );
  OAI221_X1 U24143 ( .B1(n21285), .B2(n21254), .C1(n21311), .C2(n21253), .A(
        n21315), .ZN(n21272) );
  AOI22_X1 U24144 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21318), .ZN(n21255) );
  OAI211_X1 U24145 ( .C1(n21321), .C2(n21275), .A(n21256), .B(n21255), .ZN(
        P1_U3073) );
  AOI22_X1 U24146 ( .A1(n21323), .A2(n21270), .B1(n21322), .B2(n21269), .ZN(
        n21258) );
  AOI22_X1 U24147 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21324), .ZN(n21257) );
  OAI211_X1 U24148 ( .C1(n21327), .C2(n21275), .A(n21258), .B(n21257), .ZN(
        P1_U3074) );
  AOI22_X1 U24149 ( .A1(n21329), .A2(n21270), .B1(n21328), .B2(n21269), .ZN(
        n21260) );
  AOI22_X1 U24150 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21330), .ZN(n21259) );
  OAI211_X1 U24151 ( .C1(n21333), .C2(n21275), .A(n21260), .B(n21259), .ZN(
        P1_U3075) );
  AOI22_X1 U24152 ( .A1(n21335), .A2(n21270), .B1(n21334), .B2(n21269), .ZN(
        n21262) );
  AOI22_X1 U24153 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21336), .ZN(n21261) );
  OAI211_X1 U24154 ( .C1(n21339), .C2(n21275), .A(n21262), .B(n21261), .ZN(
        P1_U3076) );
  AOI22_X1 U24155 ( .A1(n21341), .A2(n21270), .B1(n21340), .B2(n21269), .ZN(
        n21264) );
  AOI22_X1 U24156 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21342), .ZN(n21263) );
  OAI211_X1 U24157 ( .C1(n21345), .C2(n21275), .A(n21264), .B(n21263), .ZN(
        P1_U3077) );
  AOI22_X1 U24158 ( .A1(n21347), .A2(n21270), .B1(n21346), .B2(n21269), .ZN(
        n21266) );
  AOI22_X1 U24159 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21348), .ZN(n21265) );
  OAI211_X1 U24160 ( .C1(n21351), .C2(n21275), .A(n21266), .B(n21265), .ZN(
        P1_U3078) );
  AOI22_X1 U24161 ( .A1(n21353), .A2(n21270), .B1(n21352), .B2(n21269), .ZN(
        n21268) );
  AOI22_X1 U24162 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21354), .ZN(n21267) );
  OAI211_X1 U24163 ( .C1(n21357), .C2(n21275), .A(n21268), .B(n21267), .ZN(
        P1_U3079) );
  AOI22_X1 U24164 ( .A1(n21361), .A2(n21270), .B1(n21359), .B2(n21269), .ZN(
        n21274) );
  AOI22_X1 U24165 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21272), .B1(
        n21271), .B2(n21362), .ZN(n21273) );
  OAI211_X1 U24166 ( .C1(n21368), .C2(n21275), .A(n21274), .B(n21273), .ZN(
        P1_U3080) );
  OR2_X1 U24167 ( .A1(n21276), .A2(n21309), .ZN(n21278) );
  NOR2_X1 U24168 ( .A1(n21307), .A2(n21279), .ZN(n21300) );
  INV_X1 U24169 ( .A(n21300), .ZN(n21277) );
  AND2_X1 U24170 ( .A1(n21278), .A2(n21277), .ZN(n21280) );
  OAI22_X1 U24171 ( .A1(n21280), .A2(n21311), .B1(n21279), .B2(n11775), .ZN(
        n21301) );
  AOI22_X1 U24172 ( .A1(n21314), .A2(n21301), .B1(n21313), .B2(n21300), .ZN(
        n21287) );
  OAI21_X1 U24173 ( .B1(n21282), .B2(n21281), .A(n21280), .ZN(n21283) );
  OAI221_X1 U24174 ( .B1(n21285), .B2(n21284), .C1(n21311), .C2(n21283), .A(
        n21315), .ZN(n21303) );
  AOI22_X1 U24175 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21318), .ZN(n21286) );
  OAI211_X1 U24176 ( .C1(n21321), .C2(n21306), .A(n21287), .B(n21286), .ZN(
        P1_U3105) );
  AOI22_X1 U24177 ( .A1(n21323), .A2(n21301), .B1(n21322), .B2(n21300), .ZN(
        n21289) );
  AOI22_X1 U24178 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21324), .ZN(n21288) );
  OAI211_X1 U24179 ( .C1(n21327), .C2(n21306), .A(n21289), .B(n21288), .ZN(
        P1_U3106) );
  AOI22_X1 U24180 ( .A1(n21329), .A2(n21301), .B1(n21328), .B2(n21300), .ZN(
        n21291) );
  AOI22_X1 U24181 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21330), .ZN(n21290) );
  OAI211_X1 U24182 ( .C1(n21333), .C2(n21306), .A(n21291), .B(n21290), .ZN(
        P1_U3107) );
  AOI22_X1 U24183 ( .A1(n21335), .A2(n21301), .B1(n21334), .B2(n21300), .ZN(
        n21293) );
  AOI22_X1 U24184 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21336), .ZN(n21292) );
  OAI211_X1 U24185 ( .C1(n21339), .C2(n21306), .A(n21293), .B(n21292), .ZN(
        P1_U3108) );
  AOI22_X1 U24186 ( .A1(n21341), .A2(n21301), .B1(n21340), .B2(n21300), .ZN(
        n21295) );
  AOI22_X1 U24187 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21342), .ZN(n21294) );
  OAI211_X1 U24188 ( .C1(n21345), .C2(n21306), .A(n21295), .B(n21294), .ZN(
        P1_U3109) );
  AOI22_X1 U24189 ( .A1(n21347), .A2(n21301), .B1(n21346), .B2(n21300), .ZN(
        n21297) );
  AOI22_X1 U24190 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21348), .ZN(n21296) );
  OAI211_X1 U24191 ( .C1(n21351), .C2(n21306), .A(n21297), .B(n21296), .ZN(
        P1_U3110) );
  AOI22_X1 U24192 ( .A1(n21353), .A2(n21301), .B1(n21352), .B2(n21300), .ZN(
        n21299) );
  AOI22_X1 U24193 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21354), .ZN(n21298) );
  OAI211_X1 U24194 ( .C1(n21357), .C2(n21306), .A(n21299), .B(n21298), .ZN(
        P1_U3111) );
  AOI22_X1 U24195 ( .A1(n21361), .A2(n21301), .B1(n21359), .B2(n21300), .ZN(
        n21305) );
  AOI22_X1 U24196 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21303), .B1(
        n21302), .B2(n21362), .ZN(n21304) );
  OAI211_X1 U24197 ( .C1(n21368), .C2(n21306), .A(n21305), .B(n21304), .ZN(
        P1_U3112) );
  NOR2_X1 U24198 ( .A1(n21307), .A2(n21310), .ZN(n21358) );
  INV_X1 U24199 ( .A(n21358), .ZN(n21312) );
  OAI222_X1 U24200 ( .A1(n21312), .A2(n21311), .B1(n11775), .B2(n21310), .C1(
        n21309), .C2(n21308), .ZN(n21360) );
  AOI22_X1 U24201 ( .A1(n21314), .A2(n21360), .B1(n21313), .B2(n21358), .ZN(
        n21320) );
  AOI22_X1 U24202 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21318), .ZN(n21319) );
  OAI211_X1 U24203 ( .C1(n21321), .C2(n21367), .A(n21320), .B(n21319), .ZN(
        P1_U3137) );
  AOI22_X1 U24204 ( .A1(n21323), .A2(n21360), .B1(n21322), .B2(n21358), .ZN(
        n21326) );
  AOI22_X1 U24205 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21324), .ZN(n21325) );
  OAI211_X1 U24206 ( .C1(n21327), .C2(n21367), .A(n21326), .B(n21325), .ZN(
        P1_U3138) );
  AOI22_X1 U24207 ( .A1(n21329), .A2(n21360), .B1(n21328), .B2(n21358), .ZN(
        n21332) );
  AOI22_X1 U24208 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21330), .ZN(n21331) );
  OAI211_X1 U24209 ( .C1(n21333), .C2(n21367), .A(n21332), .B(n21331), .ZN(
        P1_U3139) );
  AOI22_X1 U24210 ( .A1(n21335), .A2(n21360), .B1(n21334), .B2(n21358), .ZN(
        n21338) );
  AOI22_X1 U24211 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21336), .ZN(n21337) );
  OAI211_X1 U24212 ( .C1(n21339), .C2(n21367), .A(n21338), .B(n21337), .ZN(
        P1_U3140) );
  AOI22_X1 U24213 ( .A1(n21341), .A2(n21360), .B1(n21340), .B2(n21358), .ZN(
        n21344) );
  AOI22_X1 U24214 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21342), .ZN(n21343) );
  OAI211_X1 U24215 ( .C1(n21345), .C2(n21367), .A(n21344), .B(n21343), .ZN(
        P1_U3141) );
  AOI22_X1 U24216 ( .A1(n21347), .A2(n21360), .B1(n21346), .B2(n21358), .ZN(
        n21350) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21348), .ZN(n21349) );
  OAI211_X1 U24218 ( .C1(n21351), .C2(n21367), .A(n21350), .B(n21349), .ZN(
        P1_U3142) );
  AOI22_X1 U24219 ( .A1(n21353), .A2(n21360), .B1(n21352), .B2(n21358), .ZN(
        n21356) );
  AOI22_X1 U24220 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21354), .ZN(n21355) );
  OAI211_X1 U24221 ( .C1(n21357), .C2(n21367), .A(n21356), .B(n21355), .ZN(
        P1_U3143) );
  AOI22_X1 U24222 ( .A1(n21361), .A2(n21360), .B1(n21359), .B2(n21358), .ZN(
        n21366) );
  AOI22_X1 U24223 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21364), .B1(
        n21363), .B2(n21362), .ZN(n21365) );
  OAI211_X1 U24224 ( .C1(n21368), .C2(n21367), .A(n21366), .B(n21365), .ZN(
        P1_U3144) );
  NOR2_X1 U24225 ( .A1(n21369), .A2(n13625), .ZN(n21372) );
  INV_X1 U24226 ( .A(n21370), .ZN(n21371) );
  OAI21_X1 U24227 ( .B1(n21372), .B2(n11775), .A(n21371), .ZN(P1_U3163) );
  NOR2_X1 U24228 ( .A1(n21450), .A2(n21373), .ZN(P1_U3164) );
  INV_X1 U24229 ( .A(n21450), .ZN(n21447) );
  AND2_X1 U24230 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21447), .ZN(
        P1_U3165) );
  AND2_X1 U24231 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21447), .ZN(
        P1_U3166) );
  AND2_X1 U24232 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21447), .ZN(
        P1_U3167) );
  AND2_X1 U24233 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21447), .ZN(
        P1_U3168) );
  NOR2_X1 U24234 ( .A1(n21450), .A2(n21374), .ZN(P1_U3169) );
  AND2_X1 U24235 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21447), .ZN(
        P1_U3170) );
  AND2_X1 U24236 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21447), .ZN(
        P1_U3171) );
  AND2_X1 U24237 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21447), .ZN(
        P1_U3172) );
  AND2_X1 U24238 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21447), .ZN(
        P1_U3173) );
  AND2_X1 U24239 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21447), .ZN(
        P1_U3174) );
  AND2_X1 U24240 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21447), .ZN(
        P1_U3175) );
  AND2_X1 U24241 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21447), .ZN(
        P1_U3176) );
  AND2_X1 U24242 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21447), .ZN(
        P1_U3177) );
  AND2_X1 U24243 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21447), .ZN(
        P1_U3178) );
  AND2_X1 U24244 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21447), .ZN(
        P1_U3179) );
  AND2_X1 U24245 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21447), .ZN(
        P1_U3180) );
  AND2_X1 U24246 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21447), .ZN(
        P1_U3181) );
  NOR2_X1 U24247 ( .A1(n21450), .A2(n21375), .ZN(P1_U3182) );
  AND2_X1 U24248 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21447), .ZN(
        P1_U3183) );
  AND2_X1 U24249 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21447), .ZN(
        P1_U3184) );
  AND2_X1 U24250 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21447), .ZN(
        P1_U3185) );
  AND2_X1 U24251 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21447), .ZN(P1_U3186) );
  AND2_X1 U24252 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21447), .ZN(P1_U3187) );
  AND2_X1 U24253 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21447), .ZN(P1_U3188) );
  AND2_X1 U24254 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21447), .ZN(P1_U3189) );
  AND2_X1 U24255 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21447), .ZN(P1_U3190) );
  AND2_X1 U24256 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21447), .ZN(P1_U3191) );
  NOR2_X1 U24257 ( .A1(n21450), .A2(n21376), .ZN(P1_U3192) );
  AND2_X1 U24258 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21447), .ZN(P1_U3193) );
  INV_X1 U24259 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21378) );
  NAND2_X1 U24260 ( .A1(n21378), .A2(n21377), .ZN(n21381) );
  INV_X1 U24261 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21474) );
  NOR2_X1 U24262 ( .A1(NA), .A2(n21474), .ZN(n21386) );
  INV_X1 U24263 ( .A(n21386), .ZN(n21380) );
  AOI22_X1 U24264 ( .A1(HOLD), .A2(n21381), .B1(n21380), .B2(n21379), .ZN(
        n21385) );
  AOI21_X1 U24265 ( .B1(n21383), .B2(n21467), .A(n21382), .ZN(n21384) );
  OAI21_X1 U24266 ( .B1(n21461), .B2(n21385), .A(n21384), .ZN(P1_U3194) );
  AOI21_X1 U24267 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21386), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n21395) );
  NAND2_X1 U24268 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21461), .ZN(n21433) );
  INV_X1 U24269 ( .A(n21433), .ZN(n21440) );
  AOI211_X1 U24270 ( .C1(n21390), .C2(n21388), .A(n21387), .B(n21440), .ZN(
        n21394) );
  NOR3_X1 U24271 ( .A1(NA), .A2(n21390), .A3(n21389), .ZN(n21391) );
  OAI22_X1 U24272 ( .A1(n21392), .A2(n21391), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21474), .ZN(n21393) );
  OAI22_X1 U24273 ( .A1(n21395), .A2(n21394), .B1(n19925), .B2(n21393), .ZN(
        P1_U3196) );
  AOI22_X1 U24274 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n21440), .ZN(n21396) );
  OAI21_X1 U24275 ( .B1(n21397), .B2(n21436), .A(n21396), .ZN(P1_U3197) );
  AOI22_X1 U24276 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21440), .ZN(n21398) );
  OAI21_X1 U24277 ( .B1(n21401), .B2(n21436), .A(n21398), .ZN(P1_U3198) );
  OAI222_X1 U24278 ( .A1(n21433), .A2(n21401), .B1(n21400), .B2(n21461), .C1(
        n21399), .C2(n21436), .ZN(P1_U3199) );
  AOI222_X1 U24279 ( .A1(n21439), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21440), .ZN(n21402) );
  INV_X1 U24280 ( .A(n21402), .ZN(P1_U3200) );
  AOI222_X1 U24281 ( .A1(n21440), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n21439), .ZN(n21403) );
  INV_X1 U24282 ( .A(n21403), .ZN(P1_U3201) );
  AOI222_X1 U24283 ( .A1(n21440), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n21439), .ZN(n21404) );
  INV_X1 U24284 ( .A(n21404), .ZN(P1_U3202) );
  AOI22_X1 U24285 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21439), .ZN(n21405) );
  OAI21_X1 U24286 ( .B1(n21406), .B2(n21433), .A(n21405), .ZN(P1_U3203) );
  AOI222_X1 U24287 ( .A1(n21439), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n21440), .ZN(n21407) );
  INV_X1 U24288 ( .A(n21407), .ZN(P1_U3204) );
  AOI222_X1 U24289 ( .A1(n21440), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21439), .ZN(n21408) );
  INV_X1 U24290 ( .A(n21408), .ZN(P1_U3205) );
  AOI22_X1 U24291 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n21439), .ZN(n21409) );
  OAI21_X1 U24292 ( .B1(n21410), .B2(n21433), .A(n21409), .ZN(P1_U3206) );
  AOI22_X1 U24293 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21439), .ZN(n21411) );
  OAI21_X1 U24294 ( .B1(n15230), .B2(n21433), .A(n21411), .ZN(P1_U3207) );
  AOI22_X1 U24295 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21440), .ZN(n21412) );
  OAI21_X1 U24296 ( .B1(n15210), .B2(n21436), .A(n21412), .ZN(P1_U3208) );
  AOI222_X1 U24297 ( .A1(n21440), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21439), .ZN(n21413) );
  INV_X1 U24298 ( .A(n21413), .ZN(P1_U3209) );
  AOI222_X1 U24299 ( .A1(n21439), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n21440), .ZN(n21414) );
  INV_X1 U24300 ( .A(n21414), .ZN(P1_U3210) );
  AOI222_X1 U24301 ( .A1(n21440), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n21439), .ZN(n21415) );
  INV_X1 U24302 ( .A(n21415), .ZN(P1_U3211) );
  AOI222_X1 U24303 ( .A1(n21440), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n21439), .ZN(n21416) );
  INV_X1 U24304 ( .A(n21416), .ZN(P1_U3212) );
  AOI22_X1 U24305 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21439), .ZN(n21417) );
  OAI21_X1 U24306 ( .B1(n21418), .B2(n21433), .A(n21417), .ZN(P1_U3213) );
  AOI22_X1 U24307 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n21440), .ZN(n21419) );
  OAI21_X1 U24308 ( .B1(n21420), .B2(n21436), .A(n21419), .ZN(P1_U3214) );
  AOI222_X1 U24309 ( .A1(n21439), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21440), .ZN(n21421) );
  INV_X1 U24310 ( .A(n21421), .ZN(P1_U3215) );
  AOI22_X1 U24311 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n21439), .ZN(n21422) );
  OAI21_X1 U24312 ( .B1(n21423), .B2(n21433), .A(n21422), .ZN(P1_U3216) );
  AOI22_X1 U24313 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n21439), .ZN(n21424) );
  OAI21_X1 U24314 ( .B1(n15122), .B2(n21433), .A(n21424), .ZN(P1_U3217) );
  AOI22_X1 U24315 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21476), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n21440), .ZN(n21425) );
  OAI21_X1 U24316 ( .B1(n21427), .B2(n21436), .A(n21425), .ZN(P1_U3218) );
  AOI22_X1 U24317 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n21439), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21476), .ZN(n21426) );
  OAI21_X1 U24318 ( .B1(n21427), .B2(n21433), .A(n21426), .ZN(P1_U3219) );
  AOI22_X1 U24319 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n21440), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21476), .ZN(n21428) );
  OAI21_X1 U24320 ( .B1(n21429), .B2(n21436), .A(n21428), .ZN(P1_U3220) );
  AOI222_X1 U24321 ( .A1(n21439), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n21440), .ZN(n21430) );
  INV_X1 U24322 ( .A(n21430), .ZN(P1_U3221) );
  AOI222_X1 U24323 ( .A1(n21440), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n21439), .ZN(n21431) );
  INV_X1 U24324 ( .A(n21431), .ZN(P1_U3222) );
  AOI22_X1 U24325 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21439), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21476), .ZN(n21432) );
  OAI21_X1 U24326 ( .B1(n21434), .B2(n21433), .A(n21432), .ZN(P1_U3223) );
  AOI22_X1 U24327 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21440), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21476), .ZN(n21435) );
  OAI21_X1 U24328 ( .B1(n21437), .B2(n21436), .A(n21435), .ZN(P1_U3224) );
  AOI222_X1 U24329 ( .A1(n21440), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n21439), .ZN(n21438) );
  INV_X1 U24330 ( .A(n21438), .ZN(P1_U3225) );
  AOI222_X1 U24331 ( .A1(n21440), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21476), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21439), .ZN(n21441) );
  INV_X1 U24332 ( .A(n21441), .ZN(P1_U3226) );
  OAI22_X1 U24333 ( .A1(n21476), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21461), .ZN(n21442) );
  INV_X1 U24334 ( .A(n21442), .ZN(P1_U3458) );
  OAI22_X1 U24335 ( .A1(n21476), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21461), .ZN(n21443) );
  INV_X1 U24336 ( .A(n21443), .ZN(P1_U3459) );
  OAI22_X1 U24337 ( .A1(n21476), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21461), .ZN(n21444) );
  INV_X1 U24338 ( .A(n21444), .ZN(P1_U3460) );
  OAI22_X1 U24339 ( .A1(n21476), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21461), .ZN(n21445) );
  INV_X1 U24340 ( .A(n21445), .ZN(P1_U3461) );
  INV_X1 U24341 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21452) );
  INV_X1 U24342 ( .A(n21448), .ZN(n21446) );
  AOI21_X1 U24343 ( .B1(n21452), .B2(n21447), .A(n21446), .ZN(P1_U3464) );
  INV_X1 U24344 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21449) );
  OAI21_X1 U24345 ( .B1(n21450), .B2(n21449), .A(n21448), .ZN(P1_U3465) );
  NOR3_X1 U24346 ( .A1(n21452), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n21451) );
  AOI221_X1 U24347 ( .B1(n21453), .B2(n21452), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n21451), .ZN(n21455) );
  INV_X1 U24348 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21454) );
  INV_X1 U24349 ( .A(n21459), .ZN(n21456) );
  AOI22_X1 U24350 ( .A1(n21459), .A2(n21455), .B1(n21454), .B2(n21456), .ZN(
        P1_U3481) );
  NOR2_X1 U24351 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21458) );
  INV_X1 U24352 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21457) );
  AOI22_X1 U24353 ( .A1(n21459), .A2(n21458), .B1(n21457), .B2(n21456), .ZN(
        P1_U3482) );
  AOI22_X1 U24354 ( .A1(n21461), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21460), 
        .B2(n21476), .ZN(P1_U3483) );
  INV_X1 U24355 ( .A(n21462), .ZN(n21465) );
  INV_X1 U24356 ( .A(n21463), .ZN(n21464) );
  OAI211_X1 U24357 ( .C1(n21467), .C2(n21466), .A(n21465), .B(n21464), .ZN(
        n21475) );
  NOR2_X1 U24358 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21468), .ZN(n21473) );
  OAI211_X1 U24359 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21470), .A(n21469), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21471) );
  NAND2_X1 U24360 ( .A1(n21475), .A2(n21471), .ZN(n21472) );
  OAI22_X1 U24361 ( .A1(n21475), .A2(n21474), .B1(n21473), .B2(n21472), .ZN(
        P1_U3485) );
  MUX2_X1 U24362 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n21476), .Z(P1_U3486) );
  INV_X1 U11184 ( .A(n9608), .ZN(n18258) );
  AND3_X1 U13849 ( .A1(n9733), .A2(n10616), .A3(n10615), .ZN(n10617) );
  NOR2_X2 U11158 ( .A1(n10675), .A2(n9605), .ZN(n17176) );
  CLKBUF_X1 U11053 ( .A(n12018), .Z(n12325) );
  CLKBUF_X1 U11054 ( .A(n12637), .Z(n12682) );
  NAND2_X2 U11059 ( .A1(n14299), .A2(n14542), .ZN(n12626) );
  CLKBUF_X1 U11068 ( .A(n12641), .Z(n9610) );
  CLKBUF_X1 U11089 ( .A(n11660), .Z(n14325) );
  CLKBUF_X3 U11093 ( .A(n10803), .Z(n13398) );
  CLKBUF_X1 U11123 ( .A(n11185), .Z(n9626) );
  CLKBUF_X1 U11134 ( .A(n10683), .Z(n10684) );
  CLKBUF_X1 U11140 ( .A(n14235), .Z(n9625) );
  CLKBUF_X2 U11152 ( .A(n11685), .Z(n14436) );
  CLKBUF_X1 U11165 ( .A(n12532), .Z(n15559) );
  AOI211_X1 U11170 ( .C1(n20503), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20502), .ZN(n20504) );
  INV_X2 U11178 ( .A(n19224), .ZN(n19398) );
  CLKBUF_X1 U11376 ( .A(n9605), .Z(n9615) );
  CLKBUF_X1 U11436 ( .A(n17343), .Z(n9612) );
  CLKBUF_X1 U11444 ( .A(n17787), .Z(n17799) );
  NAND2_X1 U11621 ( .A1(n13031), .A2(n14132), .ZN(n21477) );
endmodule

