

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput127,
         keyinput126, keyinput125, keyinput124, keyinput123, keyinput122,
         keyinput121, keyinput120, keyinput119, keyinput118, keyinput117,
         keyinput116, keyinput115, keyinput114, keyinput113, keyinput112,
         keyinput111, keyinput110, keyinput109, keyinput108, keyinput107,
         keyinput106, keyinput105, keyinput104, keyinput103, keyinput102,
         keyinput101, keyinput100, keyinput99, keyinput98, keyinput97,
         keyinput96, keyinput95, keyinput94, keyinput93, keyinput92,
         keyinput91, keyinput90, keyinput89, keyinput88, keyinput87,
         keyinput86, keyinput85, keyinput84, keyinput83, keyinput82,
         keyinput81, keyinput80, keyinput79, keyinput78, keyinput77,
         keyinput76, keyinput75, keyinput74, keyinput73, keyinput72,
         keyinput71, keyinput70, keyinput69, keyinput68, keyinput67,
         keyinput66, keyinput65, keyinput64, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6542, n6543, n6545, n6546, n6548, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482;

  AOI21_X2 U7290 ( .B1(n12213), .B2(n8371), .A(n6698), .ZN(n14344) );
  AND2_X1 U7291 ( .A1(n9567), .A2(n9566), .ZN(n13029) );
  NOR2_X1 U7292 ( .A1(n14656), .A2(n14657), .ZN(n14655) );
  NAND2_X1 U7293 ( .A1(n9116), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9118) );
  XNOR2_X1 U7294 ( .A(n14455), .B(n15301), .ZN(n15476) );
  NAND2_X2 U7295 ( .A1(n12031), .A2(n12030), .ZN(n15084) );
  INV_X2 U7296 ( .A(n12305), .ZN(n12366) );
  CLKBUF_X2 U7297 ( .A(n8349), .Z(n11903) );
  INV_X1 U7298 ( .A(n10685), .ZN(n10846) );
  INV_X1 U7299 ( .A(n8578), .ZN(n6546) );
  AND4_X1 U7300 ( .A1(n8340), .A2(n8339), .A3(n8338), .A4(n8337), .ZN(n11232)
         );
  CLKBUF_X1 U7302 ( .A(n7721), .Z(n8161) );
  AND2_X1 U7303 ( .A1(n14380), .A2(n8303), .ZN(n8346) );
  NAND2_X1 U7304 ( .A1(n8774), .A2(n8773), .ZN(n8779) );
  CLKBUF_X2 U7305 ( .A(n7999), .Z(n6563) );
  INV_X1 U7306 ( .A(n6566), .ZN(n8177) );
  NAND2_X1 U7307 ( .A1(n8308), .A2(n8299), .ZN(n8311) );
  BUF_X2 U7308 ( .A(n9903), .Z(n6551) );
  INV_X2 U7310 ( .A(n6906), .ZN(n9903) );
  AND2_X1 U7311 ( .A1(n7376), .A2(n7620), .ZN(n7598) );
  INV_X1 U7312 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7642) );
  INV_X1 U7313 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7679) );
  INV_X1 U7314 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7715) );
  NAND3_X1 U7315 ( .A1(n6914), .A2(n6909), .A3(n6912), .ZN(P1_U3262) );
  OR2_X2 U7316 ( .A1(n6542), .A2(n6754), .ZN(n6723) );
  AOI21_X1 U7317 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n6542) );
  NAND2_X1 U7318 ( .A1(n8769), .A2(n8770), .ZN(n8768) );
  NAND2_X1 U7319 ( .A1(n8762), .A2(n8763), .ZN(n8770) );
  INV_X1 U7320 ( .A(n6543), .ZN(n6650) );
  NOR2_X1 U7321 ( .A1(n8950), .A2(n8945), .ZN(n6543) );
  NAND3_X1 U7322 ( .A1(n8799), .A2(n8798), .A3(n6623), .ZN(n6722) );
  INV_X2 U7323 ( .A(n11752), .ZN(n11004) );
  OAI21_X1 U7324 ( .B1(n13039), .B2(n12806), .A(n12788), .ZN(n12775) );
  AND3_X1 U7325 ( .A1(n7619), .A2(n7617), .A3(n7618), .ZN(n7376) );
  OR2_X1 U7326 ( .A1(n13554), .A2(n7406), .ZN(n7403) );
  OAI21_X1 U7327 ( .B1(n12727), .B2(n12014), .A(n10611), .ZN(n10612) );
  NAND3_X1 U7328 ( .A1(n11270), .A2(n11572), .A3(n6576), .ZN(n13565) );
  NAND2_X1 U7329 ( .A1(n7688), .A2(n7687), .ZN(n10273) );
  AND2_X1 U7330 ( .A1(n7598), .A2(n7536), .ZN(n7375) );
  INV_X1 U7331 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7766) );
  INV_X1 U7332 ( .A(n11448), .ZN(n10522) );
  NAND2_X2 U7333 ( .A1(n8713), .A2(n11925), .ZN(n10282) );
  AND2_X2 U7334 ( .A1(n10613), .A2(n10612), .ZN(n12421) );
  INV_X1 U7335 ( .A(n10376), .ZN(n14941) );
  NAND2_X1 U7336 ( .A1(n9141), .A2(n9140), .ZN(n12718) );
  OAI21_X1 U7337 ( .B1(n9446), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U7338 ( .A1(n10438), .A2(n9720), .ZN(n10569) );
  CLKBUF_X2 U7339 ( .A(n13564), .Z(n9813) );
  INV_X1 U7340 ( .A(n12364), .ZN(n12343) );
  INV_X1 U7341 ( .A(n13954), .ZN(n11456) );
  AOI21_X1 U7342 ( .B1(n11214), .B2(n7346), .A(n7345), .ZN(n7344) );
  NOR2_X1 U7343 ( .A1(n11923), .A2(n11922), .ZN(n11969) );
  OAI21_X1 U7345 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n13978), .A(n13965), .ZN(
        n14678) );
  OR2_X1 U7346 ( .A1(n14547), .A2(n14546), .ZN(n7268) );
  XNOR2_X1 U7347 ( .A(n12517), .B(n12516), .ZN(n12518) );
  XNOR2_X1 U7348 ( .A(n9168), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9169) );
  XNOR2_X1 U7349 ( .A(n9219), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U7350 ( .A1(n7826), .A2(n7825), .ZN(n11277) );
  NAND2_X1 U7351 ( .A1(n7813), .A2(n7812), .ZN(n11250) );
  INV_X1 U7352 ( .A(n8979), .ZN(n8970) );
  NAND2_X1 U7353 ( .A1(n8116), .A2(n8115), .ZN(n13696) );
  NAND2_X1 U7354 ( .A1(n7923), .A2(n7922), .ZN(n13715) );
  INV_X2 U7355 ( .A(n6568), .ZN(n9902) );
  INV_X1 U7356 ( .A(n11783), .ZN(n14774) );
  AND3_X1 U7357 ( .A1(n11932), .A2(n11931), .A3(n11930), .ZN(n11976) );
  AND4_X1 U7358 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n11787)
         );
  OAI21_X1 U7359 ( .B1(n10246), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10243), .ZN(
        n10419) );
  OAI21_X1 U7360 ( .B1(n10582), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10581), .ZN(
        n10583) );
  BUF_X1 U7361 ( .A(n10728), .Z(n6552) );
  XNOR2_X1 U7362 ( .A(n8969), .B(n8968), .ZN(n13721) );
  NAND4_X1 U7363 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n9585)
         );
  AOI21_X1 U7364 ( .B1(n9632), .B2(n15039), .A(n9631), .ZN(n12386) );
  AND2_X1 U7366 ( .A1(n8981), .A2(n8980), .ZN(n13684) );
  NAND2_X1 U7367 ( .A1(n8650), .A2(n8651), .ZN(n11925) );
  INV_X1 U7369 ( .A(n9940), .ZN(n7999) );
  INV_X2 U7370 ( .A(n7808), .ZN(n7702) );
  AND2_X2 U7371 ( .A1(n10375), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10793) );
  AND2_X2 U7372 ( .A1(n6917), .A2(n6920), .ZN(n10201) );
  INV_X2 U7373 ( .A(n13292), .ZN(n9002) );
  AOI21_X2 U7374 ( .B1(n9707), .B2(n9706), .A(n6665), .ZN(n10259) );
  NAND2_X2 U7375 ( .A1(n9140), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9138) );
  NOR2_X2 U7376 ( .A1(n8311), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n8300) );
  NOR3_X2 U7377 ( .A1(n12179), .A2(n12178), .A3(n12177), .ZN(n12181) );
  INV_X1 U7379 ( .A(n8578), .ZN(n6545) );
  AOI21_X2 U7380 ( .B1(n12823), .B2(n12822), .A(n9520), .ZN(n12809) );
  OAI21_X2 U7381 ( .B1(n12836), .B2(n12114), .A(n12112), .ZN(n12823) );
  OAI21_X2 U7382 ( .B1(n12538), .B2(n12397), .A(n12399), .ZN(n12438) );
  NAND2_X2 U7383 ( .A1(n13722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7623) );
  OAI21_X2 U7384 ( .B1(n10569), .B2(n10570), .A(n9725), .ZN(n10650) );
  NAND2_X2 U7385 ( .A1(n13082), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9166) );
  OR2_X1 U7386 ( .A1(n13008), .A2(n15099), .ZN(n12021) );
  NAND2_X2 U7387 ( .A1(n6723), .A2(n7543), .ZN(n8867) );
  AOI21_X2 U7388 ( .B1(n10127), .B2(n14443), .A(n15477), .ZN(n15471) );
  AOI21_X1 U7389 ( .B1(n14034), .B2(n14033), .A(n14032), .ZN(n14251) );
  INV_X1 U7391 ( .A(n10376), .ZN(n6550) );
  NOR3_X2 U7392 ( .A1(n12124), .A2(n12123), .A3(n12789), .ZN(n12131) );
  NAND2_X2 U7393 ( .A1(n7448), .A2(n7446), .ZN(n6906) );
  OAI21_X2 U7394 ( .B1(n9272), .B2(n9090), .A(n9091), .ZN(n9286) );
  NAND2_X2 U7395 ( .A1(n9088), .A2(n9087), .ZN(n9272) );
  NOR2_X2 U7396 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10356) );
  AOI21_X2 U7397 ( .B1(n14725), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14716), .ZN(
        n14735) );
  NOR2_X2 U7398 ( .A1(n14955), .A2(n6713), .ZN(n10816) );
  NOR2_X4 U7399 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n14952), .ZN(n14436) );
  INV_X2 U7400 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14952) );
  INV_X1 U7401 ( .A(n13684), .ZN(n13311) );
  AOI22_X2 U7402 ( .A1(n13721), .A2(n7702), .B1(n8970), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n13680) );
  NAND2_X1 U7403 ( .A1(n6703), .A2(n6702), .ZN(n12471) );
  NAND2_X1 U7404 ( .A1(n8617), .A2(n8616), .ZN(n14248) );
  OR2_X1 U7405 ( .A1(n11227), .A2(n11228), .ZN(n6849) );
  NAND2_X1 U7406 ( .A1(n10787), .A2(n10786), .ZN(n11147) );
  NAND2_X1 U7407 ( .A1(n10921), .A2(n10922), .ZN(n10920) );
  XNOR2_X1 U7408 ( .A(n11212), .B(n11213), .ZN(n11227) );
  NAND2_X1 U7409 ( .A1(n7333), .A2(n6635), .ZN(n11212) );
  INV_X1 U7410 ( .A(n11782), .ZN(n13956) );
  OR2_X1 U7411 ( .A1(n13009), .A2(n14934), .ZN(n13014) );
  INV_X4 U7412 ( .A(n11921), .ZN(n11911) );
  INV_X1 U7413 ( .A(n13233), .ZN(n7221) );
  CLKBUF_X2 U7414 ( .A(P2_U3947), .Z(n6554) );
  INV_X2 U7415 ( .A(n9184), .ZN(n9369) );
  INV_X4 U7416 ( .A(n12345), .ZN(n10521) );
  INV_X2 U7418 ( .A(n6589), .ZN(n12362) );
  NAND2_X4 U7419 ( .A1(n10281), .A2(n11448), .ZN(n12345) );
  INV_X2 U7420 ( .A(n9184), .ZN(n6553) );
  CLKBUF_X2 U7421 ( .A(n9571), .Z(n6559) );
  INV_X4 U7422 ( .A(n6557), .ZN(n9555) );
  BUF_X1 U7423 ( .A(n11009), .Z(n6562) );
  NAND2_X1 U7424 ( .A1(n9170), .A2(n13090), .ZN(n9275) );
  NAND2_X1 U7426 ( .A1(n6824), .A2(n14444), .ZN(n14448) );
  AND2_X1 U7427 ( .A1(n8754), .A2(n9002), .ZN(n11114) );
  BUF_X1 U7428 ( .A(n8238), .Z(n6564) );
  XNOR2_X1 U7429 ( .A(n8189), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8238) );
  XNOR2_X1 U7430 ( .A(n8316), .B(n8317), .ZN(n10499) );
  INV_X8 U7431 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9415) );
  INV_X1 U7432 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7610) );
  INV_X2 U7433 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14371) );
  AOI21_X1 U7434 ( .B1(n7520), .B2(n7519), .A(n7515), .ZN(n12193) );
  OR2_X1 U7435 ( .A1(n12186), .A2(n15123), .ZN(n7518) );
  AOI21_X1 U7436 ( .B1(n7324), .B2(n7326), .A(n6727), .ZN(n12186) );
  OR2_X1 U7437 ( .A1(n13027), .A2(n15179), .ZN(n6970) );
  NAND2_X1 U7438 ( .A1(n13128), .A2(n13127), .ZN(n9812) );
  NAND2_X1 U7439 ( .A1(n6786), .A2(n12768), .ZN(n12947) );
  AND2_X1 U7440 ( .A1(n14236), .A2(n14238), .ZN(n14337) );
  OAI21_X1 U7441 ( .B1(n12158), .B2(n12157), .A(n12156), .ZN(n7521) );
  NAND2_X1 U7442 ( .A1(n7414), .A2(n7412), .ZN(n13128) );
  NOR2_X1 U7443 ( .A1(n8927), .A2(n8926), .ZN(n8928) );
  OR2_X1 U7444 ( .A1(n12769), .A2(n15110), .ZN(n6786) );
  AND2_X1 U7445 ( .A1(n15162), .A2(n12944), .ZN(n6971) );
  AND2_X1 U7446 ( .A1(n7563), .A2(n7564), .ZN(n6805) );
  OAI21_X1 U7447 ( .B1(n7017), .B2(n7015), .A(n7028), .ZN(n7014) );
  OAI21_X1 U7448 ( .B1(n9802), .B2(n7417), .A(n9806), .ZN(n7413) );
  NAND2_X1 U7449 ( .A1(n8661), .A2(n14522), .ZN(n7563) );
  AND2_X1 U7450 ( .A1(n7022), .A2(n7024), .ZN(n7015) );
  NAND2_X1 U7451 ( .A1(n9621), .A2(n6958), .ZN(n6961) );
  OR2_X1 U7452 ( .A1(n12782), .A2(n15110), .ZN(n6751) );
  NAND2_X1 U7453 ( .A1(n12775), .A2(n6735), .ZN(n9621) );
  NAND2_X1 U7454 ( .A1(n6894), .A2(n6891), .ZN(n13325) );
  AND2_X1 U7455 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  NOR2_X1 U7456 ( .A1(n7030), .A2(n11901), .ZN(n7027) );
  NAND2_X1 U7457 ( .A1(n12471), .A2(n12420), .ZN(n12424) );
  NOR2_X1 U7458 ( .A1(n6807), .A2(n6806), .ZN(n13339) );
  MUX2_X1 U7459 ( .A(n12371), .B(n8747), .S(n11911), .Z(n11914) );
  NAND2_X1 U7460 ( .A1(n11901), .A2(n7030), .ZN(n7026) );
  AND2_X1 U7461 ( .A1(n6893), .A2(n6892), .ZN(n6891) );
  AOI21_X2 U7462 ( .B1(n13721), .B2(n8371), .A(n11919), .ZN(n14340) );
  INV_X1 U7463 ( .A(n8664), .ZN(n6879) );
  NAND2_X1 U7464 ( .A1(n8710), .A2(n8709), .ZN(n14010) );
  XNOR2_X1 U7465 ( .A(n8978), .B(n8977), .ZN(n12213) );
  OR2_X1 U7466 ( .A1(n7264), .A2(n7262), .ZN(n6893) );
  NAND2_X1 U7467 ( .A1(n13759), .A2(n13756), .ZN(n12324) );
  NOR2_X1 U7468 ( .A1(n9562), .A2(n12141), .ZN(n12763) );
  NAND2_X1 U7469 ( .A1(n7500), .A2(n12125), .ZN(n12778) );
  AOI21_X1 U7470 ( .B1(n7361), .B2(n7363), .A(n7360), .ZN(n7359) );
  AND2_X1 U7471 ( .A1(n14070), .A2(n8595), .ZN(n7601) );
  NAND2_X1 U7472 ( .A1(n6907), .A2(n8160), .ZN(n13598) );
  XNOR2_X1 U7473 ( .A(n14551), .B(n14550), .ZN(n14549) );
  OAI21_X1 U7474 ( .B1(n13400), .B2(n7224), .A(n7222), .ZN(n8232) );
  NAND2_X1 U7475 ( .A1(n7364), .A2(n6637), .ZN(n13790) );
  NAND2_X1 U7476 ( .A1(n12129), .A2(n9539), .ZN(n12789) );
  NAND2_X1 U7477 ( .A1(n8159), .A2(n8158), .ZN(n8175) );
  CLKBUF_X1 U7478 ( .A(n12565), .Z(n6797) );
  NAND2_X1 U7479 ( .A1(n9543), .A2(n9542), .ZN(n12579) );
  NAND2_X1 U7480 ( .A1(n12843), .A2(n12104), .ZN(n9615) );
  NAND2_X1 U7481 ( .A1(n8690), .A2(n8689), .ZN(n14202) );
  NAND2_X1 U7482 ( .A1(n13419), .A2(n8227), .ZN(n13402) );
  OR2_X1 U7483 ( .A1(n13453), .A2(n7396), .ZN(n7393) );
  NAND2_X1 U7484 ( .A1(n8130), .A2(n8129), .ZN(n13361) );
  NAND2_X1 U7485 ( .A1(n12857), .A2(n9614), .ZN(n12843) );
  OR2_X1 U7486 ( .A1(n13417), .A2(n13416), .ZN(n13419) );
  NAND2_X1 U7487 ( .A1(n6823), .A2(n6822), .ZN(n7271) );
  NAND2_X1 U7488 ( .A1(n8597), .A2(n8596), .ZN(n14259) );
  AOI21_X1 U7489 ( .B1(n14108), .B2(n8572), .A(n7155), .ZN(n7154) );
  NAND2_X1 U7490 ( .A1(n13899), .A2(n13900), .ZN(n13898) );
  NAND2_X1 U7491 ( .A1(n8687), .A2(n6582), .ZN(n14332) );
  NAND2_X1 U7492 ( .A1(n12859), .A2(n12858), .ZN(n12857) );
  NAND2_X1 U7493 ( .A1(n11646), .A2(n7193), .ZN(n8687) );
  NAND2_X1 U7494 ( .A1(n12882), .A2(n6992), .ZN(n12874) );
  AND2_X1 U7495 ( .A1(n6922), .A2(n6921), .ZN(n14730) );
  NAND2_X1 U7496 ( .A1(n8096), .A2(n8095), .ZN(n13620) );
  OR2_X1 U7497 ( .A1(n14720), .A2(n6700), .ZN(n6922) );
  NAND2_X1 U7498 ( .A1(n9489), .A2(n9488), .ZN(n12848) );
  NAND2_X1 U7499 ( .A1(n8058), .A2(n8057), .ZN(n13705) );
  XNOR2_X1 U7500 ( .A(n8071), .B(n8070), .ZN(n11636) );
  NAND2_X1 U7501 ( .A1(n11524), .A2(n11947), .ZN(n11523) );
  XNOR2_X1 U7502 ( .A(n8110), .B(SI_24_), .ZN(n8107) );
  AOI21_X1 U7503 ( .B1(n8069), .B2(n8087), .A(n8068), .ZN(n8071) );
  NOR2_X2 U7504 ( .A1(n13472), .A2(n13642), .ZN(n13460) );
  AOI21_X1 U7505 ( .B1(n14597), .B2(n6619), .A(n7525), .ZN(n12916) );
  NAND2_X1 U7506 ( .A1(n7602), .A2(n9339), .ZN(n14597) );
  NAND2_X1 U7507 ( .A1(n8094), .A2(n8093), .ZN(n8110) );
  AND2_X1 U7508 ( .A1(n14478), .A2(n14477), .ZN(n14659) );
  NAND2_X1 U7509 ( .A1(n8540), .A2(n8539), .ZN(n14298) );
  CLKBUF_X1 U7510 ( .A(n14599), .Z(n6746) );
  NAND2_X1 U7511 ( .A1(n8001), .A2(n8000), .ZN(n13647) );
  NAND2_X1 U7512 ( .A1(n7141), .A2(n7140), .ZN(n7139) );
  NAND2_X1 U7513 ( .A1(n9118), .A2(n9117), .ZN(n9471) );
  AOI21_X1 U7514 ( .B1(n7006), .B2(n7005), .A(n7004), .ZN(n12621) );
  NAND2_X1 U7515 ( .A1(n6817), .A2(n6602), .ZN(n7006) );
  NAND2_X1 U7516 ( .A1(n8529), .A2(n8528), .ZN(n14304) );
  NAND2_X1 U7517 ( .A1(n6793), .A2(n6792), .ZN(n6820) );
  NAND2_X1 U7518 ( .A1(n7963), .A2(n7962), .ZN(n13656) );
  NAND2_X1 U7519 ( .A1(n7285), .A2(n7286), .ZN(n9116) );
  OR2_X1 U7520 ( .A1(n11397), .A2(n9325), .ZN(n6817) );
  OR2_X1 U7521 ( .A1(n8037), .A2(n10504), .ZN(n8038) );
  XNOR2_X1 U7522 ( .A(n8037), .B(n10504), .ZN(n8036) );
  CLKBUF_X1 U7523 ( .A(n9443), .Z(n6774) );
  NAND2_X1 U7524 ( .A1(n8023), .A2(n8022), .ZN(n8037) );
  NAND2_X1 U7525 ( .A1(n8498), .A2(n8497), .ZN(n14320) );
  OR2_X1 U7526 ( .A1(n7910), .A2(n7909), .ZN(n7485) );
  NAND2_X1 U7527 ( .A1(n7911), .A2(n7895), .ZN(n7910) );
  NAND2_X1 U7528 ( .A1(n7844), .A2(n7843), .ZN(n11479) );
  NAND2_X1 U7529 ( .A1(n9103), .A2(n9102), .ZN(n9357) );
  NAND2_X1 U7530 ( .A1(n8404), .A2(n8403), .ZN(n11806) );
  NAND2_X1 U7531 ( .A1(n7792), .A2(n7791), .ZN(n10913) );
  AND2_X1 U7532 ( .A1(n6929), .A2(n6928), .ZN(n10317) );
  INV_X2 U7533 ( .A(n15129), .ZN(n15038) );
  AND2_X1 U7534 ( .A1(n10689), .A2(n10615), .ZN(n10620) );
  NAND2_X1 U7535 ( .A1(n12042), .A2(n12041), .ZN(n15056) );
  AND2_X1 U7536 ( .A1(n12039), .A2(n12036), .ZN(n15076) );
  CLKBUF_X1 U7537 ( .A(n9331), .Z(n6773) );
  OR2_X1 U7538 ( .A1(n12609), .A2(n15078), .ZN(n12039) );
  INV_X2 U7539 ( .A(n14529), .ZN(n14224) );
  AND2_X2 U7540 ( .A1(n10981), .A2(n13573), .ZN(n13552) );
  NAND2_X1 U7541 ( .A1(n7458), .A2(n7456), .ZN(n7788) );
  INV_X2 U7542 ( .A(n12421), .ZN(n12462) );
  NAND2_X1 U7543 ( .A1(n12199), .A2(n14526), .ZN(n14529) );
  NAND4_X2 U7544 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(n15045)
         );
  NAND4_X1 U7545 ( .A1(n9188), .A2(n9186), .A3(n9187), .A4(n9185), .ZN(n13009)
         );
  NAND2_X1 U7546 ( .A1(n8332), .A2(n6745), .ZN(n13961) );
  OAI211_X1 U7547 ( .C1(n9853), .C2(n10204), .A(n8345), .B(n8344), .ZN(n10685)
         );
  NAND2_X2 U7548 ( .A1(n7061), .A2(n7060), .ZN(n11921) );
  NAND4_X1 U7549 ( .A1(n7678), .A2(n7677), .A3(n7676), .A4(n7675), .ZN(n13233)
         );
  BUF_X2 U7550 ( .A(n8760), .Z(n7655) );
  INV_X1 U7551 ( .A(n9275), .ZN(n9184) );
  AND2_X1 U7552 ( .A1(n8302), .A2(n14383), .ZN(n8347) );
  CLKBUF_X2 U7553 ( .A(n9203), .Z(n6557) );
  AND2_X1 U7554 ( .A1(n14380), .A2(n14383), .ZN(n8349) );
  INV_X1 U7555 ( .A(n11009), .ZN(n6561) );
  OAI211_X1 U7556 ( .C1(n10519), .C2(n9179), .A(n9211), .B(n9210), .ZN(n11098)
         );
  OAI211_X1 U7557 ( .C1(n10548), .C2(n9179), .A(n9202), .B(n9201), .ZN(n15099)
         );
  XNOR2_X1 U7558 ( .A(n14447), .B(n14448), .ZN(n15473) );
  AOI21_X1 U7559 ( .B1(n6899), .B2(n6901), .A(n6897), .ZN(n6896) );
  INV_X1 U7560 ( .A(n10286), .ZN(n10297) );
  OAI211_X1 U7561 ( .C1(n9853), .C2(n6548), .A(n8319), .B(n8318), .ZN(n10728)
         );
  CLKBUF_X3 U7562 ( .A(n8240), .Z(n6566) );
  INV_X1 U7563 ( .A(n7721), .ZN(n7691) );
  AND2_X2 U7564 ( .A1(n12215), .A2(n7627), .ZN(n7721) );
  AND2_X1 U7565 ( .A1(n8733), .A2(n8732), .ZN(n10286) );
  NAND2_X2 U7566 ( .A1(n9179), .A2(n6568), .ZN(n12005) );
  AND2_X1 U7567 ( .A1(n8301), .A2(n14373), .ZN(n8303) );
  AND2_X1 U7568 ( .A1(n6900), .A2(n7486), .ZN(n6899) );
  NAND2_X2 U7569 ( .A1(n13386), .A2(n9694), .ZN(n9807) );
  CLKBUF_X1 U7570 ( .A(n13386), .Z(n6794) );
  NAND2_X1 U7571 ( .A1(n8648), .A2(n7606), .ZN(n8665) );
  INV_X1 U7572 ( .A(n9169), .ZN(n13090) );
  AOI21_X1 U7573 ( .B1(n7460), .B2(n7462), .A(n7457), .ZN(n7456) );
  NAND2_X2 U7574 ( .A1(n11114), .A2(n11732), .ZN(n8994) );
  MUX2_X1 U7575 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8647), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8648) );
  AOI21_X1 U7576 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n10203), .A(n10495), .ZN(
        n10402) );
  AND2_X2 U7577 ( .A1(n8238), .A2(n11322), .ZN(n8754) );
  INV_X1 U7578 ( .A(n7627), .ZN(n7629) );
  MUX2_X1 U7579 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9139), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n9141) );
  CLKBUF_X1 U7580 ( .A(n11322), .Z(n6771) );
  AND2_X1 U7581 ( .A1(n6741), .A2(n6740), .ZN(n15479) );
  MUX2_X1 U7582 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8309), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8310) );
  NOR2_X1 U7583 ( .A1(n7838), .A2(n7489), .ZN(n7488) );
  NAND2_X1 U7584 ( .A1(n7371), .A2(n7368), .ZN(n8651) );
  NAND2_X1 U7585 ( .A1(n7057), .A2(n7059), .ZN(n8720) );
  XNOR2_X1 U7586 ( .A(n8191), .B(n8188), .ZN(n11322) );
  OR2_X1 U7587 ( .A1(n8248), .A2(n7636), .ZN(n8194) );
  NAND2_X1 U7588 ( .A1(n10537), .A2(n10536), .ZN(n10535) );
  NAND2_X1 U7589 ( .A1(n8190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U7590 ( .A1(n10560), .A2(n6591), .ZN(n10536) );
  AND2_X2 U7591 ( .A1(n9135), .A2(n9134), .ZN(n9640) );
  NAND2_X2 U7592 ( .A1(n9902), .A2(P2_U3088), .ZN(n13736) );
  NOR2_X1 U7593 ( .A1(n8192), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U7594 ( .A1(n8192), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U7595 ( .A1(n7803), .A2(SI_9_), .ZN(n7820) );
  OAI21_X1 U7596 ( .B1(n14441), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6641), .ZN(
        n7277) );
  AND2_X1 U7597 ( .A1(n8414), .A2(n8297), .ZN(n6834) );
  NAND2_X1 U7599 ( .A1(n7559), .A2(n8284), .ZN(n8354) );
  NOR2_X1 U7600 ( .A1(n7508), .A2(n9054), .ZN(n7511) );
  NAND2_X1 U7601 ( .A1(n9181), .A2(n9180), .ZN(n10568) );
  NOR2_X1 U7602 ( .A1(n8719), .A2(n8296), .ZN(n8297) );
  NAND2_X1 U7603 ( .A1(n7514), .A2(n6640), .ZN(n7508) );
  AND2_X1 U7604 ( .A1(n8293), .A2(n6676), .ZN(n7589) );
  AND2_X1 U7605 ( .A1(n9051), .A2(n9052), .ZN(n9062) );
  AND4_X1 U7606 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n8293)
         );
  NAND3_X1 U7607 ( .A1(n7766), .A2(n7809), .A3(n7610), .ZN(n7938) );
  AND2_X1 U7608 ( .A1(n7915), .A2(n7615), .ZN(n7616) );
  INV_X1 U7609 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9039) );
  INV_X1 U7610 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n15206) );
  INV_X1 U7611 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9254) );
  INV_X4 U7612 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7613 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n9041) );
  NOR2_X1 U7614 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7915) );
  INV_X4 U7615 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7616 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9043) );
  INV_X1 U7617 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9056) );
  INV_X1 U7618 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8316) );
  INV_X1 U7619 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6990) );
  INV_X1 U7620 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8368) );
  INV_X1 U7621 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8656) );
  INV_X1 U7622 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8653) );
  NOR2_X1 U7623 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8654) );
  NOR2_X1 U7624 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9051) );
  NOR2_X1 U7625 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n9052) );
  NOR2_X1 U7626 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8290) );
  AND2_X1 U7627 ( .A1(n7598), .A2(n7537), .ZN(n7534) );
  XNOR2_X1 U7628 ( .A(n8175), .B(n8174), .ZN(n13728) );
  AND2_X1 U7629 ( .A1(n10785), .A2(n10784), .ZN(n10787) );
  OR2_X1 U7630 ( .A1(n8300), .A2(n14371), .ZN(n7560) );
  INV_X2 U7631 ( .A(n8662), .ZN(n11023) );
  OAI22_X1 U7632 ( .A1(n8979), .A2(n9910), .B1(n9940), .B2(n9962), .ZN(n7373)
         );
  OAI21_X2 U7634 ( .B1(n13158), .B2(n7425), .A(n7423), .ZN(n9796) );
  INV_X1 U7635 ( .A(n12380), .ZN(n9170) );
  XNOR2_X1 U7636 ( .A(n9050), .B(n9049), .ZN(n12727) );
  NOR2_X1 U7637 ( .A1(n14572), .A2(n14573), .ZN(n14571) );
  INV_X4 U7638 ( .A(n7950), .ZN(n8182) );
  XNOR2_X1 U7639 ( .A(n7708), .B(n7710), .ZN(n9894) );
  CLKBUF_X1 U7640 ( .A(n9203), .Z(n6556) );
  NAND2_X1 U7641 ( .A1(n12380), .A2(n9169), .ZN(n9203) );
  AOI21_X2 U7642 ( .B1(n10421), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10418), .ZN(
        n10432) );
  INV_X1 U7643 ( .A(n11984), .ZN(n9571) );
  OAI211_X2 U7644 ( .C1(n10535), .C2(n10519), .A(n7133), .B(n7130), .ZN(n10601) );
  NAND2_X1 U7645 ( .A1(n13386), .A2(n9694), .ZN(n6560) );
  OAI21_X1 U7646 ( .B1(n9916), .B2(n7808), .A(n6941), .ZN(n11009) );
  AOI21_X2 U7647 ( .B1(n10406), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10400), .ZN(
        n10483) );
  NOR2_X2 U7648 ( .A1(n14735), .A2(n14736), .ZN(n14734) );
  CLKBUF_X3 U7649 ( .A(n8822), .Z(n6565) );
  BUF_X4 U7650 ( .A(n8822), .Z(n8946) );
  INV_X4 U7651 ( .A(n8822), .ZN(n8943) );
  AOI21_X2 U7652 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13984), .A(n14734), .ZN(
        n13985) );
  AND2_X1 U7654 ( .A1(n13545), .A2(n7409), .ZN(n7408) );
  NAND2_X1 U7655 ( .A1(n7908), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U7656 ( .A1(n7001), .A2(n7000), .ZN(n6999) );
  INV_X1 U7657 ( .A(n10872), .ZN(n7000) );
  NOR2_X1 U7658 ( .A1(n12763), .A2(n6959), .ZN(n6958) );
  INV_X1 U7659 ( .A(n6962), .ZN(n6959) );
  OR2_X1 U7660 ( .A1(n12986), .A2(n12900), .ZN(n12089) );
  AOI21_X1 U7661 ( .B1(n6978), .B2(n6980), .A(n6976), .ZN(n6975) );
  OR2_X1 U7662 ( .A1(n12605), .A2(n14610), .ZN(n12064) );
  AND2_X1 U7663 ( .A1(n12064), .A2(n12063), .ZN(n11593) );
  AND2_X1 U7664 ( .A1(n13447), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U7665 ( .A1(n8033), .A2(n7400), .ZN(n7399) );
  INV_X1 U7666 ( .A(n6841), .ZN(n6840) );
  NAND2_X1 U7667 ( .A1(n11304), .A2(n7152), .ZN(n11530) );
  NOR2_X1 U7668 ( .A1(n11947), .A2(n7153), .ZN(n7152) );
  INV_X1 U7669 ( .A(n8431), .ZN(n7153) );
  NAND2_X1 U7670 ( .A1(n6834), .A2(n6832), .ZN(n6833) );
  AND2_X1 U7671 ( .A1(n7589), .A2(n8313), .ZN(n6832) );
  AND3_X1 U7672 ( .A1(n9338), .A2(n9337), .A3(n9336), .ZN(n12391) );
  AND2_X1 U7673 ( .A1(n12495), .A2(n7098), .ZN(n7097) );
  NAND2_X1 U7674 ( .A1(n12428), .A2(n7104), .ZN(n7098) );
  AND2_X1 U7675 ( .A1(n12619), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7004) );
  INV_X1 U7676 ( .A(n12617), .ZN(n7005) );
  INV_X1 U7677 ( .A(n12657), .ZN(n7002) );
  INV_X1 U7678 ( .A(n7408), .ZN(n7406) );
  OAI21_X1 U7679 ( .B1(n13140), .B2(n6565), .A(n8882), .ZN(n8883) );
  AND2_X1 U7680 ( .A1(n7466), .A2(n11882), .ZN(n7464) );
  NAND2_X1 U7681 ( .A1(n7470), .A2(n7468), .ZN(n7467) );
  AOI21_X1 U7682 ( .B1(n7475), .B2(n7479), .A(n6660), .ZN(n7474) );
  INV_X1 U7683 ( .A(n7837), .ZN(n7840) );
  NOR2_X1 U7684 ( .A1(n7487), .A2(n6903), .ZN(n6902) );
  INV_X1 U7685 ( .A(n7801), .ZN(n6903) );
  INV_X1 U7686 ( .A(n7488), .ZN(n7487) );
  NAND2_X1 U7687 ( .A1(n13032), .A2(n12752), .ZN(n6960) );
  NOR2_X1 U7688 ( .A1(n9561), .A2(n12752), .ZN(n12141) );
  OR2_X1 U7689 ( .A1(n12837), .A2(n12845), .ZN(n12112) );
  OR2_X1 U7690 ( .A1(n13062), .A2(n12884), .ZN(n12095) );
  AOI21_X1 U7691 ( .B1(n7288), .B2(n7290), .A(n7287), .ZN(n7286) );
  INV_X1 U7692 ( .A(n9115), .ZN(n7287) );
  AOI21_X1 U7693 ( .B1(n7300), .B2(n7302), .A(n7299), .ZN(n7298) );
  INV_X1 U7694 ( .A(n9100), .ZN(n7299) );
  XNOR2_X1 U7695 ( .A(n6560), .B(n6561), .ZN(n9697) );
  AND2_X1 U7696 ( .A1(n11657), .A2(n9760), .ZN(n7442) );
  AND2_X1 U7697 ( .A1(n11333), .A2(n9745), .ZN(n7437) );
  NAND2_X1 U7698 ( .A1(n7387), .A2(n6592), .ZN(n7386) );
  INV_X1 U7699 ( .A(n7389), .ZN(n7387) );
  INV_X1 U7700 ( .A(n7267), .ZN(n7266) );
  XNOR2_X1 U7701 ( .A(n7221), .B(n10273), .ZN(n7220) );
  INV_X1 U7702 ( .A(n13232), .ZN(n10276) );
  INV_X1 U7703 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7638) );
  NAND4_X1 U7704 ( .A1(n7614), .A2(n7613), .A3(n7612), .A4(n7611), .ZN(n7916)
         );
  INV_X1 U7705 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7614) );
  INV_X1 U7706 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7613) );
  INV_X1 U7707 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7611) );
  INV_X1 U7708 ( .A(n6839), .ZN(n6838) );
  OAI21_X1 U7709 ( .B1(n6844), .B2(n6840), .A(n13824), .ZN(n6839) );
  INV_X1 U7710 ( .A(n7174), .ZN(n7173) );
  OAI21_X1 U7711 ( .B1(n14058), .B2(n7175), .A(n8615), .ZN(n7174) );
  AOI21_X1 U7712 ( .B1(n7166), .B2(n7164), .A(n7163), .ZN(n7162) );
  INV_X1 U7713 ( .A(n11865), .ZN(n7163) );
  INV_X1 U7714 ( .A(n14182), .ZN(n7164) );
  OAI21_X1 U7715 ( .B1(n11944), .B2(n7180), .A(n11942), .ZN(n7179) );
  NAND2_X1 U7716 ( .A1(n8662), .A2(n12212), .ZN(n11764) );
  AOI21_X1 U7717 ( .B1(n7593), .B2(n14100), .A(n6648), .ZN(n7591) );
  AND2_X1 U7718 ( .A1(n8293), .A2(n8514), .ZN(n7059) );
  AND2_X1 U7719 ( .A1(n7971), .A2(n7959), .ZN(n7969) );
  XNOR2_X1 U7720 ( .A(n7277), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14431) );
  NOR2_X1 U7721 ( .A1(n14408), .A2(n14407), .ZN(n14430) );
  NOR2_X1 U7722 ( .A1(n14456), .A2(n14457), .ZN(n14407) );
  OAI22_X1 U7723 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n14472), .B1(n14473), 
        .B2(n14417), .ZN(n14476) );
  AND2_X1 U7724 ( .A1(n6677), .A2(n7092), .ZN(n7091) );
  NAND2_X1 U7725 ( .A1(n7095), .A2(n7093), .ZN(n7092) );
  NAND2_X1 U7726 ( .A1(n12431), .A2(n12765), .ZN(n7101) );
  NAND2_X1 U7727 ( .A1(n12430), .A2(n12806), .ZN(n7102) );
  NOR2_X1 U7728 ( .A1(n6609), .A2(n6577), .ZN(n7104) );
  INV_X1 U7729 ( .A(n9478), .ZN(n9570) );
  NAND2_X1 U7730 ( .A1(n7114), .A2(n6593), .ZN(n7113) );
  NOR2_X1 U7731 ( .A1(n10819), .A2(n15307), .ZN(n10869) );
  INV_X1 U7732 ( .A(n11396), .ZN(n10871) );
  NAND2_X1 U7733 ( .A1(n7137), .A2(n7136), .ZN(n7135) );
  INV_X1 U7734 ( .A(n10856), .ZN(n7136) );
  INV_X1 U7735 ( .A(n6790), .ZN(n11543) );
  NAND2_X1 U7736 ( .A1(n7135), .A2(n7134), .ZN(n6775) );
  NAND2_X1 U7737 ( .A1(n11396), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7134) );
  XNOR2_X1 U7738 ( .A(n7139), .B(n15006), .ZN(n15014) );
  NOR2_X1 U7739 ( .A1(n15014), .A2(n9365), .ZN(n15013) );
  INV_X1 U7740 ( .A(n12710), .ZN(n7125) );
  INV_X1 U7741 ( .A(n12777), .ZN(n12752) );
  NAND2_X1 U7742 ( .A1(n7492), .A2(n7491), .ZN(n12753) );
  AOI21_X1 U7743 ( .B1(n6572), .B2(n7495), .A(n9562), .ZN(n7491) );
  AOI21_X1 U7744 ( .B1(n7498), .B2(n12126), .A(n7497), .ZN(n7496) );
  NOR2_X1 U7745 ( .A1(n12822), .A2(n6965), .ZN(n6963) );
  NOR2_X1 U7746 ( .A1(n6571), .A2(n7523), .ZN(n7522) );
  INV_X1 U7747 ( .A(n12087), .ZN(n7523) );
  INV_X1 U7748 ( .A(n12602), .ZN(n12912) );
  NOR2_X1 U7749 ( .A1(n9603), .A2(n6985), .ZN(n6981) );
  NAND2_X1 U7750 ( .A1(n9624), .A2(n12133), .ZN(n15107) );
  NAND2_X1 U7751 ( .A1(n9666), .A2(n12184), .ZN(n15039) );
  INV_X1 U7752 ( .A(n9487), .ZN(n12004) );
  INV_X1 U7753 ( .A(n12005), .ZN(n9565) );
  AND2_X1 U7754 ( .A1(n9664), .A2(n9646), .ZN(n10008) );
  OR2_X1 U7755 ( .A1(n9498), .A2(n9497), .ZN(n9122) );
  INV_X1 U7756 ( .A(n7289), .ZN(n7288) );
  OAI21_X1 U7757 ( .B1(n9442), .B2(n7290), .A(n9456), .ZN(n7289) );
  NOR2_X1 U7758 ( .A1(n9055), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n9383) );
  INV_X1 U7759 ( .A(n7301), .ZN(n7300) );
  OAI21_X1 U7760 ( .B1(n9330), .B2(n7302), .A(n9346), .ZN(n7301) );
  AND2_X1 U7761 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NOR2_X1 U7762 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9044) );
  NAND2_X1 U7763 ( .A1(n9047), .A2(n7514), .ZN(n9055) );
  INV_X1 U7764 ( .A(n7307), .ZN(n7306) );
  OAI21_X1 U7765 ( .B1(n9285), .B2(n7308), .A(n9300), .ZN(n7307) );
  NAND2_X1 U7766 ( .A1(n15351), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n15208) );
  AND3_X2 U7767 ( .A1(n6991), .A2(n6990), .A3(n9039), .ZN(n9218) );
  INV_X1 U7768 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U7769 ( .A1(n11561), .A2(n7442), .ZN(n13201) );
  INV_X1 U7770 ( .A(n9807), .ZN(n9824) );
  NAND2_X1 U7771 ( .A1(n7630), .A2(n7629), .ZN(n8240) );
  NOR2_X2 U7772 ( .A1(n6954), .A2(n13598), .ZN(n13327) );
  NAND2_X1 U7773 ( .A1(n6856), .A2(n6581), .ZN(n8124) );
  AOI21_X1 U7774 ( .B1(n7398), .B2(n7395), .A(n6646), .ZN(n7394) );
  INV_X1 U7775 ( .A(n7400), .ZN(n7395) );
  INV_X1 U7776 ( .A(n7398), .ZN(n7396) );
  OR2_X1 U7777 ( .A1(n13642), .A2(n13218), .ZN(n7400) );
  OR2_X1 U7778 ( .A1(n13495), .A2(n8219), .ZN(n7258) );
  AOI21_X1 U7779 ( .B1(n7408), .B2(n7405), .A(n6645), .ZN(n7404) );
  INV_X1 U7780 ( .A(n7410), .ZN(n7405) );
  OAI21_X1 U7781 ( .B1(n11412), .B2(n7888), .A(n7889), .ZN(n13554) );
  OR2_X1 U7782 ( .A1(n11488), .A2(n8211), .ZN(n8214) );
  NAND2_X1 U7783 ( .A1(n6944), .A2(n6947), .ZN(n6943) );
  XNOR2_X1 U7784 ( .A(n8764), .B(n6562), .ZN(n11006) );
  NAND2_X2 U7785 ( .A1(n13733), .A2(n9945), .ZN(n9940) );
  NAND2_X1 U7786 ( .A1(n8263), .A2(n8250), .ZN(n8266) );
  INV_X1 U7787 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U7788 ( .A1(n7344), .A2(n6849), .ZN(n6848) );
  NAND2_X1 U7789 ( .A1(n10658), .A2(n7341), .ZN(n7340) );
  INV_X1 U7790 ( .A(n7342), .ZN(n7338) );
  INV_X1 U7791 ( .A(n10660), .ZN(n7341) );
  NAND2_X1 U7792 ( .A1(n13856), .A2(n13855), .ZN(n7364) );
  NAND2_X1 U7793 ( .A1(n8456), .A2(n8455), .ZN(n12233) );
  NAND2_X1 U7794 ( .A1(n6843), .A2(n6842), .ZN(n6841) );
  INV_X1 U7795 ( .A(n12259), .ZN(n6842) );
  INV_X1 U7796 ( .A(n12258), .ZN(n6843) );
  XNOR2_X1 U7797 ( .A(n6850), .B(n12364), .ZN(n10660) );
  OAI21_X1 U7798 ( .B1(n8675), .B2(n6589), .A(n6851), .ZN(n6850) );
  NAND2_X1 U7799 ( .A1(n6552), .A2(n11448), .ZN(n6851) );
  INV_X1 U7800 ( .A(n7577), .ZN(n7576) );
  AOI21_X1 U7801 ( .B1(n7575), .B2(n7577), .A(n7574), .ZN(n7573) );
  INV_X1 U7802 ( .A(n8701), .ZN(n7574) );
  NAND2_X1 U7803 ( .A1(n14202), .A2(n14208), .ZN(n7561) );
  NAND2_X1 U7804 ( .A1(n11523), .A2(n7571), .ZN(n7570) );
  AOI21_X1 U7805 ( .B1(n11607), .B2(n13804), .A(n7572), .ZN(n7571) );
  INV_X1 U7806 ( .A(n8683), .ZN(n7572) );
  NAND2_X1 U7807 ( .A1(n11530), .A2(n8441), .ZN(n11515) );
  NOR2_X1 U7808 ( .A1(n6584), .A2(n8660), .ZN(n7564) );
  INV_X1 U7809 ( .A(n8356), .ZN(n8538) );
  INV_X1 U7810 ( .A(n9853), .ZN(n8537) );
  NAND2_X2 U7811 ( .A1(n9853), .A2(n6568), .ZN(n8356) );
  AND2_X1 U7812 ( .A1(n8665), .A2(n11924), .ZN(n10300) );
  NAND2_X1 U7813 ( .A1(n6833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U7814 ( .A(n8314), .B(n8313), .ZN(n14387) );
  OAI21_X1 U7815 ( .B1(n14414), .B2(n14468), .A(n14413), .ZN(n14428) );
  NOR2_X1 U7816 ( .A1(n6739), .A2(n14655), .ZN(n14478) );
  AND2_X1 U7817 ( .A1(n7269), .A2(n7268), .ZN(n14551) );
  INV_X1 U7818 ( .A(n12803), .ZN(n12833) );
  NAND2_X1 U7819 ( .A1(n6787), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6816) );
  OR2_X1 U7820 ( .A1(n12616), .A2(n12627), .ZN(n7138) );
  INV_X1 U7821 ( .A(n14719), .ZN(n14749) );
  AOI21_X1 U7822 ( .B1(n7581), .B2(n7580), .A(n7583), .ZN(n7579) );
  NOR2_X1 U7823 ( .A1(n14508), .A2(n14509), .ZN(n14469) );
  NAND2_X1 U7824 ( .A1(n6653), .A2(n8804), .ZN(n7542) );
  NAND2_X1 U7825 ( .A1(n8827), .A2(n6621), .ZN(n7540) );
  OAI21_X1 U7826 ( .B1(n8820), .B2(n8819), .A(n6631), .ZN(n7541) );
  INV_X1 U7827 ( .A(n11796), .ZN(n7052) );
  INV_X1 U7828 ( .A(n8838), .ZN(n7533) );
  OR2_X1 U7829 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  NAND2_X1 U7830 ( .A1(n11828), .A2(n11830), .ZN(n7056) );
  INV_X1 U7831 ( .A(n11845), .ZN(n7041) );
  NAND2_X1 U7832 ( .A1(n7045), .A2(n7042), .ZN(n11876) );
  NAND2_X1 U7833 ( .A1(n7044), .A2(n7043), .ZN(n7042) );
  INV_X1 U7834 ( .A(n7048), .ZN(n7043) );
  NAND2_X1 U7835 ( .A1(n6586), .A2(n7036), .ZN(n7035) );
  NAND2_X1 U7836 ( .A1(n11888), .A2(n11885), .ZN(n7036) );
  INV_X1 U7837 ( .A(n11885), .ZN(n7037) );
  NAND2_X1 U7838 ( .A1(n11884), .A2(n11883), .ZN(n11886) );
  OAI21_X1 U7839 ( .B1(n7470), .B2(n7465), .A(n7012), .ZN(n11883) );
  INV_X1 U7840 ( .A(n7035), .ZN(n7034) );
  NAND2_X1 U7841 ( .A1(n10394), .A2(n7219), .ZN(n7218) );
  NOR2_X1 U7842 ( .A1(n7220), .A2(n9017), .ZN(n7219) );
  INV_X1 U7843 ( .A(n7026), .ZN(n7020) );
  NAND2_X1 U7844 ( .A1(n13958), .A2(n14766), .ZN(n11770) );
  NAND2_X1 U7845 ( .A1(n8675), .A2(n6552), .ZN(n11771) );
  NAND2_X1 U7846 ( .A1(n8016), .A2(n8015), .ZN(n8023) );
  NAND2_X1 U7847 ( .A1(n6889), .A2(n7956), .ZN(n6888) );
  INV_X1 U7848 ( .A(n7954), .ZN(n6889) );
  INV_X1 U7849 ( .A(n7956), .ZN(n6890) );
  INV_X1 U7850 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U7851 ( .A1(n7957), .A2(n15251), .ZN(n7971) );
  INV_X1 U7852 ( .A(n7856), .ZN(n6897) );
  INV_X1 U7853 ( .A(n7820), .ZN(n7489) );
  OAI21_X1 U7854 ( .B1(n9903), .B2(n9895), .A(n6795), .ZN(n7701) );
  NAND2_X1 U7855 ( .A1(n9903), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U7856 ( .A1(n9902), .A2(n7078), .ZN(n7077) );
  INV_X1 U7857 ( .A(n9875), .ZN(n7078) );
  NAND2_X1 U7858 ( .A1(n6568), .A2(SI_1_), .ZN(n7076) );
  INV_X1 U7859 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7531) );
  AND2_X1 U7860 ( .A1(n14992), .A2(n10818), .ZN(n10867) );
  NAND2_X1 U7861 ( .A1(n6999), .A2(n6998), .ZN(n6790) );
  NAND2_X1 U7862 ( .A1(n11396), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U7863 ( .A1(n12673), .A2(n6995), .ZN(n12692) );
  NOR2_X1 U7864 ( .A1(n12653), .A2(n12918), .ZN(n6995) );
  NAND2_X1 U7865 ( .A1(n12579), .A2(n12792), .ZN(n6962) );
  NAND2_X1 U7866 ( .A1(n13036), .A2(n12765), .ZN(n6735) );
  OR2_X1 U7867 ( .A1(n12499), .A2(n12806), .ZN(n12129) );
  NOR2_X1 U7868 ( .A1(n9617), .A2(n6967), .ZN(n6966) );
  INV_X1 U7869 ( .A(n12103), .ZN(n6967) );
  INV_X1 U7870 ( .A(n7506), .ZN(n7505) );
  INV_X1 U7871 ( .A(n12039), .ZN(n7507) );
  NAND2_X1 U7872 ( .A1(n6796), .A2(n13018), .ZN(n15108) );
  NAND3_X1 U7873 ( .A1(n6986), .A2(n6987), .A3(n10614), .ZN(n12018) );
  INV_X1 U7874 ( .A(n9530), .ZN(n7282) );
  NAND2_X1 U7875 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  NAND2_X1 U7876 ( .A1(n9062), .A2(n6749), .ZN(n9054) );
  AND2_X1 U7877 ( .A1(n9053), .A2(n9061), .ZN(n6749) );
  NAND2_X1 U7878 ( .A1(n9431), .A2(n9111), .ZN(n9443) );
  AND2_X1 U7879 ( .A1(n9383), .A2(n9384), .ZN(n9400) );
  NAND2_X1 U7880 ( .A1(n9321), .A2(n9096), .ZN(n9331) );
  AND2_X1 U7881 ( .A1(n13119), .A2(n7427), .ZN(n7426) );
  INV_X1 U7882 ( .A(n13155), .ZN(n7424) );
  INV_X1 U7883 ( .A(n13186), .ZN(n7433) );
  INV_X1 U7884 ( .A(n6592), .ZN(n7388) );
  OR2_X1 U7885 ( .A1(n13361), .A2(n13696), .ZN(n6953) );
  INV_X1 U7886 ( .A(n8230), .ZN(n7224) );
  OR2_X1 U7887 ( .A1(n7227), .A2(n7224), .ZN(n7223) );
  AND2_X1 U7888 ( .A1(n8228), .A2(n13382), .ZN(n7227) );
  INV_X1 U7889 ( .A(n13545), .ZN(n7235) );
  AND2_X1 U7890 ( .A1(n7245), .A2(n7240), .ZN(n7233) );
  INV_X1 U7891 ( .A(n9014), .ZN(n7248) );
  INV_X1 U7892 ( .A(n7210), .ZN(n7209) );
  OAI21_X1 U7893 ( .B1(n9016), .B2(n7211), .A(n10908), .ZN(n7210) );
  INV_X1 U7894 ( .A(n9015), .ZN(n7211) );
  NAND2_X1 U7895 ( .A1(n8195), .A2(n13292), .ZN(n13386) );
  XNOR2_X1 U7896 ( .A(n8755), .B(n8754), .ZN(n8195) );
  INV_X1 U7897 ( .A(n8214), .ZN(n7238) );
  AND2_X1 U7898 ( .A1(n7243), .A2(n7241), .ZN(n7240) );
  NAND2_X1 U7899 ( .A1(n7242), .A2(n13222), .ZN(n7241) );
  OR2_X1 U7900 ( .A1(n8216), .A2(n7244), .ZN(n7243) );
  NAND2_X1 U7901 ( .A1(n7247), .A2(n8215), .ZN(n7244) );
  NAND2_X1 U7902 ( .A1(n9902), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7204) );
  NOR2_X1 U7903 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7537) );
  NOR2_X1 U7904 ( .A1(n8249), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8263) );
  AND2_X1 U7905 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  NOR2_X1 U7906 ( .A1(n6879), .A2(n11912), .ZN(n6878) );
  INV_X1 U7907 ( .A(n8605), .ZN(n7175) );
  NOR2_X1 U7908 ( .A1(n14284), .A2(n6866), .ZN(n6865) );
  INV_X1 U7909 ( .A(n6867), .ZN(n6866) );
  NOR2_X1 U7910 ( .A1(n14288), .A2(n14292), .ZN(n6867) );
  NOR2_X1 U7911 ( .A1(n11953), .A2(n7189), .ZN(n7188) );
  INV_X1 U7912 ( .A(n11838), .ZN(n7189) );
  INV_X1 U7913 ( .A(n8688), .ZN(n7587) );
  AND2_X1 U7914 ( .A1(n8387), .A2(n8388), .ZN(n11944) );
  NAND2_X1 U7915 ( .A1(n11764), .A2(n11761), .ZN(n7144) );
  NAND2_X1 U7916 ( .A1(n7201), .A2(n7200), .ZN(n7199) );
  INV_X1 U7917 ( .A(n11515), .ZN(n7201) );
  NAND2_X1 U7918 ( .A1(n8430), .A2(n8429), .ZN(n11304) );
  NAND2_X1 U7919 ( .A1(n10835), .A2(n11778), .ZN(n10770) );
  INV_X1 U7920 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6802) );
  INV_X1 U7921 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8299) );
  INV_X1 U7922 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U7923 ( .A1(n7932), .A2(n7484), .ZN(n7483) );
  INV_X1 U7924 ( .A(n7909), .ZN(n7484) );
  AOI21_X1 U7925 ( .B1(n7480), .B2(n7873), .A(n6654), .ZN(n7479) );
  INV_X1 U7926 ( .A(n7859), .ZN(n7480) );
  NOR2_X2 U7927 ( .A1(n8354), .A2(n8288), .ZN(n8414) );
  INV_X1 U7928 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8286) );
  INV_X1 U7929 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8285) );
  INV_X1 U7930 ( .A(n7461), .ZN(n7460) );
  OAI21_X1 U7931 ( .B1(n7761), .B2(n7462), .A(n7782), .ZN(n7461) );
  INV_X1 U7932 ( .A(n7763), .ZN(n7462) );
  NAND2_X1 U7933 ( .A1(n7737), .A2(n7736), .ZN(n7762) );
  INV_X1 U7934 ( .A(n7697), .ZN(n7698) );
  NAND2_X1 U7935 ( .A1(n6905), .A2(SI_3_), .ZN(n7700) );
  OAI21_X1 U7936 ( .B1(SI_3_), .B2(n6905), .A(n7700), .ZN(n7697) );
  NAND2_X1 U7937 ( .A1(n6779), .A2(n7686), .ZN(n7699) );
  NAND2_X1 U7938 ( .A1(n7455), .A2(n9874), .ZN(n7454) );
  NOR2_X1 U7939 ( .A1(n7646), .A2(n8333), .ZN(n7647) );
  NAND2_X1 U7940 ( .A1(n6733), .A2(n6732), .ZN(n6814) );
  NAND2_X1 U7941 ( .A1(n9863), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7942 ( .A1(n14436), .A2(n14396), .ZN(n6733) );
  OAI21_X1 U7943 ( .B1(n7091), .B2(n7089), .A(n6662), .ZN(n7088) );
  INV_X1 U7944 ( .A(n12460), .ZN(n7089) );
  INV_X1 U7945 ( .A(n12573), .ZN(n7096) );
  OR2_X1 U7946 ( .A1(n9553), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U7947 ( .A1(n9151), .A2(n9150), .ZN(n9436) );
  INV_X1 U7948 ( .A(n9421), .ZN(n9151) );
  AND2_X1 U7949 ( .A1(n11149), .A2(n11146), .ZN(n7085) );
  AND2_X1 U7950 ( .A1(n12452), .A2(n7072), .ZN(n7071) );
  NAND2_X1 U7951 ( .A1(n12564), .A2(n7073), .ZN(n7072) );
  INV_X1 U7952 ( .A(n12563), .ZN(n7073) );
  INV_X1 U7953 ( .A(n12564), .ZN(n7074) );
  INV_X1 U7954 ( .A(n12389), .ZN(n7109) );
  OR2_X1 U7955 ( .A1(n11682), .A2(n11683), .ZN(n11703) );
  NAND2_X1 U7956 ( .A1(n12390), .A2(n12389), .ZN(n12481) );
  INV_X1 U7957 ( .A(n11237), .ZN(n7082) );
  OAI21_X1 U7958 ( .B1(n7085), .B2(n7082), .A(n11461), .ZN(n7081) );
  NAND2_X1 U7959 ( .A1(n10535), .A2(n7132), .ZN(n7133) );
  AND2_X1 U7960 ( .A1(n10519), .A2(n10369), .ZN(n7132) );
  INV_X1 U7961 ( .A(n7131), .ZN(n7130) );
  OAI21_X1 U7962 ( .B1(n10369), .B2(n10519), .A(P3_REG1_REG_3__SCAN_IN), .ZN(
        n7131) );
  NAND2_X1 U7963 ( .A1(n7129), .A2(n10370), .ZN(n10599) );
  NAND2_X1 U7964 ( .A1(n10535), .A2(n10369), .ZN(n7129) );
  XNOR2_X1 U7965 ( .A(n10816), .B(n14982), .ZN(n14973) );
  NAND2_X1 U7966 ( .A1(n6772), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7114) );
  XNOR2_X1 U7967 ( .A(n10867), .B(n10868), .ZN(n10819) );
  NAND2_X1 U7968 ( .A1(n14991), .A2(n10796), .ZN(n6777) );
  XNOR2_X1 U7969 ( .A(n6790), .B(n11389), .ZN(n11397) );
  XNOR2_X1 U7970 ( .A(n12640), .B(n14566), .ZN(n14572) );
  NAND2_X1 U7971 ( .A1(n7138), .A2(n12645), .ZN(n12640) );
  NAND2_X1 U7972 ( .A1(n6815), .A2(n6604), .ZN(n6997) );
  AND2_X1 U7973 ( .A1(n6997), .A2(n6996), .ZN(n12673) );
  INV_X1 U7974 ( .A(n12663), .ZN(n6996) );
  AOI21_X1 U7975 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n12674), .A(n12671), .ZN(
        n12706) );
  NOR2_X1 U7976 ( .A1(n12675), .A2(n12905), .ZN(n12693) );
  INV_X1 U7977 ( .A(n12733), .ZN(n7123) );
  NAND2_X1 U7978 ( .A1(n7496), .A2(n7499), .ZN(n6825) );
  INV_X1 U7980 ( .A(n7496), .ZN(n7495) );
  INV_X1 U7981 ( .A(n7499), .ZN(n7498) );
  OAI21_X1 U7982 ( .B1(n12795), .B2(n12126), .A(n7500), .ZN(n7499) );
  OR2_X1 U7983 ( .A1(n9534), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9544) );
  INV_X1 U7984 ( .A(n12789), .ZN(n12795) );
  INV_X1 U7985 ( .A(n12860), .ZN(n12834) );
  AND2_X1 U7986 ( .A1(n12108), .A2(n12112), .ZN(n12835) );
  AND2_X1 U7987 ( .A1(n9612), .A2(n9611), .ZN(n6992) );
  OR2_X1 U7988 ( .A1(n9436), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9450) );
  AND4_X1 U7989 ( .A1(n9455), .A2(n9454), .A3(n9453), .A4(n9452), .ZN(n12900)
         );
  AND4_X1 U7990 ( .A1(n9427), .A2(n9426), .A3(n9425), .A4(n9424), .ZN(n12925)
         );
  AND2_X1 U7991 ( .A1(n12073), .A2(n12080), .ZN(n12928) );
  NOR2_X1 U7992 ( .A1(n9377), .A2(n7605), .ZN(n9378) );
  NOR2_X1 U7993 ( .A1(n9376), .A2(n14582), .ZN(n7605) );
  NAND2_X1 U7994 ( .A1(n14597), .A2(n9374), .ZN(n7527) );
  AOI21_X1 U7995 ( .B1(n6981), .B2(n6979), .A(n6661), .ZN(n6978) );
  INV_X1 U7996 ( .A(n6598), .ZN(n6979) );
  INV_X1 U7997 ( .A(n12055), .ZN(n7490) );
  NAND2_X1 U7998 ( .A1(n9146), .A2(n9145), .ZN(n9340) );
  INV_X1 U7999 ( .A(n9307), .ZN(n9146) );
  CLKBUF_X1 U8000 ( .A(n15077), .Z(n6783) );
  AND3_X1 U8001 ( .A1(n9260), .A2(n9259), .A3(n9258), .ZN(n15078) );
  NAND2_X1 U8002 ( .A1(n10641), .A2(n12133), .ZN(n15105) );
  NAND2_X1 U8003 ( .A1(n7291), .A2(n6701), .ZN(n12147) );
  NAND2_X1 U8004 ( .A1(n13085), .A2(n12004), .ZN(n7291) );
  AND3_X1 U8005 ( .A1(n9356), .A2(n9355), .A3(n9354), .ZN(n14610) );
  AND2_X1 U8006 ( .A1(n10633), .A2(n9851), .ZN(n10624) );
  OAI21_X1 U8007 ( .B1(n9564), .B2(n9132), .A(n9133), .ZN(n11993) );
  INV_X1 U8008 ( .A(n12718), .ZN(n10376) );
  OAI21_X1 U8009 ( .B1(n9541), .B2(n9128), .A(n9129), .ZN(n9552) );
  AND2_X1 U8010 ( .A1(n9636), .A2(n9635), .ZN(n9664) );
  XNOR2_X1 U8011 ( .A(n9125), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9521) );
  OAI21_X1 U8012 ( .B1(n7313), .B2(n9471), .A(n7312), .ZN(n9498) );
  INV_X1 U8013 ( .A(n7310), .ZN(n7312) );
  OAI21_X1 U8014 ( .B1(n9118), .B2(n7315), .A(n9120), .ZN(n7310) );
  NOR2_X1 U8015 ( .A1(n9054), .A2(n7513), .ZN(n7510) );
  NAND2_X1 U8016 ( .A1(n7514), .A2(n9056), .ZN(n7513) );
  OR2_X1 U8017 ( .A1(n9471), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9473) );
  AND2_X1 U8018 ( .A1(n9115), .A2(n9114), .ZN(n9456) );
  INV_X1 U8019 ( .A(n9113), .ZN(n7290) );
  AND2_X1 U8020 ( .A1(n9113), .A2(n9112), .ZN(n9442) );
  NAND2_X1 U8021 ( .A1(n6774), .A2(n9442), .ZN(n9445) );
  OR2_X1 U8022 ( .A1(n9432), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n9446) );
  AND2_X1 U8023 ( .A1(n9109), .A2(n9108), .ZN(n9411) );
  OAI21_X1 U8024 ( .B1(n9357), .B2(n7318), .A(n7316), .ZN(n9397) );
  NAND2_X1 U8025 ( .A1(n9379), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7318) );
  OAI21_X1 U8026 ( .B1(n9103), .B2(n7321), .A(n9105), .ZN(n7317) );
  AND2_X1 U8027 ( .A1(n9107), .A2(n9106), .ZN(n9396) );
  NAND2_X1 U8028 ( .A1(n9397), .A2(n9396), .ZN(n9399) );
  AND2_X1 U8029 ( .A1(n9100), .A2(n9099), .ZN(n9346) );
  INV_X1 U8030 ( .A(n9098), .ZN(n7302) );
  AND2_X1 U8031 ( .A1(n9098), .A2(n9097), .ZN(n9330) );
  NAND2_X1 U8032 ( .A1(n6773), .A2(n9330), .ZN(n9333) );
  AND2_X1 U8033 ( .A1(n9094), .A2(n9093), .ZN(n9300) );
  INV_X1 U8034 ( .A(n15208), .ZN(n7308) );
  AND2_X1 U8035 ( .A1(n15208), .A2(n9092), .ZN(n9285) );
  NAND2_X1 U8036 ( .A1(n9286), .A2(n9285), .ZN(n9288) );
  NOR2_X1 U8037 ( .A1(n9281), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9315) );
  OR2_X1 U8038 ( .A1(n9280), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n9281) );
  NOR2_X1 U8039 ( .A1(n9252), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U8040 ( .A1(n6767), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8041 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6767) );
  NAND2_X1 U8042 ( .A1(n7432), .A2(n9819), .ZN(n7431) );
  INV_X1 U8043 ( .A(n13095), .ZN(n7432) );
  NAND2_X1 U8044 ( .A1(n7434), .A2(n9695), .ZN(n7436) );
  AND2_X1 U8045 ( .A1(n7440), .A2(n9764), .ZN(n7439) );
  NAND2_X1 U8046 ( .A1(n7442), .A2(n11559), .ZN(n7440) );
  INV_X1 U8047 ( .A(n7442), .ZN(n7441) );
  NAND2_X1 U8048 ( .A1(n9736), .A2(n9735), .ZN(n10961) );
  AND4_X1 U8050 ( .A1(n8153), .A2(n8152), .A3(n8151), .A4(n8150), .ZN(n13189)
         );
  INV_X1 U8051 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7972) );
  AND4_X1 U8052 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n13096)
         );
  OR2_X1 U8053 ( .A1(n7264), .A2(n7261), .ZN(n6894) );
  NAND2_X1 U8054 ( .A1(n7265), .A2(n6608), .ZN(n13335) );
  NOR2_X1 U8055 ( .A1(n8137), .A2(n7390), .ZN(n7389) );
  INV_X1 U8056 ( .A(n8123), .ZN(n7390) );
  AOI21_X1 U8057 ( .B1(n13384), .B2(n6858), .A(n6624), .ZN(n6857) );
  INV_X1 U8058 ( .A(n8082), .ZN(n6858) );
  NAND2_X1 U8059 ( .A1(n6760), .A2(n13384), .ZN(n6856) );
  INV_X1 U8060 ( .A(n8083), .ZN(n6760) );
  INV_X1 U8061 ( .A(n13400), .ZN(n7226) );
  INV_X1 U8062 ( .A(n8228), .ZN(n7225) );
  NAND2_X1 U8063 ( .A1(n13400), .A2(n7227), .ZN(n13381) );
  NOR2_X1 U8064 ( .A1(n13422), .A2(n7392), .ZN(n7391) );
  INV_X1 U8065 ( .A(n7394), .ZN(n7392) );
  AND2_X1 U8066 ( .A1(n6612), .A2(n7986), .ZN(n6861) );
  NAND2_X1 U8067 ( .A1(n13498), .A2(n6862), .ZN(n13488) );
  NOR2_X1 U8068 ( .A1(n13491), .A2(n6863), .ZN(n6862) );
  INV_X1 U8069 ( .A(n7968), .ZN(n6863) );
  NAND2_X1 U8070 ( .A1(n13531), .A2(n13504), .ZN(n13506) );
  NAND2_X1 U8071 ( .A1(n13500), .A2(n13499), .ZN(n13498) );
  NAND2_X1 U8072 ( .A1(n13515), .A2(n8218), .ZN(n13495) );
  OR2_X1 U8073 ( .A1(n13513), .A2(n13512), .ZN(n13515) );
  NOR2_X1 U8074 ( .A1(n7402), .A2(n13524), .ZN(n7401) );
  INV_X1 U8075 ( .A(n7404), .ZN(n7402) );
  OR2_X1 U8076 ( .A1(n13718), .A2(n13222), .ZN(n7410) );
  OAI21_X1 U8077 ( .B1(n11483), .B2(n7871), .A(n7872), .ZN(n11412) );
  AOI21_X1 U8078 ( .B1(n7215), .B2(n7217), .A(n6617), .ZN(n7213) );
  INV_X1 U8079 ( .A(n7216), .ZN(n7215) );
  OAI21_X1 U8080 ( .B1(n11130), .B2(n7779), .A(n7780), .ZN(n10904) );
  OR2_X1 U8081 ( .A1(n10904), .A2(n10908), .ZN(n10905) );
  NAND2_X1 U8082 ( .A1(n7250), .A2(n7249), .ZN(n11118) );
  AND2_X1 U8083 ( .A1(n7253), .A2(n8206), .ZN(n7249) );
  NAND2_X1 U8084 ( .A1(n7382), .A2(n9018), .ZN(n7378) );
  INV_X1 U8085 ( .A(n7689), .ZN(n7382) );
  NAND2_X1 U8086 ( .A1(n7380), .A2(n9018), .ZN(n7379) );
  NAND2_X1 U8087 ( .A1(n10271), .A2(n7220), .ZN(n7690) );
  NAND2_X1 U8088 ( .A1(n13728), .A2(n7702), .ZN(n6907) );
  NAND2_X1 U8089 ( .A1(n7977), .A2(n7976), .ZN(n13651) );
  AND2_X1 U8090 ( .A1(n8268), .A2(n9939), .ZN(n9842) );
  INV_X1 U8091 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7536) );
  AOI21_X1 U8092 ( .B1(n13740), .B2(n12352), .A(n12361), .ZN(n7356) );
  INV_X1 U8093 ( .A(n7356), .ZN(n7354) );
  NAND2_X1 U8094 ( .A1(n11613), .A2(n11612), .ZN(n7331) );
  AND2_X1 U8095 ( .A1(n11624), .A2(n7331), .ZN(n7330) );
  INV_X1 U8096 ( .A(n7362), .ZN(n7361) );
  OAI21_X1 U8097 ( .B1(n13758), .B2(n7363), .A(n13844), .ZN(n7362) );
  NOR2_X1 U8098 ( .A1(n7366), .A2(n12258), .ZN(n6844) );
  OAI21_X1 U8099 ( .B1(n7367), .B2(n6840), .A(n6838), .ZN(n13831) );
  NAND2_X1 U8100 ( .A1(n12275), .A2(n13832), .ZN(n13835) );
  AOI21_X1 U8101 ( .B1(n6838), .B2(n6840), .A(n13833), .ZN(n6836) );
  NOR2_X1 U8102 ( .A1(n8578), .A2(n8320), .ZN(n8321) );
  AND4_X1 U8103 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n13914)
         );
  AND4_X1 U8104 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(n13817)
         );
  AND4_X1 U8105 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n8425), .ZN(n13774)
         );
  XNOR2_X1 U8106 ( .A(n10201), .B(n6826), .ZN(n9852) );
  XNOR2_X1 U8107 ( .A(n10201), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9859) );
  OR2_X1 U8108 ( .A1(n10250), .A2(n10249), .ZN(n6926) );
  NAND2_X1 U8109 ( .A1(n6926), .A2(n6925), .ZN(n6924) );
  NAND2_X1 U8110 ( .A1(n10246), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6925) );
  OR2_X1 U8111 ( .A1(n10429), .A2(n10428), .ZN(n6931) );
  AND2_X1 U8112 ( .A1(n6931), .A2(n6930), .ZN(n10213) );
  NAND2_X1 U8113 ( .A1(n10433), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6930) );
  OR2_X1 U8114 ( .A1(n10213), .A2(n10212), .ZN(n6929) );
  NOR2_X1 U8115 ( .A1(n10759), .A2(n6692), .ZN(n10763) );
  NOR2_X1 U8116 ( .A1(n14686), .A2(n14687), .ZN(n14685) );
  INV_X1 U8117 ( .A(n14732), .ZN(n6921) );
  NAND2_X1 U8118 ( .A1(n7601), .A2(n14058), .ZN(n14052) );
  NAND2_X1 U8119 ( .A1(n14080), .A2(n14270), .ZN(n14081) );
  AND2_X1 U8120 ( .A1(n14067), .A2(n8704), .ZN(n7593) );
  NAND2_X1 U8121 ( .A1(n7156), .A2(n7154), .ZN(n14090) );
  INV_X1 U8122 ( .A(n14100), .ZN(n7155) );
  OR2_X1 U8123 ( .A1(n14107), .A2(n14108), .ZN(n14105) );
  INV_X1 U8124 ( .A(n8700), .ZN(n7578) );
  NAND2_X1 U8125 ( .A1(n14145), .A2(n8663), .ZN(n14146) );
  OR2_X2 U8126 ( .A1(n14181), .A2(n8695), .ZN(n14134) );
  NAND2_X1 U8127 ( .A1(n14134), .A2(n8699), .ZN(n14137) );
  NOR2_X1 U8128 ( .A1(n11956), .A2(n8535), .ZN(n7166) );
  NAND2_X1 U8129 ( .A1(n14170), .A2(n14182), .ZN(n7167) );
  AND4_X1 U8130 ( .A1(n8502), .A2(n8501), .A3(n8500), .A4(n8499), .ZN(n14213)
         );
  AND4_X1 U8131 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n14211)
         );
  INV_X1 U8132 ( .A(n7186), .ZN(n7185) );
  OAI21_X1 U8133 ( .B1(n11953), .B2(n7187), .A(n11844), .ZN(n7186) );
  NAND2_X1 U8134 ( .A1(n7190), .A2(n11838), .ZN(n7187) );
  NAND2_X1 U8135 ( .A1(n11690), .A2(n7188), .ZN(n7184) );
  NOR2_X1 U8136 ( .A1(n14320), .A2(n6874), .ZN(n6873) );
  INV_X1 U8137 ( .A(n6875), .ZN(n6874) );
  INV_X1 U8138 ( .A(n6601), .ZN(n7190) );
  AND4_X1 U8139 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n13928)
         );
  AND4_X1 U8140 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n13929)
         );
  AND2_X1 U8141 ( .A1(n14519), .A2(n6603), .ZN(n7569) );
  OAI21_X1 U8142 ( .B1(n11515), .B2(n7194), .A(n7192), .ZN(n11647) );
  INV_X1 U8143 ( .A(n7195), .ZN(n7194) );
  AOI21_X1 U8144 ( .B1(n7195), .B2(n7197), .A(n7193), .ZN(n7192) );
  AOI21_X1 U8145 ( .B1(n7198), .B2(n8453), .A(n7196), .ZN(n7195) );
  INV_X1 U8146 ( .A(n8464), .ZN(n7196) );
  NOR2_X1 U8147 ( .A1(n11526), .A2(n13896), .ZN(n14513) );
  AND4_X1 U8148 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n12219)
         );
  NAND2_X1 U8149 ( .A1(n8436), .A2(n8435), .ZN(n13768) );
  OAI211_X1 U8150 ( .C1(n11936), .C2(n7151), .A(n7150), .B(n10775), .ZN(n10773) );
  INV_X1 U8151 ( .A(n8360), .ZN(n7151) );
  INV_X1 U8152 ( .A(n10836), .ZN(n11936) );
  INV_X1 U8153 ( .A(n14210), .ZN(n14172) );
  NAND2_X1 U8154 ( .A1(n8607), .A2(n8606), .ZN(n12347) );
  NAND2_X1 U8155 ( .A1(n8518), .A2(n8517), .ZN(n14310) );
  XNOR2_X1 U8156 ( .A(n8657), .B(n8656), .ZN(n11924) );
  OAI21_X1 U8157 ( .B1(n8720), .B2(n8655), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8657) );
  OR2_X1 U8158 ( .A1(n8651), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n7606) );
  INV_X1 U8159 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U8160 ( .A1(n6895), .A2(n6899), .ZN(n7857) );
  OR2_X1 U8161 ( .A1(n7788), .A2(n6901), .ZN(n6895) );
  OR2_X1 U8162 ( .A1(n8433), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U8163 ( .A1(n7802), .A2(n7801), .ZN(n7806) );
  NAND2_X1 U8164 ( .A1(n7806), .A2(n7805), .ZN(n7821) );
  NAND2_X1 U8165 ( .A1(n7453), .A2(n7668), .ZN(n7685) );
  NAND2_X1 U8166 ( .A1(n7454), .A2(n7647), .ZN(n7453) );
  NAND2_X1 U8167 ( .A1(n7454), .A2(n7668), .ZN(n7649) );
  XNOR2_X1 U8168 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14435) );
  XNOR2_X1 U8169 ( .A(n14398), .B(n7278), .ZN(n14441) );
  NOR2_X1 U8170 ( .A1(n14404), .A2(n14403), .ZN(n14453) );
  NOR2_X1 U8171 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14445), .ZN(n14403) );
  AOI21_X1 U8172 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15003), .A(n14409), .ZN(
        n14462) );
  AOI22_X1 U8173 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n14416), .B1(n14428), 
        .B2(n14415), .ZN(n14473) );
  NAND2_X1 U8174 ( .A1(n10620), .A2(n10618), .ZN(n10690) );
  AND4_X1 U8175 ( .A1(n9441), .A2(n9440), .A3(n9439), .A4(n9438), .ZN(n12913)
         );
  AND2_X1 U8176 ( .A1(n12583), .A2(n12404), .ZN(n12504) );
  NAND2_X1 U8177 ( .A1(n9435), .A2(n9434), .ZN(n12903) );
  AND2_X1 U8178 ( .A1(n7103), .A2(n7102), .ZN(n12572) );
  OAI211_X1 U8179 ( .C1(n9369), .C2(n9519), .A(n9518), .B(n9517), .ZN(n12803)
         );
  NAND2_X1 U8180 ( .A1(n7113), .A2(n7112), .ZN(n14991) );
  INV_X1 U8181 ( .A(n14988), .ZN(n7112) );
  INV_X1 U8182 ( .A(n7001), .ZN(n10873) );
  INV_X1 U8183 ( .A(n7006), .ZN(n12618) );
  INV_X1 U8184 ( .A(n6775), .ZN(n11537) );
  INV_X1 U8185 ( .A(n7003), .ZN(n12658) );
  INV_X1 U8186 ( .A(n7139), .ZN(n12614) );
  OR2_X1 U8187 ( .A1(n14564), .A2(n14565), .ZN(n6815) );
  INV_X1 U8188 ( .A(n7124), .ZN(n12734) );
  OR2_X1 U8189 ( .A1(n12731), .A2(n12730), .ZN(n6818) );
  INV_X1 U8190 ( .A(n12176), .ZN(n6784) );
  NOR2_X1 U8191 ( .A1(n12155), .A2(n9579), .ZN(n6785) );
  NAND2_X1 U8192 ( .A1(n12751), .A2(n6972), .ZN(n12943) );
  NOR2_X1 U8193 ( .A1(n6684), .A2(n6973), .ZN(n6972) );
  NOR2_X1 U8194 ( .A1(n12752), .A2(n15107), .ZN(n6973) );
  NAND2_X1 U8195 ( .A1(n12780), .A2(n6629), .ZN(n12951) );
  NOR2_X1 U8196 ( .A1(n10974), .A2(n15098), .ZN(n12889) );
  NAND2_X1 U8197 ( .A1(n9462), .A2(n9461), .ZN(n13062) );
  OR2_X1 U8198 ( .A1(n15169), .A2(n15098), .ZN(n13074) );
  CLKBUF_X1 U8199 ( .A(n9350), .Z(n9351) );
  OR3_X1 U8200 ( .A1(n9850), .A2(n11674), .A3(n9849), .ZN(n9943) );
  AND2_X1 U8201 ( .A1(n11561), .A2(n9760), .ZN(n11658) );
  NAND2_X1 U8202 ( .A1(n10961), .A2(n7438), .ZN(n11192) );
  AND2_X1 U8203 ( .A1(n11193), .A2(n9739), .ZN(n7438) );
  NAND2_X1 U8204 ( .A1(n8040), .A2(n8039), .ZN(n13636) );
  NAND2_X1 U8205 ( .A1(n8025), .A2(n8024), .ZN(n13642) );
  AND2_X1 U8206 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  XNOR2_X1 U8207 ( .A(n13385), .B(n13384), .ZN(n13623) );
  INV_X1 U8208 ( .A(n6942), .ZN(n6941) );
  NAND2_X1 U8209 ( .A1(n14929), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U8210 ( .A1(n8247), .A2(n6860), .ZN(n13595) );
  AND2_X1 U8211 ( .A1(n13322), .A2(n13318), .ZN(n6860) );
  OR2_X1 U8212 ( .A1(n11446), .A2(n11447), .ZN(n6845) );
  NAND2_X1 U8213 ( .A1(n8482), .A2(n8481), .ZN(n14329) );
  NAND2_X1 U8214 ( .A1(n13898), .A2(n12287), .ZN(n13783) );
  AND2_X1 U8215 ( .A1(n13802), .A2(n13800), .ZN(n6744) );
  XNOR2_X1 U8216 ( .A(n10660), .B(n10659), .ZN(n10661) );
  OR2_X1 U8217 ( .A1(n10304), .A2(n10293), .ZN(n13938) );
  AND2_X1 U8218 ( .A1(n11928), .A2(n10047), .ZN(n14174) );
  INV_X1 U8219 ( .A(n12219), .ZN(n13950) );
  NOR2_X1 U8220 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  NAND2_X1 U8221 ( .A1(n13991), .A2(n14749), .ZN(n6911) );
  AOI21_X1 U8222 ( .B1(n13989), .B2(n14753), .A(n14726), .ZN(n6916) );
  OAI21_X1 U8223 ( .B1(n13995), .B2(n14761), .A(n13994), .ZN(n6913) );
  NAND2_X1 U8224 ( .A1(n8645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8536) );
  OR2_X1 U8225 ( .A1(n8525), .A2(n6595), .ZN(n8645) );
  NAND2_X1 U8226 ( .A1(n14517), .A2(n10746), .ZN(n14233) );
  NAND2_X1 U8227 ( .A1(n6578), .A2(n6805), .ZN(n7170) );
  NAND2_X1 U8228 ( .A1(n9853), .A2(n6622), .ZN(n8328) );
  INV_X1 U8229 ( .A(n14498), .ZN(n6740) );
  OR2_X1 U8230 ( .A1(n14497), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n6741) );
  INV_X1 U8231 ( .A(n14653), .ZN(n6792) );
  INV_X1 U8232 ( .A(n14671), .ZN(n6822) );
  NAND2_X1 U8233 ( .A1(n6708), .A2(n6707), .ZN(n8786) );
  INV_X1 U8234 ( .A(n8785), .ZN(n6708) );
  INV_X1 U8235 ( .A(n8784), .ZN(n6707) );
  INV_X1 U8236 ( .A(n8796), .ZN(n6761) );
  INV_X1 U8237 ( .A(n11763), .ZN(n11766) );
  NAND2_X1 U8238 ( .A1(n8815), .A2(n8814), .ZN(n8820) );
  NAND2_X1 U8239 ( .A1(n11786), .A2(n7599), .ZN(n11792) );
  OR2_X1 U8240 ( .A1(n11785), .A2(n11784), .ZN(n7599) );
  OR2_X1 U8241 ( .A1(n11798), .A2(n11796), .ZN(n7051) );
  NAND2_X1 U8242 ( .A1(n6725), .A2(n6724), .ZN(n7604) );
  INV_X1 U8243 ( .A(n8832), .ZN(n6724) );
  NAND2_X1 U8244 ( .A1(n6600), .A2(n8850), .ZN(n7543) );
  AND2_X1 U8245 ( .A1(n7064), .A2(n11808), .ZN(n7063) );
  INV_X1 U8246 ( .A(n11807), .ZN(n7064) );
  NAND2_X1 U8247 ( .A1(n11819), .A2(n11821), .ZN(n7054) );
  INV_X1 U8248 ( .A(n8893), .ZN(n7539) );
  NAND2_X1 U8249 ( .A1(n8897), .A2(n8896), .ZN(n8900) );
  OR2_X1 U8250 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U8251 ( .A1(n7550), .A2(n7551), .ZN(n7549) );
  INV_X1 U8252 ( .A(n8911), .ZN(n7550) );
  OAI21_X1 U8253 ( .B1(n11834), .B2(n11833), .A(n11832), .ZN(n11837) );
  AND2_X1 U8254 ( .A1(n7040), .A2(n11851), .ZN(n7039) );
  OR2_X1 U8255 ( .A1(n11842), .A2(n7041), .ZN(n7040) );
  OAI21_X1 U8256 ( .B1(n13122), .B2(n6565), .A(n8914), .ZN(n8915) );
  NOR2_X1 U8257 ( .A1(n11872), .A2(n11870), .ZN(n7048) );
  OAI21_X1 U8258 ( .B1(n11862), .B2(n11861), .A(n11860), .ZN(n11864) );
  NOR2_X1 U8259 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  INV_X1 U8260 ( .A(n7450), .ZN(n7047) );
  AOI21_X1 U8261 ( .B1(n11869), .B2(n11868), .A(n7451), .ZN(n7450) );
  INV_X1 U8262 ( .A(n11867), .ZN(n7451) );
  INV_X1 U8263 ( .A(n7049), .ZN(n7044) );
  AOI21_X1 U8264 ( .B1(n11870), .B2(n11872), .A(n6663), .ZN(n7049) );
  NAND2_X1 U8265 ( .A1(n7469), .A2(n11879), .ZN(n7468) );
  INV_X1 U8266 ( .A(n11878), .ZN(n7469) );
  NAND2_X1 U8267 ( .A1(n6652), .A2(n8934), .ZN(n7547) );
  NAND2_X1 U8268 ( .A1(n7463), .A2(n11878), .ZN(n7466) );
  OR2_X1 U8269 ( .A1(n11874), .A2(n11877), .ZN(n7470) );
  AND2_X1 U8270 ( .A1(n7468), .A2(n7013), .ZN(n7012) );
  INV_X1 U8271 ( .A(n11882), .ZN(n7013) );
  INV_X1 U8272 ( .A(n8942), .ZN(n7556) );
  INV_X1 U8273 ( .A(n7890), .ZN(n7891) );
  NOR2_X1 U8274 ( .A1(n7478), .A2(n7892), .ZN(n7477) );
  INV_X1 U8275 ( .A(n7479), .ZN(n7478) );
  NOR2_X1 U8276 ( .A1(n7873), .A2(n7892), .ZN(n7475) );
  INV_X1 U8277 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7509) );
  INV_X1 U8278 ( .A(n7378), .ZN(n6853) );
  NOR2_X1 U8279 ( .A1(n11277), .A2(n11479), .ZN(n6956) );
  INV_X1 U8280 ( .A(n7033), .ZN(n7032) );
  OAI21_X1 U8281 ( .B1(n7035), .B2(n6585), .A(n6570), .ZN(n7033) );
  INV_X1 U8282 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15377) );
  INV_X1 U8283 ( .A(n7104), .ZN(n7093) );
  OR2_X1 U8284 ( .A1(n12573), .A2(n7102), .ZN(n7100) );
  NAND2_X1 U8285 ( .A1(n10531), .A2(n6633), .ZN(n10359) );
  XNOR2_X1 U8286 ( .A(n7128), .B(n10383), .ZN(n10375) );
  NOR2_X1 U8287 ( .A1(n10815), .A2(n9243), .ZN(n6713) );
  AOI21_X1 U8288 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n14962), .A(n14959), .ZN(
        n10794) );
  NAND2_X1 U8289 ( .A1(n9155), .A2(n9154), .ZN(n9515) );
  NAND2_X1 U8290 ( .A1(n12021), .A2(n12022), .ZN(n9580) );
  AND2_X1 U8291 ( .A1(n6615), .A2(n7530), .ZN(n7529) );
  NOR2_X1 U8292 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7530) );
  INV_X1 U8293 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9137) );
  AND2_X1 U8294 ( .A1(n9640), .A2(n9136), .ZN(n9637) );
  INV_X1 U8295 ( .A(n9107), .ZN(n7295) );
  NAND2_X1 U8296 ( .A1(n9906), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n15210) );
  AND2_X1 U8297 ( .A1(n7828), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7846) );
  NOR2_X1 U8298 ( .A1(n7814), .A2(n10072), .ZN(n7828) );
  NOR2_X1 U8299 ( .A1(n7901), .A2(n7900), .ZN(n7925) );
  AOI22_X1 U8300 ( .A1(n13311), .A2(n8943), .B1(n8946), .B2(n13208), .ZN(n8993) );
  NOR2_X1 U8301 ( .A1(n11115), .A2(n7218), .ZN(n9019) );
  OR2_X1 U8302 ( .A1(n8181), .A2(n11740), .ZN(n7654) );
  OR2_X1 U8303 ( .A1(n7660), .A2(n11737), .ZN(n7652) );
  INV_X1 U8304 ( .A(n8233), .ZN(n7262) );
  NOR2_X1 U8305 ( .A1(n13330), .A2(n7263), .ZN(n6892) );
  INV_X1 U8306 ( .A(n8234), .ZN(n7263) );
  NOR2_X1 U8307 ( .A1(n13436), .A2(n13705), .ZN(n6940) );
  AND2_X1 U8308 ( .A1(n7978), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U8309 ( .A1(n7255), .A2(n7254), .ZN(n13444) );
  NOR2_X1 U8310 ( .A1(n7256), .A2(n6630), .ZN(n7254) );
  INV_X1 U8311 ( .A(n8210), .ZN(n7217) );
  NOR2_X1 U8312 ( .A1(n8205), .A2(n7252), .ZN(n7251) );
  INV_X1 U8313 ( .A(n8203), .ZN(n7252) );
  NAND2_X1 U8314 ( .A1(n11270), .A2(n6956), .ZN(n11484) );
  NAND2_X1 U8315 ( .A1(n11270), .A2(n11269), .ZN(n11349) );
  NOR2_X1 U8316 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7428) );
  AND2_X1 U8317 ( .A1(n7810), .A2(n7809), .ZN(n7919) );
  NAND4_X1 U8318 ( .A1(n7715), .A2(n7679), .A3(n7713), .A4(n7740), .ZN(n7742)
         );
  AOI21_X1 U8319 ( .B1(n7330), .B2(n7328), .A(n11711), .ZN(n7327) );
  INV_X1 U8320 ( .A(n7330), .ZN(n7329) );
  INV_X1 U8321 ( .A(n11614), .ZN(n7328) );
  INV_X1 U8323 ( .A(n7062), .ZN(n7061) );
  OAI21_X1 U8324 ( .B1(n11908), .B2(n8713), .A(n10282), .ZN(n7062) );
  NAND2_X1 U8325 ( .A1(n7026), .A2(n7025), .ZN(n7024) );
  NAND2_X1 U8326 ( .A1(n11915), .A2(n11916), .ZN(n7029) );
  NAND2_X1 U8327 ( .A1(n6718), .A2(n7019), .ZN(n6738) );
  INV_X1 U8328 ( .A(n7022), .ZN(n6718) );
  OR2_X1 U8329 ( .A1(n14320), .A2(n14213), .ZN(n11844) );
  NOR2_X1 U8330 ( .A1(n14329), .A2(n13868), .ZN(n6875) );
  AND2_X1 U8331 ( .A1(n8457), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8472) );
  AND2_X1 U8332 ( .A1(n11162), .A2(n11632), .ZN(n11161) );
  NOR2_X1 U8333 ( .A1(n11795), .A2(n11789), .ZN(n6870) );
  NAND2_X1 U8334 ( .A1(n11033), .A2(n11944), .ZN(n11032) );
  NAND2_X1 U8335 ( .A1(n10300), .A2(n11925), .ZN(n10281) );
  OAI21_X1 U8336 ( .B1(n11033), .B2(n7178), .A(n7177), .ZN(n11160) );
  NAND2_X1 U8337 ( .A1(n8388), .A2(n8400), .ZN(n7178) );
  NAND2_X1 U8338 ( .A1(n7179), .A2(n8400), .ZN(n7177) );
  AND3_X1 U8339 ( .A1(n10840), .A2(n6870), .A3(n6869), .ZN(n11162) );
  INV_X1 U8340 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8298) );
  INV_X1 U8341 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U8342 ( .A1(n6886), .A2(n6884), .ZN(n8016) );
  AOI21_X1 U8343 ( .B1(n6606), .B2(n6890), .A(n6885), .ZN(n6884) );
  INV_X1 U8344 ( .A(n7971), .ZN(n6885) );
  XNOR2_X1 U8345 ( .A(n8016), .B(SI_18_), .ZN(n7988) );
  AOI21_X1 U8346 ( .B1(n7804), .B2(n7488), .A(n6659), .ZN(n7486) );
  NAND2_X1 U8347 ( .A1(n6902), .A2(n7786), .ZN(n6900) );
  INV_X1 U8348 ( .A(n6902), .ZN(n6901) );
  OAI21_X1 U8349 ( .B1(n9903), .B2(n9869), .A(n6780), .ZN(n7669) );
  NAND2_X1 U8350 ( .A1(n9903), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6780) );
  AOI21_X1 U8351 ( .B1(n6814), .B2(n6813), .A(n6812), .ZN(n14398) );
  AND2_X1 U8352 ( .A1(n14397), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6812) );
  INV_X1 U8353 ( .A(n14434), .ZN(n6813) );
  INV_X1 U8354 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14397) );
  INV_X1 U8355 ( .A(n6734), .ZN(n14402) );
  OAI21_X1 U8356 ( .B1(n14431), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6658), .ZN(
        n6734) );
  INV_X1 U8357 ( .A(n7277), .ZN(n14400) );
  INV_X1 U8358 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14401) );
  XNOR2_X1 U8359 ( .A(n14402), .B(n14401), .ZN(n14445) );
  INV_X1 U8360 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U8361 ( .A1(n9158), .A2(n12574), .ZN(n9553) );
  NAND2_X1 U8362 ( .A1(n9179), .A2(n7075), .ZN(n7079) );
  NAND2_X1 U8363 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  INV_X1 U8364 ( .A(n12474), .ZN(n6702) );
  OR2_X1 U8365 ( .A1(n9404), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9421) );
  NOR2_X1 U8366 ( .A1(n12586), .A2(n7066), .ZN(n7065) );
  INV_X1 U8367 ( .A(n12402), .ZN(n7066) );
  NAND2_X1 U8368 ( .A1(n9640), .A2(n7528), .ZN(n9635) );
  AND2_X1 U8369 ( .A1(n6615), .A2(n9136), .ZN(n7528) );
  OR2_X1 U8370 ( .A1(n12178), .A2(n12152), .ZN(n12157) );
  NAND2_X1 U8371 ( .A1(n12156), .A2(n7323), .ZN(n6727) );
  NAND2_X1 U8372 ( .A1(n12179), .A2(n12743), .ZN(n7323) );
  INV_X1 U8373 ( .A(n12157), .ZN(n7326) );
  NOR2_X1 U8374 ( .A1(n12182), .A2(n12183), .ZN(n7517) );
  OAI22_X1 U8375 ( .A1(n11984), .A2(n9176), .B1(n6556), .B2(n10557), .ZN(n6988) );
  OR2_X1 U8376 ( .A1(n9423), .A2(n6736), .ZN(n6989) );
  OAI21_X1 U8377 ( .B1(n10548), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6721), .ZN(
        n10537) );
  NAND2_X1 U8378 ( .A1(n10548), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6721) );
  INV_X1 U8379 ( .A(n6994), .ZN(n10812) );
  NOR2_X1 U8380 ( .A1(n10793), .A2(n7127), .ZN(n14961) );
  AND2_X1 U8381 ( .A1(n7128), .A2(n10814), .ZN(n7127) );
  AND2_X1 U8382 ( .A1(n6994), .A2(n6993), .ZN(n14957) );
  NAND2_X1 U8383 ( .A1(n10813), .A2(n10814), .ZN(n6993) );
  OR2_X1 U8384 ( .A1(n14973), .A2(n9265), .ZN(n7009) );
  OR2_X1 U8385 ( .A1(n10869), .A2(n10870), .ZN(n7001) );
  INV_X1 U8386 ( .A(n6999), .ZN(n11395) );
  OR2_X1 U8387 ( .A1(n10854), .A2(n10855), .ZN(n7137) );
  INV_X1 U8388 ( .A(n6777), .ZN(n10853) );
  OR3_X1 U8389 ( .A1(n15010), .A2(n12629), .A3(n12628), .ZN(n12647) );
  NAND2_X1 U8390 ( .A1(n6816), .A2(n6610), .ZN(n7003) );
  NAND2_X1 U8391 ( .A1(n12619), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7140) );
  AND2_X1 U8392 ( .A1(n12694), .A2(n12695), .ZN(n6788) );
  OR2_X1 U8393 ( .A1(n12735), .A2(n7126), .ZN(n7121) );
  AND2_X1 U8394 ( .A1(n12735), .A2(n7126), .ZN(n7120) );
  NOR2_X1 U8395 ( .A1(n12753), .A2(n9578), .ZN(n12155) );
  NAND2_X1 U8396 ( .A1(n6961), .A2(n6627), .ZN(n12748) );
  AND2_X1 U8397 ( .A1(n6961), .A2(n6960), .ZN(n12749) );
  NAND2_X1 U8398 ( .A1(n12146), .A2(n12139), .ZN(n12754) );
  NAND2_X1 U8399 ( .A1(n9621), .A2(n6962), .ZN(n12761) );
  NAND2_X1 U8400 ( .A1(n12120), .A2(n12121), .ZN(n12807) );
  NAND2_X1 U8401 ( .A1(n12802), .A2(n12807), .ZN(n12801) );
  AND3_X1 U8402 ( .A1(n9528), .A2(n9527), .A3(n9526), .ZN(n12821) );
  AND2_X1 U8403 ( .A1(n6964), .A2(n9616), .ZN(n12817) );
  AND2_X1 U8404 ( .A1(n12104), .A2(n12103), .ZN(n12846) );
  AOI21_X1 U8405 ( .B1(n9470), .B2(n12094), .A(n9469), .ZN(n12856) );
  INV_X1 U8406 ( .A(n12871), .ZN(n9612) );
  INV_X1 U8407 ( .A(n9450), .ZN(n9152) );
  OAI21_X1 U8408 ( .B1(n6574), .B2(n7526), .A(n12073), .ZN(n7525) );
  INV_X1 U8409 ( .A(n9410), .ZN(n7526) );
  INV_X1 U8410 ( .A(n6978), .ZN(n6977) );
  NAND2_X1 U8411 ( .A1(n9148), .A2(n9147), .ZN(n9389) );
  NAND2_X1 U8412 ( .A1(n9149), .A2(n15366), .ZN(n9404) );
  INV_X1 U8413 ( .A(n9389), .ZN(n9149) );
  OR2_X1 U8414 ( .A1(n9375), .A2(n11593), .ZN(n14582) );
  OR3_X1 U8415 ( .A1(n9340), .A2(P3_REG3_REG_11__SCAN_IN), .A3(
        P3_REG3_REG_12__SCAN_IN), .ZN(n9366) );
  OR2_X1 U8416 ( .A1(n12606), .A2(n14603), .ZN(n12059) );
  NAND2_X1 U8417 ( .A1(n6982), .A2(n6984), .ZN(n11594) );
  NAND2_X1 U8418 ( .A1(n6983), .A2(n6598), .ZN(n6982) );
  INV_X1 U8419 ( .A(n6746), .ZN(n6983) );
  OAI21_X1 U8420 ( .B1(n15051), .B2(n9306), .A(n12051), .ZN(n15026) );
  NAND2_X1 U8421 ( .A1(n9263), .A2(n9262), .ZN(n9292) );
  AOI21_X1 U8422 ( .B1(n7505), .B2(n7507), .A(n7503), .ZN(n7502) );
  INV_X1 U8423 ( .A(n12042), .ZN(n7503) );
  AND2_X1 U8424 ( .A1(n9227), .A2(n9226), .ZN(n9241) );
  AND2_X1 U8425 ( .A1(n9241), .A2(n15331), .ZN(n9263) );
  NOR2_X1 U8426 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9227) );
  NAND2_X1 U8427 ( .A1(n10617), .A2(n12018), .ZN(n15097) );
  INV_X1 U8428 ( .A(n11591), .ZN(n15115) );
  NOR2_X1 U8429 ( .A1(n9679), .A2(n9670), .ZN(n10643) );
  NAND2_X1 U8430 ( .A1(n7322), .A2(n9131), .ZN(n9564) );
  OR2_X1 U8431 ( .A1(n9552), .A2(n9130), .ZN(n7322) );
  INV_X1 U8432 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9161) );
  AND2_X1 U8433 ( .A1(n9126), .A2(n7282), .ZN(n7281) );
  OR2_X1 U8434 ( .A1(n9125), .A2(n15371), .ZN(n9126) );
  XNOR2_X1 U8435 ( .A(n9067), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12014) );
  NOR2_X1 U8436 ( .A1(n9054), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U8437 ( .A1(n9473), .A2(n9118), .ZN(n9484) );
  OR2_X1 U8438 ( .A1(n9116), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9117) );
  OAI21_X1 U8439 ( .B1(n9399), .B2(n7296), .A(n7293), .ZN(n9429) );
  INV_X1 U8440 ( .A(n9411), .ZN(n7296) );
  AOI21_X1 U8441 ( .B1(n9411), .B2(n7295), .A(n7294), .ZN(n7293) );
  INV_X1 U8442 ( .A(n9109), .ZN(n7294) );
  AND2_X1 U8443 ( .A1(n9111), .A2(n9110), .ZN(n9428) );
  AND2_X1 U8444 ( .A1(n9400), .A2(n9048), .ZN(n9416) );
  INV_X1 U8445 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U8446 ( .A1(n9359), .A2(n9103), .ZN(n9380) );
  OR2_X1 U8447 ( .A1(n9101), .A2(n10157), .ZN(n9102) );
  OR2_X1 U8448 ( .A1(n9357), .A2(n10158), .ZN(n9359) );
  AOI21_X1 U8449 ( .B1(n7306), .B2(n7308), .A(n7305), .ZN(n7304) );
  INV_X1 U8450 ( .A(n9094), .ZN(n7305) );
  AND2_X1 U8451 ( .A1(n9091), .A2(n9089), .ZN(n9271) );
  AND2_X1 U8452 ( .A1(n9084), .A2(n9083), .ZN(n9236) );
  OR2_X1 U8453 ( .A1(n9234), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9252) );
  AND2_X1 U8454 ( .A1(n9081), .A2(n9080), .ZN(n9220) );
  AND2_X1 U8455 ( .A1(n9077), .A2(n9076), .ZN(n9199) );
  OAI211_X1 U8456 ( .C1(n7142), .C2(n10356), .A(n6715), .B(n7143), .ZN(n6714)
         );
  NAND2_X1 U8457 ( .A1(n9415), .A2(n9039), .ZN(n7143) );
  INV_X1 U8458 ( .A(n9218), .ZN(n6715) );
  XNOR2_X1 U8459 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9178) );
  NAND2_X1 U8460 ( .A1(n9073), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9191) );
  INV_X1 U8461 ( .A(n7430), .ZN(n7429) );
  OAI22_X1 U8462 ( .A1(n6597), .A2(n7431), .B1(n9822), .B2(n9823), .ZN(n7430)
         );
  NAND2_X1 U8463 ( .A1(n7846), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7865) );
  OR2_X1 U8464 ( .A1(n7865), .A2(n10149), .ZN(n7882) );
  INV_X1 U8465 ( .A(n13147), .ZN(n7417) );
  NOR2_X1 U8466 ( .A1(n7417), .A2(n7416), .ZN(n7415) );
  INV_X1 U8467 ( .A(n13103), .ZN(n7416) );
  AOI21_X1 U8468 ( .B1(n7426), .B2(n7424), .A(n6620), .ZN(n7423) );
  INV_X1 U8469 ( .A(n7426), .ZN(n7425) );
  AND2_X1 U8470 ( .A1(n7435), .A2(n9699), .ZN(n6706) );
  NAND2_X1 U8471 ( .A1(n9812), .A2(n6597), .ZN(n13184) );
  INV_X1 U8472 ( .A(n8754), .ZN(n9694) );
  NAND2_X1 U8473 ( .A1(n7384), .A2(n7383), .ZN(n13331) );
  NAND2_X1 U8474 ( .A1(n8124), .A2(n6573), .ZN(n7384) );
  AOI21_X1 U8475 ( .B1(n6573), .B2(n7388), .A(n6647), .ZN(n7383) );
  NOR2_X1 U8476 ( .A1(n13347), .A2(n6953), .ZN(n6951) );
  NOR2_X1 U8477 ( .A1(n13390), .A2(n6953), .ZN(n13364) );
  AND2_X1 U8478 ( .A1(n7223), .A2(n13372), .ZN(n7222) );
  NAND2_X1 U8479 ( .A1(n6940), .A2(n6939), .ZN(n13406) );
  INV_X1 U8480 ( .A(n6940), .ZN(n13426) );
  NAND2_X1 U8481 ( .A1(n13460), .A2(n13442), .ZN(n13436) );
  NAND2_X1 U8482 ( .A1(n8002), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8043) );
  AND2_X1 U8483 ( .A1(n13444), .A2(n13443), .ZN(n13455) );
  NAND2_X1 U8484 ( .A1(n7234), .A2(n7232), .ZN(n13513) );
  AOI21_X1 U8485 ( .B1(n7233), .B2(n7235), .A(n6616), .ZN(n7232) );
  NAND2_X1 U8486 ( .A1(n8214), .A2(n6638), .ZN(n7234) );
  INV_X1 U8487 ( .A(n13188), .ZN(n13516) );
  AND2_X1 U8488 ( .A1(n9938), .A2(n6944), .ZN(n13518) );
  AOI21_X1 U8489 ( .B1(n11176), .B2(n6855), .A(n6636), .ZN(n6854) );
  INV_X1 U8490 ( .A(n7800), .ZN(n6855) );
  AOI21_X1 U8491 ( .B1(n7209), .B2(n7211), .A(n6634), .ZN(n7207) );
  AND2_X1 U8492 ( .A1(n11137), .A2(n11107), .ZN(n11185) );
  NOR2_X1 U8493 ( .A1(n11138), .A2(n14917), .ZN(n11137) );
  NAND2_X1 U8494 ( .A1(n6937), .A2(n6936), .ZN(n11138) );
  INV_X1 U8495 ( .A(n11125), .ZN(n6937) );
  NAND2_X1 U8496 ( .A1(n7250), .A2(n8206), .ZN(n11116) );
  NAND2_X1 U8497 ( .A1(n6697), .A2(n6938), .ZN(n11125) );
  INV_X1 U8498 ( .A(n7220), .ZN(n10274) );
  NAND2_X1 U8499 ( .A1(n9940), .A2(n6568), .ZN(n7808) );
  NAND2_X1 U8500 ( .A1(n7236), .A2(n7240), .ZN(n13539) );
  NAND2_X1 U8501 ( .A1(n7238), .A2(n7237), .ZN(n7236) );
  NOR2_X1 U8502 ( .A1(n7999), .A2(n7204), .ZN(n7205) );
  INV_X1 U8503 ( .A(n14902), .ZN(n14918) );
  INV_X1 U8504 ( .A(n14905), .ZN(n14921) );
  INV_X1 U8505 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U8506 ( .A1(n7535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7639) );
  NOR2_X1 U8507 ( .A1(n8260), .A2(n8259), .ZN(n8279) );
  CLKBUF_X1 U8508 ( .A(n7916), .Z(n7917) );
  NOR2_X1 U8509 ( .A1(n7744), .A2(n7743), .ZN(n7941) );
  CLKBUF_X1 U8510 ( .A(n7742), .Z(n7743) );
  OR2_X1 U8511 ( .A1(n7666), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n7744) );
  INV_X1 U8512 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9073) );
  INV_X1 U8513 ( .A(n10661), .ZN(n7339) );
  NOR2_X1 U8514 ( .A1(n8394), .A2(n8393), .ZN(n8405) );
  AND2_X1 U8515 ( .A1(n12340), .A2(n12338), .ZN(n13813) );
  AND2_X1 U8516 ( .A1(n13812), .A2(n12331), .ZN(n13844) );
  OR2_X1 U8517 ( .A1(n8423), .A2(n8422), .ZN(n8447) );
  NOR2_X1 U8518 ( .A1(n7347), .A2(n7349), .ZN(n7345) );
  INV_X1 U8519 ( .A(n11369), .ZN(n7349) );
  INV_X1 U8520 ( .A(n11368), .ZN(n7347) );
  NAND2_X1 U8521 ( .A1(n7367), .A2(n7365), .ZN(n13923) );
  AND2_X1 U8522 ( .A1(n8713), .A2(n14393), .ZN(n11928) );
  AND4_X1 U8523 ( .A1(n8643), .A2(n8642), .A3(n8641), .A4(n8640), .ZN(n12371)
         );
  AND4_X1 U8524 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n13804)
         );
  NAND2_X1 U8525 ( .A1(n10315), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6928) );
  NOR2_X1 U8526 ( .A1(n10762), .A2(n10763), .ZN(n10942) );
  NOR2_X1 U8527 ( .A1(n10942), .A2(n6934), .ZN(n10943) );
  AND2_X1 U8528 ( .A1(n10952), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8529 ( .A1(n10943), .A2(n10944), .ZN(n13965) );
  AOI21_X1 U8530 ( .B1(n14681), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14673), .ZN(
        n14690) );
  NOR2_X1 U8531 ( .A1(n14676), .A2(n6933), .ZN(n14686) );
  AND2_X1 U8532 ( .A1(n14681), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6933) );
  INV_X1 U8533 ( .A(n13967), .ZN(n13968) );
  XNOR2_X1 U8534 ( .A(n14710), .B(n13982), .ZN(n14706) );
  NOR2_X1 U8535 ( .A1(n14685), .A2(n6932), .ZN(n13967) );
  AND2_X1 U8536 ( .A1(n13980), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U8537 ( .A1(n11933), .A2(n6877), .ZN(n6876) );
  INV_X1 U8538 ( .A(n6878), .ZN(n6877) );
  AND4_X1 U8539 ( .A1(n8633), .A2(n8632), .A3(n8631), .A4(n8630), .ZN(n13741)
         );
  AND2_X1 U8540 ( .A1(n14034), .A2(n8708), .ZN(n7581) );
  INV_X1 U8541 ( .A(n8710), .ZN(n7583) );
  AOI21_X1 U8542 ( .B1(n7173), .B2(n7175), .A(n6639), .ZN(n7172) );
  AND2_X1 U8543 ( .A1(n14145), .A2(n6588), .ZN(n14080) );
  NAND2_X1 U8544 ( .A1(n14145), .A2(n6865), .ZN(n14112) );
  NAND2_X1 U8545 ( .A1(n8566), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8575) );
  AND2_X1 U8546 ( .A1(n8557), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U8547 ( .A1(n7157), .A2(n7158), .ZN(n14119) );
  AOI21_X1 U8548 ( .B1(n6569), .B2(n7165), .A(n6655), .ZN(n7158) );
  NAND2_X1 U8549 ( .A1(n7160), .A2(n7162), .ZN(n14138) );
  NAND2_X1 U8550 ( .A1(n7161), .A2(n7166), .ZN(n7160) );
  INV_X1 U8551 ( .A(n14170), .ZN(n7161) );
  NAND2_X1 U8552 ( .A1(n6587), .A2(n6596), .ZN(n7182) );
  NOR2_X1 U8553 ( .A1(n14206), .A2(n6872), .ZN(n6871) );
  INV_X1 U8554 ( .A(n6873), .ZN(n6872) );
  NAND2_X1 U8555 ( .A1(n14332), .A2(n7586), .ZN(n8690) );
  NOR2_X1 U8556 ( .A1(n14228), .A2(n7587), .ZN(n7586) );
  NAND2_X1 U8557 ( .A1(n14514), .A2(n6875), .ZN(n14220) );
  NAND2_X1 U8558 ( .A1(n14514), .A2(n14645), .ZN(n11693) );
  AND2_X1 U8559 ( .A1(n14513), .A2(n14538), .ZN(n14514) );
  AND4_X1 U8560 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(n12231)
         );
  OR2_X1 U8561 ( .A1(n11525), .A2(n13768), .ZN(n11526) );
  NAND2_X1 U8562 ( .A1(n11032), .A2(n8388), .ZN(n11050) );
  OAI21_X1 U8563 ( .B1(n11033), .B2(n7180), .A(n7176), .ZN(n11049) );
  INV_X1 U8564 ( .A(n7179), .ZN(n7176) );
  AND4_X1 U8565 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n11719)
         );
  NAND2_X1 U8566 ( .A1(n10840), .A2(n6870), .ZN(n11054) );
  AND2_X1 U8567 ( .A1(n8375), .A2(n8374), .ZN(n10775) );
  NAND2_X1 U8568 ( .A1(n10832), .A2(n8360), .ZN(n10774) );
  NAND2_X1 U8569 ( .A1(n10840), .A2(n11788), .ZN(n11039) );
  AND2_X1 U8570 ( .A1(n10838), .A2(n14774), .ZN(n10840) );
  NAND2_X1 U8571 ( .A1(n10679), .A2(n11777), .ZN(n10833) );
  NAND2_X1 U8572 ( .A1(n10833), .A2(n11936), .ZN(n10832) );
  NAND2_X1 U8573 ( .A1(n8359), .A2(n8360), .ZN(n10836) );
  NAND2_X1 U8574 ( .A1(n10837), .A2(n10836), .ZN(n10835) );
  NAND2_X1 U8575 ( .A1(n11763), .A2(n7144), .ZN(n10709) );
  INV_X1 U8576 ( .A(n13961), .ZN(n8672) );
  NAND2_X1 U8577 ( .A1(n7199), .A2(n7198), .ZN(n14523) );
  NAND2_X1 U8578 ( .A1(n7199), .A2(n7202), .ZN(n14520) );
  NAND2_X1 U8579 ( .A1(n11304), .A2(n8431), .ZN(n11532) );
  AND2_X1 U8580 ( .A1(n8381), .A2(n8380), .ZN(n14779) );
  INV_X1 U8581 ( .A(n14512), .ZN(n14252) );
  NOR2_X1 U8582 ( .A1(n10291), .A2(n8744), .ZN(n10719) );
  OAI21_X1 U8583 ( .B1(n8978), .B2(n8976), .A(n8966), .ZN(n8969) );
  NAND2_X1 U8584 ( .A1(n6803), .A2(n6801), .ZN(n8301) );
  NAND2_X1 U8585 ( .A1(n6802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U8586 ( .A1(n6804), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6803) );
  XNOR2_X1 U8587 ( .A(n8724), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8731) );
  XNOR2_X1 U8588 ( .A(n8139), .B(n8128), .ZN(n13735) );
  XNOR2_X1 U8589 ( .A(n8729), .B(n8728), .ZN(n10296) );
  OAI21_X1 U8590 ( .B1(n7606), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8729) );
  NOR2_X1 U8591 ( .A1(n6595), .A2(n7369), .ZN(n7368) );
  NAND2_X1 U8592 ( .A1(n8646), .A2(n7370), .ZN(n7369) );
  AND2_X1 U8593 ( .A1(n8417), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U8594 ( .A1(n6887), .A2(n7956), .ZN(n7970) );
  NAND2_X1 U8595 ( .A1(n7955), .A2(n7954), .ZN(n6887) );
  OR2_X1 U8596 ( .A1(n8454), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U8597 ( .A1(n7911), .A2(n7485), .ZN(n7933) );
  OAI21_X1 U8598 ( .B1(n7860), .B2(n7481), .A(n7479), .ZN(n7893) );
  NAND2_X1 U8599 ( .A1(n7860), .A2(n7859), .ZN(n7874) );
  NAND2_X1 U8600 ( .A1(n7821), .A2(n7820), .ZN(n7839) );
  INV_X1 U8601 ( .A(n7784), .ZN(n7457) );
  NAND2_X1 U8602 ( .A1(n7788), .A2(n7787), .ZN(n7802) );
  OR2_X1 U8603 ( .A1(n8389), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U8604 ( .A1(n7459), .A2(n7763), .ZN(n7783) );
  NAND2_X1 U8605 ( .A1(n7762), .A2(n7761), .ZN(n7459) );
  NAND2_X1 U8606 ( .A1(n7471), .A2(n7700), .ZN(n7710) );
  NAND2_X1 U8607 ( .A1(n7699), .A2(n7698), .ZN(n7471) );
  XNOR2_X1 U8608 ( .A(n7699), .B(n7697), .ZN(n8343) );
  INV_X1 U8609 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8284) );
  INV_X1 U8610 ( .A(n8315), .ZN(n6920) );
  NAND2_X1 U8611 ( .A1(n15481), .A2(n15482), .ZN(n6827) );
  INV_X1 U8612 ( .A(n6814), .ZN(n14433) );
  XNOR2_X1 U8613 ( .A(n14431), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14432) );
  XNOR2_X1 U8614 ( .A(n14445), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U8615 ( .A1(n14501), .A2(n14500), .ZN(n7275) );
  OAI21_X1 U8616 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14411), .A(n14410), .ZN(
        n14466) );
  AOI22_X1 U8617 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14684), .B1(n14476), 
        .B2(n14418), .ZN(n14480) );
  INV_X1 U8618 ( .A(n12597), .ZN(n12766) );
  NAND2_X1 U8619 ( .A1(n9512), .A2(n9511), .ZN(n12824) );
  NAND2_X1 U8620 ( .A1(n11703), .A2(n7110), .ZN(n12390) );
  AND2_X1 U8621 ( .A1(n11703), .A2(n11702), .ZN(n11705) );
  NAND2_X1 U8622 ( .A1(n7070), .A2(n12564), .ZN(n12453) );
  NAND2_X1 U8623 ( .A1(n6797), .A2(n12563), .ZN(n7070) );
  OAI21_X1 U8624 ( .B1(n6797), .B2(n7074), .A(n7071), .ZN(n12451) );
  INV_X1 U8625 ( .A(n7086), .ZN(n12464) );
  NAND2_X1 U8626 ( .A1(n7095), .A2(n12460), .ZN(n7090) );
  INV_X1 U8627 ( .A(n7088), .ZN(n7087) );
  NAND2_X1 U8628 ( .A1(n9533), .A2(n9532), .ZN(n12499) );
  NAND2_X1 U8629 ( .A1(n11238), .A2(n11237), .ZN(n11462) );
  NAND2_X1 U8630 ( .A1(n12502), .A2(n12408), .ZN(n12510) );
  AND3_X1 U8631 ( .A1(n9538), .A2(n9537), .A3(n9536), .ZN(n12806) );
  NAND2_X1 U8632 ( .A1(n9523), .A2(n9522), .ZN(n12810) );
  NAND2_X1 U8633 ( .A1(n11147), .A2(n7085), .ZN(n11238) );
  NOR2_X1 U8634 ( .A1(n7084), .A2(n7083), .ZN(n11148) );
  INV_X1 U8635 ( .A(n11146), .ZN(n7083) );
  INV_X1 U8636 ( .A(n11147), .ZN(n7084) );
  AOI21_X1 U8637 ( .B1(n7071), .B2(n7074), .A(n6685), .ZN(n7069) );
  AOI21_X1 U8638 ( .B1(n7111), .B2(n7107), .A(n7106), .ZN(n7105) );
  INV_X1 U8639 ( .A(n12395), .ZN(n7106) );
  NAND2_X1 U8640 ( .A1(n9501), .A2(n9500), .ZN(n12837) );
  INV_X1 U8641 ( .A(n12391), .ZN(n14603) );
  NAND2_X1 U8642 ( .A1(n10625), .A2(n10932), .ZN(n14935) );
  INV_X1 U8643 ( .A(n7081), .ZN(n7080) );
  NAND2_X1 U8644 ( .A1(n10638), .A2(n10637), .ZN(n12578) );
  NAND2_X1 U8645 ( .A1(n7067), .A2(n12402), .ZN(n12585) );
  INV_X1 U8646 ( .A(n12184), .ZN(n7519) );
  NAND2_X1 U8647 ( .A1(n9560), .A2(n9559), .ZN(n12777) );
  INV_X1 U8648 ( .A(n12821), .ZN(n12791) );
  INV_X1 U8649 ( .A(n12872), .ZN(n12599) );
  INV_X1 U8650 ( .A(n12913), .ZN(n12883) );
  INV_X1 U8651 ( .A(n14591), .ZN(n12603) );
  NAND4_X1 U8652 ( .A1(n9312), .A2(n9311), .A3(n9310), .A4(n9309), .ZN(n15044)
         );
  OR2_X1 U8653 ( .A1(n9423), .A2(n14947), .ZN(n9186) );
  OR2_X1 U8654 ( .A1(n9275), .A2(n14942), .ZN(n9185) );
  OR2_X1 U8655 ( .A1(n10550), .A2(n10330), .ZN(n10552) );
  NAND2_X1 U8656 ( .A1(n7133), .A2(n10599), .ZN(n10512) );
  INV_X1 U8657 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15003) );
  INV_X1 U8658 ( .A(n7113), .ZN(n14989) );
  XNOR2_X1 U8659 ( .A(n6777), .B(n6776), .ZN(n10797) );
  NOR2_X1 U8660 ( .A1(n15236), .A2(n10797), .ZN(n10854) );
  INV_X1 U8661 ( .A(n7135), .ZN(n11382) );
  INV_X1 U8662 ( .A(n7137), .ZN(n10857) );
  INV_X1 U8663 ( .A(n6817), .ZN(n11544) );
  XNOR2_X1 U8664 ( .A(n6775), .B(n11389), .ZN(n11383) );
  NOR2_X1 U8665 ( .A1(n14571), .A2(n12641), .ZN(n12644) );
  INV_X1 U8666 ( .A(n6997), .ZN(n12664) );
  NOR2_X1 U8667 ( .A1(n12693), .A2(n6769), .ZN(n12678) );
  AND2_X1 U8668 ( .A1(n12675), .A2(n12905), .ZN(n6769) );
  XOR2_X1 U8669 ( .A(n12754), .B(n12753), .Z(n12944) );
  OAI21_X1 U8670 ( .B1(n12764), .B2(n12763), .A(n12762), .ZN(n12948) );
  OAI21_X1 U8671 ( .B1(n12796), .B2(n7495), .A(n6572), .ZN(n12762) );
  NAND2_X1 U8672 ( .A1(n12796), .A2(n7498), .ZN(n7493) );
  AOI21_X1 U8673 ( .B1(n12796), .B2(n12795), .A(n12126), .ZN(n12779) );
  NAND2_X1 U8674 ( .A1(n9615), .A2(n12103), .ZN(n12831) );
  NAND2_X1 U8675 ( .A1(n9475), .A2(n9474), .ZN(n12866) );
  NAND2_X1 U8676 ( .A1(n12882), .A2(n9611), .ZN(n12870) );
  NAND2_X1 U8677 ( .A1(n7524), .A2(n12087), .ZN(n12892) );
  NAND2_X1 U8678 ( .A1(n9449), .A2(n9448), .ZN(n12986) );
  NAND2_X1 U8679 ( .A1(n7527), .A2(n6574), .ZN(n12927) );
  INV_X1 U8680 ( .A(n12889), .ZN(n12934) );
  NAND2_X1 U8681 ( .A1(n7527), .A2(n9378), .ZN(n11668) );
  NAND2_X1 U8682 ( .A1(n6974), .A2(n6978), .ZN(n11664) );
  NAND2_X1 U8683 ( .A1(n6746), .A2(n6981), .ZN(n6974) );
  NAND2_X1 U8684 ( .A1(n7504), .A2(n12039), .ZN(n11285) );
  NAND2_X1 U8685 ( .A1(n6783), .A2(n15076), .ZN(n7504) );
  NAND2_X1 U8686 ( .A1(n10920), .A2(n9590), .ZN(n15071) );
  INV_X1 U8687 ( .A(n15123), .ZN(n15102) );
  AND2_X1 U8688 ( .A1(n10932), .A2(n15102), .ZN(n15125) );
  INV_X1 U8689 ( .A(n12147), .ZN(n13023) );
  AND2_X1 U8690 ( .A1(n12007), .A2(n12006), .ZN(n13026) );
  NOR2_X1 U8691 ( .A1(n12951), .A2(n6750), .ZN(n13033) );
  AND2_X1 U8692 ( .A1(n12952), .A2(n15168), .ZN(n6750) );
  INV_X1 U8693 ( .A(n12499), .ZN(n13039) );
  AND2_X1 U8694 ( .A1(n9652), .A2(n9651), .ZN(n13077) );
  AND2_X1 U8695 ( .A1(n9649), .A2(n9648), .ZN(n13079) );
  INV_X1 U8696 ( .A(n9851), .ZN(n13078) );
  XNOR2_X1 U8697 ( .A(n7292), .B(n12001), .ZN(n13085) );
  NAND2_X1 U8698 ( .A1(n11999), .A2(n11998), .ZN(n7292) );
  INV_X1 U8699 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9165) );
  INV_X1 U8700 ( .A(n9664), .ZN(n11504) );
  NAND2_X1 U8701 ( .A1(n9047), .A2(n7510), .ZN(n9058) );
  INV_X1 U8702 ( .A(SI_20_), .ZN(n10504) );
  XNOR2_X1 U8703 ( .A(n9065), .B(n9064), .ZN(n10611) );
  OAI21_X1 U8704 ( .B1(n6774), .B2(n7290), .A(n7288), .ZN(n9459) );
  NAND2_X1 U8705 ( .A1(n9445), .A2(n9113), .ZN(n9457) );
  INV_X1 U8706 ( .A(SI_17_), .ZN(n15251) );
  NAND2_X1 U8707 ( .A1(n9412), .A2(n9411), .ZN(n9414) );
  NAND2_X1 U8708 ( .A1(n9399), .A2(n9107), .ZN(n9412) );
  INV_X1 U8709 ( .A(SI_16_), .ZN(n15337) );
  INV_X1 U8710 ( .A(SI_15_), .ZN(n15383) );
  OAI21_X1 U8711 ( .B1(n6773), .B2(n7302), .A(n7300), .ZN(n9349) );
  NAND2_X1 U8712 ( .A1(n9333), .A2(n9098), .ZN(n9347) );
  INV_X1 U8713 ( .A(SI_11_), .ZN(n9898) );
  XNOR2_X1 U8714 ( .A(n9317), .B(n9316), .ZN(n11396) );
  INV_X1 U8715 ( .A(SI_10_), .ZN(n15445) );
  OAI21_X1 U8716 ( .B1(n9286), .B2(n7308), .A(n7306), .ZN(n9303) );
  NAND2_X1 U8717 ( .A1(n9288), .A2(n15208), .ZN(n9301) );
  NAND2_X1 U8718 ( .A1(n9284), .A2(n9283), .ZN(n14995) );
  XNOR2_X1 U8719 ( .A(n9270), .B(P3_IR_REG_7__SCAN_IN), .ZN(n14982) );
  INV_X1 U8720 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7010) );
  NOR2_X1 U8721 ( .A1(n9218), .A2(n9415), .ZN(n7011) );
  INV_X2 U8722 ( .A(n6714), .ZN(n10548) );
  NAND2_X1 U8723 ( .A1(n6768), .A2(n6766), .ZN(n9181) );
  NAND2_X1 U8724 ( .A1(n6990), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8725 ( .A1(n13184), .A2(n9819), .ZN(n13094) );
  NOR2_X1 U8726 ( .A1(n7422), .A2(n13202), .ZN(n7420) );
  NAND2_X1 U8727 ( .A1(n13598), .A2(n14638), .ZN(n7419) );
  NAND2_X1 U8728 ( .A1(n7436), .A2(n9699), .ZN(n10162) );
  OR2_X1 U8729 ( .A1(n14626), .A2(n13203), .ZN(n9765) );
  AND2_X1 U8730 ( .A1(n9720), .A2(n9719), .ZN(n10440) );
  NAND2_X1 U8731 ( .A1(n7418), .A2(n9802), .ZN(n13148) );
  NAND2_X1 U8732 ( .A1(n13104), .A2(n13103), .ZN(n7418) );
  NAND2_X1 U8733 ( .A1(n9759), .A2(n9758), .ZN(n11561) );
  AND2_X1 U8734 ( .A1(n11192), .A2(n9745), .ZN(n11334) );
  OR2_X1 U8735 ( .A1(n9836), .A2(n9835), .ZN(n13178) );
  AND2_X1 U8736 ( .A1(n9781), .A2(n9775), .ZN(n7443) );
  INV_X1 U8737 ( .A(n13172), .ZN(n9781) );
  NAND2_X1 U8738 ( .A1(n13135), .A2(n9775), .ZN(n13173) );
  INV_X1 U8739 ( .A(n13178), .ZN(n14635) );
  NAND2_X1 U8740 ( .A1(n9812), .A2(n9811), .ZN(n13187) );
  OR3_X1 U8741 ( .A1(n8974), .A2(n8973), .A3(n8972), .ZN(n13302) );
  NAND2_X1 U8742 ( .A1(n7721), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7633) );
  OR2_X1 U8743 ( .A1(n8240), .A2(n7631), .ZN(n7632) );
  INV_X2 U8744 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7656) );
  AND2_X1 U8745 ( .A1(n14835), .A2(n14834), .ZN(n14840) );
  CLKBUF_X1 U8746 ( .A(n7993), .Z(n7974) );
  INV_X1 U8747 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U8748 ( .A1(n13335), .A2(n8234), .ZN(n13323) );
  NAND2_X1 U8749 ( .A1(n7385), .A2(n6592), .ZN(n13340) );
  NAND2_X1 U8750 ( .A1(n8124), .A2(n7389), .ZN(n7385) );
  NAND2_X1 U8751 ( .A1(n8124), .A2(n8123), .ZN(n13352) );
  NAND2_X1 U8752 ( .A1(n6856), .A2(n6857), .ZN(n13373) );
  NAND2_X1 U8753 ( .A1(n13381), .A2(n8230), .ZN(n13369) );
  NOR2_X1 U8754 ( .A1(n7226), .A2(n7225), .ZN(n13383) );
  NAND2_X1 U8755 ( .A1(n7393), .A2(n7394), .ZN(n13423) );
  NAND2_X1 U8756 ( .A1(n7397), .A2(n7400), .ZN(n13435) );
  OR2_X1 U8757 ( .A1(n13453), .A2(n8033), .ZN(n7397) );
  AND2_X1 U8758 ( .A1(n7255), .A2(n7257), .ZN(n13469) );
  NAND2_X1 U8759 ( .A1(n13488), .A2(n7986), .ZN(n13467) );
  NAND2_X1 U8760 ( .A1(n13498), .A2(n7968), .ZN(n13490) );
  NAND2_X1 U8761 ( .A1(n7258), .A2(n7259), .ZN(n13480) );
  NAND2_X1 U8762 ( .A1(n7403), .A2(n7404), .ZN(n13525) );
  NAND2_X1 U8763 ( .A1(n7407), .A2(n7410), .ZN(n13546) );
  OR2_X1 U8764 ( .A1(n13554), .A2(n7908), .ZN(n7407) );
  NAND2_X1 U8765 ( .A1(n7239), .A2(n8215), .ZN(n13560) );
  NAND2_X1 U8766 ( .A1(n8214), .A2(n7246), .ZN(n7239) );
  NAND2_X1 U8767 ( .A1(n8214), .A2(n8213), .ZN(n11410) );
  NAND2_X1 U8768 ( .A1(n7214), .A2(n8210), .ZN(n11341) );
  NAND2_X1 U8769 ( .A1(n11259), .A2(n11258), .ZN(n7214) );
  NAND2_X1 U8770 ( .A1(n11177), .A2(n11176), .ZN(n11179) );
  NAND2_X1 U8771 ( .A1(n10905), .A2(n7800), .ZN(n11177) );
  NAND2_X1 U8772 ( .A1(n7208), .A2(n9015), .ZN(n10909) );
  NAND2_X1 U8773 ( .A1(n11132), .A2(n9016), .ZN(n7208) );
  NAND2_X1 U8774 ( .A1(n8204), .A2(n8203), .ZN(n10992) );
  NAND2_X1 U8775 ( .A1(n7379), .A2(n7377), .ZN(n10984) );
  AND2_X1 U8776 ( .A1(n7378), .A2(n7707), .ZN(n7377) );
  NAND2_X1 U8777 ( .A1(n7690), .A2(n7689), .ZN(n10390) );
  AND2_X1 U8778 ( .A1(n13557), .A2(n10983), .ZN(n13579) );
  AND2_X1 U8779 ( .A1(n13557), .A2(n10986), .ZN(n13577) );
  INV_X1 U8780 ( .A(n13549), .ZN(n13581) );
  NAND2_X1 U8781 ( .A1(n7946), .A2(n7945), .ZN(n14637) );
  NOR2_X1 U8782 ( .A1(n14863), .A2(n14893), .ZN(n14884) );
  CLKBUF_X1 U8783 ( .A(n14884), .Z(n14888) );
  AND2_X1 U8784 ( .A1(n9842), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14891) );
  INV_X1 U8785 ( .A(n14891), .ZN(n14893) );
  INV_X1 U8786 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13723) );
  XNOR2_X1 U8787 ( .A(n8254), .B(n8253), .ZN(n11674) );
  OAI21_X1 U8788 ( .B1(n8266), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8254) );
  XNOR2_X1 U8789 ( .A(n8251), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11641) );
  INV_X1 U8790 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10831) );
  INV_X1 U8791 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10704) );
  INV_X1 U8792 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10671) );
  INV_X1 U8793 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10137) );
  INV_X1 U8794 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10090) );
  INV_X1 U8795 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9935) );
  INV_X1 U8796 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9932) );
  INV_X1 U8797 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9925) );
  INV_X1 U8798 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9922) );
  INV_X1 U8799 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9909) );
  AND2_X1 U8800 ( .A1(n7718), .A2(n7739), .ZN(n9986) );
  INV_X1 U8801 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9913) );
  INV_X1 U8802 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9906) );
  INV_X1 U8803 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9910) );
  CLKBUF_X1 U8804 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n6810) );
  AND2_X1 U8805 ( .A1(n8638), .A2(n8621), .ZN(n14028) );
  XNOR2_X1 U8806 ( .A(n6831), .B(n13740), .ZN(n6830) );
  NAND2_X1 U8807 ( .A1(n13909), .A2(n12353), .ZN(n6831) );
  NAND2_X1 U8808 ( .A1(n7367), .A2(n12245), .ZN(n13747) );
  INV_X1 U8809 ( .A(n7333), .ZN(n11208) );
  NOR2_X1 U8810 ( .A1(n12369), .A2(n7354), .ZN(n7351) );
  OAI22_X1 U8811 ( .A1(n7354), .A2(n7353), .B1(n12369), .B2(n7356), .ZN(n7352)
         );
  NOR2_X1 U8812 ( .A1(n13740), .A2(n12369), .ZN(n7353) );
  INV_X1 U8813 ( .A(n12369), .ZN(n7355) );
  NAND2_X1 U8814 ( .A1(n7332), .A2(n7330), .ZN(n11712) );
  NAND2_X1 U8815 ( .A1(n11615), .A2(n11614), .ZN(n7332) );
  NAND2_X1 U8816 ( .A1(n7364), .A2(n12297), .ZN(n13792) );
  NAND2_X1 U8817 ( .A1(n8556), .A2(n8555), .ZN(n14288) );
  OAI21_X1 U8818 ( .B1(n12324), .B2(n7363), .A(n7361), .ZN(n13845) );
  NAND2_X1 U8819 ( .A1(n6837), .A2(n6841), .ZN(n13823) );
  NAND2_X1 U8820 ( .A1(n7367), .A2(n6844), .ZN(n6837) );
  NAND2_X1 U8821 ( .A1(n12324), .A2(n13758), .ZN(n13760) );
  NAND2_X1 U8822 ( .A1(n8587), .A2(n8586), .ZN(n14266) );
  INV_X1 U8823 ( .A(n6849), .ZN(n11226) );
  NAND2_X1 U8824 ( .A1(n13783), .A2(n12290), .ZN(n13856) );
  NAND2_X1 U8825 ( .A1(n13801), .A2(n12239), .ZN(n13863) );
  NAND2_X1 U8826 ( .A1(n7344), .A2(n7343), .ZN(n11445) );
  NAND2_X1 U8827 ( .A1(n11226), .A2(n7346), .ZN(n7343) );
  INV_X1 U8828 ( .A(n13938), .ZN(n13912) );
  INV_X1 U8829 ( .A(n13741), .ZN(n13942) );
  INV_X1 U8830 ( .A(n8675), .ZN(n13958) );
  AND3_X1 U8831 ( .A1(n9852), .A2(P1_REG1_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n10189) );
  AOI21_X1 U8832 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(n10201), .A(n10189), .ZN(
        n10497) );
  NOR2_X1 U8833 ( .A1(n10484), .A2(n6927), .ZN(n10250) );
  NOR2_X1 U8834 ( .A1(n10488), .A2(n10207), .ZN(n6927) );
  INV_X1 U8835 ( .A(n6926), .ZN(n10248) );
  AOI21_X1 U8836 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n10209), .A(n10481), .ZN(
        n10244) );
  INV_X1 U8837 ( .A(n10416), .ZN(n6923) );
  INV_X1 U8838 ( .A(n6924), .ZN(n10417) );
  INV_X1 U8839 ( .A(n6931), .ZN(n10427) );
  AOI21_X1 U8840 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10433), .A(n10430), .ZN(
        n10197) );
  INV_X1 U8841 ( .A(n6929), .ZN(n10314) );
  NAND2_X1 U8842 ( .A1(n10951), .A2(n6720), .ZN(n10953) );
  OR2_X1 U8843 ( .A1(n10952), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6720) );
  INV_X1 U8844 ( .A(n6922), .ZN(n14731) );
  AND2_X1 U8845 ( .A1(n10051), .A2(n6705), .ZN(n14753) );
  NAND2_X1 U8846 ( .A1(n14031), .A2(n7584), .ZN(n14013) );
  NAND2_X1 U8847 ( .A1(n14031), .A2(n8708), .ZN(n14011) );
  NAND2_X1 U8848 ( .A1(n14052), .A2(n8605), .ZN(n14042) );
  NAND2_X1 U8849 ( .A1(n14278), .A2(n7593), .ZN(n14075) );
  NAND2_X1 U8850 ( .A1(n14278), .A2(n8704), .ZN(n14073) );
  OR2_X1 U8851 ( .A1(n14101), .A2(n14100), .ZN(n14278) );
  NAND2_X1 U8852 ( .A1(n14105), .A2(n8572), .ZN(n14091) );
  NAND2_X1 U8853 ( .A1(n14137), .A2(n8700), .ZN(n14128) );
  AND2_X1 U8854 ( .A1(n7167), .A2(n8534), .ZN(n14162) );
  NAND2_X1 U8855 ( .A1(n7167), .A2(n7166), .ZN(n14160) );
  NAND2_X1 U8856 ( .A1(n7184), .A2(n7185), .ZN(n14209) );
  OAI21_X1 U8857 ( .B1(n11690), .B2(n7190), .A(n11838), .ZN(n14229) );
  NAND2_X1 U8858 ( .A1(n14332), .A2(n8688), .ZN(n14219) );
  NAND2_X1 U8859 ( .A1(n8687), .A2(n8686), .ZN(n11697) );
  NAND2_X1 U8860 ( .A1(n7191), .A2(n7195), .ZN(n11648) );
  NAND2_X1 U8861 ( .A1(n11515), .A2(n7198), .ZN(n7191) );
  NAND2_X1 U8862 ( .A1(n11523), .A2(n8683), .ZN(n11514) );
  NAND2_X1 U8863 ( .A1(n11979), .A2(n10302), .ZN(n14526) );
  INV_X1 U8864 ( .A(n14779), .ZN(n11795) );
  OR2_X1 U8865 ( .A1(n8356), .A2(n9869), .ZN(n8319) );
  INV_X1 U8866 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U8867 ( .A1(n8444), .A2(n8443), .ZN(n13896) );
  NAND2_X1 U8868 ( .A1(n8421), .A2(n8420), .ZN(n11810) );
  INV_X1 U8869 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7169) );
  INV_X1 U8870 ( .A(n12347), .ZN(n14350) );
  OR2_X1 U8871 ( .A1(n14297), .A2(n14296), .ZN(n14358) );
  INV_X1 U8872 ( .A(n13896), .ZN(n11607) );
  INV_X1 U8873 ( .A(n8302), .ZN(n14380) );
  INV_X1 U8874 ( .A(n8303), .ZN(n14383) );
  CLKBUF_X1 U8875 ( .A(n14387), .Z(n6705) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n15248) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11202) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10702) );
  AND2_X1 U8879 ( .A1(n8417), .A2(n8293), .ZN(n8515) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10672) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10463) );
  INV_X1 U8882 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10135) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10130) );
  INV_X1 U8884 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10091) );
  AND2_X1 U8885 ( .A1(n8434), .A2(n8454), .ZN(n10760) );
  INV_X1 U8886 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9936) );
  OR2_X1 U8887 ( .A1(n8419), .A2(n8418), .ZN(n10308) );
  INV_X1 U8888 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n15351) );
  INV_X1 U8889 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9926) );
  INV_X1 U8890 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9919) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9901) );
  INV_X1 U8892 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n15396) );
  NAND2_X1 U8893 ( .A1(n6950), .A2(n7668), .ZN(n6949) );
  INV_X1 U8894 ( .A(n7453), .ZN(n6950) );
  INV_X1 U8895 ( .A(n10201), .ZN(n9870) );
  XNOR2_X1 U8896 ( .A(n14437), .B(n6742), .ZN(n15481) );
  AND2_X1 U8897 ( .A1(n14440), .A2(n14439), .ZN(n14497) );
  XNOR2_X1 U8898 ( .A(n14432), .B(n6791), .ZN(n15472) );
  XNOR2_X1 U8899 ( .A(n14451), .B(n7276), .ZN(n14501) );
  INV_X1 U8900 ( .A(n7274), .ZN(n14505) );
  OAI21_X1 U8901 ( .B1(n14502), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6613), .ZN(
        n7274) );
  INV_X1 U8902 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6728) );
  INV_X1 U8903 ( .A(n14659), .ZN(n6729) );
  AND2_X1 U8904 ( .A1(n14486), .A2(n14487), .ZN(n14666) );
  AND2_X1 U8905 ( .A1(n12581), .A2(n12580), .ZN(n6704) );
  INV_X1 U8906 ( .A(n7141), .ZN(n12613) );
  INV_X1 U8907 ( .A(n6816), .ZN(n15004) );
  INV_X1 U8908 ( .A(n7138), .ZN(n12639) );
  INV_X1 U8909 ( .A(n6815), .ZN(n14563) );
  AOI21_X1 U8910 ( .B1(n12716), .B2(n14981), .A(n12703), .ZN(n12713) );
  AOI21_X1 U8911 ( .B1(n12385), .B2(n12889), .A(n12384), .ZN(n6743) );
  INV_X1 U8912 ( .A(n6969), .ZN(n6968) );
  OAI22_X1 U8913 ( .A1(n13029), .A2(n13001), .B1(n15181), .B2(n12945), .ZN(
        n6969) );
  OAI21_X1 U8914 ( .B1(n9674), .B2(n13074), .A(n9673), .ZN(n9675) );
  OAI21_X1 U8915 ( .B1(n13027), .B2(n15169), .A(n6752), .ZN(P3_U3455) );
  INV_X1 U8916 ( .A(n6753), .ZN(n6752) );
  OAI22_X1 U8917 ( .A1(n13029), .A2(n13074), .B1(n15170), .B2(n13028), .ZN(
        n6753) );
  INV_X1 U8918 ( .A(n7229), .ZN(n7228) );
  NAND2_X1 U8919 ( .A1(n13595), .A2(n14931), .ZN(n7231) );
  OAI21_X1 U8920 ( .B1(n13596), .B2(n13629), .A(n7230), .ZN(n7229) );
  AND2_X1 U8921 ( .A1(n8283), .A2(n6691), .ZN(n6904) );
  NAND2_X1 U8922 ( .A1(n13595), .A2(n14908), .ZN(n6859) );
  NOR2_X1 U8923 ( .A1(n10524), .A2(n7342), .ZN(n10662) );
  INV_X1 U8924 ( .A(n6913), .ZN(n6912) );
  AND2_X1 U8925 ( .A1(n7568), .A2(n7563), .ZN(n12195) );
  INV_X1 U8926 ( .A(n6747), .ZN(n14036) );
  OAI21_X1 U8927 ( .B1(n14251), .B2(n14201), .A(n6748), .ZN(n6747) );
  AOI21_X1 U8928 ( .B1(n14247), .B2(n14194), .A(n14035), .ZN(n6748) );
  NAND2_X1 U8929 ( .A1(n7567), .A2(n7565), .ZN(n8748) );
  NAND2_X1 U8930 ( .A1(n14800), .A2(n7566), .ZN(n7565) );
  NAND2_X1 U8931 ( .A1(n7170), .A2(n7168), .ZN(n8753) );
  NAND2_X1 U8932 ( .A1(n14794), .A2(n7169), .ZN(n7168) );
  OAI21_X1 U8933 ( .B1(n11727), .B2(n14390), .A(n7147), .ZN(P1_U3327) );
  NOR2_X1 U8934 ( .A1(n14384), .A2(n11726), .ZN(n7148) );
  INV_X1 U8935 ( .A(n6820), .ZN(n14651) );
  INV_X1 U8936 ( .A(n7271), .ZN(n14669) );
  INV_X1 U8937 ( .A(n7268), .ZN(n14545) );
  NOR2_X1 U8938 ( .A1(n14553), .A2(n14552), .ZN(n14562) );
  INV_X1 U8939 ( .A(n13598), .ZN(n7422) );
  AND2_X1 U8940 ( .A1(n7162), .A2(n7159), .ZN(n6569) );
  NAND2_X1 U8941 ( .A1(n11889), .A2(n11891), .ZN(n6570) );
  CLKBUF_X3 U8942 ( .A(n8181), .Z(n8149) );
  NAND2_X1 U8944 ( .A1(n12089), .A2(n12088), .ZN(n6571) );
  NAND2_X2 U8945 ( .A1(n7998), .A2(n8190), .ZN(n13292) );
  AND2_X1 U8946 ( .A1(n6825), .A2(n12763), .ZN(n6572) );
  AND2_X1 U8947 ( .A1(n13341), .A2(n7386), .ZN(n6573) );
  AND2_X1 U8948 ( .A1(n6976), .A2(n9378), .ZN(n6574) );
  INV_X1 U8949 ( .A(n8534), .ZN(n8535) );
  OR2_X1 U8950 ( .A1(n12144), .A2(n12133), .ZN(n6575) );
  AND2_X1 U8951 ( .A1(n6956), .A2(n6955), .ZN(n6576) );
  NAND2_X1 U8952 ( .A1(n14392), .A2(n9853), .ZN(n13882) );
  AND3_X1 U8953 ( .A1(n12426), .A2(n12833), .A3(n12821), .ZN(n6577) );
  AND2_X1 U8954 ( .A1(n7562), .A2(n14796), .ZN(n6578) );
  INV_X1 U8955 ( .A(n7313), .ZN(n7314) );
  NOR2_X1 U8956 ( .A1(n8220), .A2(n7260), .ZN(n6579) );
  AND2_X1 U8957 ( .A1(n14137), .A2(n7577), .ZN(n6580) );
  AND2_X1 U8958 ( .A1(n6857), .A2(n6632), .ZN(n6581) );
  NAND2_X1 U8959 ( .A1(n9182), .A2(n7079), .ZN(n10614) );
  AND2_X1 U8960 ( .A1(n7588), .A2(n8686), .ZN(n6582) );
  OR2_X1 U8961 ( .A1(n6643), .A2(n8792), .ZN(n6583) );
  INV_X1 U8962 ( .A(n7166), .ZN(n7165) );
  NAND2_X1 U8963 ( .A1(n12203), .A2(n12198), .ZN(n6584) );
  INV_X1 U8964 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U8965 ( .A1(n11887), .A2(n7037), .ZN(n6585) );
  NAND2_X1 U8966 ( .A1(n11890), .A2(n7449), .ZN(n6586) );
  INV_X1 U8967 ( .A(n11889), .ZN(n7449) );
  NAND2_X1 U8968 ( .A1(n12579), .A2(n12765), .ZN(n12125) );
  INV_X1 U8969 ( .A(n12125), .ZN(n7497) );
  NAND2_X1 U8970 ( .A1(n7185), .A2(n7183), .ZN(n6587) );
  AND2_X1 U8971 ( .A1(n6864), .A2(n6865), .ZN(n6588) );
  INV_X1 U8972 ( .A(n11957), .ZN(n7159) );
  INV_X1 U8973 ( .A(n13843), .ZN(n7363) );
  INV_X1 U8974 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10158) );
  INV_X1 U8975 ( .A(n10989), .ZN(n6938) );
  INV_X1 U8976 ( .A(n8346), .ZN(n8363) );
  OR2_X2 U8977 ( .A1(n10282), .A2(n10286), .ZN(n6589) );
  OR2_X1 U8978 ( .A1(n10816), .A2(n14982), .ZN(n6590) );
  OR3_X1 U8979 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10366), .ZN(n6591) );
  OR2_X1 U8980 ( .A1(n13693), .A2(n9011), .ZN(n6592) );
  INV_X1 U8981 ( .A(n11835), .ZN(n7588) );
  INV_X1 U8982 ( .A(n11951), .ZN(n7193) );
  NAND2_X1 U8983 ( .A1(n9637), .A2(n9137), .ZN(n9633) );
  OR2_X1 U8984 ( .A1(n14982), .A2(n10794), .ZN(n6593) );
  NOR2_X1 U8985 ( .A1(n14010), .A2(n7585), .ZN(n7584) );
  OR2_X1 U8986 ( .A1(n13566), .A2(n13715), .ZN(n6594) );
  NAND2_X1 U8987 ( .A1(n8652), .A2(n7058), .ZN(n6595) );
  NAND2_X1 U8988 ( .A1(n14206), .A2(n13928), .ZN(n6596) );
  INV_X1 U8989 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7514) );
  AND2_X1 U8990 ( .A1(n7433), .A2(n9811), .ZN(n6597) );
  NAND2_X1 U8991 ( .A1(n12606), .A2(n12391), .ZN(n6598) );
  AND3_X1 U8992 ( .A1(n7663), .A2(n7662), .A3(n7661), .ZN(n6599) );
  AND2_X1 U8993 ( .A1(n8848), .A2(n8847), .ZN(n6600) );
  OR2_X1 U8994 ( .A1(n14329), .A2(n13929), .ZN(n6601) );
  OR2_X1 U8995 ( .A1(n11549), .A2(n11543), .ZN(n6602) );
  OR2_X1 U8996 ( .A1(n11607), .A2(n13804), .ZN(n6603) );
  OR2_X1 U8997 ( .A1(n12660), .A2(n12661), .ZN(n6604) );
  AND2_X1 U8998 ( .A1(n8941), .A2(n8940), .ZN(n6605) );
  AND2_X1 U8999 ( .A1(n7969), .A2(n6888), .ZN(n6606) );
  INV_X1 U9000 ( .A(n12168), .ZN(n6976) );
  INV_X1 U9001 ( .A(n13740), .ZN(n7357) );
  NOR2_X1 U9002 ( .A1(n14592), .A2(n12604), .ZN(n6607) );
  OR2_X1 U9003 ( .A1(n13357), .A2(n8233), .ZN(n6608) );
  INV_X1 U9004 ( .A(n10036), .ZN(n6946) );
  INV_X1 U9005 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14399) );
  INV_X1 U9006 ( .A(n7873), .ZN(n7481) );
  AND2_X1 U9007 ( .A1(n12519), .A2(n12427), .ZN(n6609) );
  INV_X1 U9008 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7278) );
  NAND2_X1 U9009 ( .A1(n8471), .A2(n8470), .ZN(n13868) );
  OR2_X1 U9010 ( .A1(n9257), .A2(n9256), .ZN(n14962) );
  AOI21_X1 U9011 ( .B1(n9103), .B2(n10158), .A(n7321), .ZN(n7320) );
  OR2_X1 U9012 ( .A1(n12620), .A2(n12621), .ZN(n6610) );
  OR3_X1 U9013 ( .A1(n8525), .A2(P1_IR_REG_19__SCAN_IN), .A3(n6595), .ZN(n6611) );
  NAND2_X1 U9014 ( .A1(n8505), .A2(n8504), .ZN(n14206) );
  OR2_X1 U9015 ( .A1(n13647), .A2(n13219), .ZN(n6612) );
  OR2_X1 U9016 ( .A1(n14461), .A2(n14460), .ZN(n6613) );
  OR2_X1 U9017 ( .A1(n13390), .A2(n13696), .ZN(n6614) );
  INV_X1 U9018 ( .A(n7265), .ZN(n7264) );
  AND2_X1 U9019 ( .A1(n9137), .A2(n7531), .ZN(n6615) );
  AND2_X1 U9020 ( .A1(n13715), .A2(n8217), .ZN(n6616) );
  AND2_X1 U9021 ( .A1(n11479), .A2(n11438), .ZN(n6617) );
  AND2_X1 U9022 ( .A1(n6924), .A2(n6923), .ZN(n6618) );
  INV_X1 U9023 ( .A(n8453), .ZN(n7200) );
  NAND2_X1 U9024 ( .A1(n8550), .A2(n8549), .ZN(n14292) );
  AND2_X1 U9025 ( .A1(n9410), .A2(n9374), .ZN(n6619) );
  AND2_X1 U9026 ( .A1(n9793), .A2(n9792), .ZN(n6620) );
  AND2_X1 U9027 ( .A1(n8824), .A2(n8823), .ZN(n6621) );
  AND2_X1 U9028 ( .A1(n6568), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6622) );
  OR2_X1 U9029 ( .A1(n6653), .A2(n8804), .ZN(n6623) );
  AND2_X1 U9030 ( .A1(n13620), .A2(n13214), .ZN(n6624) );
  OR2_X1 U9031 ( .A1(n8993), .A2(n8992), .ZN(n6625) );
  INV_X1 U9032 ( .A(n6954), .ZN(n13343) );
  NAND2_X1 U9033 ( .A1(n6952), .A2(n6951), .ZN(n6954) );
  OR2_X1 U9034 ( .A1(n8716), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n6626) );
  AND2_X1 U9035 ( .A1(n12754), .A2(n6960), .ZN(n6627) );
  AND2_X1 U9036 ( .A1(n7027), .A2(n7026), .ZN(n6628) );
  AND2_X1 U9037 ( .A1(n6751), .A2(n12781), .ZN(n6629) );
  INV_X1 U9038 ( .A(n12579), .ZN(n13036) );
  NOR2_X1 U9039 ( .A1(n13647), .A2(n13177), .ZN(n6630) );
  OR2_X1 U9040 ( .A1(n8827), .A2(n6621), .ZN(n6631) );
  NAND2_X1 U9041 ( .A1(n13696), .A2(n13213), .ZN(n6632) );
  OR2_X1 U9042 ( .A1(n10548), .A2(n15120), .ZN(n6633) );
  AND2_X1 U9043 ( .A1(n10913), .A2(n10966), .ZN(n6634) );
  NAND2_X1 U9044 ( .A1(n11207), .A2(n11206), .ZN(n6635) );
  AND2_X1 U9045 ( .A1(n11250), .A2(n13227), .ZN(n6636) );
  AND2_X1 U9046 ( .A1(n12304), .A2(n12297), .ZN(n6637) );
  AND2_X1 U9047 ( .A1(n7235), .A2(n7240), .ZN(n6638) );
  AND2_X1 U9048 ( .A1(n12347), .A2(n13818), .ZN(n6639) );
  AND2_X1 U9049 ( .A1(n9056), .A2(n7509), .ZN(n6640) );
  OR2_X1 U9050 ( .A1(n14398), .A2(n7278), .ZN(n6641) );
  NAND2_X1 U9051 ( .A1(n6906), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6642) );
  AND2_X1 U9052 ( .A1(n8791), .A2(n8790), .ZN(n6643) );
  INV_X1 U9053 ( .A(n8665), .ZN(n8713) );
  OR2_X1 U9054 ( .A1(n13406), .A2(n13620), .ZN(n13390) );
  INV_X1 U9055 ( .A(n13390), .ZN(n6952) );
  INV_X1 U9056 ( .A(n6985), .ZN(n6984) );
  NOR2_X1 U9057 ( .A1(n12391), .A2(n12606), .ZN(n6985) );
  NOR2_X1 U9058 ( .A1(n13651), .A2(n13140), .ZN(n6644) );
  NOR2_X1 U9059 ( .A1(n13715), .A2(n13519), .ZN(n6645) );
  NOR2_X1 U9060 ( .A1(n13636), .A2(n13217), .ZN(n6646) );
  NOR2_X1 U9061 ( .A1(n13689), .A2(n13189), .ZN(n6647) );
  NOR2_X1 U9062 ( .A1(n14266), .A2(n14093), .ZN(n6648) );
  NOR2_X1 U9063 ( .A1(n8706), .A2(n14041), .ZN(n6649) );
  INV_X1 U9064 ( .A(n8347), .ZN(n8581) );
  INV_X1 U9065 ( .A(n7366), .ZN(n7365) );
  NAND2_X1 U9066 ( .A1(n12252), .A2(n12245), .ZN(n7366) );
  INV_X1 U9067 ( .A(n7203), .ZN(n7202) );
  NOR2_X1 U9068 ( .A1(n11607), .A2(n13949), .ZN(n7203) );
  INV_X1 U9069 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7996) );
  INV_X1 U9070 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U9071 ( .A1(n9047), .A2(n7512), .ZN(n6651) );
  AND2_X1 U9072 ( .A1(n8931), .A2(n8930), .ZN(n6652) );
  INV_X1 U9073 ( .A(n8388), .ZN(n7180) );
  NAND2_X1 U9074 ( .A1(n7880), .A2(n7879), .ZN(n11575) );
  AND2_X1 U9075 ( .A1(n8801), .A2(n8800), .ZN(n6653) );
  AND2_X1 U9076 ( .A1(n7875), .A2(n9915), .ZN(n6654) );
  NOR2_X1 U9077 ( .A1(n14292), .A2(n13785), .ZN(n6655) );
  XOR2_X1 U9078 ( .A(n7685), .B(n7683), .Z(n6656) );
  OR2_X1 U9079 ( .A1(n8939), .A2(n8938), .ZN(n6657) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9869) );
  INV_X1 U9081 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9895) );
  OR2_X1 U9082 ( .A1(n14400), .A2(n14399), .ZN(n6658) );
  AND2_X1 U9083 ( .A1(n7840), .A2(n15445), .ZN(n6659) );
  AND2_X1 U9084 ( .A1(n7891), .A2(SI_13_), .ZN(n6660) );
  NAND2_X1 U9085 ( .A1(n9605), .A2(n9604), .ZN(n6661) );
  NAND2_X1 U9086 ( .A1(n12314), .A2(n13872), .ZN(n13759) );
  NAND2_X1 U9087 ( .A1(n12459), .A2(n12752), .ZN(n6662) );
  INV_X1 U9088 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U9089 ( .A1(n11702), .A2(n11704), .ZN(n7111) );
  NOR2_X1 U9090 ( .A1(n11869), .A2(n11868), .ZN(n6663) );
  AND2_X1 U9091 ( .A1(n12265), .A2(n12264), .ZN(n13833) );
  NAND2_X1 U9092 ( .A1(n8754), .A2(n8756), .ZN(n7411) );
  INV_X1 U9093 ( .A(n7095), .ZN(n7094) );
  AND2_X1 U9094 ( .A1(n7097), .A2(n7096), .ZN(n7095) );
  INV_X1 U9095 ( .A(n7247), .ZN(n7246) );
  NAND2_X1 U9096 ( .A1(n8213), .A2(n7248), .ZN(n7247) );
  AND2_X1 U9097 ( .A1(n11845), .A2(n11835), .ZN(n6664) );
  AND2_X1 U9098 ( .A1(n9709), .A2(n9708), .ZN(n6665) );
  OR2_X1 U9099 ( .A1(n12383), .A2(n12869), .ZN(n6666) );
  OR2_X1 U9100 ( .A1(n6600), .A2(n8850), .ZN(n6667) );
  INV_X1 U9101 ( .A(n13347), .ZN(n13689) );
  NAND2_X1 U9102 ( .A1(n8144), .A2(n8143), .ZN(n13347) );
  OR2_X1 U9103 ( .A1(n8838), .A2(n8840), .ZN(n6668) );
  AND2_X1 U9104 ( .A1(n12948), .A2(n15168), .ZN(n6669) );
  AND2_X1 U9105 ( .A1(n7188), .A2(n6596), .ZN(n6670) );
  OR2_X1 U9106 ( .A1(n7381), .A2(n7730), .ZN(n6671) );
  INV_X1 U9107 ( .A(n8708), .ZN(n7585) );
  INV_X1 U9108 ( .A(n7260), .ZN(n7259) );
  NOR2_X1 U9109 ( .A1(n13504), .A2(n13517), .ZN(n7260) );
  INV_X1 U9110 ( .A(n7348), .ZN(n7346) );
  NOR2_X1 U9111 ( .A1(n11368), .A2(n11369), .ZN(n7348) );
  OR2_X1 U9112 ( .A1(n8893), .A2(n8895), .ZN(n6672) );
  OR2_X1 U9113 ( .A1(n7539), .A2(n8894), .ZN(n6673) );
  OR2_X1 U9114 ( .A1(n7533), .A2(n8839), .ZN(n6674) );
  OR2_X1 U9115 ( .A1(n11819), .A2(n11821), .ZN(n6675) );
  AND2_X1 U9116 ( .A1(n8298), .A2(n7590), .ZN(n6676) );
  AND2_X1 U9117 ( .A1(n7100), .A2(n7101), .ZN(n6677) );
  OR2_X1 U9118 ( .A1(n11797), .A2(n7052), .ZN(n6678) );
  AND2_X1 U9119 ( .A1(n7419), .A2(n7596), .ZN(n6679) );
  NAND2_X1 U9120 ( .A1(n8910), .A2(n8911), .ZN(n6680) );
  INV_X1 U9121 ( .A(n7700), .ZN(n7473) );
  INV_X1 U9122 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8313) );
  INV_X1 U9123 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7058) );
  AND2_X1 U9124 ( .A1(n7934), .A2(n7914), .ZN(n7932) );
  INV_X1 U9125 ( .A(n7245), .ZN(n7237) );
  OR2_X1 U9126 ( .A1(n8216), .A2(n9013), .ZN(n7245) );
  OR2_X1 U9127 ( .A1(n8934), .A2(n6652), .ZN(n6681) );
  INV_X1 U9128 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U9129 ( .A1(n9902), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6948) );
  INV_X1 U9130 ( .A(n7108), .ZN(n7107) );
  OR2_X1 U9131 ( .A1(n12396), .A2(n7109), .ZN(n7108) );
  OR2_X1 U9132 ( .A1(n7357), .A2(n7355), .ZN(n6682) );
  INV_X2 U9133 ( .A(n7660), .ZN(n7950) );
  INV_X1 U9134 ( .A(n10868), .ZN(n6776) );
  INV_X1 U9135 ( .A(n14208), .ZN(n7183) );
  NAND2_X1 U9136 ( .A1(n8073), .A2(n8072), .ZN(n13408) );
  INV_X1 U9137 ( .A(n13408), .ZN(n6939) );
  XNOR2_X1 U9138 ( .A(n10276), .B(n10393), .ZN(n9018) );
  INV_X1 U9139 ( .A(n14276), .ZN(n6864) );
  OR2_X1 U9140 ( .A1(n10315), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6683) );
  INV_X1 U9141 ( .A(n13812), .ZN(n7360) );
  AND2_X1 U9142 ( .A1(n12750), .A2(n15043), .ZN(n6684) );
  INV_X1 U9143 ( .A(n7621), .ZN(n7960) );
  NOR2_X1 U9144 ( .A1(n14129), .A2(n7578), .ZN(n7577) );
  NOR2_X1 U9145 ( .A1(n14176), .A2(n14298), .ZN(n14145) );
  INV_X1 U9146 ( .A(n12792), .ZN(n12765) );
  NAND2_X1 U9147 ( .A1(n9550), .A2(n9549), .ZN(n12792) );
  NAND2_X1 U9148 ( .A1(n7598), .A2(n7973), .ZN(n8256) );
  AND2_X1 U9149 ( .A1(n12415), .A2(n12884), .ZN(n6685) );
  NOR2_X1 U9150 ( .A1(n15060), .A2(n15061), .ZN(n6686) );
  NAND2_X1 U9151 ( .A1(n14145), .A2(n6867), .ZN(n6868) );
  OR2_X1 U9152 ( .A1(n13032), .A2(n13001), .ZN(n6687) );
  INV_X1 U9153 ( .A(n6935), .ZN(n13483) );
  NOR2_X1 U9154 ( .A1(n13506), .A2(n13651), .ZN(n6935) );
  OR2_X1 U9155 ( .A1(n13032), .A2(n13074), .ZN(n6688) );
  INV_X1 U9156 ( .A(n8660), .ZN(n7568) );
  INV_X1 U9157 ( .A(n9379), .ZN(n7321) );
  AND2_X1 U9158 ( .A1(n7570), .A2(n6603), .ZN(n6689) );
  INV_X1 U9159 ( .A(n7257), .ZN(n7256) );
  AOI21_X1 U9160 ( .B1(n6579), .B2(n8219), .A(n6644), .ZN(n7257) );
  OR2_X1 U9161 ( .A1(n11830), .A2(n11828), .ZN(n6690) );
  INV_X1 U9162 ( .A(n9616), .ZN(n6965) );
  NAND2_X1 U9163 ( .A1(n10387), .A2(n10386), .ZN(n14929) );
  AND2_X2 U9164 ( .A1(n8751), .A2(n10719), .ZN(n14796) );
  OR2_X1 U9165 ( .A1(n9836), .A2(n9830), .ZN(n13202) );
  INV_X1 U9166 ( .A(n14803), .ZN(n14800) );
  OR2_X1 U9167 ( .A1(n14908), .A2(n8178), .ZN(n6691) );
  NAND2_X1 U9168 ( .A1(n9833), .A2(n13573), .ZN(n14638) );
  INV_X1 U9169 ( .A(n7198), .ZN(n7197) );
  NOR2_X1 U9170 ( .A1(n14519), .A2(n7203), .ZN(n7198) );
  INV_X1 U9171 ( .A(n6981), .ZN(n6980) );
  NAND2_X1 U9172 ( .A1(n11270), .A2(n6576), .ZN(n6957) );
  AND2_X1 U9173 ( .A1(n10760), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6692) );
  INV_X2 U9174 ( .A(n8363), .ZN(n8668) );
  AND2_X1 U9175 ( .A1(n14514), .A2(n6873), .ZN(n6693) );
  AND2_X1 U9176 ( .A1(n7332), .A2(n7331), .ZN(n6694) );
  AND2_X1 U9177 ( .A1(n7009), .A2(n6590), .ZN(n6695) );
  AND2_X1 U9178 ( .A1(n10961), .A2(n9739), .ZN(n6696) );
  INV_X1 U9179 ( .A(n9483), .ZN(n7315) );
  INV_X1 U9180 ( .A(n7146), .ZN(n10047) );
  INV_X1 U9181 ( .A(n6555), .ZN(n12180) );
  INV_X1 U9182 ( .A(n14910), .ZN(n6936) );
  NAND2_X1 U9183 ( .A1(n7864), .A2(n7863), .ZN(n13578) );
  INV_X1 U9184 ( .A(n13578), .ZN(n6955) );
  AND2_X1 U9185 ( .A1(n10391), .A2(n11062), .ZN(n6697) );
  INV_X1 U9186 ( .A(n12133), .ZN(n12143) );
  AND2_X1 U9187 ( .A1(n12190), .A2(n12014), .ZN(n12133) );
  NOR2_X1 U9188 ( .A1(n8356), .A2(n14378), .ZN(n6698) );
  NAND2_X1 U9189 ( .A1(n7899), .A2(n7898), .ZN(n13718) );
  INV_X1 U9190 ( .A(n13718), .ZN(n7242) );
  AND2_X1 U9191 ( .A1(n13984), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U9192 ( .A1(n8392), .A2(n8391), .ZN(n11799) );
  INV_X1 U9193 ( .A(n11799), .ZN(n6869) );
  AND2_X1 U9194 ( .A1(n14725), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6700) );
  INV_X1 U9195 ( .A(n15104), .ZN(n6796) );
  INV_X1 U9196 ( .A(n9945), .ZN(n6944) );
  OR2_X1 U9197 ( .A1(n12005), .A2(n13080), .ZN(n6701) );
  INV_X1 U9198 ( .A(n7707), .ZN(n7381) );
  INV_X1 U9199 ( .A(n11760), .ZN(n13992) );
  INV_X1 U9200 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n6736) );
  INV_X1 U9201 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7276) );
  INV_X1 U9202 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6791) );
  INV_X1 U9203 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6742) );
  INV_X1 U9204 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6826) );
  AOI21_X1 U9205 ( .B1(n8246), .B2(n13540), .A(n8245), .ZN(n13322) );
  AOI211_X1 U9206 ( .C1(n13540), .C2(n13389), .A(n13388), .B(n13387), .ZN(
        n13622) );
  NAND2_X2 U9207 ( .A1(n6551), .A2(P3_U3151), .ZN(n13092) );
  OAI21_X1 U9208 ( .B1(n11147), .B2(n7082), .A(n7080), .ZN(n11465) );
  NAND2_X1 U9209 ( .A1(n12529), .A2(n12528), .ZN(n12527) );
  INV_X1 U9210 ( .A(n12473), .ZN(n6703) );
  NAND2_X1 U9211 ( .A1(n11467), .A2(n11466), .ZN(n11507) );
  NAND2_X1 U9212 ( .A1(n12438), .A2(n12437), .ZN(n7067) );
  OAI21_X1 U9213 ( .B1(n12582), .B2(n12594), .A(n6704), .ZN(P3_U3180) );
  NAND2_X1 U9214 ( .A1(n7068), .A2(n7069), .ZN(n12529) );
  NAND2_X1 U9215 ( .A1(n12412), .A2(n12411), .ZN(n12565) );
  NAND2_X1 U9216 ( .A1(n9416), .A2(n9417), .ZN(n9432) );
  NAND2_X1 U9217 ( .A1(n7099), .A2(n7097), .ZN(n7103) );
  NAND2_X1 U9218 ( .A1(n13814), .A2(n12340), .ZN(n13910) );
  NAND2_X1 U9219 ( .A1(n13892), .A2(n6744), .ZN(n13801) );
  NOR2_X1 U9220 ( .A1(n7337), .A2(n10664), .ZN(n7334) );
  OR2_X1 U9221 ( .A1(n12145), .A2(n12143), .ZN(n7325) );
  XNOR2_X1 U9222 ( .A(n8157), .B(n8142), .ZN(n13732) );
  NAND2_X1 U9223 ( .A1(n8141), .A2(n8140), .ZN(n8157) );
  NAND2_X1 U9224 ( .A1(n6898), .A2(n6896), .ZN(n7860) );
  NAND2_X1 U9225 ( .A1(n7231), .A2(n7228), .ZN(P2_U3528) );
  NAND2_X1 U9226 ( .A1(n15104), .A2(n13018), .ZN(n12017) );
  NAND2_X2 U9227 ( .A1(n6986), .A2(n6987), .ZN(n15104) );
  NAND2_X1 U9228 ( .A1(n6859), .A2(n6904), .ZN(P2_U3496) );
  AOI21_X1 U9229 ( .B1(n12058), .B2(n12057), .A(n14598), .ZN(n12067) );
  OAI21_X1 U9230 ( .B1(n12116), .B2(n12115), .A(n12822), .ZN(n12118) );
  AOI211_X1 U9231 ( .C1(n12086), .C2(n12085), .A(n12896), .B(n6571), .ZN(
        n12098) );
  AOI211_X1 U9232 ( .C1(n12143), .C2(n12035), .A(n12040), .B(n12034), .ZN(
        n12045) );
  NAND2_X1 U9233 ( .A1(n10678), .A2(n10677), .ZN(n10676) );
  NAND2_X1 U9234 ( .A1(n10706), .A2(n11934), .ZN(n10708) );
  OAI21_X2 U9235 ( .B1(n14186), .B2(n8692), .A(n8693), .ZN(n14181) );
  NAND2_X1 U9236 ( .A1(n12914), .A2(n12081), .ZN(n12902) );
  NAND2_X1 U9237 ( .A1(n15096), .A2(n12021), .ZN(n11087) );
  NAND2_X1 U9238 ( .A1(n9224), .A2(n12031), .ZN(n10919) );
  NAND2_X1 U9239 ( .A1(n14630), .A2(n9771), .ZN(n13136) );
  NAND2_X1 U9240 ( .A1(n10220), .A2(n9705), .ZN(n10323) );
  INV_X1 U9241 ( .A(n10963), .ZN(n9736) );
  NAND2_X1 U9242 ( .A1(n8674), .A2(n8673), .ZN(n10706) );
  NAND2_X1 U9243 ( .A1(n7436), .A2(n6706), .ZN(n10160) );
  NAND2_X1 U9244 ( .A1(n9193), .A2(n12017), .ZN(n10617) );
  NAND2_X2 U9245 ( .A1(n11763), .A2(n11764), .ZN(n11759) );
  NAND2_X2 U9246 ( .A1(n13960), .A2(n11023), .ZN(n11763) );
  NAND2_X1 U9247 ( .A1(n11031), .A2(n8679), .ZN(n11048) );
  NAND2_X1 U9248 ( .A1(n11156), .A2(n8681), .ZN(n11303) );
  NOR2_X1 U9249 ( .A1(n12943), .A2(n6971), .ZN(n13027) );
  NAND2_X1 U9250 ( .A1(n10439), .A2(n10440), .ZN(n10438) );
  INV_X1 U9251 ( .A(n11560), .ZN(n9759) );
  NAND2_X1 U9252 ( .A1(n6970), .A2(n6968), .ZN(P3_U3487) );
  NAND2_X1 U9253 ( .A1(n6726), .A2(n8998), .ZN(n9035) );
  AOI21_X1 U9254 ( .B1(n6756), .B2(n8975), .A(n9010), .ZN(n8991) );
  AOI21_X1 U9255 ( .B1(n8833), .B2(n8832), .A(n8830), .ZN(n8831) );
  NAND2_X1 U9256 ( .A1(n6717), .A2(n6716), .ZN(n7600) );
  AOI21_X1 U9257 ( .B1(n8950), .B2(n8945), .A(n8949), .ZN(n8951) );
  OAI21_X1 U9258 ( .B1(n7541), .B2(n8821), .A(n7540), .ZN(n8833) );
  OR2_X1 U9259 ( .A1(n7691), .A2(n7658), .ZN(n7664) );
  NAND2_X1 U9260 ( .A1(n7544), .A2(n6583), .ZN(n8797) );
  INV_X1 U9261 ( .A(n8797), .ZN(n6762) );
  INV_X1 U9262 ( .A(n8783), .ZN(n6711) );
  INV_X1 U9263 ( .A(n8925), .ZN(n6758) );
  AOI22_X1 U9264 ( .A1(n13578), .A2(n8946), .B1(n13224), .B2(n8943), .ZN(n8843) );
  NAND2_X1 U9265 ( .A1(n6710), .A2(n6709), .ZN(n8780) );
  INV_X1 U9266 ( .A(n8777), .ZN(n6709) );
  NAND2_X1 U9267 ( .A1(n8779), .A2(n8778), .ZN(n6710) );
  NAND2_X1 U9268 ( .A1(n6712), .A2(n6711), .ZN(n8787) );
  NAND2_X1 U9269 ( .A1(n8785), .A2(n8784), .ZN(n6712) );
  NAND2_X1 U9270 ( .A1(n6829), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6994) );
  XNOR2_X1 U9271 ( .A(n12621), .B(n12620), .ZN(n15005) );
  NOR2_X1 U9272 ( .A1(n12693), .A2(n6788), .ZN(n12698) );
  XNOR2_X1 U9273 ( .A(n10813), .B(n10814), .ZN(n10362) );
  NAND3_X1 U9274 ( .A1(n8952), .A2(n6650), .A3(n8953), .ZN(n6756) );
  INV_X1 U9275 ( .A(n8778), .ZN(n6716) );
  INV_X1 U9276 ( .A(n8779), .ZN(n6717) );
  NAND2_X1 U9277 ( .A1(n7759), .A2(n7758), .ZN(n11130) );
  NAND2_X1 U9278 ( .A1(n7855), .A2(n7854), .ZN(n11483) );
  NAND2_X1 U9279 ( .A1(n13425), .A2(n8067), .ZN(n13399) );
  NOR2_X1 U9280 ( .A1(n6853), .A2(n6671), .ZN(n6852) );
  INV_X1 U9281 ( .A(n7027), .ZN(n7021) );
  OAI21_X2 U9282 ( .B1(n8126), .B2(n8125), .A(n8127), .ZN(n8139) );
  NAND2_X1 U9283 ( .A1(n6908), .A2(n8111), .ZN(n8126) );
  NAND2_X1 U9284 ( .A1(n8964), .A2(n8963), .ZN(n8978) );
  OAI21_X2 U9285 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8961) );
  NAND2_X1 U9286 ( .A1(n6719), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U9287 ( .A1(n13990), .A2(n14753), .ZN(n6719) );
  NAND2_X1 U9288 ( .A1(n10953), .A2(n10954), .ZN(n13977) );
  NOR2_X1 U9289 ( .A1(n14751), .A2(n15249), .ZN(n14750) );
  XNOR2_X1 U9290 ( .A(n13985), .B(n14756), .ZN(n14751) );
  AOI21_X2 U9291 ( .B1(n10760), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10754), .ZN(
        n10757) );
  NAND2_X1 U9292 ( .A1(n10603), .A2(n10374), .ZN(n7128) );
  INV_X1 U9293 ( .A(n14971), .ZN(n6772) );
  NOR2_X1 U9294 ( .A1(n9324), .A2(n11383), .ZN(n11538) );
  NAND2_X1 U9295 ( .A1(n10310), .A2(n6683), .ZN(n10311) );
  NOR2_X1 U9296 ( .A1(n12615), .A2(n15013), .ZN(n12616) );
  NOR2_X1 U9297 ( .A1(n14961), .A2(n14960), .ZN(n14959) );
  NAND2_X1 U9298 ( .A1(n6722), .A2(n7542), .ZN(n8810) );
  INV_X1 U9299 ( .A(n8833), .ZN(n6725) );
  INV_X1 U9300 ( .A(n7411), .ZN(n8759) );
  OAI21_X2 U9301 ( .B1(n8991), .B2(n8990), .A(n6625), .ZN(n6726) );
  NOR2_X1 U9302 ( .A1(n12137), .A2(n12136), .ZN(n12142) );
  AOI21_X2 U9303 ( .B1(n6729), .B2(n6728), .A(n14660), .ZN(n14663) );
  INV_X1 U9304 ( .A(n14652), .ZN(n6793) );
  AND2_X2 U9305 ( .A1(n6731), .A2(n6730), .ZN(n14508) );
  NAND2_X1 U9306 ( .A1(n14464), .A2(n14465), .ZN(n6730) );
  INV_X1 U9307 ( .A(n14503), .ZN(n6731) );
  INV_X1 U9308 ( .A(n8335), .ZN(n11934) );
  NAND2_X1 U9309 ( .A1(n6834), .A2(n7589), .ZN(n8312) );
  NAND2_X1 U9310 ( .A1(n11093), .A2(n9587), .ZN(n15085) );
  OAI21_X1 U9311 ( .B1(n12766), .B2(n13029), .A(n12748), .ZN(n9622) );
  NAND2_X1 U9312 ( .A1(n6737), .A2(n9602), .ZN(n14599) );
  AOI21_X1 U9313 ( .B1(n11282), .B2(n9598), .A(n9597), .ZN(n15042) );
  OAI21_X1 U9314 ( .B1(n14611), .B2(n12383), .A(n12386), .ZN(n9691) );
  OAI22_X2 U9315 ( .A1(n12923), .A2(n9608), .B1(n12930), .B2(n12602), .ZN(
        n12910) );
  NAND2_X1 U9316 ( .A1(n15028), .A2(n15027), .ZN(n6737) );
  NAND3_X1 U9317 ( .A1(n7028), .A2(n11900), .A3(n6738), .ZN(n7016) );
  NAND2_X1 U9318 ( .A1(n11918), .A2(n11917), .ZN(n7028) );
  NAND2_X1 U9319 ( .A1(n6811), .A2(n6642), .ZN(n7645) );
  OAI21_X2 U9320 ( .B1(n12910), .B2(n12915), .A(n9609), .ZN(n12897) );
  AOI21_X1 U9321 ( .B1(n14656), .B2(n14657), .A(P2_ADDR_REG_12__SCAN_IN), .ZN(
        n6739) );
  NAND2_X1 U9323 ( .A1(n14652), .A2(n14653), .ZN(n14470) );
  OAI21_X1 U9324 ( .B1(n7698), .B2(n7473), .A(n7709), .ZN(n7472) );
  NAND2_X1 U9325 ( .A1(n9212), .A2(n12026), .ZN(n15083) );
  XNOR2_X1 U9326 ( .A(n7521), .B(n12180), .ZN(n7520) );
  NAND2_X1 U9327 ( .A1(n12902), .A2(n12901), .ZN(n7524) );
  XNOR2_X1 U9328 ( .A(n6785), .B(n6784), .ZN(n12383) );
  OAI211_X1 U9329 ( .C1(n12386), .C2(n15038), .A(n6666), .B(n6743), .ZN(
        P3_U3204) );
  NOR2_X2 U9331 ( .A1(n10287), .A2(n10288), .ZN(n10524) );
  AND2_X1 U9332 ( .A1(n8331), .A2(n8330), .ZN(n6745) );
  NAND3_X1 U9333 ( .A1(n9046), .A2(n9045), .A3(n9218), .ZN(n9350) );
  AOI21_X2 U9334 ( .B1(n15085), .B2(n15084), .A(n9589), .ZN(n10922) );
  NAND2_X2 U9335 ( .A1(n9798), .A2(n9797), .ZN(n9801) );
  NAND3_X1 U9336 ( .A1(n10920), .A2(n9590), .A3(n9591), .ZN(n11282) );
  NAND2_X1 U9337 ( .A1(n7546), .A2(n7547), .ZN(n8939) );
  OAI21_X1 U9338 ( .B1(n8845), .B2(n8844), .A(n6667), .ZN(n6754) );
  AND2_X4 U9339 ( .A1(n11744), .A2(n6771), .ZN(n13528) );
  AND2_X2 U9340 ( .A1(n11732), .A2(n11406), .ZN(n11744) );
  AND4_X4 U9341 ( .A1(n8323), .A2(n8324), .A3(n8325), .A4(n8322), .ZN(n12212)
         );
  INV_X1 U9342 ( .A(n15084), .ZN(n15082) );
  NAND2_X1 U9343 ( .A1(n7476), .A2(n7474), .ZN(n7894) );
  OAI21_X1 U9344 ( .B1(n7472), .B2(n7700), .A(n7711), .ZN(n6882) );
  OAI21_X1 U9345 ( .B1(n8139), .B2(n11502), .A(n8138), .ZN(n8141) );
  NAND2_X1 U9346 ( .A1(n8939), .A2(n8938), .ZN(n6809) );
  OR2_X1 U9347 ( .A1(n6906), .A2(n8333), .ZN(n7657) );
  OAI21_X2 U9348 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(n8885) );
  NAND2_X1 U9349 ( .A1(n8922), .A2(n8921), .ZN(n8927) );
  NAND2_X2 U9350 ( .A1(n7628), .A2(n7627), .ZN(n7660) );
  NAND3_X1 U9351 ( .A1(n6755), .A2(n9006), .A3(n9005), .ZN(n9038) );
  NAND2_X1 U9352 ( .A1(n9001), .A2(n9000), .ZN(n6755) );
  NAND2_X1 U9353 ( .A1(n7538), .A2(n6673), .ZN(n8901) );
  NAND2_X1 U9354 ( .A1(n7548), .A2(n7549), .ZN(n8917) );
  NAND2_X1 U9355 ( .A1(n6763), .A2(n8761), .ZN(n8769) );
  NAND2_X1 U9356 ( .A1(n7553), .A2(n7552), .ZN(n8950) );
  NAND2_X1 U9357 ( .A1(n8780), .A2(n7600), .ZN(n8785) );
  NAND2_X1 U9358 ( .A1(n6759), .A2(n6758), .ZN(n6757) );
  NAND3_X1 U9359 ( .A1(n6657), .A2(n7555), .A3(n7554), .ZN(n7553) );
  NAND3_X1 U9360 ( .A1(n8929), .A2(n6757), .A3(n6681), .ZN(n7546) );
  AOI211_X1 U9361 ( .C1(n6564), .C2(n13292), .A(n9007), .B(n8999), .ZN(n9000)
         );
  NAND2_X1 U9362 ( .A1(n8927), .A2(n8926), .ZN(n6759) );
  NAND2_X1 U9363 ( .A1(n6762), .A2(n6761), .ZN(n8798) );
  AND2_X2 U9364 ( .A1(n6821), .A2(n6820), .ZN(n14656) );
  NOR2_X1 U9365 ( .A1(n14549), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14553) );
  NAND2_X1 U9366 ( .A1(n7379), .A2(n6852), .ZN(n7732) );
  NAND2_X1 U9367 ( .A1(n11263), .A2(n11262), .ZN(n11265) );
  AOI211_X1 U9368 ( .C1(n14905), .C2(n13605), .A(n13604), .B(n13603), .ZN(
        n13686) );
  NAND2_X1 U9369 ( .A1(n8755), .A2(n8196), .ZN(n8756) );
  NAND2_X1 U9370 ( .A1(n8757), .A2(n8758), .ZN(n6763) );
  NAND2_X1 U9371 ( .A1(n8810), .A2(n8811), .ZN(n8809) );
  NAND4_X4 U9372 ( .A1(n7635), .A2(n7633), .A3(n7632), .A4(n7634), .ZN(n8764)
         );
  NAND2_X1 U9373 ( .A1(n12874), .A2(n9613), .ZN(n12859) );
  NAND2_X1 U9374 ( .A1(n12816), .A2(n9619), .ZN(n12802) );
  NAND2_X1 U9375 ( .A1(n12801), .A2(n9620), .ZN(n12790) );
  NAND2_X1 U9376 ( .A1(n6765), .A2(n11431), .ZN(n11434) );
  NAND2_X1 U9377 ( .A1(n10221), .A2(n10222), .ZN(n10220) );
  NAND2_X1 U9378 ( .A1(n6764), .A2(n10733), .ZN(n10963) );
  NAND2_X1 U9379 ( .A1(n10735), .A2(n10734), .ZN(n6764) );
  NAND2_X1 U9380 ( .A1(n6964), .A2(n6963), .ZN(n12816) );
  NAND2_X1 U9381 ( .A1(n10257), .A2(n9713), .ZN(n10439) );
  NAND2_X1 U9382 ( .A1(n11332), .A2(n11430), .ZN(n6765) );
  INV_X1 U9383 ( .A(n7413), .ZN(n7412) );
  NAND2_X1 U9384 ( .A1(n12897), .A2(n12896), .ZN(n12895) );
  INV_X1 U9385 ( .A(n10362), .ZN(n6829) );
  INV_X1 U9386 ( .A(n15005), .ZN(n6787) );
  NOR2_X1 U9387 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  INV_X1 U9388 ( .A(n10359), .ZN(n6789) );
  AOI21_X1 U9389 ( .B1(n6590), .B2(n9265), .A(n14994), .ZN(n7007) );
  OAI21_X1 U9390 ( .B1(n10595), .B2(n10593), .A(n10594), .ZN(n10597) );
  CLKBUF_X2 U9391 ( .A(n8994), .Z(n6770) );
  OR2_X1 U9392 ( .A1(n12611), .A2(n15090), .ZN(n12031) );
  NAND2_X1 U9393 ( .A1(n9240), .A2(n12009), .ZN(n15077) );
  NAND2_X1 U9394 ( .A1(n7493), .A2(n7496), .ZN(n12764) );
  NOR2_X1 U9395 ( .A1(n12947), .A2(n6669), .ZN(n13030) );
  AOI21_X1 U9396 ( .B1(n15026), .B2(n12159), .A(n7490), .ZN(n7602) );
  OR2_X1 U9397 ( .A1(n7019), .A2(n7026), .ZN(n7018) );
  NAND2_X1 U9398 ( .A1(n7955), .A2(n6606), .ZN(n6886) );
  INV_X1 U9399 ( .A(n7645), .ZN(n7455) );
  INV_X1 U9400 ( .A(n11902), .ZN(n7030) );
  NAND2_X1 U9401 ( .A1(n10371), .A2(n10598), .ZN(n10603) );
  NAND2_X1 U9402 ( .A1(n9510), .A2(n9509), .ZN(n9124) );
  NAND2_X1 U9403 ( .A1(n9085), .A2(n9084), .ZN(n9251) );
  OAI211_X2 U9404 ( .C1(n7910), .C2(n7483), .A(n7934), .B(n6778), .ZN(n7955)
         );
  NAND2_X1 U9405 ( .A1(n7482), .A2(n7932), .ZN(n6778) );
  NAND2_X1 U9406 ( .A1(n7684), .A2(n7685), .ZN(n6779) );
  INV_X1 U9407 ( .A(n11914), .ZN(n7025) );
  NAND2_X1 U9408 ( .A1(n11157), .A2(n11158), .ZN(n11156) );
  NAND2_X1 U9409 ( .A1(n10770), .A2(n11940), .ZN(n10769) );
  INV_X2 U9410 ( .A(n12212), .ZN(n13960) );
  NAND2_X1 U9411 ( .A1(n8917), .A2(n8918), .ZN(n8916) );
  NAND2_X1 U9412 ( .A1(n8901), .A2(n8900), .ZN(n8905) );
  INV_X1 U9413 ( .A(n8937), .ZN(n6808) );
  NAND2_X1 U9414 ( .A1(n6643), .A2(n8792), .ZN(n7545) );
  NAND3_X1 U9415 ( .A1(n6782), .A2(n6781), .A3(n6672), .ZN(n7538) );
  NAND2_X1 U9416 ( .A1(n8888), .A2(n8887), .ZN(n6781) );
  NAND2_X1 U9417 ( .A1(n8884), .A2(n8883), .ZN(n6782) );
  NAND2_X1 U9418 ( .A1(n15097), .A2(n15109), .ZN(n15096) );
  NAND2_X1 U9419 ( .A1(n13031), .A2(n6688), .ZN(P3_U3454) );
  NAND2_X1 U9420 ( .A1(n12950), .A2(n6687), .ZN(P3_U3486) );
  NOR2_X2 U9421 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n9061) );
  NAND2_X1 U9422 ( .A1(n9291), .A2(n12048), .ZN(n15051) );
  NOR2_X1 U9423 ( .A1(n10511), .A2(n10341), .ZN(n10595) );
  OAI21_X1 U9424 ( .B1(n10373), .B2(n10361), .A(n10597), .ZN(n10813) );
  NAND2_X1 U9425 ( .A1(n6789), .A2(n10519), .ZN(n6828) );
  NAND2_X1 U9426 ( .A1(n14470), .A2(n14471), .ZN(n6821) );
  NOR2_X1 U9427 ( .A1(n14663), .A2(n14664), .ZN(n14662) );
  NOR2_X1 U9428 ( .A1(n14666), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n14488) );
  XNOR2_X2 U9429 ( .A(n9801), .B(n9799), .ZN(n13104) );
  INV_X1 U9430 ( .A(n6882), .ZN(n6881) );
  NAND2_X1 U9431 ( .A1(n9730), .A2(n9729), .ZN(n10735) );
  BUF_X4 U9432 ( .A(n8755), .Z(n11732) );
  NAND2_X1 U9433 ( .A1(n10259), .A2(n10258), .ZN(n10257) );
  NAND2_X1 U9434 ( .A1(n11192), .A2(n7437), .ZN(n11332) );
  NAND2_X1 U9435 ( .A1(n10311), .A2(n10312), .ZN(n10581) );
  NAND2_X1 U9436 ( .A1(n7557), .A2(n14371), .ZN(n6919) );
  NOR2_X1 U9437 ( .A1(n14717), .A2(n14718), .ZN(n14716) );
  INV_X1 U9438 ( .A(n6918), .ZN(n6917) );
  NAND2_X1 U9439 ( .A1(n6910), .A2(n13992), .ZN(n6909) );
  XNOR2_X1 U9440 ( .A(n13988), .B(n13987), .ZN(n13989) );
  INV_X1 U9441 ( .A(n13989), .ZN(n13990) );
  AND2_X2 U9442 ( .A1(n6989), .A2(n9177), .ZN(n6986) );
  AOI21_X4 U9443 ( .B1(n12547), .B2(n12845), .A(n12425), .ZN(n12517) );
  NAND2_X1 U9444 ( .A1(n6799), .A2(n6798), .ZN(n8799) );
  INV_X1 U9445 ( .A(n8795), .ZN(n6798) );
  NAND2_X1 U9446 ( .A1(n8797), .A2(n8796), .ZN(n6799) );
  OAI211_X1 U9447 ( .C1(n9834), .C2(n7421), .A(n6800), .B(n6679), .ZN(P2_U3192) );
  NAND2_X1 U9448 ( .A1(n9834), .A2(n7420), .ZN(n6800) );
  XNOR2_X1 U9449 ( .A(n9796), .B(n9794), .ZN(n13165) );
  INV_X1 U9450 ( .A(n10163), .ZN(n7435) );
  NAND2_X1 U9451 ( .A1(n9615), .A2(n6966), .ZN(n6964) );
  NOR2_X1 U9452 ( .A1(n12162), .A2(n9583), .ZN(n9584) );
  XNOR2_X2 U9453 ( .A(n9166), .B(n9165), .ZN(n12380) );
  NAND2_X1 U9454 ( .A1(n7297), .A2(n7298), .ZN(n9101) );
  NAND2_X1 U9455 ( .A1(n7518), .A2(n7516), .ZN(n7515) );
  AND2_X1 U9456 ( .A1(n11212), .A2(n11213), .ZN(n11214) );
  OR2_X1 U9457 ( .A1(n8413), .A2(n9905), .ZN(n8344) );
  NAND2_X1 U9458 ( .A1(n6830), .A2(n13912), .ZN(n13745) );
  MUX2_X1 U9459 ( .A(n9073), .B(n9189), .S(n6906), .Z(n7646) );
  XNOR2_X1 U9460 ( .A(n12218), .B(n12216), .ZN(n11715) );
  NAND2_X1 U9461 ( .A1(n7344), .A2(n7348), .ZN(n6847) );
  NAND2_X1 U9462 ( .A1(n8311), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6804) );
  INV_X1 U9463 ( .A(n6833), .ZN(n8308) );
  NAND2_X1 U9464 ( .A1(n8685), .A2(n8684), .ZN(n11646) );
  NAND2_X1 U9465 ( .A1(n7592), .A2(n7591), .ZN(n14059) );
  NAND2_X1 U9466 ( .A1(n6915), .A2(n11760), .ZN(n6914) );
  AND2_X1 U9467 ( .A1(n13336), .A2(n13341), .ZN(n6806) );
  INV_X1 U9468 ( .A(n13335), .ZN(n6807) );
  NOR2_X1 U9469 ( .A1(n13341), .A2(n7266), .ZN(n7265) );
  NAND2_X1 U9470 ( .A1(n8056), .A2(n8055), .ZN(n8086) );
  NAND2_X1 U9471 ( .A1(n6881), .A2(n6880), .ZN(n7735) );
  NAND2_X1 U9472 ( .A1(n8109), .A2(n8108), .ZN(n6908) );
  NOR3_X1 U9473 ( .A1(n11977), .A2(n11976), .A3(n11975), .ZN(n11983) );
  NAND3_X1 U9474 ( .A1(n8834), .A2(n7604), .A3(n6668), .ZN(n7532) );
  NAND2_X1 U9475 ( .A1(n6809), .A2(n6808), .ZN(n7555) );
  INV_X2 U9476 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U9477 ( .A1(n7997), .A2(n7996), .ZN(n8190) );
  NAND2_X1 U9478 ( .A1(n7532), .A2(n6674), .ZN(n8845) );
  NAND2_X1 U9479 ( .A1(n9903), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6811) );
  INV_X1 U9480 ( .A(n9580), .ZN(n15109) );
  NAND2_X2 U9481 ( .A1(n12808), .A2(n12121), .ZN(n12796) );
  INV_X2 U9482 ( .A(n9350), .ZN(n9047) );
  NAND2_X1 U9483 ( .A1(n7018), .A2(n7029), .ZN(n7017) );
  NAND2_X1 U9484 ( .A1(n6883), .A2(n7699), .ZN(n6880) );
  NAND2_X1 U9485 ( .A1(n7016), .A2(n7014), .ZN(n11932) );
  NAND2_X1 U9486 ( .A1(n8139), .A2(n11502), .ZN(n8140) );
  NAND2_X1 U9487 ( .A1(n8053), .A2(n8052), .ZN(n8056) );
  NAND2_X1 U9488 ( .A1(n7273), .A2(n14492), .ZN(n7272) );
  NOR2_X1 U9489 ( .A1(n14505), .A2(n14504), .ZN(n14503) );
  INV_X1 U9490 ( .A(n14670), .ZN(n6823) );
  OAI21_X2 U9491 ( .B1(n14469), .B2(n14832), .A(n14507), .ZN(n14652) );
  NAND2_X1 U9492 ( .A1(n10360), .A2(n6828), .ZN(n10511) );
  AOI21_X1 U9493 ( .B1(n6819), .B2(n12732), .A(n6818), .ZN(n12740) );
  XNOR2_X1 U9494 ( .A(n12726), .B(n12725), .ZN(n6819) );
  NOR2_X2 U9495 ( .A1(n14488), .A2(n14667), .ZN(n14670) );
  NAND2_X1 U9496 ( .A1(n15472), .A2(n15471), .ZN(n6824) );
  NAND2_X1 U9497 ( .A1(n9082), .A2(n9081), .ZN(n9237) );
  NAND2_X1 U9498 ( .A1(n9319), .A2(n9318), .ZN(n9321) );
  NAND2_X1 U9499 ( .A1(n7280), .A2(n9075), .ZN(n9200) );
  NAND2_X1 U9500 ( .A1(n9122), .A2(n9121), .ZN(n9510) );
  NAND2_X1 U9501 ( .A1(n7279), .A2(n9077), .ZN(n9209) );
  NAND2_X1 U9502 ( .A1(n7309), .A2(n9483), .ZN(n7313) );
  NAND2_X1 U9503 ( .A1(n9429), .A2(n9428), .ZN(n9431) );
  INV_X1 U9504 ( .A(n7317), .ZN(n7316) );
  NAND2_X1 U9505 ( .A1(n7283), .A2(n9126), .ZN(n9531) );
  OAI21_X1 U9506 ( .B1(n13991), .B2(n14719), .A(n6916), .ZN(n6915) );
  OAI21_X1 U9507 ( .B1(n8326), .B2(n7557), .A(n6919), .ZN(n6918) );
  NAND2_X1 U9508 ( .A1(n6827), .A2(n14438), .ZN(n14439) );
  NAND2_X1 U9509 ( .A1(n14670), .A2(n14671), .ZN(n7273) );
  AOI21_X2 U9510 ( .B1(n14847), .B2(n14482), .A(n14662), .ZN(n14486) );
  NAND2_X1 U9511 ( .A1(n14547), .A2(n14546), .ZN(n7270) );
  NAND2_X1 U9512 ( .A1(n7270), .A2(n14494), .ZN(n7269) );
  NAND2_X1 U9513 ( .A1(n7008), .A2(n7007), .ZN(n14992) );
  NAND2_X2 U9514 ( .A1(n13910), .A2(n13911), .ZN(n13909) );
  NAND2_X4 U9515 ( .A1(n7146), .A2(n14387), .ZN(n9853) );
  NAND2_X1 U9516 ( .A1(n8310), .A2(n8311), .ZN(n7146) );
  NAND2_X1 U9517 ( .A1(n7367), .A2(n6838), .ZN(n6835) );
  NAND2_X1 U9518 ( .A1(n6835), .A2(n6836), .ZN(n12275) );
  OAI21_X2 U9519 ( .B1(n11615), .B2(n7329), .A(n7327), .ZN(n12218) );
  NAND2_X2 U9520 ( .A1(n6846), .A2(n6845), .ZN(n11615) );
  NAND3_X1 U9521 ( .A1(n6848), .A2(n6847), .A3(n11444), .ZN(n6846) );
  INV_X1 U9522 ( .A(n10728), .ZN(n14766) );
  OAI21_X1 U9523 ( .B1(n10905), .B2(n11180), .A(n6854), .ZN(n11263) );
  NAND2_X1 U9524 ( .A1(n8083), .A2(n8082), .ZN(n13385) );
  NAND2_X1 U9525 ( .A1(n13488), .A2(n6861), .ZN(n8012) );
  NAND2_X2 U9526 ( .A1(n9940), .A2(n9902), .ZN(n8979) );
  XNOR2_X2 U9527 ( .A(n7639), .B(n7638), .ZN(n9945) );
  XNOR2_X2 U9528 ( .A(n7641), .B(n7640), .ZN(n13733) );
  INV_X1 U9529 ( .A(n6868), .ZN(n14123) );
  NAND2_X1 U9530 ( .A1(n14514), .A2(n6871), .ZN(n14203) );
  NAND2_X1 U9531 ( .A1(n14017), .A2(n6878), .ZN(n13996) );
  NAND2_X1 U9532 ( .A1(n14017), .A2(n6876), .ZN(n14002) );
  NAND2_X1 U9533 ( .A1(n14017), .A2(n8664), .ZN(n14018) );
  INV_X1 U9534 ( .A(n13996), .ZN(n14003) );
  NAND2_X1 U9535 ( .A1(n7735), .A2(n7734), .ZN(n7737) );
  INV_X1 U9536 ( .A(n7472), .ZN(n6883) );
  NAND2_X1 U9537 ( .A1(n7788), .A2(n6899), .ZN(n6898) );
  MUX2_X1 U9538 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6906), .Z(n6905) );
  OAI21_X2 U9539 ( .B1(n8036), .B2(n8035), .A(n8038), .ZN(n8053) );
  NOR2_X2 U9540 ( .A1(n14730), .A2(n6699), .ZN(n13973) );
  NOR2_X2 U9541 ( .A1(n6594), .A2(n14637), .ZN(n13531) );
  OAI211_X1 U9542 ( .C1(n13733), .C2(n6948), .A(n6945), .B(n6943), .ZN(n6942)
         );
  NAND3_X1 U9543 ( .A1(n13733), .A2(n9945), .A3(n6946), .ZN(n6945) );
  NAND2_X1 U9544 ( .A1(n7650), .A2(n6949), .ZN(n9916) );
  INV_X1 U9545 ( .A(n6957), .ZN(n11487) );
  INV_X1 U9546 ( .A(n6961), .ZN(n12760) );
  OAI21_X1 U9547 ( .B1(n14599), .B2(n6977), .A(n6975), .ZN(n9607) );
  INV_X1 U9548 ( .A(n6988), .ZN(n6987) );
  INV_X1 U9549 ( .A(n10614), .ZN(n13018) );
  NAND2_X2 U9550 ( .A1(n12017), .A2(n12018), .ZN(n13015) );
  AND2_X2 U9551 ( .A1(n12895), .A2(n9610), .ZN(n7597) );
  AOI21_X2 U9552 ( .B1(n7003), .B2(n7002), .A(n12659), .ZN(n12661) );
  NAND2_X1 U9553 ( .A1(n6590), .A2(n14973), .ZN(n7008) );
  INV_X1 U9554 ( .A(n7009), .ZN(n14972) );
  XNOR2_X2 U9555 ( .A(n7011), .B(n7010), .ZN(n10519) );
  AOI21_X1 U9557 ( .B1(n6628), .B2(n7025), .A(n7023), .ZN(n7022) );
  INV_X1 U9558 ( .A(n11913), .ZN(n7023) );
  NAND2_X1 U9559 ( .A1(n11886), .A2(n7034), .ZN(n7031) );
  NAND2_X1 U9560 ( .A1(n7031), .A2(n7032), .ZN(n11894) );
  NAND2_X1 U9561 ( .A1(n7038), .A2(n7039), .ZN(n11859) );
  NAND3_X1 U9562 ( .A1(n11837), .A2(n6664), .A3(n11836), .ZN(n7038) );
  NAND2_X1 U9563 ( .A1(n7452), .A2(n7046), .ZN(n7045) );
  NAND2_X1 U9564 ( .A1(n7050), .A2(n6678), .ZN(n11803) );
  NAND3_X1 U9565 ( .A1(n11794), .A2(n11793), .A3(n7051), .ZN(n7050) );
  NAND3_X1 U9566 ( .A1(n11818), .A2(n11817), .A3(n6675), .ZN(n7053) );
  NAND2_X1 U9567 ( .A1(n7053), .A2(n7054), .ZN(n11825) );
  NAND3_X1 U9568 ( .A1(n11827), .A2(n11826), .A3(n6690), .ZN(n7055) );
  NAND2_X1 U9569 ( .A1(n7055), .A2(n7056), .ZN(n11834) );
  NAND2_X1 U9570 ( .A1(n7059), .A2(n8417), .ZN(n8525) );
  NAND2_X1 U9571 ( .A1(n11908), .A2(n11929), .ZN(n7060) );
  OAI22_X1 U9572 ( .A1(n11809), .A2(n7063), .B1(n11808), .B2(n7064), .ZN(
        n11813) );
  INV_X1 U9573 ( .A(n11813), .ZN(n11816) );
  AND2_X2 U9574 ( .A1(n7511), .A2(n9047), .ZN(n9135) );
  NAND2_X1 U9575 ( .A1(n7067), .A2(n7065), .ZN(n12583) );
  NAND2_X1 U9576 ( .A1(n12565), .A2(n7071), .ZN(n7068) );
  NAND2_X2 U9577 ( .A1(n9179), .A2(n9902), .ZN(n9487) );
  OAI21_X1 U9578 ( .B1(n12517), .B2(n7094), .A(n7091), .ZN(n12461) );
  OAI21_X1 U9579 ( .B1(n12517), .B2(n7090), .A(n7087), .ZN(n7086) );
  NAND2_X1 U9580 ( .A1(n12517), .A2(n7104), .ZN(n7099) );
  OAI21_X1 U9581 ( .B1(n12517), .B2(n12428), .A(n7104), .ZN(n12494) );
  OAI21_X1 U9582 ( .B1(n11703), .B2(n7108), .A(n7105), .ZN(n12538) );
  INV_X1 U9583 ( .A(n7114), .ZN(n14970) );
  XNOR2_X1 U9584 ( .A(n10794), .B(n14982), .ZN(n14971) );
  NAND3_X1 U9585 ( .A1(n7118), .A2(n7116), .A3(n7115), .ZN(n12738) );
  NAND2_X1 U9586 ( .A1(n12704), .A2(n7120), .ZN(n7115) );
  OAI21_X1 U9587 ( .B1(n7122), .B2(n12735), .A(n7117), .ZN(n7116) );
  NAND2_X1 U9588 ( .A1(n7122), .A2(n7121), .ZN(n7117) );
  NAND3_X1 U9589 ( .A1(n7119), .A2(n7122), .A3(n12736), .ZN(n7118) );
  INV_X1 U9590 ( .A(n12704), .ZN(n7119) );
  AOI21_X2 U9591 ( .B1(n7125), .B2(n7126), .A(n7123), .ZN(n7122) );
  OAI21_X1 U9592 ( .B1(n12704), .B2(n7125), .A(n7126), .ZN(n7124) );
  INV_X1 U9593 ( .A(n12709), .ZN(n7126) );
  OR2_X2 U9594 ( .A1(n11542), .A2(n11541), .ZN(n7141) );
  NAND2_X1 U9595 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7142) );
  NAND3_X1 U9596 ( .A1(n8335), .A2(n11763), .A3(n7144), .ZN(n10711) );
  AND2_X1 U9597 ( .A1(n11770), .A2(n11771), .ZN(n8335) );
  NAND2_X1 U9598 ( .A1(n10047), .A2(n7145), .ZN(n9858) );
  INV_X1 U9599 ( .A(n6705), .ZN(n7145) );
  NAND2_X1 U9600 ( .A1(n11928), .A2(n7146), .ZN(n14210) );
  NOR2_X1 U9601 ( .A1(n10477), .A2(n7146), .ZN(n10478) );
  AOI21_X1 U9602 ( .B1(n10047), .B2(P1_STATE_REG_SCAN_IN), .A(n7148), .ZN(
        n7147) );
  NAND2_X1 U9603 ( .A1(n10679), .A2(n7149), .ZN(n7150) );
  AND2_X1 U9604 ( .A1(n11777), .A2(n8360), .ZN(n7149) );
  NAND2_X1 U9605 ( .A1(n14107), .A2(n8572), .ZN(n7156) );
  NAND2_X1 U9606 ( .A1(n14170), .A2(n6569), .ZN(n7157) );
  NAND2_X1 U9607 ( .A1(n7601), .A2(n7173), .ZN(n7171) );
  NAND2_X1 U9608 ( .A1(n7171), .A2(n7172), .ZN(n14024) );
  NAND2_X1 U9609 ( .A1(n11690), .A2(n6670), .ZN(n7181) );
  NAND2_X1 U9610 ( .A1(n7181), .A2(n7182), .ZN(n14188) );
  NOR2_X1 U9611 ( .A1(n12644), .A2(n12643), .ZN(n12671) );
  NOR2_X1 U9612 ( .A1(n11539), .A2(n11538), .ZN(n11542) );
  NOR2_X2 U9613 ( .A1(n12992), .A2(n12672), .ZN(n12704) );
  OR2_X2 U9614 ( .A1(n13718), .A2(n13565), .ZN(n13566) );
  NOR2_X2 U9615 ( .A1(n10268), .A2(n10273), .ZN(n10391) );
  AOI21_X1 U9616 ( .B1(n6563), .B2(n10120), .A(n7205), .ZN(n7688) );
  NAND2_X1 U9617 ( .A1(n11132), .A2(n7209), .ZN(n7206) );
  NAND2_X1 U9618 ( .A1(n7206), .A2(n7207), .ZN(n11181) );
  NAND2_X1 U9619 ( .A1(n11259), .A2(n7215), .ZN(n7212) );
  NAND2_X1 U9620 ( .A1(n7212), .A2(n7213), .ZN(n11488) );
  OAI21_X1 U9621 ( .B1(n11258), .B2(n7217), .A(n11345), .ZN(n7216) );
  INV_X1 U9622 ( .A(n11115), .ZN(n7253) );
  NAND2_X1 U9623 ( .A1(n8204), .A2(n7251), .ZN(n7250) );
  NAND2_X1 U9624 ( .A1(n13495), .A2(n6579), .ZN(n7255) );
  INV_X1 U9625 ( .A(n13357), .ZN(n7261) );
  NAND2_X1 U9626 ( .A1(n6608), .A2(n7267), .ZN(n13336) );
  OR2_X1 U9627 ( .A1(n13361), .A2(n9011), .ZN(n7267) );
  AND2_X2 U9628 ( .A1(n7272), .A2(n7271), .ZN(n14547) );
  NOR2_X2 U9631 ( .A1(n14449), .A2(n14450), .ZN(n14451) );
  NAND2_X1 U9632 ( .A1(n9200), .A2(n9199), .ZN(n7279) );
  NAND2_X1 U9633 ( .A1(n9074), .A2(n9178), .ZN(n7280) );
  NAND2_X1 U9634 ( .A1(n9521), .A2(n11643), .ZN(n7283) );
  NAND2_X1 U9635 ( .A1(n7283), .A2(n7281), .ZN(n7284) );
  NAND2_X1 U9636 ( .A1(n7284), .A2(n9127), .ZN(n9541) );
  NAND2_X1 U9637 ( .A1(n9443), .A2(n7288), .ZN(n7285) );
  NAND2_X1 U9638 ( .A1(n9331), .A2(n7300), .ZN(n7297) );
  NAND2_X1 U9639 ( .A1(n9286), .A2(n7306), .ZN(n7303) );
  NAND2_X1 U9640 ( .A1(n7303), .A2(n7304), .ZN(n9319) );
  NAND2_X1 U9641 ( .A1(n9118), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7309) );
  NAND2_X1 U9642 ( .A1(n7311), .A2(n7314), .ZN(n9486) );
  NAND2_X1 U9643 ( .A1(n9471), .A2(n9118), .ZN(n7311) );
  NAND2_X1 U9644 ( .A1(n7319), .A2(n7320), .ZN(n9382) );
  NAND2_X1 U9645 ( .A1(n9357), .A2(n9103), .ZN(n7319) );
  NAND3_X1 U9646 ( .A1(n7325), .A2(n12153), .A3(n6575), .ZN(n7324) );
  OAI21_X1 U9647 ( .B1(n10661), .B2(n7338), .A(n7340), .ZN(n7337) );
  NAND2_X1 U9648 ( .A1(n7334), .A2(n7336), .ZN(n7333) );
  NAND2_X1 U9649 ( .A1(n7335), .A2(n7336), .ZN(n10663) );
  INV_X1 U9650 ( .A(n7337), .ZN(n7335) );
  NAND2_X1 U9651 ( .A1(n7339), .A2(n10524), .ZN(n7336) );
  AND2_X1 U9652 ( .A1(n10525), .A2(n10526), .ZN(n7342) );
  NOR2_X1 U9653 ( .A1(n11226), .A2(n11214), .ZN(n11370) );
  OAI22_X1 U9654 ( .A1(n6589), .A2(n12212), .B1(n11023), .B2(n10522), .ZN(
        n10283) );
  AND2_X2 U9655 ( .A1(n10282), .A2(n10297), .ZN(n11448) );
  NAND2_X1 U9656 ( .A1(n13909), .A2(n7351), .ZN(n7350) );
  OAI211_X1 U9657 ( .C1(n13909), .C2(n6682), .A(n7352), .B(n7350), .ZN(n12376)
         );
  NAND2_X1 U9658 ( .A1(n7358), .A2(n7359), .ZN(n12339) );
  NAND2_X1 U9659 ( .A1(n12324), .A2(n7361), .ZN(n7358) );
  NAND2_X2 U9660 ( .A1(n13863), .A2(n13862), .ZN(n7367) );
  INV_X1 U9661 ( .A(n8525), .ZN(n7371) );
  XNOR2_X1 U9662 ( .A(n13234), .B(n7671), .ZN(n10183) );
  NAND2_X2 U9663 ( .A1(n7374), .A2(n7372), .ZN(n7671) );
  INV_X1 U9664 ( .A(n7373), .ZN(n7372) );
  OR2_X1 U9665 ( .A1(n7808), .A2(n6656), .ZN(n7374) );
  AND2_X2 U9666 ( .A1(n7621), .A2(n7375), .ZN(n8259) );
  AND3_X2 U9667 ( .A1(n7444), .A2(n7616), .A3(n7445), .ZN(n7621) );
  INV_X1 U9668 ( .A(n7690), .ZN(n7380) );
  NAND2_X1 U9669 ( .A1(n7393), .A2(n7391), .ZN(n13425) );
  NAND2_X1 U9670 ( .A1(n7403), .A2(n7401), .ZN(n13527) );
  NAND2_X1 U9671 ( .A1(n13104), .A2(n7415), .ZN(n7414) );
  NAND2_X1 U9672 ( .A1(n7422), .A2(n14633), .ZN(n7421) );
  OAI21_X1 U9673 ( .B1(n13158), .B2(n13154), .A(n13155), .ZN(n13120) );
  NAND2_X1 U9674 ( .A1(n13154), .A2(n13155), .ZN(n7427) );
  NAND2_X1 U9675 ( .A1(n7997), .A2(n7428), .ZN(n8192) );
  OAI21_X2 U9676 ( .B1(n9812), .B2(n7431), .A(n7429), .ZN(n9827) );
  NAND2_X1 U9677 ( .A1(n9697), .A2(n9696), .ZN(n9699) );
  INV_X1 U9678 ( .A(n9697), .ZN(n7434) );
  OAI21_X1 U9679 ( .B1(n9759), .B2(n7441), .A(n7439), .ZN(n9767) );
  NAND2_X1 U9680 ( .A1(n13135), .A2(n7443), .ZN(n13174) );
  AND2_X2 U9681 ( .A1(n13174), .A2(n9782), .ZN(n13113) );
  NAND4_X1 U9682 ( .A1(n7444), .A2(n7445), .A3(n7616), .A4(n7972), .ZN(n7993)
         );
  INV_X1 U9683 ( .A(n7960), .ZN(n7973) );
  NOR2_X2 U9684 ( .A1(n7742), .A2(n7666), .ZN(n7444) );
  NOR2_X2 U9685 ( .A1(n7916), .A2(n7938), .ZN(n7445) );
  INV_X1 U9686 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12729) );
  INV_X1 U9687 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15392) );
  INV_X1 U9688 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13995) );
  INV_X1 U9689 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7447) );
  NAND4_X1 U9690 ( .A1(n12729), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n7447), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7446) );
  NAND4_X1 U9691 ( .A1(n13297), .A2(n15392), .A3(n13995), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U9692 ( .A1(n11894), .A2(n11895), .ZN(n11893) );
  NAND3_X1 U9693 ( .A1(n11864), .A2(n14161), .A3(n11863), .ZN(n7452) );
  NAND2_X1 U9694 ( .A1(n7762), .A2(n7460), .ZN(n7458) );
  INV_X1 U9695 ( .A(n11879), .ZN(n7463) );
  INV_X1 U9696 ( .A(n7466), .ZN(n7465) );
  NAND2_X1 U9697 ( .A1(n7464), .A2(n7467), .ZN(n11881) );
  NAND2_X1 U9698 ( .A1(n7860), .A2(n7477), .ZN(n7476) );
  INV_X1 U9699 ( .A(n7911), .ZN(n7482) );
  NAND2_X1 U9700 ( .A1(n12796), .A2(n6572), .ZN(n7492) );
  INV_X1 U9701 ( .A(n12127), .ZN(n7500) );
  NAND2_X1 U9702 ( .A1(n15077), .A2(n7505), .ZN(n7501) );
  NAND2_X1 U9703 ( .A1(n7501), .A2(n7502), .ZN(n15055) );
  OAI21_X1 U9704 ( .B1(n15076), .B2(n7507), .A(n11284), .ZN(n7506) );
  AOI21_X2 U9705 ( .B1(n12186), .B2(n12185), .A(n7517), .ZN(n7516) );
  NAND2_X1 U9706 ( .A1(n7524), .A2(n7522), .ZN(n12890) );
  OAI21_X2 U9707 ( .B1(n12847), .B2(n12106), .A(n12105), .ZN(n12836) );
  AND2_X2 U9708 ( .A1(n9640), .A2(n7529), .ZN(n9162) );
  NAND2_X1 U9709 ( .A1(n7621), .A2(n7534), .ZN(n7535) );
  INV_X1 U9710 ( .A(n7535), .ZN(n7637) );
  AOI21_X1 U9711 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8878) );
  NAND3_X1 U9712 ( .A1(n8787), .A2(n8786), .A3(n7545), .ZN(n7544) );
  NAND3_X1 U9713 ( .A1(n8906), .A2(n8907), .A3(n6680), .ZN(n7548) );
  INV_X1 U9714 ( .A(n8910), .ZN(n7551) );
  NAND2_X1 U9715 ( .A1(n6605), .A2(n7556), .ZN(n7552) );
  OR2_X1 U9716 ( .A1(n6605), .A2(n7556), .ZN(n7554) );
  INV_X1 U9717 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7557) );
  INV_X1 U9718 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7558) );
  NOR2_X1 U9719 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8315) );
  NAND3_X1 U9720 ( .A1(n8316), .A2(n7558), .A3(n7557), .ZN(n8341) );
  INV_X1 U9721 ( .A(n8341), .ZN(n7559) );
  NAND2_X2 U9722 ( .A1(n8302), .A2(n8303), .ZN(n8578) );
  XNOR2_X2 U9723 ( .A(n7560), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8302) );
  NAND2_X2 U9724 ( .A1(n7561), .A2(n8691), .ZN(n14186) );
  NAND2_X1 U9725 ( .A1(n12205), .A2(n14793), .ZN(n7562) );
  NAND4_X1 U9726 ( .A1(n7562), .A2(n7564), .A3(n7563), .A4(n14803), .ZN(n7567)
         );
  NAND2_X1 U9727 ( .A1(n7570), .A2(n7569), .ZN(n8685) );
  INV_X1 U9728 ( .A(n8699), .ZN(n7575) );
  OAI21_X2 U9729 ( .B1(n14134), .B2(n7576), .A(n7573), .ZN(n14104) );
  NAND2_X1 U9730 ( .A1(n14033), .A2(n7584), .ZN(n7582) );
  INV_X1 U9731 ( .A(n14010), .ZN(n7580) );
  NAND2_X1 U9732 ( .A1(n7582), .A2(n7579), .ZN(n8712) );
  OR2_X2 U9733 ( .A1(n14033), .A2(n14034), .ZN(n14031) );
  NAND3_X1 U9734 ( .A1(n8414), .A2(n8297), .A3(n8293), .ZN(n8716) );
  NAND2_X1 U9735 ( .A1(n14101), .A2(n7593), .ZN(n7592) );
  XNOR2_X2 U9736 ( .A(n15045), .B(n15066), .ZN(n15061) );
  CLKBUF_X1 U9737 ( .A(n11332), .Z(n11429) );
  INV_X1 U9738 ( .A(n11509), .ZN(n11467) );
  OAI21_X1 U9739 ( .B1(n9691), .B2(n15179), .A(n9690), .ZN(n9693) );
  CLKBUF_X1 U9740 ( .A(P3_IR_REG_9__SCAN_IN), .Z(n9313) );
  NAND2_X1 U9741 ( .A1(n9167), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U9742 ( .A1(n9162), .A2(n9161), .ZN(n9167) );
  OR2_X1 U9743 ( .A1(n10675), .A2(n9487), .ZN(n9489) );
  OR2_X1 U9744 ( .A1(n10505), .A2(n9487), .ZN(n9475) );
  NAND4_X2 U9745 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), .ZN(n13008)
         );
  INV_X2 U9746 ( .A(n9179), .ZN(n9460) );
  NAND2_X2 U9747 ( .A1(n13111), .A2(n9786), .ZN(n13158) );
  AOI22_X1 U9748 ( .A1(n13960), .A2(n10521), .B1(n12362), .B2(n8662), .ZN(
        n10526) );
  INV_X1 U9749 ( .A(n8810), .ZN(n8813) );
  NAND2_X1 U9750 ( .A1(n11764), .A2(n11911), .ZN(n11765) );
  NAND2_X1 U9751 ( .A1(n9035), .A2(n9004), .ZN(n9005) );
  AND2_X1 U9752 ( .A1(n14803), .A2(n14330), .ZN(n14235) );
  INV_X1 U9753 ( .A(n15181), .ZN(n15179) );
  NAND2_X1 U9754 ( .A1(n10387), .A2(n14890), .ZN(n14924) );
  OR2_X1 U9755 ( .A1(n8747), .A2(n14327), .ZN(n7594) );
  OR2_X1 U9756 ( .A1(n8747), .A2(n8752), .ZN(n7595) );
  AND2_X1 U9757 ( .A1(n9848), .A2(n9847), .ZN(n7596) );
  INV_X1 U9758 ( .A(n14598), .ZN(n9339) );
  INV_X1 U9759 ( .A(n13702), .ZN(n8282) );
  INV_X1 U9760 ( .A(n13328), .ZN(n9846) );
  INV_X1 U9761 ( .A(n11158), .ZN(n8411) );
  INV_X1 U9762 ( .A(n15076), .ZN(n9591) );
  AND2_X1 U9763 ( .A1(n13771), .A2(n13770), .ZN(n7603) );
  INV_X1 U9764 ( .A(n12822), .ZN(n9618) );
  INV_X1 U9765 ( .A(n14108), .ZN(n8571) );
  AND2_X1 U9766 ( .A1(n8347), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7607) );
  AND2_X1 U9767 ( .A1(n11774), .A2(n11937), .ZN(n7608) );
  AND2_X1 U9768 ( .A1(n6545), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9769 ( .A1(n8764), .A2(n8994), .ZN(n8762) );
  NAND2_X1 U9770 ( .A1(n13234), .A2(n8822), .ZN(n8776) );
  OAI21_X1 U9771 ( .B1(n11911), .B2(n11766), .A(n11765), .ZN(n11767) );
  OAI21_X1 U9772 ( .B1(n8803), .B2(n8946), .A(n8802), .ZN(n8804) );
  INV_X1 U9773 ( .A(n8811), .ZN(n8812) );
  OAI211_X1 U9774 ( .C1(n8867), .C2(n8866), .A(n8876), .B(n8864), .ZN(n8879)
         );
  AOI22_X1 U9775 ( .A1(n13636), .A2(n8943), .B1(n8946), .B2(n13217), .ZN(n8910) );
  NAND2_X1 U9776 ( .A1(n8913), .A2(n8912), .ZN(n8918) );
  INV_X1 U9777 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9040) );
  NOR2_X1 U9778 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n9053) );
  INV_X1 U9779 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8295) );
  INV_X1 U9780 ( .A(n9524), .ZN(n9157) );
  NAND2_X1 U9781 ( .A1(n13015), .A2(n13007), .ZN(n13006) );
  INV_X1 U9782 ( .A(n8051), .ZN(n8052) );
  INV_X1 U9783 ( .A(n12604), .ZN(n12439) );
  INV_X1 U9784 ( .A(n9502), .ZN(n9155) );
  INV_X1 U9785 ( .A(n10519), .ZN(n10370) );
  NAND2_X1 U9786 ( .A1(n9157), .A2(n9156), .ZN(n9534) );
  INV_X1 U9787 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15273) );
  INV_X1 U9788 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15366) );
  INV_X1 U9789 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9134) );
  NOR2_X1 U9790 ( .A1(n7964), .A2(n13141), .ZN(n7978) );
  INV_X1 U9791 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10072) );
  OAI22_X1 U9792 ( .A1(n14007), .A2(n8634), .B1(n13741), .B2(n6879), .ZN(n8644) );
  INV_X1 U9793 ( .A(n14067), .ZN(n8593) );
  OR2_X1 U9794 ( .A1(n8484), .A2(n8483), .ZN(n8508) );
  INV_X1 U9795 ( .A(n14243), .ZN(n8664) );
  NAND2_X1 U9796 ( .A1(n8086), .A2(n8085), .ZN(n8094) );
  INV_X1 U9797 ( .A(n8034), .ZN(n8035) );
  INV_X1 U9798 ( .A(n11510), .ZN(n11466) );
  INV_X1 U9799 ( .A(n9490), .ZN(n9153) );
  INV_X1 U9800 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9226) );
  MUX2_X1 U9801 ( .A(n12018), .B(n15108), .S(n12421), .Z(n10689) );
  OR2_X1 U9802 ( .A1(n9515), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9524) );
  INV_X1 U9803 ( .A(n10383), .ZN(n10814) );
  AND2_X1 U9804 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  INV_X1 U9805 ( .A(n12807), .ZN(n9529) );
  AND2_X1 U9806 ( .A1(n12837), .A2(n12845), .ZN(n12114) );
  OR2_X1 U9807 ( .A1(n9463), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U9808 ( .A1(n9152), .A2(n15273), .ZN(n9463) );
  INV_X1 U9809 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15331) );
  AND2_X1 U9810 ( .A1(n9096), .A2(n9095), .ZN(n9318) );
  INV_X1 U9811 ( .A(n14643), .ZN(n9845) );
  AND2_X1 U9812 ( .A1(n14631), .A2(n9765), .ZN(n9766) );
  INV_X1 U9813 ( .A(n10964), .ZN(n9735) );
  INV_X1 U9814 ( .A(n13528), .ZN(n9714) );
  NOR2_X1 U9815 ( .A1(n8099), .A2(n8098), .ZN(n8118) );
  OR2_X1 U9816 ( .A1(n8043), .A2(n8042), .ZN(n8059) );
  OR2_X1 U9817 ( .A1(n7882), .A2(n11563), .ZN(n7901) );
  INV_X1 U9818 ( .A(n8131), .ZN(n8132) );
  OR2_X1 U9819 ( .A1(n7794), .A2(n10739), .ZN(n7814) );
  AND2_X1 U9820 ( .A1(n9009), .A2(n6564), .ZN(n9938) );
  OR2_X1 U9821 ( .A1(n7841), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7861) );
  NOR2_X1 U9822 ( .A1(n15336), .A2(n8575), .ZN(n8588) );
  INV_X1 U9823 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8422) );
  NOR2_X1 U9824 ( .A1(n8447), .A2(n8446), .ZN(n8457) );
  NOR2_X1 U9825 ( .A1(n8508), .A2(n8507), .ZN(n8519) );
  INV_X1 U9826 ( .A(n14017), .ZN(n14027) );
  INV_X1 U9827 ( .A(n14080), .ZN(n14095) );
  INV_X1 U9828 ( .A(n14292), .ZN(n8663) );
  NAND2_X1 U9829 ( .A1(n8961), .A2(n8960), .ZN(n8964) );
  OR2_X1 U9830 ( .A1(n8157), .A2(n11589), .ZN(n8158) );
  NOR2_X1 U9831 ( .A1(n14430), .A2(n14429), .ZN(n14409) );
  INV_X1 U9832 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U9833 ( .A1(n9153), .A2(n15291), .ZN(n9502) );
  OR2_X1 U9834 ( .A1(n9476), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9490) );
  INV_X1 U9835 ( .A(n12555), .ZN(n12587) );
  INV_X1 U9836 ( .A(n9423), .ZN(n9175) );
  INV_X1 U9837 ( .A(n12818), .ZN(n12845) );
  AND2_X1 U9838 ( .A1(n12095), .A2(n12094), .ZN(n12871) );
  AND2_X1 U9839 ( .A1(n12074), .A2(n12081), .ZN(n12915) );
  OR2_X1 U9840 ( .A1(n9292), .A2(n9144), .ZN(n9307) );
  INV_X1 U9841 ( .A(n13077), .ZN(n9686) );
  NAND2_X1 U9842 ( .A1(n15169), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9673) );
  INV_X1 U9843 ( .A(n12190), .ZN(n12012) );
  INV_X1 U9844 ( .A(n15039), .ZN(n15110) );
  AND2_X1 U9845 ( .A1(n9105), .A2(n9104), .ZN(n9379) );
  AND2_X1 U9846 ( .A1(n15210), .A2(n9078), .ZN(n9208) );
  INV_X1 U9847 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11563) );
  INV_X1 U9848 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7750) );
  OR2_X1 U9849 ( .A1(n9836), .A2(n10985), .ZN(n9833) );
  NOR2_X1 U9850 ( .A1(n8059), .A2(n13167), .ZN(n8074) );
  OR2_X1 U9851 ( .A1(n10231), .A2(n10232), .ZN(n10882) );
  INV_X1 U9852 ( .A(n9840), .ZN(n9832) );
  INV_X1 U9853 ( .A(n13518), .ZN(n13190) );
  INV_X1 U9854 ( .A(n9023), .ZN(n13499) );
  INV_X1 U9855 ( .A(n13540), .ZN(n13562) );
  AND2_X1 U9856 ( .A1(n7941), .A2(n7766), .ZN(n7810) );
  AND2_X1 U9857 ( .A1(n13843), .A2(n12323), .ZN(n13758) );
  OR3_X1 U9858 ( .A1(n8543), .A2(n8542), .A3(n8541), .ZN(n8551) );
  AND2_X1 U9859 ( .A1(n13756), .A2(n12313), .ZN(n13872) );
  NAND2_X1 U9860 ( .A1(n10665), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13887) );
  NOR2_X1 U9861 ( .A1(n8551), .A2(n15252), .ZN(n8557) );
  INV_X1 U9862 ( .A(n10308), .ZN(n10582) );
  INV_X1 U9863 ( .A(n11953), .ZN(n14228) );
  INV_X1 U9864 ( .A(n11789), .ZN(n11788) );
  NAND2_X1 U9865 ( .A1(n14529), .A2(n10720), .ZN(n14525) );
  XNOR2_X1 U9866 ( .A(n14248), .B(n13943), .ZN(n14034) );
  INV_X1 U9867 ( .A(n13868), .ZN(n14645) );
  INV_X1 U9868 ( .A(n14174), .ZN(n14212) );
  INV_X1 U9869 ( .A(n14522), .ZN(n14110) );
  INV_X1 U9870 ( .A(n14330), .ZN(n14788) );
  AND2_X1 U9871 ( .A1(n10300), .A2(n8746), .ZN(n14330) );
  INV_X1 U9872 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8646) );
  AND2_X1 U9873 ( .A1(n7956), .A2(n7937), .ZN(n7954) );
  XNOR2_X1 U9874 ( .A(n7875), .B(SI_12_), .ZN(n7873) );
  OAI21_X1 U9875 ( .B1(n7669), .B2(SI_2_), .A(n7686), .ZN(n7683) );
  OAI22_X1 U9876 ( .A1(n14453), .A2(n14405), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14969), .ZN(n14406) );
  INV_X1 U9877 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15304) );
  AND2_X1 U9878 ( .A1(n10643), .A2(n10642), .ZN(n12555) );
  AND2_X1 U9879 ( .A1(n10624), .A2(n15065), .ZN(n10932) );
  INV_X1 U9880 ( .A(n12594), .ZN(n14938) );
  INV_X1 U9881 ( .A(n14935), .ZN(n12592) );
  OR2_X1 U9882 ( .A1(n12381), .A2(n9478), .ZN(n11990) );
  AND4_X1 U9883 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n12872)
         );
  AND4_X1 U9884 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(n14591)
         );
  OR2_X1 U9885 ( .A1(n10364), .A2(n10363), .ZN(n10377) );
  INV_X1 U9886 ( .A(n15017), .ZN(n14999) );
  INV_X1 U9887 ( .A(n15007), .ZN(n14981) );
  INV_X1 U9888 ( .A(n15107), .ZN(n15046) );
  INV_X1 U9889 ( .A(n12869), .ZN(n15079) );
  INV_X1 U9890 ( .A(n15125), .ZN(n15101) );
  AND3_X1 U9891 ( .A1(n9681), .A2(n9680), .A3(n9679), .ZN(n10931) );
  NAND2_X1 U9892 ( .A1(n12012), .A2(n10934), .ZN(n15098) );
  INV_X1 U9893 ( .A(n14611), .ZN(n15162) );
  INV_X1 U9894 ( .A(n12946), .ZN(n15168) );
  INV_X1 U9895 ( .A(n15105), .ZN(n15043) );
  OR2_X1 U9896 ( .A1(n10008), .A2(n13078), .ZN(n15466) );
  AND2_X1 U9897 ( .A1(n10353), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9851) );
  AND2_X1 U9898 ( .A1(n9060), .A2(n9059), .ZN(n12190) );
  INV_X1 U9899 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9417) );
  OR2_X1 U9900 ( .A1(n7948), .A2(n7947), .ZN(n7964) );
  INV_X1 U9901 ( .A(n13202), .ZN(n14633) );
  INV_X1 U9902 ( .A(n14850), .ZN(n14833) );
  INV_X1 U9903 ( .A(n14862), .ZN(n14838) );
  NAND2_X1 U9904 ( .A1(n14891), .A2(n9832), .ZN(n13573) );
  INV_X1 U9905 ( .A(n13629), .ZN(n13675) );
  AND2_X1 U9906 ( .A1(n8261), .A2(n8279), .ZN(n14863) );
  AND3_X1 U9907 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n11920) );
  AND4_X1 U9908 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n13818)
         );
  AND4_X1 U9909 ( .A1(n8548), .A2(n8547), .A3(n8546), .A4(n8545), .ZN(n13902)
         );
  OR2_X1 U9910 ( .A1(n9860), .A2(n10047), .ZN(n14757) );
  INV_X1 U9911 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15395) );
  INV_X1 U9912 ( .A(n14753), .ZN(n14715) );
  OR2_X1 U9913 ( .A1(n9860), .A2(n9858), .ZN(n14719) );
  INV_X1 U9914 ( .A(n14757), .ZN(n14726) );
  INV_X1 U9915 ( .A(n10281), .ZN(n14512) );
  INV_X1 U9916 ( .A(n11850), .ZN(n14189) );
  INV_X1 U9917 ( .A(n14516), .ZN(n14194) );
  INV_X1 U9918 ( .A(n14525), .ZN(n14225) );
  INV_X1 U9919 ( .A(n14793), .ZN(n14313) );
  NAND2_X1 U9920 ( .A1(n14524), .A2(n10768), .ZN(n14793) );
  AND2_X1 U9921 ( .A1(n14796), .A2(n14330), .ZN(n11173) );
  NAND2_X1 U9922 ( .A1(n10296), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10080) );
  AND2_X1 U9923 ( .A1(n8469), .A2(n8479), .ZN(n14681) );
  NAND2_X1 U9924 ( .A1(n9664), .A2(n9663), .ZN(n10633) );
  INV_X1 U9925 ( .A(n12578), .ZN(n12590) );
  NAND2_X1 U9926 ( .A1(n10623), .A2(n10624), .ZN(n12594) );
  AND2_X1 U9927 ( .A1(n11990), .A2(n9629), .ZN(n12148) );
  INV_X1 U9928 ( .A(P3_U3897), .ZN(n12598) );
  INV_X1 U9929 ( .A(n12925), .ZN(n12601) );
  INV_X1 U9930 ( .A(n14978), .ZN(n15008) );
  INV_X1 U9931 ( .A(n12732), .ZN(n15023) );
  INV_X1 U9932 ( .A(n12737), .ZN(n15015) );
  NAND2_X1 U9933 ( .A1(n10935), .A2(n15101), .ZN(n15129) );
  NAND2_X1 U9934 ( .A1(n12385), .A2(n12938), .ZN(n9692) );
  INV_X1 U9935 ( .A(n12938), .ZN(n13001) );
  AND2_X2 U9936 ( .A1(n10931), .A2(n9688), .ZN(n15181) );
  NAND2_X1 U9937 ( .A1(n9691), .A2(n15170), .ZN(n9677) );
  INV_X2 U9938 ( .A(n15169), .ZN(n15170) );
  AND2_X1 U9939 ( .A1(n9672), .A2(n9671), .ZN(n15169) );
  INV_X2 U9940 ( .A(n15466), .ZN(n10034) );
  INV_X1 U9941 ( .A(n12014), .ZN(n10934) );
  INV_X1 U9942 ( .A(SI_18_), .ZN(n15448) );
  INV_X1 U9943 ( .A(SI_12_), .ZN(n9915) );
  INV_X1 U9944 ( .A(n13656), .ZN(n13504) );
  INV_X1 U9945 ( .A(n14638), .ZN(n13183) );
  NAND2_X1 U9946 ( .A1(n10164), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14643) );
  INV_X1 U9947 ( .A(n9837), .ZN(n13209) );
  OR3_X1 U9948 ( .A1(n7931), .A2(n7930), .A3(n7929), .ZN(n13519) );
  INV_X1 U9949 ( .A(n14855), .ZN(n14848) );
  INV_X1 U9950 ( .A(n13577), .ZN(n13486) );
  INV_X1 U9951 ( .A(n13579), .ZN(n13509) );
  INV_X2 U9952 ( .A(n14929), .ZN(n14931) );
  NAND2_X1 U9953 ( .A1(n8281), .A2(n8280), .ZN(n14890) );
  INV_X1 U9954 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11676) );
  INV_X1 U9955 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11204) );
  INV_X1 U9956 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n15303) );
  OR3_X1 U9957 ( .A1(n13891), .A2(n13772), .A3(n13938), .ZN(n13779) );
  INV_X1 U9958 ( .A(n12233), .ZN(n14538) );
  INV_X1 U9959 ( .A(n11810), .ZN(n11725) );
  INV_X1 U9960 ( .A(n13936), .ZN(n13921) );
  INV_X1 U9961 ( .A(n11920), .ZN(n13999) );
  INV_X1 U9962 ( .A(n13804), .ZN(n13949) );
  NAND2_X1 U9963 ( .A1(n9862), .A2(n9861), .ZN(n14761) );
  OR2_X1 U9964 ( .A1(n12199), .A2(n11760), .ZN(n14516) );
  INV_X1 U9965 ( .A(n14233), .ZN(n14201) );
  INV_X1 U9966 ( .A(n14235), .ZN(n14327) );
  AND2_X2 U9967 ( .A1(n8745), .A2(n10719), .ZN(n14803) );
  INV_X1 U9968 ( .A(n14206), .ZN(n14365) );
  INV_X1 U9969 ( .A(n14796), .ZN(n14794) );
  INV_X1 U9970 ( .A(n14764), .ZN(n14763) );
  NAND2_X1 U9971 ( .A1(n11979), .A2(n10079), .ZN(n14764) );
  INV_X1 U9972 ( .A(n11924), .ZN(n14393) );
  INV_X1 U9973 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10829) );
  INV_X1 U9974 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10157) );
  NOR2_X2 U9975 ( .A1(n10633), .A2(n13078), .ZN(P3_U3897) );
  NAND2_X1 U9976 ( .A1(n9677), .A2(n9676), .ZN(P3_U3456) );
  NOR2_X1 U9977 ( .A1(P2_U3088), .A2(n9943), .ZN(P2_U3947) );
  INV_X1 U9978 ( .A(n13959), .ZN(P1_U4016) );
  INV_X2 U9979 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7713) );
  INV_X2 U9980 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7740) );
  INV_X2 U9981 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7612) );
  NAND2_X2 U9982 ( .A1(n7656), .A2(n7642), .ZN(n7666) );
  NOR2_X1 U9983 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7615) );
  NOR3_X1 U9984 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n7620) );
  NOR2_X1 U9985 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7619) );
  NOR2_X1 U9986 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n7618) );
  NOR2_X1 U9987 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n7617) );
  NAND2_X1 U9988 ( .A1(n7637), .A2(n7638), .ZN(n7624) );
  INV_X1 U9989 ( .A(n7624), .ZN(n7622) );
  NAND2_X1 U9990 ( .A1(n7622), .A2(n7625), .ZN(n13722) );
  XNOR2_X2 U9991 ( .A(n7623), .B(n13723), .ZN(n7630) );
  INV_X2 U9992 ( .A(n7630), .ZN(n7628) );
  NAND2_X1 U9993 ( .A1(n7624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7626) );
  XNOR2_X2 U9994 ( .A(n7626), .B(n7625), .ZN(n7627) );
  NAND2_X4 U9995 ( .A1(n7628), .A2(n7629), .ZN(n8181) );
  INV_X1 U9996 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11007) );
  OR2_X1 U9997 ( .A1(n8181), .A2(n11007), .ZN(n7635) );
  INV_X1 U9998 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9963) );
  OR2_X1 U9999 ( .A1(n7660), .A2(n9963), .ZN(n7634) );
  BUF_X2 U10000 ( .A(n7630), .Z(n12215) );
  INV_X1 U10001 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7631) );
  INV_X1 U10002 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7636) );
  OR2_X2 U10003 ( .A1(n8259), .A2(n7636), .ZN(n7641) );
  NAND2_X1 U10004 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6810), .ZN(n7643) );
  MUX2_X1 U10005 ( .A(n7643), .B(P2_IR_REG_31__SCAN_IN), .S(n7642), .Z(n7644)
         );
  NAND2_X1 U10006 ( .A1(n7644), .A2(n7666), .ZN(n10036) );
  NAND2_X1 U10007 ( .A1(n7645), .A2(SI_1_), .ZN(n7668) );
  INV_X1 U10008 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9189) );
  INV_X1 U10009 ( .A(SI_0_), .ZN(n8333) );
  INV_X1 U10010 ( .A(n7647), .ZN(n7648) );
  NAND2_X1 U10011 ( .A1(n7649), .A2(n7648), .ZN(n7650) );
  INV_X1 U10012 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9917) );
  INV_X1 U10013 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11740) );
  INV_X1 U10014 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11736) );
  OR2_X1 U10015 ( .A1(n8240), .A2(n11736), .ZN(n7653) );
  INV_X1 U10016 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11737) );
  NAND2_X1 U10017 ( .A1(n7721), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7651) );
  NAND4_X1 U10018 ( .A1(n7654), .A2(n7651), .A3(n7653), .A4(n7652), .ZN(n8760)
         );
  XNOR2_X1 U10019 ( .A(n7657), .B(n9073), .ZN(n13738) );
  MUX2_X2 U10020 ( .A(n7656), .B(n13738), .S(n9940), .Z(n11752) );
  NAND2_X1 U10021 ( .A1(n7655), .A2(n11004), .ZN(n9698) );
  INV_X1 U10022 ( .A(n9698), .ZN(n11005) );
  OAI22_X1 U10023 ( .A1(n11006), .A2(n11005), .B1(n6562), .B2(n8764), .ZN(
        n10181) );
  INV_X1 U10024 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7658) );
  INV_X1 U10025 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11070) );
  OR2_X1 U10026 ( .A1(n8181), .A2(n11070), .ZN(n7663) );
  INV_X1 U10027 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7659) );
  OR2_X1 U10028 ( .A1(n8240), .A2(n7659), .ZN(n7662) );
  NAND2_X1 U10029 ( .A1(n7950), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7661) );
  NAND2_X2 U10030 ( .A1(n7664), .A2(n6599), .ZN(n13234) );
  NAND2_X1 U10031 ( .A1(n7666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7665) );
  MUX2_X1 U10032 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7665), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7667) );
  NAND2_X1 U10033 ( .A1(n7667), .A2(n7744), .ZN(n9962) );
  NAND2_X1 U10034 ( .A1(n7669), .A2(SI_2_), .ZN(n7686) );
  INV_X1 U10035 ( .A(n10183), .ZN(n7670) );
  NAND2_X1 U10036 ( .A1(n10181), .A2(n7670), .ZN(n7673) );
  INV_X1 U10037 ( .A(n13234), .ZN(n10277) );
  INV_X1 U10038 ( .A(n7671), .ZN(n11071) );
  NAND2_X1 U10039 ( .A1(n10277), .A2(n11071), .ZN(n7672) );
  NAND2_X1 U10040 ( .A1(n7673), .A2(n7672), .ZN(n10271) );
  NAND2_X1 U10041 ( .A1(n8177), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7678) );
  OR2_X1 U10042 ( .A1(n8149), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7677) );
  INV_X1 U10043 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11083) );
  OR2_X1 U10044 ( .A1(n8182), .A2(n11083), .ZN(n7676) );
  INV_X1 U10045 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7674) );
  OR2_X1 U10046 ( .A1(n7691), .A2(n7674), .ZN(n7675) );
  NAND2_X1 U10047 ( .A1(n7744), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7680) );
  MUX2_X1 U10048 ( .A(n7680), .B(P2_IR_REG_31__SCAN_IN), .S(n7679), .Z(n7681)
         );
  INV_X1 U10049 ( .A(n7681), .ZN(n7682) );
  NOR2_X1 U10050 ( .A1(n7744), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7714) );
  NOR2_X1 U10051 ( .A1(n7682), .A2(n7714), .ZN(n10120) );
  INV_X1 U10052 ( .A(n7683), .ZN(n7684) );
  NAND2_X1 U10053 ( .A1(n8343), .A2(n7702), .ZN(n7687) );
  INV_X1 U10054 ( .A(n10273), .ZN(n11079) );
  NAND2_X1 U10055 ( .A1(n7221), .A2(n11079), .ZN(n7689) );
  NAND2_X1 U10056 ( .A1(n8177), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7696) );
  INV_X1 U10057 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7692) );
  OR2_X1 U10058 ( .A1(n7691), .A2(n7692), .ZN(n7695) );
  AND2_X1 U10059 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7722) );
  INV_X1 U10060 ( .A(n7722), .ZN(n7724) );
  OAI21_X1 U10061 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7724), .ZN(n11061) );
  OR2_X1 U10062 ( .A1(n8181), .A2(n11061), .ZN(n7694) );
  INV_X1 U10063 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11066) );
  OR2_X1 U10064 ( .A1(n8182), .A2(n11066), .ZN(n7693) );
  NAND4_X1 U10065 ( .A1(n7696), .A2(n7695), .A3(n7694), .A4(n7693), .ZN(n13232) );
  NAND2_X1 U10066 ( .A1(n7701), .A2(SI_4_), .ZN(n7711) );
  OAI21_X1 U10067 ( .B1(n7701), .B2(SI_4_), .A(n7711), .ZN(n7708) );
  NAND2_X1 U10068 ( .A1(n9894), .A2(n7702), .ZN(n7706) );
  INV_X1 U10069 ( .A(n7714), .ZN(n7703) );
  NAND2_X1 U10070 ( .A1(n7703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7704) );
  XNOR2_X1 U10071 ( .A(n7704), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U10072 ( .A1(n8970), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6563), .B2(
        n10001), .ZN(n7705) );
  NAND2_X1 U10073 ( .A1(n7706), .A2(n7705), .ZN(n10393) );
  OR2_X1 U10074 ( .A1(n13232), .A2(n10393), .ZN(n7707) );
  INV_X1 U10075 ( .A(n7708), .ZN(n7709) );
  MUX2_X1 U10076 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6568), .Z(n7712) );
  NAND2_X1 U10077 ( .A1(n7712), .A2(SI_5_), .ZN(n7736) );
  OAI21_X1 U10078 ( .B1(n7712), .B2(SI_5_), .A(n7736), .ZN(n7733) );
  XNOR2_X1 U10079 ( .A(n7735), .B(n7733), .ZN(n9899) );
  NAND2_X1 U10080 ( .A1(n9899), .A2(n7702), .ZN(n7720) );
  NAND2_X1 U10081 ( .A1(n7714), .A2(n7713), .ZN(n7717) );
  NAND2_X1 U10082 ( .A1(n7717), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7716) );
  MUX2_X1 U10083 ( .A(n7716), .B(P2_IR_REG_31__SCAN_IN), .S(n7715), .Z(n7718)
         );
  OR2_X1 U10084 ( .A1(n7717), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7739) );
  AOI22_X1 U10085 ( .A1(n8970), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6563), .B2(
        n9986), .ZN(n7719) );
  NAND2_X1 U10086 ( .A1(n7720), .A2(n7719), .ZN(n10989) );
  NAND2_X1 U10087 ( .A1(n8161), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7729) );
  INV_X1 U10088 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9948) );
  OR2_X1 U10089 ( .A1(n6566), .A2(n9948), .ZN(n7728) );
  NAND2_X1 U10090 ( .A1(n7722), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7751) );
  INV_X1 U10091 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10092 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  NAND2_X1 U10093 ( .A1(n7751), .A2(n7725), .ZN(n10987) );
  OR2_X1 U10094 ( .A1(n8149), .A2(n10987), .ZN(n7727) );
  INV_X1 U10095 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9971) );
  OR2_X1 U10096 ( .A1(n8182), .A2(n9971), .ZN(n7726) );
  NAND4_X1 U10097 ( .A1(n7729), .A2(n7728), .A3(n7727), .A4(n7726), .ZN(n13231) );
  NOR2_X1 U10098 ( .A1(n10989), .A2(n13231), .ZN(n7730) );
  NAND2_X1 U10099 ( .A1(n10989), .A2(n13231), .ZN(n7731) );
  NAND2_X1 U10100 ( .A1(n7732), .A2(n7731), .ZN(n11113) );
  INV_X1 U10101 ( .A(n7733), .ZN(n7734) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6551), .Z(n7738) );
  NAND2_X1 U10103 ( .A1(n7738), .A2(SI_6_), .ZN(n7763) );
  OAI21_X1 U10104 ( .B1(n7738), .B2(SI_6_), .A(n7763), .ZN(n7760) );
  XNOR2_X1 U10105 ( .A(n7762), .B(n7760), .ZN(n9918) );
  NAND2_X1 U10106 ( .A1(n9918), .A2(n7702), .ZN(n7748) );
  NAND2_X1 U10107 ( .A1(n7739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7741) );
  MUX2_X1 U10108 ( .A(n7741), .B(P2_IR_REG_31__SCAN_IN), .S(n7740), .Z(n7746)
         );
  INV_X1 U10109 ( .A(n7941), .ZN(n7745) );
  NAND2_X1 U10110 ( .A1(n7746), .A2(n7745), .ZN(n9989) );
  INV_X1 U10111 ( .A(n9989), .ZN(n10061) );
  AOI22_X1 U10112 ( .A1(n8970), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6563), .B2(
        n10061), .ZN(n7747) );
  NAND2_X1 U10113 ( .A1(n7748), .A2(n7747), .ZN(n14910) );
  NAND2_X1 U10114 ( .A1(n8161), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7756) );
  INV_X1 U10115 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7749) );
  OR2_X1 U10116 ( .A1(n6566), .A2(n7749), .ZN(n7755) );
  NOR2_X1 U10117 ( .A1(n7751), .A2(n7750), .ZN(n7771) );
  INV_X1 U10118 ( .A(n7771), .ZN(n7773) );
  NAND2_X1 U10119 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U10120 ( .A1(n7773), .A2(n7752), .ZN(n11126) );
  OR2_X1 U10121 ( .A1(n8149), .A2(n11126), .ZN(n7754) );
  INV_X1 U10122 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11123) );
  OR2_X1 U10123 ( .A1(n8182), .A2(n11123), .ZN(n7753) );
  NAND4_X1 U10124 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n13230) );
  INV_X1 U10125 ( .A(n13230), .ZN(n8803) );
  NAND2_X1 U10126 ( .A1(n14910), .A2(n8803), .ZN(n8207) );
  OR2_X1 U10127 ( .A1(n14910), .A2(n8803), .ZN(n7757) );
  NAND2_X1 U10128 ( .A1(n8207), .A2(n7757), .ZN(n11115) );
  NAND2_X1 U10129 ( .A1(n11113), .A2(n11115), .ZN(n7759) );
  NAND2_X1 U10130 ( .A1(n14910), .A2(n13230), .ZN(n7758) );
  INV_X1 U10131 ( .A(n7760), .ZN(n7761) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6568), .Z(n7764) );
  NAND2_X1 U10133 ( .A1(n7764), .A2(SI_7_), .ZN(n7784) );
  OAI21_X1 U10134 ( .B1(n7764), .B2(SI_7_), .A(n7784), .ZN(n7781) );
  XNOR2_X1 U10135 ( .A(n7783), .B(n7781), .ZN(n9923) );
  NAND2_X1 U10136 ( .A1(n9923), .A2(n7702), .ZN(n7769) );
  NOR2_X1 U10137 ( .A1(n7941), .A2(n7636), .ZN(n7765) );
  MUX2_X1 U10138 ( .A(n7636), .B(n7765), .S(P2_IR_REG_7__SCAN_IN), .Z(n7767)
         );
  NOR2_X1 U10139 ( .A1(n7767), .A2(n7810), .ZN(n13240) );
  AOI22_X1 U10140 ( .A1(n8970), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6563), .B2(
        n13240), .ZN(n7768) );
  NAND2_X1 U10141 ( .A1(n7769), .A2(n7768), .ZN(n14917) );
  NAND2_X1 U10142 ( .A1(n8161), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7778) );
  INV_X1 U10143 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7770) );
  OR2_X1 U10144 ( .A1(n6566), .A2(n7770), .ZN(n7777) );
  NAND2_X1 U10145 ( .A1(n7771), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7794) );
  INV_X1 U10146 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10147 ( .A1(n7773), .A2(n7772), .ZN(n7774) );
  NAND2_X1 U10148 ( .A1(n7794), .A2(n7774), .ZN(n11139) );
  OR2_X1 U10149 ( .A1(n8181), .A2(n11139), .ZN(n7776) );
  INV_X1 U10150 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11136) );
  OR2_X1 U10151 ( .A1(n8182), .A2(n11136), .ZN(n7775) );
  NAND4_X1 U10152 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .ZN(n13229) );
  AND2_X1 U10153 ( .A1(n14917), .A2(n13229), .ZN(n7779) );
  OR2_X1 U10154 ( .A1(n14917), .A2(n13229), .ZN(n7780) );
  INV_X1 U10155 ( .A(n7781), .ZN(n7782) );
  MUX2_X1 U10156 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6568), .Z(n7785) );
  NAND2_X1 U10157 ( .A1(n7785), .A2(SI_8_), .ZN(n7801) );
  OAI21_X1 U10158 ( .B1(n7785), .B2(SI_8_), .A(n7801), .ZN(n7786) );
  INV_X1 U10159 ( .A(n7786), .ZN(n7787) );
  OR2_X1 U10160 ( .A1(n7788), .A2(n7787), .ZN(n7789) );
  NAND2_X1 U10161 ( .A1(n7802), .A2(n7789), .ZN(n9931) );
  OR2_X1 U10162 ( .A1(n9931), .A2(n7808), .ZN(n7792) );
  OR2_X1 U10163 ( .A1(n7810), .A2(n7636), .ZN(n7790) );
  XNOR2_X1 U10164 ( .A(n7790), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U10165 ( .A1(n8970), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6563), .B2(
        n13258), .ZN(n7791) );
  NAND2_X1 U10166 ( .A1(n8177), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7799) );
  INV_X1 U10167 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7793) );
  OR2_X1 U10168 ( .A1(n7691), .A2(n7793), .ZN(n7798) );
  INV_X1 U10169 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U10170 ( .A1(n7794), .A2(n10739), .ZN(n7795) );
  NAND2_X1 U10171 ( .A1(n7814), .A2(n7795), .ZN(n11106) );
  OR2_X1 U10172 ( .A1(n8149), .A2(n11106), .ZN(n7797) );
  INV_X1 U10173 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11105) );
  OR2_X1 U10174 ( .A1(n8182), .A2(n11105), .ZN(n7796) );
  NAND4_X1 U10175 ( .A1(n7799), .A2(n7798), .A3(n7797), .A4(n7796), .ZN(n13228) );
  XNOR2_X1 U10176 ( .A(n10913), .B(n13228), .ZN(n10908) );
  NAND2_X1 U10177 ( .A1(n10913), .A2(n13228), .ZN(n7800) );
  MUX2_X1 U10178 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9903), .Z(n7803) );
  OAI21_X1 U10179 ( .B1(n7803), .B2(SI_9_), .A(n7820), .ZN(n7804) );
  INV_X1 U10180 ( .A(n7804), .ZN(n7805) );
  OR2_X1 U10181 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U10182 ( .A1(n7821), .A2(n7807), .ZN(n9937) );
  OR2_X1 U10183 ( .A1(n9937), .A2(n7808), .ZN(n7813) );
  OR2_X1 U10184 ( .A1(n7919), .A2(n7636), .ZN(n7811) );
  XNOR2_X1 U10185 ( .A(n7811), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U10186 ( .A1(n8970), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6563), .B2(
        n10067), .ZN(n7812) );
  NAND2_X1 U10187 ( .A1(n8161), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7819) );
  INV_X1 U10188 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10104) );
  OR2_X1 U10189 ( .A1(n6566), .A2(n10104), .ZN(n7818) );
  INV_X1 U10190 ( .A(n7828), .ZN(n7830) );
  NAND2_X1 U10191 ( .A1(n7814), .A2(n10072), .ZN(n7815) );
  NAND2_X1 U10192 ( .A1(n7830), .A2(n7815), .ZN(n11247) );
  OR2_X1 U10193 ( .A1(n8149), .A2(n11247), .ZN(n7817) );
  INV_X1 U10194 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11248) );
  OR2_X1 U10195 ( .A1(n8182), .A2(n11248), .ZN(n7816) );
  NAND4_X1 U10196 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n13227) );
  INV_X1 U10197 ( .A(n13227), .ZN(n8826) );
  XNOR2_X1 U10198 ( .A(n11250), .B(n8826), .ZN(n11176) );
  MUX2_X1 U10199 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9903), .Z(n7837) );
  XNOR2_X1 U10200 ( .A(n7837), .B(SI_10_), .ZN(n7822) );
  XNOR2_X1 U10201 ( .A(n7839), .B(n7822), .ZN(n10088) );
  NAND2_X1 U10202 ( .A1(n10088), .A2(n7702), .ZN(n7826) );
  INV_X1 U10203 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10204 ( .A1(n7919), .A2(n7823), .ZN(n7841) );
  NAND2_X1 U10205 ( .A1(n7841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7824) );
  XNOR2_X1 U10206 ( .A(n7824), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U10207 ( .A1(n8970), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6563), 
        .B2(n14824), .ZN(n7825) );
  NAND2_X1 U10208 ( .A1(n8177), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7835) );
  INV_X1 U10209 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7827) );
  OR2_X1 U10210 ( .A1(n7691), .A2(n7827), .ZN(n7834) );
  INV_X1 U10211 ( .A(n7846), .ZN(n7847) );
  INV_X1 U10212 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10213 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U10214 ( .A1(n7847), .A2(n7831), .ZN(n11266) );
  OR2_X1 U10215 ( .A1(n8149), .A2(n11266), .ZN(n7833) );
  INV_X1 U10216 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11267) );
  OR2_X1 U10217 ( .A1(n8182), .A2(n11267), .ZN(n7832) );
  NAND4_X1 U10218 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n13226) );
  INV_X1 U10219 ( .A(n13226), .ZN(n10965) );
  XNOR2_X1 U10220 ( .A(n11277), .B(n10965), .ZN(n11262) );
  NAND2_X1 U10221 ( .A1(n11277), .A2(n13226), .ZN(n7836) );
  NAND2_X1 U10222 ( .A1(n11265), .A2(n7836), .ZN(n11344) );
  NOR2_X1 U10223 ( .A1(n7840), .A2(n15445), .ZN(n7838) );
  MUX2_X1 U10224 ( .A(n10130), .B(n15303), .S(n6568), .Z(n7858) );
  XNOR2_X1 U10225 ( .A(n7858), .B(SI_11_), .ZN(n7856) );
  XNOR2_X1 U10226 ( .A(n7857), .B(n7856), .ZN(n10129) );
  NAND2_X1 U10227 ( .A1(n10129), .A2(n7702), .ZN(n7844) );
  NAND2_X1 U10228 ( .A1(n7861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7842) );
  XNOR2_X1 U10229 ( .A(n7842), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U10230 ( .A1(n8970), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6563), 
        .B2(n10138), .ZN(n7843) );
  NAND2_X1 U10231 ( .A1(n8177), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7852) );
  INV_X1 U10232 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7845) );
  OR2_X1 U10233 ( .A1(n7691), .A2(n7845), .ZN(n7851) );
  INV_X1 U10234 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U10235 ( .A1(n7847), .A2(n15348), .ZN(n7848) );
  NAND2_X1 U10236 ( .A1(n7865), .A2(n7848), .ZN(n11346) );
  OR2_X1 U10237 ( .A1(n8149), .A2(n11346), .ZN(n7850) );
  INV_X1 U10238 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11347) );
  OR2_X1 U10239 ( .A1(n8182), .A2(n11347), .ZN(n7849) );
  NAND4_X1 U10240 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n13225) );
  OR2_X1 U10241 ( .A1(n11479), .A2(n13225), .ZN(n7853) );
  NAND2_X1 U10242 ( .A1(n11344), .A2(n7853), .ZN(n7855) );
  NAND2_X1 U10243 ( .A1(n11479), .A2(n13225), .ZN(n7854) );
  NAND2_X1 U10244 ( .A1(n7858), .A2(n9898), .ZN(n7859) );
  MUX2_X1 U10245 ( .A(n10135), .B(n10137), .S(n6568), .Z(n7875) );
  XNOR2_X1 U10246 ( .A(n7874), .B(n7873), .ZN(n10134) );
  NAND2_X1 U10247 ( .A1(n10134), .A2(n7702), .ZN(n7864) );
  NOR2_X1 U10248 ( .A1(n7861), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n7877) );
  OR2_X1 U10249 ( .A1(n7877), .A2(n7636), .ZN(n7862) );
  XNOR2_X1 U10250 ( .A(n7862), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U10251 ( .A1(n6563), .A2(n10144), .B1(n8970), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10252 ( .A1(n8161), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7870) );
  INV_X1 U10253 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10227) );
  OR2_X1 U10254 ( .A1(n6566), .A2(n10227), .ZN(n7869) );
  INV_X1 U10255 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U10256 ( .A1(n7865), .A2(n10149), .ZN(n7866) );
  NAND2_X1 U10257 ( .A1(n7882), .A2(n7866), .ZN(n13574) );
  OR2_X1 U10258 ( .A1(n8149), .A2(n13574), .ZN(n7868) );
  INV_X1 U10259 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n13575) );
  OR2_X1 U10260 ( .A1(n8182), .A2(n13575), .ZN(n7867) );
  NAND4_X1 U10261 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n13224) );
  AND2_X1 U10262 ( .A1(n13578), .A2(n13224), .ZN(n7871) );
  OR2_X1 U10263 ( .A1(n13578), .A2(n13224), .ZN(n7872) );
  MUX2_X1 U10264 ( .A(n10157), .B(n10158), .S(n6568), .Z(n7890) );
  XNOR2_X1 U10265 ( .A(n7890), .B(SI_13_), .ZN(n7876) );
  XNOR2_X1 U10266 ( .A(n7893), .B(n7876), .ZN(n10155) );
  NAND2_X1 U10267 ( .A1(n10155), .A2(n7702), .ZN(n7880) );
  NAND2_X1 U10268 ( .A1(n7877), .A2(n7612), .ZN(n7896) );
  NAND2_X1 U10269 ( .A1(n7896), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7878) );
  XNOR2_X1 U10270 ( .A(n7878), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U10271 ( .A1(n10880), .A2(n6563), .B1(n8970), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10272 ( .A1(n8177), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7887) );
  INV_X1 U10273 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7881) );
  OR2_X1 U10274 ( .A1(n7691), .A2(n7881), .ZN(n7886) );
  NAND2_X1 U10275 ( .A1(n7882), .A2(n11563), .ZN(n7883) );
  NAND2_X1 U10276 ( .A1(n7901), .A2(n7883), .ZN(n11415) );
  OR2_X1 U10277 ( .A1(n8149), .A2(n11415), .ZN(n7885) );
  INV_X1 U10278 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10235) );
  OR2_X1 U10279 ( .A1(n8182), .A2(n10235), .ZN(n7884) );
  NAND4_X1 U10280 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n13223) );
  NOR2_X1 U10281 ( .A1(n11575), .A2(n13223), .ZN(n7888) );
  NAND2_X1 U10282 ( .A1(n11575), .A2(n13223), .ZN(n7889) );
  NOR2_X1 U10283 ( .A1(n7891), .A2(SI_13_), .ZN(n7892) );
  OR2_X2 U10284 ( .A1(n7894), .A2(SI_14_), .ZN(n7911) );
  NAND2_X1 U10285 ( .A1(n7894), .A2(SI_14_), .ZN(n7895) );
  MUX2_X1 U10286 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6568), .Z(n7909) );
  XNOR2_X1 U10287 ( .A(n7910), .B(n7909), .ZN(n10462) );
  NAND2_X1 U10288 ( .A1(n10462), .A2(n7702), .ZN(n7899) );
  OAI21_X1 U10289 ( .B1(n7896), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7897) );
  XNOR2_X1 U10290 ( .A(n7897), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14837) );
  AOI22_X1 U10291 ( .A1(n14837), .A2(n6563), .B1(n8970), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n7898) );
  INV_X1 U10292 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7900) );
  INV_X1 U10293 ( .A(n7925), .ZN(n7927) );
  NAND2_X1 U10294 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  NAND2_X1 U10295 ( .A1(n7927), .A2(n7902), .ZN(n13555) );
  OR2_X1 U10296 ( .A1(n13555), .A2(n8149), .ZN(n7907) );
  INV_X1 U10297 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7903) );
  OR2_X1 U10298 ( .A1(n7691), .A2(n7903), .ZN(n7906) );
  INV_X1 U10299 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13556) );
  OR2_X1 U10300 ( .A1(n8182), .A2(n13556), .ZN(n7905) );
  INV_X1 U10301 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10883) );
  OR2_X1 U10302 ( .A1(n6566), .A2(n10883), .ZN(n7904) );
  NAND4_X1 U10303 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), .ZN(n13222) );
  AND2_X1 U10304 ( .A1(n13718), .A2(n13222), .ZN(n7908) );
  MUX2_X1 U10305 ( .A(n10672), .B(n10671), .S(n6551), .Z(n7912) );
  NAND2_X1 U10306 ( .A1(n7912), .A2(n15383), .ZN(n7934) );
  INV_X1 U10307 ( .A(n7912), .ZN(n7913) );
  NAND2_X1 U10308 ( .A1(n7913), .A2(SI_15_), .ZN(n7914) );
  XNOR2_X1 U10309 ( .A(n7933), .B(n7932), .ZN(n10670) );
  NAND2_X1 U10310 ( .A1(n10670), .A2(n7702), .ZN(n7923) );
  INV_X1 U10311 ( .A(n7915), .ZN(n7918) );
  NOR2_X1 U10312 ( .A1(n7918), .A2(n7917), .ZN(n7939) );
  NAND2_X1 U10313 ( .A1(n7919), .A2(n7939), .ZN(n7920) );
  NAND2_X1 U10314 ( .A1(n7920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7921) );
  XNOR2_X1 U10315 ( .A(n7921), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U10316 ( .A1(n8970), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6563), 
        .B2(n10893), .ZN(n7922) );
  INV_X1 U10317 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15235) );
  NAND2_X1 U10318 ( .A1(n8161), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7924) );
  OAI21_X1 U10319 ( .B1(n15235), .B2(n6566), .A(n7924), .ZN(n7931) );
  NAND2_X1 U10320 ( .A1(n7925), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7948) );
  INV_X1 U10321 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U10322 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NAND2_X1 U10323 ( .A1(n7948), .A2(n7928), .ZN(n13538) );
  NOR2_X1 U10324 ( .A1(n13538), .A2(n8149), .ZN(n7930) );
  INV_X1 U10325 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U10326 ( .A1(n8182), .A2(n15363), .ZN(n7929) );
  INV_X1 U10327 ( .A(n13519), .ZN(n8217) );
  XNOR2_X1 U10328 ( .A(n13715), .B(n8217), .ZN(n13545) );
  MUX2_X1 U10329 ( .A(n10702), .B(n10704), .S(n6568), .Z(n7935) );
  NAND2_X1 U10330 ( .A1(n7935), .A2(n15337), .ZN(n7956) );
  INV_X1 U10331 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U10332 ( .A1(n7936), .A2(SI_16_), .ZN(n7937) );
  XNOR2_X1 U10333 ( .A(n7955), .B(n7954), .ZN(n10701) );
  NAND2_X1 U10334 ( .A1(n10701), .A2(n7702), .ZN(n7946) );
  INV_X1 U10335 ( .A(n7938), .ZN(n7940) );
  NAND3_X1 U10336 ( .A1(n7941), .A2(n7940), .A3(n7939), .ZN(n7942) );
  NAND2_X1 U10337 ( .A1(n7942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7943) );
  MUX2_X1 U10338 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7943), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n7944) );
  NAND2_X1 U10339 ( .A1(n7944), .A2(n7960), .ZN(n11357) );
  INV_X1 U10340 ( .A(n11357), .ZN(n11359) );
  AOI22_X1 U10341 ( .A1(n8970), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6563), 
        .B2(n11359), .ZN(n7945) );
  INV_X1 U10342 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U10343 ( .A1(n7948), .A2(n7947), .ZN(n7949) );
  NAND2_X1 U10344 ( .A1(n7964), .A2(n7949), .ZN(n14642) );
  AOI22_X1 U10345 ( .A1(n8177), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n7950), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10346 ( .A1(n8161), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7951) );
  OAI211_X1 U10347 ( .C1(n14642), .C2(n8149), .A(n7952), .B(n7951), .ZN(n13221) );
  INV_X1 U10348 ( .A(n13221), .ZN(n13139) );
  XNOR2_X1 U10349 ( .A(n14637), .B(n13139), .ZN(n13512) );
  INV_X1 U10350 ( .A(n13512), .ZN(n13524) );
  NAND2_X1 U10351 ( .A1(n14637), .A2(n13221), .ZN(n7953) );
  NAND2_X1 U10352 ( .A1(n13527), .A2(n7953), .ZN(n13500) );
  MUX2_X1 U10353 ( .A(n10829), .B(n10831), .S(n6551), .Z(n7957) );
  INV_X1 U10354 ( .A(n7957), .ZN(n7958) );
  NAND2_X1 U10355 ( .A1(n7958), .A2(SI_17_), .ZN(n7959) );
  XNOR2_X1 U10356 ( .A(n7970), .B(n7969), .ZN(n10828) );
  NAND2_X1 U10357 ( .A1(n10828), .A2(n7702), .ZN(n7963) );
  OR2_X1 U10358 ( .A1(n7973), .A2(n7636), .ZN(n7961) );
  XNOR2_X1 U10359 ( .A(n7961), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U10360 ( .A1(n8970), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6563), 
        .B2(n13270), .ZN(n7962) );
  INV_X1 U10361 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13502) );
  INV_X1 U10362 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13141) );
  INV_X1 U10363 ( .A(n7978), .ZN(n7979) );
  NAND2_X1 U10364 ( .A1(n7964), .A2(n13141), .ZN(n7965) );
  NAND2_X1 U10365 ( .A1(n7979), .A2(n7965), .ZN(n13501) );
  OR2_X1 U10366 ( .A1(n13501), .A2(n8149), .ZN(n7967) );
  AOI22_X1 U10367 ( .A1(n8177), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8161), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n7966) );
  OAI211_X1 U10368 ( .C1(n8182), .C2(n13502), .A(n7967), .B(n7966), .ZN(n13517) );
  XNOR2_X1 U10369 ( .A(n13656), .B(n13517), .ZN(n9023) );
  NAND2_X1 U10370 ( .A1(n13656), .A2(n13517), .ZN(n7968) );
  MUX2_X1 U10371 ( .A(n11202), .B(n11204), .S(n6551), .Z(n8013) );
  XNOR2_X1 U10372 ( .A(n7988), .B(n8013), .ZN(n11201) );
  NAND2_X1 U10373 ( .A1(n11201), .A2(n7702), .ZN(n7977) );
  NAND2_X1 U10374 ( .A1(n7974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7975) );
  XNOR2_X1 U10375 ( .A(n7975), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U10376 ( .A1(n8970), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6563), 
        .B2(n13283), .ZN(n7976) );
  INV_X1 U10377 ( .A(n8002), .ZN(n8004) );
  INV_X1 U10378 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n15292) );
  NAND2_X1 U10379 ( .A1(n7979), .A2(n15292), .ZN(n7980) );
  AND2_X1 U10380 ( .A1(n8004), .A2(n7980), .ZN(n13484) );
  INV_X1 U10381 ( .A(n8149), .ZN(n8026) );
  NAND2_X1 U10382 ( .A1(n13484), .A2(n8026), .ZN(n7985) );
  INV_X1 U10383 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n15350) );
  NAND2_X1 U10384 ( .A1(n7950), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10385 ( .A1(n8161), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7981) );
  OAI211_X1 U10386 ( .C1(n6566), .C2(n15350), .A(n7982), .B(n7981), .ZN(n7983)
         );
  INV_X1 U10387 ( .A(n7983), .ZN(n7984) );
  NAND2_X1 U10388 ( .A1(n7985), .A2(n7984), .ZN(n13220) );
  XNOR2_X1 U10389 ( .A(n13651), .B(n13220), .ZN(n13491) );
  OR2_X1 U10390 ( .A1(n13651), .A2(n13220), .ZN(n7986) );
  INV_X1 U10391 ( .A(n8013), .ZN(n8017) );
  NOR2_X1 U10392 ( .A1(n8016), .A2(n15448), .ZN(n7987) );
  AOI21_X1 U10393 ( .B1(n7988), .B2(n8017), .A(n7987), .ZN(n7992) );
  MUX2_X1 U10394 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n6551), .Z(n7989) );
  NAND2_X1 U10395 ( .A1(n7989), .A2(SI_19_), .ZN(n8020) );
  INV_X1 U10396 ( .A(n7989), .ZN(n7990) );
  INV_X1 U10397 ( .A(SI_19_), .ZN(n10255) );
  NAND2_X1 U10398 ( .A1(n7990), .A2(n10255), .ZN(n8018) );
  AND2_X1 U10399 ( .A1(n8020), .A2(n8018), .ZN(n7991) );
  XNOR2_X1 U10400 ( .A(n7992), .B(n7991), .ZN(n11296) );
  NAND2_X1 U10401 ( .A1(n11296), .A2(n7702), .ZN(n8001) );
  NOR2_X2 U10402 ( .A1(n7993), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n7997) );
  INV_X1 U10403 ( .A(n7997), .ZN(n7994) );
  NAND2_X1 U10404 ( .A1(n7994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7995) );
  MUX2_X1 U10405 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7995), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n7998) );
  AOI22_X1 U10406 ( .A1(n8970), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6563), 
        .B2(n9002), .ZN(n8000) );
  INV_X1 U10407 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10408 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  NAND2_X1 U10409 ( .A1(n8043), .A2(n8005), .ZN(n13115) );
  OR2_X1 U10410 ( .A1(n13115), .A2(n8181), .ZN(n8010) );
  INV_X1 U10411 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U10412 ( .A1(n7950), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10413 ( .A1(n8161), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8006) );
  OAI211_X1 U10414 ( .C1(n6566), .C2(n15450), .A(n8007), .B(n8006), .ZN(n8008)
         );
  INV_X1 U10415 ( .A(n8008), .ZN(n8009) );
  NAND2_X1 U10416 ( .A1(n8010), .A2(n8009), .ZN(n13219) );
  NAND2_X1 U10417 ( .A1(n13647), .A2(n13219), .ZN(n8011) );
  NAND2_X1 U10418 ( .A1(n8012), .A2(n8011), .ZN(n13453) );
  OAI21_X1 U10419 ( .B1(n8013), .B2(n15448), .A(n8020), .ZN(n8014) );
  INV_X1 U10420 ( .A(n8014), .ZN(n8015) );
  NOR2_X1 U10421 ( .A1(n8017), .A2(SI_18_), .ZN(n8021) );
  INV_X1 U10422 ( .A(n8018), .ZN(n8019) );
  AOI21_X1 U10423 ( .B1(n8021), .B2(n8020), .A(n8019), .ZN(n8022) );
  MUX2_X1 U10424 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n6551), .Z(n8034) );
  XNOR2_X1 U10425 ( .A(n8036), .B(n8034), .ZN(n11300) );
  NAND2_X1 U10426 ( .A1(n11300), .A2(n7702), .ZN(n8025) );
  INV_X1 U10427 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11323) );
  OR2_X1 U10428 ( .A1(n8979), .A2(n11323), .ZN(n8024) );
  XNOR2_X1 U10429 ( .A(n8043), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U10430 ( .A1(n13461), .A2(n8026), .ZN(n8032) );
  INV_X1 U10431 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10432 ( .A1(n7950), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10433 ( .A1(n8161), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8027) );
  OAI211_X1 U10434 ( .C1(n6566), .C2(n8029), .A(n8028), .B(n8027), .ZN(n8030)
         );
  INV_X1 U10435 ( .A(n8030), .ZN(n8031) );
  NAND2_X1 U10436 ( .A1(n8032), .A2(n8031), .ZN(n13218) );
  AND2_X1 U10437 ( .A1(n13642), .A2(n13218), .ZN(n8033) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6568), .Z(n8054) );
  XNOR2_X1 U10439 ( .A(n8054), .B(SI_21_), .ZN(n8051) );
  XNOR2_X1 U10440 ( .A(n8053), .B(n8051), .ZN(n11405) );
  NAND2_X1 U10441 ( .A1(n11405), .A2(n7702), .ZN(n8040) );
  INV_X1 U10442 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11407) );
  OR2_X1 U10443 ( .A1(n8979), .A2(n11407), .ZN(n8039) );
  INV_X1 U10444 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13159) );
  INV_X1 U10445 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8041) );
  OAI21_X1 U10446 ( .B1(n8043), .B2(n13159), .A(n8041), .ZN(n8044) );
  NAND2_X1 U10447 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8042) );
  NAND2_X1 U10448 ( .A1(n8044), .A2(n8059), .ZN(n13439) );
  OR2_X1 U10449 ( .A1(n13439), .A2(n8181), .ZN(n8050) );
  INV_X1 U10450 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10451 ( .A1(n8161), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10452 ( .A1(n7950), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8045) );
  OAI211_X1 U10453 ( .C1(n6566), .C2(n8047), .A(n8046), .B(n8045), .ZN(n8048)
         );
  INV_X1 U10454 ( .A(n8048), .ZN(n8049) );
  NAND2_X1 U10455 ( .A1(n8050), .A2(n8049), .ZN(n13217) );
  INV_X1 U10456 ( .A(n13217), .ZN(n8224) );
  XNOR2_X1 U10457 ( .A(n13636), .B(n8224), .ZN(n13447) );
  NAND2_X1 U10458 ( .A1(n8054), .A2(SI_21_), .ZN(n8055) );
  XNOR2_X1 U10459 ( .A(n8086), .B(SI_22_), .ZN(n8564) );
  MUX2_X1 U10460 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6551), .Z(n8087) );
  XNOR2_X1 U10461 ( .A(n8564), .B(n8087), .ZN(n11731) );
  NAND2_X1 U10462 ( .A1(n11731), .A2(n7702), .ZN(n8058) );
  INV_X1 U10463 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11734) );
  OR2_X1 U10464 ( .A1(n8979), .A2(n11734), .ZN(n8057) );
  INV_X1 U10465 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13167) );
  AND2_X1 U10466 ( .A1(n8059), .A2(n13167), .ZN(n8060) );
  OR2_X1 U10467 ( .A1(n8060), .A2(n8074), .ZN(n13429) );
  INV_X1 U10468 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U10469 ( .A1(n8161), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10470 ( .A1(n7950), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8061) );
  OAI211_X1 U10471 ( .C1(n8063), .C2(n6566), .A(n8062), .B(n8061), .ZN(n8064)
         );
  INV_X1 U10472 ( .A(n8064), .ZN(n8065) );
  OAI21_X1 U10473 ( .B1(n13429), .B2(n8149), .A(n8065), .ZN(n13216) );
  INV_X1 U10474 ( .A(n13216), .ZN(n13122) );
  OR2_X1 U10475 ( .A1(n13705), .A2(n13122), .ZN(n8227) );
  NAND2_X1 U10476 ( .A1(n13705), .A2(n13122), .ZN(n8066) );
  NAND2_X1 U10477 ( .A1(n8227), .A2(n8066), .ZN(n13416) );
  INV_X1 U10478 ( .A(n13416), .ZN(n13422) );
  NAND2_X1 U10479 ( .A1(n13705), .A2(n13216), .ZN(n8067) );
  INV_X1 U10480 ( .A(n8564), .ZN(n8069) );
  AND2_X1 U10481 ( .A1(n8086), .A2(SI_22_), .ZN(n8068) );
  INV_X1 U10482 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11635) );
  INV_X1 U10483 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11639) );
  MUX2_X1 U10484 ( .A(n11635), .B(n11639), .S(n6568), .Z(n8089) );
  XNOR2_X1 U10485 ( .A(n8089), .B(SI_23_), .ZN(n8070) );
  NAND2_X1 U10486 ( .A1(n11636), .A2(n7702), .ZN(n8073) );
  OR2_X1 U10487 ( .A1(n8979), .A2(n11639), .ZN(n8072) );
  OR2_X1 U10488 ( .A1(n8074), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U10489 ( .A1(n8074), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10490 ( .A1(n8075), .A2(n8099), .ZN(n13409) );
  OR2_X1 U10491 ( .A1(n13409), .A2(n8149), .ZN(n8080) );
  INV_X1 U10492 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U10493 ( .A1(n8161), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10494 ( .A1(n7950), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8076) );
  OAI211_X1 U10495 ( .C1(n6566), .C2(n13627), .A(n8077), .B(n8076), .ZN(n8078)
         );
  INV_X1 U10496 ( .A(n8078), .ZN(n8079) );
  NAND2_X1 U10497 ( .A1(n8080), .A2(n8079), .ZN(n13215) );
  OR2_X1 U10498 ( .A1(n13408), .A2(n13215), .ZN(n8081) );
  NAND2_X1 U10499 ( .A1(n13399), .A2(n8081), .ZN(n8083) );
  NAND2_X1 U10500 ( .A1(n13408), .A2(n13215), .ZN(n8082) );
  INV_X1 U10501 ( .A(SI_23_), .ZN(n10960) );
  NAND2_X1 U10502 ( .A1(n8089), .A2(n10960), .ZN(n8091) );
  OAI21_X1 U10503 ( .B1(n8087), .B2(SI_22_), .A(n8091), .ZN(n8084) );
  INV_X1 U10504 ( .A(n8084), .ZN(n8085) );
  INV_X1 U10505 ( .A(n8087), .ZN(n8088) );
  INV_X1 U10506 ( .A(SI_22_), .ZN(n9499) );
  NOR2_X1 U10507 ( .A1(n8088), .A2(n9499), .ZN(n8092) );
  INV_X1 U10508 ( .A(n8089), .ZN(n8090) );
  AOI22_X1 U10509 ( .A1(n8092), .A2(n8091), .B1(n8090), .B2(SI_23_), .ZN(n8093) );
  MUX2_X1 U10510 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6551), .Z(n8108) );
  XNOR2_X1 U10511 ( .A(n8107), .B(n8108), .ZN(n11640) );
  NAND2_X1 U10512 ( .A1(n11640), .A2(n7702), .ZN(n8096) );
  INV_X1 U10513 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15371) );
  OR2_X1 U10514 ( .A1(n8979), .A2(n15371), .ZN(n8095) );
  NAND2_X1 U10515 ( .A1(n8161), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8106) );
  INV_X1 U10516 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8097) );
  OR2_X1 U10517 ( .A1(n8182), .A2(n8097), .ZN(n8105) );
  INV_X1 U10518 ( .A(n8099), .ZN(n8101) );
  INV_X1 U10519 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8098) );
  INV_X1 U10520 ( .A(n8118), .ZN(n8100) );
  OAI21_X1 U10521 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(n8101), .A(n8100), .ZN(
        n13391) );
  OR2_X1 U10522 ( .A1(n8149), .A2(n13391), .ZN(n8104) );
  INV_X1 U10523 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8102) );
  OR2_X1 U10524 ( .A1(n6566), .A2(n8102), .ZN(n8103) );
  NAND4_X1 U10525 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n13214) );
  XNOR2_X1 U10526 ( .A(n13620), .B(n13214), .ZN(n13382) );
  INV_X1 U10527 ( .A(n13382), .ZN(n13384) );
  INV_X1 U10528 ( .A(n8107), .ZN(n8109) );
  NAND2_X1 U10529 ( .A1(n8110), .A2(SI_24_), .ZN(n8111) );
  INV_X1 U10530 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11672) );
  MUX2_X1 U10531 ( .A(n11672), .B(n11676), .S(n6568), .Z(n8112) );
  INV_X1 U10532 ( .A(SI_25_), .ZN(n15435) );
  NAND2_X1 U10533 ( .A1(n8112), .A2(n15435), .ZN(n8127) );
  INV_X1 U10534 ( .A(n8112), .ZN(n8113) );
  NAND2_X1 U10535 ( .A1(n8113), .A2(SI_25_), .ZN(n8114) );
  NAND2_X1 U10536 ( .A1(n8127), .A2(n8114), .ZN(n8125) );
  XNOR2_X1 U10537 ( .A(n8126), .B(n8125), .ZN(n11671) );
  NAND2_X1 U10538 ( .A1(n11671), .A2(n7702), .ZN(n8116) );
  OR2_X1 U10539 ( .A1(n8979), .A2(n11676), .ZN(n8115) );
  NAND2_X1 U10540 ( .A1(n8177), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8122) );
  INV_X1 U10541 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8117) );
  OR2_X1 U10542 ( .A1(n7691), .A2(n8117), .ZN(n8121) );
  NAND2_X1 U10543 ( .A1(n8118), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8131) );
  OAI21_X1 U10544 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8118), .A(n8131), .ZN(
        n13375) );
  OR2_X1 U10545 ( .A1(n8149), .A2(n13375), .ZN(n8120) );
  INV_X1 U10546 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13376) );
  OR2_X1 U10547 ( .A1(n8182), .A2(n13376), .ZN(n8119) );
  NAND4_X1 U10548 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n13213) );
  OR2_X1 U10549 ( .A1(n13696), .A2(n13213), .ZN(n8123) );
  INV_X1 U10550 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14388) );
  INV_X1 U10551 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15264) );
  MUX2_X1 U10552 ( .A(n14388), .B(n15264), .S(n6568), .Z(n8138) );
  XNOR2_X1 U10553 ( .A(n8138), .B(SI_26_), .ZN(n8128) );
  NAND2_X1 U10554 ( .A1(n13735), .A2(n7702), .ZN(n8130) );
  OR2_X1 U10555 ( .A1(n8979), .A2(n15264), .ZN(n8129) );
  NAND2_X1 U10556 ( .A1(n8161), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8136) );
  INV_X1 U10557 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13354) );
  OR2_X1 U10558 ( .A1(n8182), .A2(n13354), .ZN(n8135) );
  NAND2_X1 U10559 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8132), .ZN(n8147) );
  OAI21_X1 U10560 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8132), .A(n8147), .ZN(
        n13353) );
  OR2_X1 U10561 ( .A1(n8149), .A2(n13353), .ZN(n8134) );
  INV_X1 U10562 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13611) );
  OR2_X1 U10563 ( .A1(n6566), .A2(n13611), .ZN(n8133) );
  NAND4_X1 U10564 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n13212) );
  NOR2_X1 U10565 ( .A1(n13361), .A2(n13212), .ZN(n8137) );
  INV_X1 U10566 ( .A(n13361), .ZN(n13693) );
  INV_X1 U10567 ( .A(n13212), .ZN(n9011) );
  INV_X1 U10568 ( .A(SI_26_), .ZN(n11502) );
  INV_X1 U10569 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14385) );
  INV_X1 U10570 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13734) );
  MUX2_X1 U10571 ( .A(n14385), .B(n13734), .S(n6551), .Z(n8154) );
  XNOR2_X1 U10572 ( .A(n8154), .B(SI_27_), .ZN(n8142) );
  NAND2_X1 U10573 ( .A1(n13732), .A2(n7702), .ZN(n8144) );
  OR2_X1 U10574 ( .A1(n8979), .A2(n13734), .ZN(n8143) );
  NAND2_X1 U10575 ( .A1(n8177), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8153) );
  INV_X1 U10576 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13687) );
  OR2_X1 U10577 ( .A1(n7691), .A2(n13687), .ZN(n8152) );
  INV_X1 U10578 ( .A(n8147), .ZN(n8145) );
  NAND2_X1 U10579 ( .A1(n8145), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8179) );
  INV_X1 U10580 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10581 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  NAND2_X1 U10582 ( .A1(n8179), .A2(n8148), .ZN(n13344) );
  OR2_X1 U10583 ( .A1(n8149), .A2(n13344), .ZN(n8151) );
  INV_X1 U10584 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13345) );
  OR2_X1 U10585 ( .A1(n8182), .A2(n13345), .ZN(n8150) );
  XNOR2_X1 U10586 ( .A(n13347), .B(n13189), .ZN(n13341) );
  INV_X1 U10587 ( .A(SI_27_), .ZN(n11589) );
  NAND2_X1 U10588 ( .A1(n8157), .A2(n11589), .ZN(n8156) );
  INV_X1 U10589 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U10590 ( .A1(n8156), .A2(n8155), .ZN(n8159) );
  MUX2_X1 U10591 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6551), .Z(n8171) );
  XNOR2_X1 U10592 ( .A(n8171), .B(SI_28_), .ZN(n8174) );
  INV_X1 U10593 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13731) );
  OR2_X1 U10594 ( .A1(n8979), .A2(n13731), .ZN(n8160) );
  NAND2_X1 U10595 ( .A1(n8161), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8168) );
  INV_X1 U10596 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8162) );
  OR2_X1 U10597 ( .A1(n8182), .A2(n8162), .ZN(n8167) );
  INV_X1 U10598 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10599 ( .A(n8179), .B(n8163), .ZN(n13328) );
  OR2_X1 U10600 ( .A1(n8149), .A2(n13328), .ZN(n8166) );
  INV_X1 U10601 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8164) );
  OR2_X1 U10602 ( .A1(n6566), .A2(n8164), .ZN(n8165) );
  XNOR2_X2 U10603 ( .A(n13598), .B(n13096), .ZN(n13330) );
  NAND2_X1 U10604 ( .A1(n13331), .A2(n13330), .ZN(n8170) );
  OR2_X1 U10605 ( .A1(n7422), .A2(n13096), .ZN(n8169) );
  NAND2_X1 U10606 ( .A1(n8170), .A2(n8169), .ZN(n8187) );
  INV_X1 U10607 ( .A(n8171), .ZN(n8172) );
  INV_X1 U10608 ( .A(SI_28_), .ZN(n11730) );
  NAND2_X1 U10609 ( .A1(n8172), .A2(n11730), .ZN(n8173) );
  INV_X1 U10610 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14381) );
  INV_X1 U10611 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n15334) );
  MUX2_X1 U10612 ( .A(n14381), .B(n15334), .S(n6551), .Z(n8962) );
  XNOR2_X1 U10613 ( .A(n8962), .B(SI_29_), .ZN(n8960) );
  NOR2_X1 U10615 ( .A1(n8979), .A2(n15334), .ZN(n8176) );
  AOI21_X2 U10616 ( .B1(n12194), .B2(n7702), .A(n8176), .ZN(n13596) );
  INV_X1 U10617 ( .A(n13596), .ZN(n13316) );
  NAND2_X1 U10618 ( .A1(n8177), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8186) );
  INV_X1 U10619 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8178) );
  OR2_X1 U10620 ( .A1(n7691), .A2(n8178), .ZN(n8185) );
  INV_X1 U10621 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U10622 ( .A1(n8180), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13313) );
  OR2_X1 U10623 ( .A1(n8181), .A2(n13313), .ZN(n8184) );
  INV_X1 U10624 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13314) );
  OR2_X1 U10625 ( .A1(n8182), .A2(n13314), .ZN(n8183) );
  AND4_X1 U10626 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n9837)
         );
  XNOR2_X1 U10627 ( .A(n13316), .B(n13209), .ZN(n9028) );
  XNOR2_X1 U10628 ( .A(n8187), .B(n9028), .ZN(n13320) );
  INV_X1 U10629 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8188) );
  INV_X1 U10630 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8193) );
  XNOR2_X2 U10631 ( .A(n8194), .B(n8193), .ZN(n8755) );
  AND2_X1 U10632 ( .A1(n9002), .A2(n11322), .ZN(n8196) );
  NAND2_X1 U10633 ( .A1(n6794), .A2(n8756), .ZN(n14905) );
  NAND2_X1 U10634 ( .A1(n13320), .A2(n14905), .ZN(n8247) );
  NOR2_X1 U10635 ( .A1(n7655), .A2(n11752), .ZN(n10999) );
  NAND2_X1 U10636 ( .A1(n11006), .A2(n10999), .ZN(n8198) );
  INV_X1 U10637 ( .A(n8764), .ZN(n10185) );
  NAND2_X1 U10638 ( .A1(n10185), .A2(n6562), .ZN(n8197) );
  NAND2_X1 U10639 ( .A1(n8198), .A2(n8197), .ZN(n10184) );
  NAND2_X1 U10640 ( .A1(n10184), .A2(n10183), .ZN(n8200) );
  NAND2_X1 U10641 ( .A1(n10277), .A2(n7671), .ZN(n8199) );
  NAND2_X1 U10642 ( .A1(n8200), .A2(n8199), .ZN(n10275) );
  NAND2_X1 U10643 ( .A1(n10275), .A2(n10274), .ZN(n8202) );
  NAND2_X1 U10644 ( .A1(n7221), .A2(n10273), .ZN(n8201) );
  NAND2_X1 U10645 ( .A1(n8202), .A2(n8201), .ZN(n10395) );
  INV_X1 U10646 ( .A(n9018), .ZN(n10394) );
  NAND2_X1 U10647 ( .A1(n10395), .A2(n10394), .ZN(n8204) );
  NAND2_X1 U10648 ( .A1(n10276), .A2(n10393), .ZN(n8203) );
  INV_X1 U10649 ( .A(n13231), .ZN(n10573) );
  AND2_X1 U10650 ( .A1(n10989), .A2(n10573), .ZN(n8205) );
  OR2_X1 U10651 ( .A1(n10989), .A2(n10573), .ZN(n8206) );
  NAND2_X1 U10652 ( .A1(n11118), .A2(n8207), .ZN(n11132) );
  INV_X1 U10653 ( .A(n13229), .ZN(n10572) );
  OR2_X1 U10654 ( .A1(n14917), .A2(n10572), .ZN(n9016) );
  NAND2_X1 U10655 ( .A1(n14917), .A2(n10572), .ZN(n9015) );
  INV_X1 U10656 ( .A(n13228), .ZN(n10966) );
  INV_X1 U10657 ( .A(n11176), .ZN(n11180) );
  NAND2_X1 U10658 ( .A1(n11181), .A2(n11180), .ZN(n8209) );
  NAND2_X1 U10659 ( .A1(n11250), .A2(n8826), .ZN(n8208) );
  NAND2_X1 U10660 ( .A1(n8209), .A2(n8208), .ZN(n11259) );
  INV_X1 U10661 ( .A(n11262), .ZN(n11258) );
  NAND2_X1 U10662 ( .A1(n11277), .A2(n10965), .ZN(n8210) );
  XNOR2_X1 U10663 ( .A(n11479), .B(n13225), .ZN(n11345) );
  INV_X1 U10664 ( .A(n13225), .ZN(n11438) );
  INV_X1 U10665 ( .A(n13224), .ZN(n8212) );
  AND2_X1 U10666 ( .A1(n13578), .A2(n8212), .ZN(n8211) );
  OR2_X1 U10667 ( .A1(n13578), .A2(n8212), .ZN(n8213) );
  INV_X1 U10668 ( .A(n13223), .ZN(n11437) );
  NOR2_X1 U10669 ( .A1(n11575), .A2(n11437), .ZN(n9014) );
  AND2_X1 U10670 ( .A1(n11575), .A2(n11437), .ZN(n9013) );
  INV_X1 U10671 ( .A(n9013), .ZN(n8215) );
  INV_X1 U10672 ( .A(n13222), .ZN(n9012) );
  AND2_X1 U10673 ( .A1(n13718), .A2(n9012), .ZN(n8216) );
  OR2_X1 U10674 ( .A1(n14637), .A2(n13139), .ZN(n8218) );
  INV_X1 U10675 ( .A(n13517), .ZN(n13176) );
  NOR2_X1 U10676 ( .A1(n13656), .A2(n13176), .ZN(n8219) );
  INV_X1 U10677 ( .A(n13220), .ZN(n13140) );
  AND2_X1 U10678 ( .A1(n13651), .A2(n13140), .ZN(n8220) );
  INV_X1 U10679 ( .A(n13219), .ZN(n13177) );
  NAND2_X1 U10680 ( .A1(n13647), .A2(n13177), .ZN(n13443) );
  INV_X1 U10681 ( .A(n13218), .ZN(n13121) );
  NAND2_X1 U10682 ( .A1(n13642), .A2(n13121), .ZN(n13445) );
  NAND3_X1 U10683 ( .A1(n13444), .A2(n13443), .A3(n13445), .ZN(n8223) );
  OAI22_X1 U10684 ( .A1(n13636), .A2(n8224), .B1(n13121), .B2(n13642), .ZN(
        n8221) );
  INV_X1 U10685 ( .A(n8221), .ZN(n8222) );
  NAND2_X1 U10686 ( .A1(n8223), .A2(n8222), .ZN(n8226) );
  NAND2_X1 U10687 ( .A1(n13636), .A2(n8224), .ZN(n8225) );
  NAND2_X1 U10688 ( .A1(n8226), .A2(n8225), .ZN(n13417) );
  XNOR2_X1 U10689 ( .A(n13408), .B(n13215), .ZN(n13401) );
  NAND2_X1 U10690 ( .A1(n13402), .A2(n13401), .ZN(n13400) );
  INV_X1 U10691 ( .A(n13215), .ZN(n13149) );
  OR2_X1 U10692 ( .A1(n13408), .A2(n13149), .ZN(n8228) );
  INV_X1 U10693 ( .A(n13214), .ZN(n8229) );
  NAND2_X1 U10694 ( .A1(n13620), .A2(n8229), .ZN(n8230) );
  XNOR2_X1 U10695 ( .A(n13696), .B(n13213), .ZN(n13372) );
  INV_X1 U10696 ( .A(n13213), .ZN(n13191) );
  NAND2_X1 U10697 ( .A1(n13696), .A2(n13191), .ZN(n8231) );
  NAND2_X1 U10698 ( .A1(n8232), .A2(n8231), .ZN(n13357) );
  AND2_X1 U10699 ( .A1(n13361), .A2(n9011), .ZN(n8233) );
  INV_X1 U10700 ( .A(n13189), .ZN(n13211) );
  OR2_X1 U10701 ( .A1(n13689), .A2(n13211), .ZN(n8234) );
  INV_X1 U10702 ( .A(n13096), .ZN(n13210) );
  NAND2_X1 U10703 ( .A1(n7422), .A2(n13210), .ZN(n8235) );
  NAND2_X1 U10704 ( .A1(n13325), .A2(n8235), .ZN(n8237) );
  INV_X1 U10705 ( .A(n9028), .ZN(n8236) );
  XNOR2_X1 U10706 ( .A(n8237), .B(n8236), .ZN(n8246) );
  INV_X1 U10707 ( .A(n6771), .ZN(n9831) );
  NAND2_X1 U10708 ( .A1(n6564), .A2(n9831), .ZN(n8239) );
  OAI21_X2 U10709 ( .B1(n11732), .B2(n13292), .A(n8239), .ZN(n13540) );
  INV_X1 U10710 ( .A(n11732), .ZN(n9009) );
  INV_X1 U10711 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13593) );
  OR2_X1 U10712 ( .A1(n6566), .A2(n13593), .ZN(n8243) );
  INV_X1 U10713 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13308) );
  OR2_X1 U10714 ( .A1(n8182), .A2(n13308), .ZN(n8242) );
  INV_X1 U10715 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13682) );
  OR2_X1 U10716 ( .A1(n7691), .A2(n13682), .ZN(n8241) );
  AND3_X1 U10717 ( .A1(n8243), .A2(n8242), .A3(n8241), .ZN(n8984) );
  NAND2_X1 U10718 ( .A1(n9938), .A2(n9945), .ZN(n13188) );
  INV_X1 U10719 ( .A(n13733), .ZN(n9946) );
  NAND2_X1 U10720 ( .A1(n9946), .A2(P2_B_REG_SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10721 ( .A1(n13516), .A2(n8244), .ZN(n13301) );
  OAI22_X1 U10722 ( .A1(n13096), .A2(n13190), .B1(n8984), .B2(n13301), .ZN(
        n8245) );
  INV_X1 U10723 ( .A(n11575), .ZN(n11572) );
  INV_X1 U10724 ( .A(n11277), .ZN(n11269) );
  NAND2_X1 U10725 ( .A1(n6561), .A2(n11752), .ZN(n11002) );
  OR2_X1 U10726 ( .A1(n11002), .A2(n7671), .ZN(n10268) );
  INV_X1 U10727 ( .A(n10393), .ZN(n11062) );
  INV_X1 U10728 ( .A(n10913), .ZN(n11107) );
  INV_X1 U10729 ( .A(n11250), .ZN(n11184) );
  AND2_X2 U10730 ( .A1(n11185), .A2(n11184), .ZN(n11270) );
  OR2_X2 U10731 ( .A1(n13647), .A2(n13483), .ZN(n13472) );
  INV_X1 U10732 ( .A(n13636), .ZN(n13442) );
  INV_X1 U10733 ( .A(n6564), .ZN(n11406) );
  NAND2_X1 U10734 ( .A1(n13596), .A2(n13327), .ZN(n13298) );
  OAI211_X1 U10735 ( .C1(n13596), .C2(n13327), .A(n13528), .B(n13298), .ZN(
        n13318) );
  INV_X1 U10736 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U10737 ( .A1(n8266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8251) );
  INV_X1 U10738 ( .A(P2_B_REG_SCAN_IN), .ZN(n8252) );
  XNOR2_X1 U10739 ( .A(n11641), .B(n8252), .ZN(n8255) );
  INV_X1 U10740 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8253) );
  NAND2_X1 U10741 ( .A1(n8255), .A2(n11674), .ZN(n8261) );
  NAND2_X1 U10742 ( .A1(n8256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8257) );
  MUX2_X1 U10743 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8257), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8258) );
  INV_X1 U10744 ( .A(n8258), .ZN(n8260) );
  INV_X1 U10745 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15401) );
  INV_X1 U10746 ( .A(n8279), .ZN(n13737) );
  AND2_X1 U10747 ( .A1(n11674), .A2(n13737), .ZN(n8262) );
  AOI21_X1 U10748 ( .B1(n14863), .B2(n15401), .A(n8262), .ZN(n10980) );
  NAND2_X1 U10749 ( .A1(n11641), .A2(n8279), .ZN(n9850) );
  OR2_X1 U10750 ( .A1(n9850), .A2(n11674), .ZN(n8268) );
  INV_X1 U10751 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U10752 ( .A1(n8264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8265) );
  MUX2_X1 U10753 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8265), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8267) );
  NAND2_X1 U10754 ( .A1(n8267), .A2(n8266), .ZN(n9939) );
  NOR2_X1 U10755 ( .A1(n10980), .A2(n14893), .ZN(n14892) );
  NOR4_X1 U10756 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8272) );
  NOR4_X1 U10757 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8271) );
  NOR4_X1 U10758 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n8270) );
  NOR4_X1 U10759 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8269) );
  NAND4_X1 U10760 ( .A1(n8272), .A2(n8271), .A3(n8270), .A4(n8269), .ZN(n8277)
         );
  NOR2_X1 U10761 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .ZN(
        n15213) );
  NOR4_X1 U10762 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n8275) );
  NOR4_X1 U10763 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8274) );
  NOR4_X1 U10764 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8273) );
  NAND4_X1 U10765 ( .A1(n15213), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(n8276) );
  OAI21_X1 U10766 ( .B1(n8277), .B2(n8276), .A(n14863), .ZN(n10978) );
  NAND2_X1 U10767 ( .A1(n13528), .A2(n9002), .ZN(n9840) );
  NAND2_X1 U10768 ( .A1(n6771), .A2(n13292), .ZN(n9835) );
  NAND2_X1 U10769 ( .A1(n9938), .A2(n9835), .ZN(n10977) );
  AND3_X1 U10770 ( .A1(n10978), .A2(n9840), .A3(n10977), .ZN(n8278) );
  AND2_X1 U10771 ( .A1(n14892), .A2(n8278), .ZN(n10387) );
  INV_X1 U10772 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14889) );
  NAND2_X1 U10773 ( .A1(n14863), .A2(n14889), .ZN(n8281) );
  OR2_X1 U10774 ( .A1(n11641), .A2(n8279), .ZN(n8280) );
  INV_X2 U10775 ( .A(n14924), .ZN(n14908) );
  NAND2_X1 U10776 ( .A1(n11744), .A2(n9835), .ZN(n14902) );
  NAND2_X1 U10777 ( .A1(n14908), .A2(n14918), .ZN(n13702) );
  NAND2_X1 U10778 ( .A1(n13316), .A2(n8282), .ZN(n8283) );
  NOR2_X1 U10779 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8287) );
  NAND4_X1 U10780 ( .A1(n8287), .A2(n8286), .A3(n8368), .A4(n8285), .ZN(n8288)
         );
  NOR2_X1 U10781 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8292) );
  NOR2_X1 U10782 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n8291) );
  NOR2_X1 U10783 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8294) );
  NAND4_X1 U10784 ( .A1(n8654), .A2(n8294), .A3(n8653), .A4(n8656), .ZN(n8719)
         );
  NAND3_X1 U10785 ( .A1(n7058), .A2(n8514), .A3(n8295), .ZN(n8296) );
  INV_X1 U10786 ( .A(n8300), .ZN(n14373) );
  NAND2_X1 U10787 ( .A1(n6545), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10788 ( .A1(n8347), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10789 ( .A1(n8349), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U10790 ( .A1(n8346), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8304) );
  AND4_X2 U10791 ( .A1(n8307), .A2(n8306), .A3(n8305), .A4(n8304), .ZN(n8675)
         );
  NAND2_X1 U10792 ( .A1(n8312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8314) );
  OR2_X1 U10793 ( .A1(n8315), .A2(n14371), .ZN(n8317) );
  NAND2_X2 U10794 ( .A1(n9853), .A2(n9902), .ZN(n8413) );
  OR2_X1 U10795 ( .A1(n8413), .A2(n6656), .ZN(n8318) );
  NAND2_X1 U10796 ( .A1(n8347), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8325) );
  NAND2_X1 U10797 ( .A1(n8346), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U10798 ( .A1(n8349), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8323) );
  INV_X1 U10799 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8320) );
  INV_X1 U10800 ( .A(n8321), .ZN(n8322) );
  NAND2_X1 U10801 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8326) );
  INV_X1 U10802 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9871) );
  OR2_X1 U10803 ( .A1(n8413), .A2(n9916), .ZN(n8327) );
  OAI211_X1 U10804 ( .C1(n9853), .C2(n9870), .A(n8328), .B(n8327), .ZN(n8662)
         );
  NOR2_X1 U10805 ( .A1(n7607), .A2(n7609), .ZN(n8332) );
  NAND2_X1 U10806 ( .A1(n8349), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10807 ( .A1(n8346), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8330) );
  NOR2_X1 U10808 ( .A1(n6568), .A2(n8333), .ZN(n8334) );
  XNOR2_X1 U10809 ( .A(n8334), .B(n9189), .ZN(n14394) );
  MUX2_X1 U10810 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14394), .S(n9853), .Z(n12209)
         );
  NAND2_X1 U10811 ( .A1(n8672), .A2(n12209), .ZN(n11761) );
  NAND2_X1 U10812 ( .A1(n10711), .A2(n11771), .ZN(n10680) );
  INV_X1 U10813 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10814 ( .A1(n6545), .A2(n8336), .ZN(n8340) );
  NAND2_X1 U10815 ( .A1(n8347), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U10816 ( .A1(n8349), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10817 ( .A1(n8346), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10818 ( .A1(n8341), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8342) );
  XNOR2_X1 U10819 ( .A(n8342), .B(n8284), .ZN(n10204) );
  OR2_X1 U10820 ( .A1(n8356), .A2(n15396), .ZN(n8345) );
  INV_X1 U10821 ( .A(n8343), .ZN(n9905) );
  NAND2_X1 U10822 ( .A1(n11232), .A2(n10685), .ZN(n11777) );
  INV_X1 U10823 ( .A(n11232), .ZN(n13957) );
  NAND2_X1 U10824 ( .A1(n13957), .A2(n10846), .ZN(n11776) );
  AND2_X1 U10825 ( .A1(n11777), .A2(n11776), .ZN(n11937) );
  NAND2_X1 U10826 ( .A1(n10680), .A2(n11937), .ZN(n10679) );
  NAND2_X1 U10827 ( .A1(n8668), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10828 ( .A1(n8669), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8352) );
  AND2_X1 U10829 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8361) );
  NOR2_X1 U10830 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8348) );
  NOR2_X1 U10831 ( .A1(n8361), .A2(n8348), .ZN(n11229) );
  NAND2_X1 U10832 ( .A1(n6546), .A2(n11229), .ZN(n8351) );
  NAND2_X1 U10833 ( .A1(n11903), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8350) );
  AND4_X2 U10834 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n11782)
         );
  NAND2_X1 U10835 ( .A1(n8354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8355) );
  XNOR2_X1 U10836 ( .A(n8355), .B(n8368), .ZN(n10488) );
  INV_X2 U10837 ( .A(n8413), .ZN(n8371) );
  NAND2_X1 U10838 ( .A1(n8371), .A2(n9894), .ZN(n8358) );
  OR2_X1 U10839 ( .A1(n8356), .A2(n9895), .ZN(n8357) );
  OAI211_X1 U10840 ( .C1(n9853), .C2(n10488), .A(n8358), .B(n8357), .ZN(n11783) );
  NAND2_X1 U10841 ( .A1(n11782), .A2(n11783), .ZN(n8360) );
  NAND2_X1 U10842 ( .A1(n13956), .A2(n14774), .ZN(n8359) );
  NAND2_X1 U10843 ( .A1(n8669), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10844 ( .A1(n11903), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8366) );
  AND2_X1 U10845 ( .A1(n8361), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8382) );
  NOR2_X1 U10846 ( .A1(n8361), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8362) );
  NOR2_X1 U10847 ( .A1(n8382), .A2(n8362), .ZN(n11219) );
  NAND2_X1 U10848 ( .A1(n6546), .A2(n11219), .ZN(n8365) );
  NAND2_X1 U10849 ( .A1(n8668), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8364) );
  INV_X1 U10850 ( .A(n8354), .ZN(n8369) );
  NAND2_X1 U10851 ( .A1(n8369), .A2(n8368), .ZN(n8376) );
  NAND2_X1 U10852 ( .A1(n8376), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8370) );
  XNOR2_X1 U10853 ( .A(n8370), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U10854 ( .A1(n8538), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8537), .B2(
        n10246), .ZN(n8373) );
  NAND2_X1 U10855 ( .A1(n9899), .A2(n8371), .ZN(n8372) );
  NAND2_X1 U10856 ( .A1(n8373), .A2(n8372), .ZN(n11789) );
  NAND2_X1 U10857 ( .A1(n11787), .A2(n11789), .ZN(n8375) );
  INV_X1 U10858 ( .A(n11787), .ZN(n13955) );
  NAND2_X1 U10859 ( .A1(n13955), .A2(n11788), .ZN(n8374) );
  NAND2_X1 U10860 ( .A1(n10773), .A2(n8375), .ZN(n11033) );
  NAND2_X1 U10861 ( .A1(n9918), .A2(n8371), .ZN(n8381) );
  INV_X1 U10862 ( .A(n8376), .ZN(n8378) );
  INV_X1 U10863 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10864 ( .A1(n8378), .A2(n8377), .ZN(n8389) );
  NAND2_X1 U10865 ( .A1(n8389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U10866 ( .A(n8379), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U10867 ( .A1(n8538), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8537), .B2(
        n10421), .ZN(n8380) );
  NAND2_X1 U10868 ( .A1(n8668), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8386) );
  INV_X2 U10869 ( .A(n8581), .ZN(n8669) );
  NAND2_X1 U10870 ( .A1(n8669), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10871 ( .A1(n8382), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8394) );
  OAI21_X1 U10872 ( .B1(n8382), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8394), .ZN(
        n11376) );
  INV_X1 U10873 ( .A(n11376), .ZN(n11041) );
  NAND2_X1 U10874 ( .A1(n6546), .A2(n11041), .ZN(n8384) );
  NAND2_X1 U10875 ( .A1(n11903), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8383) );
  NAND4_X1 U10876 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n13954) );
  NAND2_X1 U10877 ( .A1(n14779), .A2(n13954), .ZN(n8387) );
  NAND2_X1 U10878 ( .A1(n11456), .A2(n11795), .ZN(n8388) );
  NAND2_X1 U10879 ( .A1(n9923), .A2(n8371), .ZN(n8392) );
  NAND2_X1 U10880 ( .A1(n8401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10881 ( .A(n8390), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U10882 ( .A1(n8538), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8537), .B2(
        n10433), .ZN(n8391) );
  NAND2_X1 U10883 ( .A1(n8668), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U10884 ( .A1(n8669), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8398) );
  INV_X1 U10885 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8393) );
  AND2_X1 U10886 ( .A1(n8394), .A2(n8393), .ZN(n8395) );
  NOR2_X1 U10887 ( .A1(n8405), .A2(n8395), .ZN(n11453) );
  NAND2_X1 U10888 ( .A1(n6546), .A2(n11453), .ZN(n8397) );
  NAND2_X1 U10889 ( .A1(n11903), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8396) );
  NAND4_X1 U10890 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8396), .ZN(n13953) );
  XNOR2_X1 U10891 ( .A(n11799), .B(n13953), .ZN(n11942) );
  INV_X1 U10892 ( .A(n13953), .ZN(n11377) );
  NAND2_X1 U10893 ( .A1(n11799), .A2(n11377), .ZN(n8400) );
  OR2_X1 U10894 ( .A1(n9931), .A2(n8413), .ZN(n8404) );
  OAI21_X1 U10895 ( .B1(n8401), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8402) );
  XNOR2_X1 U10896 ( .A(n8402), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U10897 ( .A1(n8538), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8537), .B2(
        n10315), .ZN(n8403) );
  NAND2_X1 U10898 ( .A1(n8668), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10899 ( .A1(n8669), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10900 ( .A1(n8405), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10901 ( .A1(n8405), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8406) );
  AND2_X1 U10902 ( .A1(n8423), .A2(n8406), .ZN(n11629) );
  NAND2_X1 U10903 ( .A1(n6546), .A2(n11629), .ZN(n8408) );
  NAND2_X1 U10904 ( .A1(n11903), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8407) );
  XNOR2_X1 U10905 ( .A(n11806), .B(n11719), .ZN(n11158) );
  NAND2_X1 U10906 ( .A1(n11160), .A2(n8411), .ZN(n11159) );
  OR2_X1 U10907 ( .A1(n11806), .A2(n11719), .ZN(n8412) );
  NAND2_X1 U10908 ( .A1(n11159), .A2(n8412), .ZN(n11306) );
  INV_X1 U10909 ( .A(n11306), .ZN(n8430) );
  OR2_X1 U10910 ( .A1(n9937), .A2(n8413), .ZN(n8421) );
  NOR2_X1 U10911 ( .A1(n8417), .A2(n14371), .ZN(n8415) );
  MUX2_X1 U10912 ( .A(n14371), .B(n8415), .S(P1_IR_REG_9__SCAN_IN), .Z(n8419)
         );
  INV_X1 U10913 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10914 ( .A1(n8417), .A2(n8416), .ZN(n8433) );
  INV_X1 U10915 ( .A(n8433), .ZN(n8418) );
  AOI22_X1 U10916 ( .A1(n8538), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8537), .B2(
        n10582), .ZN(n8420) );
  NAND2_X1 U10917 ( .A1(n8669), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10918 ( .A1(n11903), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U10919 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  AND2_X1 U10920 ( .A1(n8447), .A2(n8424), .ZN(n11722) );
  NAND2_X1 U10921 ( .A1(n6546), .A2(n11722), .ZN(n8426) );
  NAND2_X1 U10922 ( .A1(n8668), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8425) );
  XNOR2_X1 U10923 ( .A(n11810), .B(n13774), .ZN(n11946) );
  INV_X1 U10924 ( .A(n11946), .ZN(n8429) );
  NAND2_X1 U10925 ( .A1(n11810), .A2(n13774), .ZN(n8431) );
  NAND2_X1 U10926 ( .A1(n10088), .A2(n8371), .ZN(n8436) );
  NAND2_X1 U10927 ( .A1(n8433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8432) );
  MUX2_X1 U10928 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8432), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n8434) );
  AOI22_X1 U10929 ( .A1(n8538), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8537), 
        .B2(n10760), .ZN(n8435) );
  XNOR2_X1 U10930 ( .A(n8447), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n13777) );
  NAND2_X1 U10931 ( .A1(n6546), .A2(n13777), .ZN(n8440) );
  NAND2_X1 U10932 ( .A1(n8669), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10933 ( .A1(n11903), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10934 ( .A1(n8668), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8437) );
  XNOR2_X1 U10935 ( .A(n13768), .B(n12219), .ZN(n11947) );
  OR2_X1 U10936 ( .A1(n13768), .A2(n12219), .ZN(n8441) );
  NAND2_X1 U10937 ( .A1(n10129), .A2(n8371), .ZN(n8444) );
  NAND2_X1 U10938 ( .A1(n8454), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8442) );
  XNOR2_X1 U10939 ( .A(n8442), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U10940 ( .A1(n8538), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8537), 
        .B2(n10952), .ZN(n8443) );
  NAND2_X1 U10941 ( .A1(n8668), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10942 ( .A1(n8669), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8451) );
  INV_X1 U10943 ( .A(n8447), .ZN(n8445) );
  AOI21_X1 U10944 ( .B1(n8445), .B2(P1_REG3_REG_10__SCAN_IN), .A(
        P1_REG3_REG_11__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U10945 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8446) );
  OR2_X1 U10946 ( .A1(n8448), .A2(n8457), .ZN(n13888) );
  INV_X1 U10947 ( .A(n13888), .ZN(n11517) );
  NAND2_X1 U10948 ( .A1(n6546), .A2(n11517), .ZN(n8450) );
  NAND2_X1 U10949 ( .A1(n11903), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8449) );
  NOR2_X1 U10950 ( .A1(n13896), .A2(n13804), .ZN(n8453) );
  NAND2_X1 U10951 ( .A1(n10134), .A2(n8371), .ZN(n8456) );
  NAND2_X1 U10952 ( .A1(n8494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8465) );
  XNOR2_X1 U10953 ( .A(n8465), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U10954 ( .A1(n8538), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8537), 
        .B2(n13978), .ZN(n8455) );
  NAND2_X1 U10955 ( .A1(n8669), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10956 ( .A1(n8668), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8461) );
  NOR2_X1 U10957 ( .A1(n8457), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8458) );
  OR2_X1 U10958 ( .A1(n8472), .A2(n8458), .ZN(n14527) );
  INV_X1 U10959 ( .A(n14527), .ZN(n13809) );
  NAND2_X1 U10960 ( .A1(n6546), .A2(n13809), .ZN(n8460) );
  NAND2_X1 U10961 ( .A1(n11903), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8459) );
  OR2_X1 U10962 ( .A1(n12233), .A2(n12231), .ZN(n8464) );
  NAND2_X1 U10963 ( .A1(n12233), .A2(n12231), .ZN(n8463) );
  NAND2_X1 U10964 ( .A1(n8464), .A2(n8463), .ZN(n14519) );
  NAND2_X1 U10965 ( .A1(n10155), .A2(n8371), .ZN(n8471) );
  INV_X1 U10966 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U10967 ( .A1(n8465), .A2(n8491), .ZN(n8466) );
  NAND2_X1 U10968 ( .A1(n8466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8468) );
  INV_X1 U10969 ( .A(n8468), .ZN(n8467) );
  NAND2_X1 U10970 ( .A1(n8467), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n8469) );
  INV_X1 U10971 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U10972 ( .A1(n8468), .A2(n8492), .ZN(n8479) );
  AOI22_X1 U10973 ( .A1(n8538), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8537), 
        .B2(n14681), .ZN(n8470) );
  NAND2_X1 U10974 ( .A1(n8669), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U10975 ( .A1(n11903), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10976 ( .A1(n8472), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8484) );
  OR2_X1 U10977 ( .A1(n8472), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8473) );
  AND2_X1 U10978 ( .A1(n8484), .A2(n8473), .ZN(n13864) );
  NAND2_X1 U10979 ( .A1(n6546), .A2(n13864), .ZN(n8475) );
  NAND2_X1 U10980 ( .A1(n8668), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8474) );
  NAND4_X1 U10981 ( .A1(n8477), .A2(n8476), .A3(n8475), .A4(n8474), .ZN(n13947) );
  XNOR2_X1 U10982 ( .A(n13868), .B(n13947), .ZN(n11951) );
  INV_X1 U10983 ( .A(n13947), .ZN(n13751) );
  OR2_X1 U10984 ( .A1(n13868), .A2(n13751), .ZN(n8478) );
  NAND2_X1 U10985 ( .A1(n11647), .A2(n8478), .ZN(n11690) );
  NAND2_X1 U10986 ( .A1(n10462), .A2(n8371), .ZN(n8482) );
  NAND2_X1 U10987 ( .A1(n8479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U10988 ( .A(n8480), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U10989 ( .A1(n8538), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8537), 
        .B2(n13980), .ZN(n8481) );
  NAND2_X1 U10990 ( .A1(n8668), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10991 ( .A1(n8669), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8488) );
  INV_X1 U10992 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10993 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  AND2_X1 U10994 ( .A1(n8508), .A2(n8485), .ZN(n13749) );
  NAND2_X1 U10995 ( .A1(n6546), .A2(n13749), .ZN(n8487) );
  NAND2_X1 U10996 ( .A1(n11903), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10997 ( .A1(n14329), .A2(n13929), .ZN(n11838) );
  NAND2_X1 U10998 ( .A1(n10670), .A2(n8371), .ZN(n8498) );
  INV_X1 U10999 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8490) );
  NAND3_X1 U11000 ( .A1(n8492), .A2(n8491), .A3(n8490), .ZN(n8493) );
  OAI21_X1 U11001 ( .B1(n8494), .B2(n8493), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8495) );
  INV_X1 U11002 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n15309) );
  XNOR2_X1 U11003 ( .A(n8495), .B(n15309), .ZN(n14710) );
  INV_X1 U11004 ( .A(n14710), .ZN(n8496) );
  AOI22_X1 U11005 ( .A1(n8538), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8537), 
        .B2(n8496), .ZN(n8497) );
  NAND2_X1 U11006 ( .A1(n8668), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U11007 ( .A1(n8669), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8501) );
  XNOR2_X1 U11008 ( .A(n8508), .B(P1_REG3_REG_15__SCAN_IN), .ZN(n14223) );
  NAND2_X1 U11009 ( .A1(n6546), .A2(n14223), .ZN(n8500) );
  NAND2_X1 U11010 ( .A1(n11903), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U11011 ( .A1(n14320), .A2(n14213), .ZN(n11843) );
  NAND2_X1 U11012 ( .A1(n11844), .A2(n11843), .ZN(n11953) );
  NAND2_X1 U11013 ( .A1(n10701), .A2(n8371), .ZN(n8505) );
  OR2_X1 U11014 ( .A1(n8515), .A2(n14371), .ZN(n8503) );
  XNOR2_X1 U11015 ( .A(n8503), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14725) );
  AOI22_X1 U11016 ( .A1(n8538), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8537), 
        .B2(n14725), .ZN(n8504) );
  NAND2_X1 U11017 ( .A1(n8668), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U11018 ( .A1(n8669), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8512) );
  INV_X1 U11019 ( .A(n8508), .ZN(n8506) );
  AOI21_X1 U11020 ( .B1(n8506), .B2(P1_REG3_REG_15__SCAN_IN), .A(
        P1_REG3_REG_16__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U11021 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n8507) );
  OR2_X1 U11022 ( .A1(n8509), .A2(n8519), .ZN(n14204) );
  INV_X1 U11023 ( .A(n14204), .ZN(n13828) );
  NAND2_X1 U11024 ( .A1(n6546), .A2(n13828), .ZN(n8511) );
  NAND2_X1 U11025 ( .A1(n11903), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8510) );
  XNOR2_X1 U11026 ( .A(n14206), .B(n13928), .ZN(n14208) );
  NAND2_X1 U11027 ( .A1(n10828), .A2(n8371), .ZN(n8518) );
  NAND2_X1 U11028 ( .A1(n8525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8516) );
  XNOR2_X1 U11029 ( .A(n8516), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U11030 ( .A1(n8538), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8537), 
        .B2(n13984), .ZN(n8517) );
  NAND2_X1 U11031 ( .A1(n8668), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U11032 ( .A1(n8669), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U11033 ( .A1(n8519), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8543) );
  OR2_X1 U11034 ( .A1(n8519), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8520) );
  AND2_X1 U11035 ( .A1(n8543), .A2(n8520), .ZN(n14195) );
  NAND2_X1 U11036 ( .A1(n6546), .A2(n14195), .ZN(n8522) );
  NAND2_X1 U11037 ( .A1(n11903), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8521) );
  XNOR2_X1 U11038 ( .A(n14310), .B(n14211), .ZN(n11850) );
  NAND2_X1 U11039 ( .A1(n14188), .A2(n14189), .ZN(n14187) );
  OR2_X1 U11040 ( .A1(n14310), .A2(n14211), .ZN(n11849) );
  NAND2_X1 U11041 ( .A1(n14187), .A2(n11849), .ZN(n14170) );
  NAND2_X1 U11042 ( .A1(n11201), .A2(n8371), .ZN(n8529) );
  NAND2_X1 U11043 ( .A1(n8720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8526) );
  INV_X1 U11044 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8652) );
  XNOR2_X1 U11045 ( .A(n8526), .B(n8652), .ZN(n14756) );
  INV_X1 U11046 ( .A(n14756), .ZN(n8527) );
  AOI22_X1 U11047 ( .A1(n8538), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8537), 
        .B2(n8527), .ZN(n8528) );
  NAND2_X1 U11048 ( .A1(n8668), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11049 ( .A1(n8669), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8532) );
  XNOR2_X1 U11050 ( .A(n8543), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U11051 ( .A1(n6546), .A2(n14178), .ZN(n8531) );
  NAND2_X1 U11052 ( .A1(n11903), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8530) );
  NAND4_X1 U11053 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n14163) );
  XNOR2_X1 U11054 ( .A(n14304), .B(n14163), .ZN(n14182) );
  INV_X1 U11055 ( .A(n14163), .ZN(n13786) );
  OR2_X1 U11056 ( .A1(n14304), .A2(n13786), .ZN(n8534) );
  NAND2_X1 U11057 ( .A1(n11296), .A2(n8371), .ZN(n8540) );
  XNOR2_X2 U11058 ( .A(n8536), .B(P1_IR_REG_19__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U11059 ( .A1(n8538), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11760), 
        .B2(n8537), .ZN(n8539) );
  INV_X1 U11060 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8542) );
  INV_X1 U11061 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8541) );
  OAI21_X1 U11062 ( .B1(n8543), .B2(n8542), .A(n8541), .ZN(n8544) );
  AND2_X1 U11063 ( .A1(n8544), .A2(n8551), .ZN(n14157) );
  NAND2_X1 U11064 ( .A1(n14157), .A2(n6546), .ZN(n8548) );
  NAND2_X1 U11065 ( .A1(n8669), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U11066 ( .A1(n11903), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11067 ( .A1(n8668), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8545) );
  XNOR2_X1 U11068 ( .A(n14298), .B(n13902), .ZN(n11956) );
  INV_X1 U11069 ( .A(n11956), .ZN(n14161) );
  NAND2_X1 U11070 ( .A1(n14298), .A2(n13902), .ZN(n11865) );
  NAND2_X1 U11071 ( .A1(n11300), .A2(n8371), .ZN(n8550) );
  INV_X1 U11072 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11301) );
  OR2_X1 U11073 ( .A1(n8356), .A2(n11301), .ZN(n8549) );
  INV_X1 U11074 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n15252) );
  AND2_X1 U11075 ( .A1(n8551), .A2(n15252), .ZN(n8552) );
  OR2_X1 U11076 ( .A1(n8552), .A2(n8557), .ZN(n14143) );
  AOI22_X1 U11077 ( .A1(n8669), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n11903), 
        .B2(P1_REG0_REG_20__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U11078 ( .A1(n8668), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8553) );
  OAI211_X1 U11079 ( .C1(n14143), .C2(n8578), .A(n8554), .B(n8553), .ZN(n14164) );
  INV_X1 U11080 ( .A(n14164), .ZN(n13785) );
  XNOR2_X1 U11081 ( .A(n14292), .B(n13785), .ZN(n11957) );
  NAND2_X1 U11082 ( .A1(n11405), .A2(n8371), .ZN(n8556) );
  INV_X1 U11083 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11408) );
  OR2_X1 U11084 ( .A1(n8356), .A2(n11408), .ZN(n8555) );
  NOR2_X1 U11085 ( .A1(n8557), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8558) );
  OR2_X1 U11086 ( .A1(n8566), .A2(n8558), .ZN(n14124) );
  AOI22_X1 U11087 ( .A1(n8668), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n8669), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U11088 ( .A1(n11903), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8559) );
  OAI211_X1 U11089 ( .C1(n14124), .C2(n8578), .A(n8560), .B(n8559), .ZN(n14140) );
  OR2_X1 U11090 ( .A1(n14288), .A2(n14140), .ZN(n8701) );
  NAND2_X1 U11091 ( .A1(n14288), .A2(n14140), .ZN(n8561) );
  NAND2_X1 U11092 ( .A1(n8701), .A2(n8561), .ZN(n14129) );
  NAND2_X1 U11093 ( .A1(n14119), .A2(n14129), .ZN(n8563) );
  INV_X1 U11094 ( .A(n14140), .ZN(n13857) );
  OR2_X1 U11095 ( .A1(n14288), .A2(n13857), .ZN(n8562) );
  NAND2_X1 U11096 ( .A1(n8563), .A2(n8562), .ZN(n14107) );
  OR2_X1 U11097 ( .A1(n8564), .A2(n6568), .ZN(n8565) );
  XNOR2_X1 U11098 ( .A(n8565), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14392) );
  OR2_X1 U11099 ( .A1(n8566), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U11100 ( .A1(n8575), .A2(n8567), .ZN(n14114) );
  AOI22_X1 U11101 ( .A1(n8668), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n8669), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U11102 ( .A1(n11903), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U11103 ( .C1(n14114), .C2(n8578), .A(n8569), .B(n8568), .ZN(n14092) );
  OR2_X1 U11104 ( .A1(n13882), .A2(n14092), .ZN(n8572) );
  NAND2_X1 U11105 ( .A1(n13882), .A2(n14092), .ZN(n8570) );
  NAND2_X1 U11106 ( .A1(n8572), .A2(n8570), .ZN(n14108) );
  NAND2_X1 U11107 ( .A1(n11636), .A2(n8371), .ZN(n8574) );
  OR2_X1 U11108 ( .A1(n8356), .A2(n11635), .ZN(n8573) );
  NAND2_X2 U11109 ( .A1(n8574), .A2(n8573), .ZN(n14276) );
  INV_X1 U11110 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15336) );
  NAND2_X1 U11111 ( .A1(n8575), .A2(n15336), .ZN(n8577) );
  INV_X1 U11112 ( .A(n8588), .ZN(n8576) );
  NAND2_X1 U11113 ( .A1(n8577), .A2(n8576), .ZN(n14096) );
  OR2_X1 U11114 ( .A1(n14096), .A2(n8578), .ZN(n8584) );
  INV_X1 U11115 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14097) );
  NAND2_X1 U11116 ( .A1(n11903), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U11117 ( .A1(n8668), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8579) );
  OAI211_X1 U11118 ( .C1(n8581), .C2(n14097), .A(n8580), .B(n8579), .ZN(n8582)
         );
  INV_X1 U11119 ( .A(n8582), .ZN(n8583) );
  NAND2_X1 U11120 ( .A1(n8584), .A2(n8583), .ZN(n14072) );
  XNOR2_X1 U11121 ( .A(n14276), .B(n14072), .ZN(n14100) );
  INV_X1 U11122 ( .A(n14072), .ZN(n13850) );
  NAND2_X1 U11123 ( .A1(n14276), .A2(n13850), .ZN(n8585) );
  NAND2_X1 U11124 ( .A1(n14090), .A2(n8585), .ZN(n14068) );
  INV_X1 U11125 ( .A(n14068), .ZN(n8594) );
  NAND2_X1 U11126 ( .A1(n11640), .A2(n8371), .ZN(n8587) );
  INV_X1 U11127 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11643) );
  OR2_X1 U11128 ( .A1(n8356), .A2(n11643), .ZN(n8586) );
  NAND2_X1 U11129 ( .A1(n8668), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11130 ( .A1(n8669), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11131 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n8588), .ZN(n8598) );
  OAI21_X1 U11132 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8588), .A(n8598), .ZN(
        n13849) );
  INV_X1 U11133 ( .A(n13849), .ZN(n14083) );
  NAND2_X1 U11134 ( .A1(n6546), .A2(n14083), .ZN(n8590) );
  NAND2_X1 U11135 ( .A1(n11903), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U11136 ( .A(n14266), .B(n13817), .ZN(n14067) );
  NAND2_X1 U11137 ( .A1(n8594), .A2(n8593), .ZN(n14070) );
  OR2_X1 U11138 ( .A1(n14266), .A2(n13817), .ZN(n8595) );
  NAND2_X1 U11139 ( .A1(n11671), .A2(n8371), .ZN(n8597) );
  OR2_X1 U11140 ( .A1(n8356), .A2(n11672), .ZN(n8596) );
  NAND2_X1 U11141 ( .A1(n8669), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11142 ( .A1(n11903), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8603) );
  INV_X1 U11143 ( .A(n8598), .ZN(n8599) );
  NAND2_X1 U11144 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8599), .ZN(n8609) );
  OAI21_X1 U11145 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8599), .A(n8609), .ZN(
        n14060) );
  INV_X1 U11146 ( .A(n14060), .ZN(n8600) );
  NAND2_X1 U11147 ( .A1(n6546), .A2(n8600), .ZN(n8602) );
  NAND2_X1 U11148 ( .A1(n8668), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U11149 ( .A(n14259), .B(n13914), .ZN(n11960) );
  NAND2_X1 U11150 ( .A1(n14259), .A2(n13914), .ZN(n8605) );
  NAND2_X1 U11151 ( .A1(n13735), .A2(n8371), .ZN(n8607) );
  OR2_X1 U11152 ( .A1(n8356), .A2(n14388), .ZN(n8606) );
  NAND2_X1 U11153 ( .A1(n8668), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11154 ( .A1(n8669), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8613) );
  INV_X1 U11155 ( .A(n8609), .ZN(n8608) );
  NAND2_X1 U11156 ( .A1(n8608), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8620) );
  INV_X1 U11157 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13917) );
  NAND2_X1 U11158 ( .A1(n8609), .A2(n13917), .ZN(n8610) );
  AND2_X1 U11159 ( .A1(n8620), .A2(n8610), .ZN(n14046) );
  NAND2_X1 U11160 ( .A1(n6545), .A2(n14046), .ZN(n8612) );
  NAND2_X1 U11161 ( .A1(n11903), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8611) );
  OR2_X1 U11162 ( .A1(n12347), .A2(n13818), .ZN(n8615) );
  NAND2_X1 U11163 ( .A1(n13732), .A2(n8371), .ZN(n8617) );
  OR2_X1 U11164 ( .A1(n8356), .A2(n14385), .ZN(n8616) );
  NAND2_X1 U11165 ( .A1(n8668), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11166 ( .A1(n8669), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8624) );
  INV_X1 U11167 ( .A(n8620), .ZN(n8618) );
  NAND2_X1 U11168 ( .A1(n8618), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8638) );
  INV_X1 U11169 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11170 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NAND2_X1 U11171 ( .A1(n6546), .A2(n14028), .ZN(n8623) );
  NAND2_X1 U11172 ( .A1(n11903), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8622) );
  NAND4_X1 U11173 ( .A1(n8625), .A2(n8624), .A3(n8623), .A4(n8622), .ZN(n13943) );
  NAND2_X1 U11174 ( .A1(n14024), .A2(n14034), .ZN(n8627) );
  INV_X1 U11175 ( .A(n13943), .ZN(n12372) );
  NAND2_X1 U11176 ( .A1(n14248), .A2(n12372), .ZN(n8626) );
  NAND2_X1 U11177 ( .A1(n8627), .A2(n8626), .ZN(n14007) );
  NAND2_X1 U11178 ( .A1(n13728), .A2(n8371), .ZN(n8629) );
  INV_X1 U11179 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11726) );
  OR2_X1 U11180 ( .A1(n8356), .A2(n11726), .ZN(n8628) );
  NAND2_X2 U11181 ( .A1(n8629), .A2(n8628), .ZN(n14243) );
  NAND2_X1 U11182 ( .A1(n8668), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11183 ( .A1(n8669), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8632) );
  XNOR2_X1 U11184 ( .A(n8638), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U11185 ( .A1(n6546), .A2(n12370), .ZN(n8631) );
  NAND2_X1 U11186 ( .A1(n11903), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8630) );
  AND2_X1 U11187 ( .A1(n14243), .A2(n13741), .ZN(n8634) );
  NAND2_X1 U11188 ( .A1(n12194), .A2(n8371), .ZN(n8636) );
  OR2_X1 U11189 ( .A1(n8356), .A2(n14381), .ZN(n8635) );
  NAND2_X2 U11190 ( .A1(n8636), .A2(n8635), .ZN(n11912) );
  NAND2_X1 U11191 ( .A1(n8668), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11192 ( .A1(n8669), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8642) );
  INV_X1 U11193 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8637) );
  NOR2_X1 U11194 ( .A1(n8638), .A2(n8637), .ZN(n12196) );
  NAND2_X1 U11195 ( .A1(n6546), .A2(n12196), .ZN(n8641) );
  NAND2_X1 U11196 ( .A1(n11903), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8640) );
  XNOR2_X1 U11197 ( .A(n11912), .B(n12371), .ZN(n8711) );
  XNOR2_X1 U11198 ( .A(n8644), .B(n8711), .ZN(n8661) );
  NAND2_X1 U11199 ( .A1(n8651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U11200 ( .A1(n6611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8649) );
  MUX2_X1 U11201 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8649), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8650) );
  INV_X1 U11202 ( .A(n11925), .ZN(n11929) );
  NAND2_X1 U11203 ( .A1(n8713), .A2(n11929), .ZN(n8659) );
  NAND3_X1 U11204 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n8655) );
  NAND2_X1 U11205 ( .A1(n11760), .A2(n14393), .ZN(n8658) );
  NAND2_X2 U11206 ( .A1(n8659), .A2(n8658), .ZN(n14522) );
  AND2_X1 U11207 ( .A1(n13942), .A2(n14174), .ZN(n8660) );
  OR2_X1 U11208 ( .A1(n8662), .A2(n12209), .ZN(n10723) );
  NOR2_X1 U11209 ( .A1(n10723), .A2(n6552), .ZN(n10722) );
  AND2_X1 U11210 ( .A1(n10722), .A2(n10846), .ZN(n10838) );
  INV_X1 U11211 ( .A(n11806), .ZN(n11632) );
  NAND2_X1 U11212 ( .A1(n11161), .A2(n11725), .ZN(n11525) );
  OR2_X1 U11213 ( .A1(n14310), .A2(n14203), .ZN(n14192) );
  OR2_X1 U11214 ( .A1(n14304), .A2(n14192), .ZN(n14176) );
  NOR2_X1 U11215 ( .A1(n14081), .A2(n14259), .ZN(n14056) );
  NAND2_X1 U11216 ( .A1(n14056), .A2(n14350), .ZN(n14045) );
  NOR2_X2 U11217 ( .A1(n14045), .A2(n14248), .ZN(n14017) );
  AOI21_X1 U11218 ( .B1(n11912), .B2(n14018), .A(n14252), .ZN(n8666) );
  NAND2_X1 U11219 ( .A1(n8666), .A2(n13996), .ZN(n12203) );
  AND2_X1 U11220 ( .A1(n7145), .A2(P1_B_REG_SCAN_IN), .ZN(n8667) );
  NOR2_X1 U11221 ( .A1(n14210), .A2(n8667), .ZN(n13998) );
  INV_X1 U11222 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U11223 ( .A1(n8669), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11224 ( .A1(n11903), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8670) );
  OAI211_X1 U11225 ( .C1(n8363), .C2(n14240), .A(n8671), .B(n8670), .ZN(n13940) );
  NAND2_X1 U11226 ( .A1(n13998), .A2(n13940), .ZN(n12198) );
  NAND2_X1 U11227 ( .A1(n13961), .A2(n12209), .ZN(n10454) );
  NAND2_X1 U11228 ( .A1(n11759), .A2(n10454), .ZN(n8674) );
  NAND2_X1 U11229 ( .A1(n12212), .A2(n11023), .ZN(n8673) );
  NAND2_X1 U11230 ( .A1(n8675), .A2(n14766), .ZN(n8676) );
  NAND2_X1 U11231 ( .A1(n10708), .A2(n8676), .ZN(n10678) );
  INV_X1 U11232 ( .A(n11937), .ZN(n10677) );
  NAND2_X1 U11233 ( .A1(n11232), .A2(n10846), .ZN(n8677) );
  NAND2_X1 U11234 ( .A1(n10676), .A2(n8677), .ZN(n10837) );
  NAND2_X1 U11235 ( .A1(n11782), .A2(n14774), .ZN(n11778) );
  INV_X1 U11236 ( .A(n10775), .ZN(n11940) );
  NAND2_X1 U11237 ( .A1(n11787), .A2(n11788), .ZN(n8678) );
  NAND2_X1 U11238 ( .A1(n10769), .A2(n8678), .ZN(n11029) );
  INV_X1 U11239 ( .A(n11944), .ZN(n11028) );
  NAND2_X1 U11240 ( .A1(n11029), .A2(n11028), .ZN(n11031) );
  NAND2_X1 U11241 ( .A1(n14779), .A2(n11456), .ZN(n8679) );
  INV_X1 U11242 ( .A(n11942), .ZN(n11047) );
  NAND2_X1 U11243 ( .A1(n11048), .A2(n11047), .ZN(n11046) );
  OR2_X1 U11244 ( .A1(n11799), .A2(n13953), .ZN(n8680) );
  NAND2_X1 U11245 ( .A1(n11046), .A2(n8680), .ZN(n11157) );
  INV_X1 U11246 ( .A(n11719), .ZN(n13952) );
  OR2_X1 U11247 ( .A1(n11806), .A2(n13952), .ZN(n8681) );
  NAND2_X1 U11248 ( .A1(n11303), .A2(n11946), .ZN(n11302) );
  INV_X1 U11249 ( .A(n13774), .ZN(n13951) );
  OR2_X1 U11250 ( .A1(n11810), .A2(n13951), .ZN(n8682) );
  NAND2_X1 U11251 ( .A1(n11302), .A2(n8682), .ZN(n11524) );
  OR2_X1 U11252 ( .A1(n13768), .A2(n13950), .ZN(n8683) );
  INV_X1 U11253 ( .A(n12231), .ZN(n13948) );
  OR2_X1 U11254 ( .A1(n12233), .A2(n13948), .ZN(n8684) );
  OR2_X1 U11255 ( .A1(n13868), .A2(n13947), .ZN(n8686) );
  INV_X1 U11256 ( .A(n13929), .ZN(n13946) );
  XNOR2_X1 U11257 ( .A(n14329), .B(n13946), .ZN(n11835) );
  NAND2_X1 U11258 ( .A1(n14329), .A2(n13946), .ZN(n8688) );
  INV_X1 U11259 ( .A(n14213), .ZN(n13945) );
  OR2_X1 U11260 ( .A1(n14320), .A2(n13945), .ZN(n8689) );
  INV_X1 U11261 ( .A(n13928), .ZN(n13944) );
  OR2_X1 U11262 ( .A1(n14206), .A2(n13944), .ZN(n8691) );
  INV_X1 U11263 ( .A(n14211), .ZN(n14175) );
  NOR2_X1 U11264 ( .A1(n14310), .A2(n14175), .ZN(n8692) );
  NAND2_X1 U11265 ( .A1(n14310), .A2(n14175), .ZN(n8693) );
  AND2_X1 U11266 ( .A1(n14304), .A2(n14163), .ZN(n14152) );
  INV_X1 U11267 ( .A(n13902), .ZN(n14173) );
  OR2_X1 U11268 ( .A1(n14298), .A2(n14173), .ZN(n8696) );
  INV_X1 U11269 ( .A(n8696), .ZN(n8694) );
  NOR2_X1 U11270 ( .A1(n8694), .A2(n11956), .ZN(n8698) );
  OR2_X1 U11271 ( .A1(n14152), .A2(n8698), .ZN(n8695) );
  OR2_X1 U11272 ( .A1(n14304), .A2(n14163), .ZN(n14153) );
  AND2_X1 U11273 ( .A1(n14153), .A2(n8696), .ZN(n8697) );
  OR2_X1 U11274 ( .A1(n8698), .A2(n8697), .ZN(n14133) );
  AND2_X1 U11275 ( .A1(n11957), .A2(n14133), .ZN(n8699) );
  NAND2_X1 U11276 ( .A1(n14292), .A2(n14164), .ZN(n8700) );
  NAND2_X1 U11277 ( .A1(n14104), .A2(n14108), .ZN(n8703) );
  INV_X1 U11278 ( .A(n14092), .ZN(n13763) );
  NAND2_X1 U11279 ( .A1(n13882), .A2(n13763), .ZN(n8702) );
  NAND2_X1 U11280 ( .A1(n8703), .A2(n8702), .ZN(n14101) );
  NAND2_X1 U11281 ( .A1(n14276), .A2(n14072), .ZN(n8704) );
  INV_X1 U11282 ( .A(n13817), .ZN(n14093) );
  INV_X1 U11283 ( .A(n11960), .ZN(n14058) );
  OR2_X2 U11284 ( .A1(n14059), .A2(n14058), .ZN(n14261) );
  INV_X1 U11285 ( .A(n13914), .ZN(n14071) );
  NAND2_X1 U11286 ( .A1(n14259), .A2(n14071), .ZN(n14037) );
  INV_X1 U11287 ( .A(n13818), .ZN(n14053) );
  NAND2_X1 U11288 ( .A1(n12347), .A2(n14053), .ZN(n8705) );
  AND2_X1 U11289 ( .A1(n14037), .A2(n8705), .ZN(n8707) );
  INV_X1 U11290 ( .A(n8705), .ZN(n8706) );
  XNOR2_X1 U11291 ( .A(n12347), .B(n13818), .ZN(n14041) );
  AOI21_X2 U11292 ( .B1(n14261), .B2(n8707), .A(n6649), .ZN(n14033) );
  OR2_X1 U11293 ( .A1(n14248), .A2(n13943), .ZN(n8708) );
  NAND2_X1 U11294 ( .A1(n14243), .A2(n13942), .ZN(n8710) );
  OR2_X1 U11295 ( .A1(n14243), .A2(n13942), .ZN(n8709) );
  INV_X1 U11296 ( .A(n8711), .ZN(n11962) );
  XNOR2_X1 U11297 ( .A(n8712), .B(n11962), .ZN(n12205) );
  NAND2_X1 U11298 ( .A1(n13992), .A2(n14393), .ZN(n8714) );
  NAND2_X2 U11299 ( .A1(n10282), .A2(n8714), .ZN(n12364) );
  OAI211_X1 U11300 ( .C1(n10282), .C2(n11924), .A(n13992), .B(n12364), .ZN(
        n14524) );
  AND2_X1 U11301 ( .A1(n11760), .A2(n11924), .ZN(n8715) );
  NAND2_X1 U11302 ( .A1(n11925), .A2(n8715), .ZN(n10768) );
  NAND2_X1 U11303 ( .A1(n14512), .A2(n11760), .ZN(n10301) );
  NAND2_X1 U11304 ( .A1(n8716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U11305 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8717), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8718) );
  NAND2_X1 U11306 ( .A1(n8718), .A2(n6626), .ZN(n11673) );
  NAND2_X1 U11307 ( .A1(n11673), .A2(P1_B_REG_SCAN_IN), .ZN(n8723) );
  OAI21_X1 U11308 ( .B1(n8720), .B2(n8719), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8721) );
  MUX2_X1 U11309 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8721), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8722) );
  NAND2_X1 U11310 ( .A1(n8722), .A2(n8716), .ZN(n11645) );
  MUX2_X1 U11311 ( .A(P1_B_REG_SCAN_IN), .B(n8723), .S(n11645), .Z(n8725) );
  NAND2_X1 U11312 ( .A1(n6626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8724) );
  AND2_X1 U11313 ( .A1(n8725), .A2(n8731), .ZN(n10078) );
  INV_X1 U11314 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U11315 ( .A1(n10078), .A2(n10087), .ZN(n8726) );
  INV_X1 U11316 ( .A(n8731), .ZN(n14391) );
  NAND2_X1 U11317 ( .A1(n14391), .A2(n11673), .ZN(n10084) );
  NAND2_X1 U11318 ( .A1(n8726), .A2(n10084), .ZN(n10716) );
  NAND2_X1 U11319 ( .A1(n10301), .A2(n10716), .ZN(n8750) );
  INV_X1 U11320 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U11321 ( .A1(n10078), .A2(n10083), .ZN(n8727) );
  NAND2_X1 U11322 ( .A1(n11645), .A2(n14391), .ZN(n10081) );
  NAND2_X1 U11323 ( .A1(n8727), .A2(n10081), .ZN(n8749) );
  NOR2_X1 U11324 ( .A1(n8750), .A2(n8749), .ZN(n8745) );
  INV_X1 U11325 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8728) );
  INV_X1 U11326 ( .A(n11645), .ZN(n8733) );
  INV_X1 U11327 ( .A(n11673), .ZN(n8730) );
  OR2_X1 U11328 ( .A1(n10080), .A2(n10286), .ZN(n10291) );
  NAND2_X1 U11329 ( .A1(n11925), .A2(n13992), .ZN(n8746) );
  NAND2_X1 U11330 ( .A1(n11928), .A2(n8746), .ZN(n11978) );
  NOR4_X1 U11331 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n8737) );
  NOR4_X1 U11332 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n8736) );
  NOR4_X1 U11333 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n8735) );
  NOR4_X1 U11334 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n8734) );
  NAND4_X1 U11335 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n8743)
         );
  NOR2_X1 U11336 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .ZN(
        n8741) );
  NOR4_X1 U11337 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8740) );
  NOR4_X1 U11338 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8739) );
  NOR4_X1 U11339 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8738) );
  NAND4_X1 U11340 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n8742)
         );
  OAI21_X1 U11341 ( .B1(n8743), .B2(n8742), .A(n10078), .ZN(n10289) );
  NAND2_X1 U11342 ( .A1(n11978), .A2(n10289), .ZN(n8744) );
  INV_X1 U11343 ( .A(n11912), .ZN(n8747) );
  NAND2_X1 U11344 ( .A1(n8748), .A2(n7594), .ZN(P1_U3557) );
  INV_X1 U11345 ( .A(n8749), .ZN(n10717) );
  NOR2_X1 U11346 ( .A1(n8750), .A2(n10717), .ZN(n8751) );
  INV_X1 U11347 ( .A(n11173), .ZN(n8752) );
  NAND2_X1 U11348 ( .A1(n8753), .A2(n7595), .ZN(P1_U3525) );
  AOI21_X1 U11349 ( .B1(n11004), .B2(n8994), .A(n8759), .ZN(n8758) );
  NAND2_X1 U11350 ( .A1(n8760), .A2(n11752), .ZN(n8757) );
  OAI211_X1 U11351 ( .C1(n11752), .C2(n7411), .A(n8760), .B(n8994), .ZN(n8761)
         );
  INV_X4 U11352 ( .A(n8994), .ZN(n8822) );
  NAND2_X1 U11353 ( .A1(n8822), .A2(n6562), .ZN(n8763) );
  NAND2_X1 U11354 ( .A1(n8764), .A2(n8822), .ZN(n8766) );
  NAND2_X1 U11355 ( .A1(n6770), .A2(n6562), .ZN(n8765) );
  NAND2_X1 U11356 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  NAND2_X1 U11357 ( .A1(n8768), .A2(n8767), .ZN(n8774) );
  INV_X1 U11358 ( .A(n8769), .ZN(n8772) );
  INV_X1 U11359 ( .A(n8770), .ZN(n8771) );
  NAND2_X1 U11360 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U11361 ( .A1(n6770), .A2(n7671), .ZN(n8775) );
  NAND2_X1 U11362 ( .A1(n8776), .A2(n8775), .ZN(n8778) );
  AOI22_X1 U11363 ( .A1(n13234), .A2(n6770), .B1(n6565), .B2(n7671), .ZN(n8777) );
  NAND2_X1 U11364 ( .A1(n13233), .A2(n6770), .ZN(n8782) );
  NAND2_X1 U11365 ( .A1(n8946), .A2(n10273), .ZN(n8781) );
  NAND2_X1 U11366 ( .A1(n8782), .A2(n8781), .ZN(n8784) );
  AOI22_X1 U11367 ( .A1(n13233), .A2(n8946), .B1(n10273), .B2(n6770), .ZN(
        n8783) );
  NAND2_X1 U11368 ( .A1(n10393), .A2(n6770), .ZN(n8789) );
  NAND2_X1 U11369 ( .A1(n13232), .A2(n8946), .ZN(n8788) );
  NAND2_X1 U11370 ( .A1(n8789), .A2(n8788), .ZN(n8792) );
  NAND2_X1 U11371 ( .A1(n10393), .A2(n8946), .ZN(n8791) );
  NAND2_X1 U11372 ( .A1(n13232), .A2(n6770), .ZN(n8790) );
  NAND2_X1 U11373 ( .A1(n10989), .A2(n8946), .ZN(n8794) );
  NAND2_X1 U11374 ( .A1(n13231), .A2(n6770), .ZN(n8793) );
  NAND2_X1 U11375 ( .A1(n8794), .A2(n8793), .ZN(n8796) );
  AOI22_X1 U11376 ( .A1(n10989), .A2(n6770), .B1(n8946), .B2(n13231), .ZN(
        n8795) );
  NAND2_X1 U11377 ( .A1(n14910), .A2(n6770), .ZN(n8801) );
  NAND2_X1 U11378 ( .A1(n13230), .A2(n8946), .ZN(n8800) );
  NAND2_X1 U11379 ( .A1(n14910), .A2(n8946), .ZN(n8802) );
  NAND2_X1 U11380 ( .A1(n14917), .A2(n8946), .ZN(n8806) );
  NAND2_X1 U11381 ( .A1(n13229), .A2(n6770), .ZN(n8805) );
  NAND2_X1 U11382 ( .A1(n8806), .A2(n8805), .ZN(n8811) );
  AOI22_X1 U11383 ( .A1(n14917), .A2(n6770), .B1(n8946), .B2(n13229), .ZN(
        n8807) );
  INV_X1 U11384 ( .A(n8807), .ZN(n8808) );
  NAND2_X1 U11385 ( .A1(n8809), .A2(n8808), .ZN(n8815) );
  NAND2_X1 U11386 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  NAND2_X1 U11387 ( .A1(n10913), .A2(n8943), .ZN(n8817) );
  NAND2_X1 U11388 ( .A1(n13228), .A2(n8946), .ZN(n8816) );
  NAND2_X1 U11389 ( .A1(n8817), .A2(n8816), .ZN(n8819) );
  AOI22_X1 U11390 ( .A1(n10913), .A2(n8946), .B1(n13228), .B2(n8943), .ZN(
        n8818) );
  AOI21_X1 U11391 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  NAND2_X1 U11392 ( .A1(n11250), .A2(n8946), .ZN(n8824) );
  NAND2_X1 U11393 ( .A1(n13227), .A2(n8943), .ZN(n8823) );
  NAND2_X1 U11394 ( .A1(n11250), .A2(n8943), .ZN(n8825) );
  OAI21_X1 U11395 ( .B1(n8826), .B2(n8943), .A(n8825), .ZN(n8827) );
  NAND2_X1 U11396 ( .A1(n11277), .A2(n8943), .ZN(n8829) );
  NAND2_X1 U11397 ( .A1(n13226), .A2(n8946), .ZN(n8828) );
  NAND2_X1 U11398 ( .A1(n8829), .A2(n8828), .ZN(n8832) );
  AOI22_X1 U11399 ( .A1(n11277), .A2(n8946), .B1(n13226), .B2(n8943), .ZN(
        n8830) );
  INV_X1 U11400 ( .A(n8831), .ZN(n8834) );
  NAND2_X1 U11401 ( .A1(n11479), .A2(n6565), .ZN(n8836) );
  NAND2_X1 U11402 ( .A1(n13225), .A2(n8943), .ZN(n8835) );
  NAND2_X1 U11403 ( .A1(n8836), .A2(n8835), .ZN(n8839) );
  NAND2_X1 U11404 ( .A1(n11479), .A2(n8943), .ZN(n8837) );
  OAI21_X1 U11405 ( .B1(n11438), .B2(n8943), .A(n8837), .ZN(n8838) );
  INV_X1 U11406 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U11407 ( .A1(n13578), .A2(n8943), .ZN(n8842) );
  NAND2_X1 U11408 ( .A1(n13224), .A2(n6565), .ZN(n8841) );
  NAND2_X1 U11409 ( .A1(n8842), .A2(n8841), .ZN(n8844) );
  NAND2_X1 U11410 ( .A1(n11575), .A2(n6565), .ZN(n8848) );
  NAND2_X1 U11411 ( .A1(n13223), .A2(n8943), .ZN(n8847) );
  NAND2_X1 U11412 ( .A1(n11575), .A2(n8943), .ZN(n8849) );
  OAI21_X1 U11413 ( .B1(n11437), .B2(n8943), .A(n8849), .ZN(n8850) );
  NAND2_X1 U11414 ( .A1(n13718), .A2(n8943), .ZN(n8852) );
  NAND2_X1 U11415 ( .A1(n13222), .A2(n6565), .ZN(n8851) );
  NAND2_X1 U11416 ( .A1(n8852), .A2(n8851), .ZN(n8866) );
  AOI22_X1 U11417 ( .A1(n13656), .A2(n8943), .B1(n6565), .B2(n13517), .ZN(
        n8855) );
  NAND2_X1 U11418 ( .A1(n13656), .A2(n8946), .ZN(n8854) );
  NAND2_X1 U11419 ( .A1(n13517), .A2(n8943), .ZN(n8853) );
  NAND2_X1 U11420 ( .A1(n8854), .A2(n8853), .ZN(n8873) );
  NAND2_X1 U11421 ( .A1(n8855), .A2(n8873), .ZN(n8860) );
  AND2_X1 U11422 ( .A1(n13221), .A2(n8946), .ZN(n8856) );
  AOI21_X1 U11423 ( .B1(n14637), .B2(n8943), .A(n8856), .ZN(n8871) );
  NAND2_X1 U11424 ( .A1(n14637), .A2(n6565), .ZN(n8858) );
  NAND2_X1 U11425 ( .A1(n13221), .A2(n8943), .ZN(n8857) );
  NAND2_X1 U11426 ( .A1(n8858), .A2(n8857), .ZN(n8870) );
  NAND2_X1 U11427 ( .A1(n8871), .A2(n8870), .ZN(n8859) );
  AND2_X1 U11428 ( .A1(n8860), .A2(n8859), .ZN(n8876) );
  AND2_X1 U11429 ( .A1(n13519), .A2(n6565), .ZN(n8861) );
  AOI21_X1 U11430 ( .B1(n13715), .B2(n8943), .A(n8861), .ZN(n8869) );
  NAND2_X1 U11431 ( .A1(n13715), .A2(n8946), .ZN(n8863) );
  NAND2_X1 U11432 ( .A1(n13519), .A2(n8943), .ZN(n8862) );
  NAND2_X1 U11433 ( .A1(n8863), .A2(n8862), .ZN(n8868) );
  NAND2_X1 U11434 ( .A1(n8869), .A2(n8868), .ZN(n8864) );
  AOI22_X1 U11435 ( .A1(n13718), .A2(n6565), .B1(n13222), .B2(n8943), .ZN(
        n8865) );
  OAI22_X1 U11436 ( .A1(n8871), .A2(n8870), .B1(n8869), .B2(n8868), .ZN(n8875)
         );
  NOR2_X1 U11437 ( .A1(n13656), .A2(n13517), .ZN(n8872) );
  NOR2_X1 U11438 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  AOI21_X1 U11439 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n8877) );
  NAND2_X1 U11440 ( .A1(n13651), .A2(n8943), .ZN(n8881) );
  NAND2_X1 U11441 ( .A1(n13220), .A2(n6565), .ZN(n8880) );
  NAND2_X1 U11442 ( .A1(n8881), .A2(n8880), .ZN(n8886) );
  NAND2_X1 U11443 ( .A1(n8885), .A2(n8886), .ZN(n8884) );
  NAND2_X1 U11444 ( .A1(n13651), .A2(n8946), .ZN(n8882) );
  INV_X1 U11445 ( .A(n8885), .ZN(n8888) );
  INV_X1 U11446 ( .A(n8886), .ZN(n8887) );
  NAND2_X1 U11447 ( .A1(n13647), .A2(n8946), .ZN(n8890) );
  NAND2_X1 U11448 ( .A1(n13219), .A2(n8943), .ZN(n8889) );
  NAND2_X1 U11449 ( .A1(n8890), .A2(n8889), .ZN(n8894) );
  NAND2_X1 U11450 ( .A1(n13647), .A2(n8943), .ZN(n8892) );
  NAND2_X1 U11451 ( .A1(n13219), .A2(n6565), .ZN(n8891) );
  NAND2_X1 U11452 ( .A1(n8892), .A2(n8891), .ZN(n8893) );
  INV_X1 U11453 ( .A(n8894), .ZN(n8895) );
  INV_X1 U11454 ( .A(n8901), .ZN(n8899) );
  NAND2_X1 U11455 ( .A1(n13642), .A2(n8943), .ZN(n8897) );
  NAND2_X1 U11456 ( .A1(n13218), .A2(n6565), .ZN(n8896) );
  INV_X1 U11457 ( .A(n8900), .ZN(n8898) );
  NAND2_X1 U11458 ( .A1(n8899), .A2(n8898), .ZN(n8907) );
  NAND2_X1 U11459 ( .A1(n13642), .A2(n6565), .ZN(n8903) );
  NAND2_X1 U11460 ( .A1(n13218), .A2(n8943), .ZN(n8902) );
  NAND2_X1 U11461 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U11462 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  NAND2_X1 U11463 ( .A1(n13636), .A2(n8946), .ZN(n8909) );
  NAND2_X1 U11464 ( .A1(n13217), .A2(n8943), .ZN(n8908) );
  NAND2_X1 U11465 ( .A1(n8909), .A2(n8908), .ZN(n8911) );
  NAND2_X1 U11466 ( .A1(n13705), .A2(n8943), .ZN(n8913) );
  NAND2_X1 U11467 ( .A1(n13216), .A2(n8946), .ZN(n8912) );
  NAND2_X1 U11468 ( .A1(n13705), .A2(n8946), .ZN(n8914) );
  NAND2_X1 U11469 ( .A1(n8916), .A2(n8915), .ZN(n8922) );
  INV_X1 U11470 ( .A(n8917), .ZN(n8920) );
  INV_X1 U11471 ( .A(n8918), .ZN(n8919) );
  NAND2_X1 U11472 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  NAND2_X1 U11473 ( .A1(n13408), .A2(n8946), .ZN(n8924) );
  NAND2_X1 U11474 ( .A1(n13215), .A2(n8943), .ZN(n8923) );
  NAND2_X1 U11475 ( .A1(n8924), .A2(n8923), .ZN(n8926) );
  AOI22_X1 U11476 ( .A1(n13408), .A2(n8943), .B1(n6565), .B2(n13215), .ZN(
        n8925) );
  INV_X1 U11477 ( .A(n8928), .ZN(n8929) );
  NAND2_X1 U11478 ( .A1(n13620), .A2(n8943), .ZN(n8931) );
  NAND2_X1 U11479 ( .A1(n13214), .A2(n6565), .ZN(n8930) );
  NAND2_X1 U11480 ( .A1(n13620), .A2(n8946), .ZN(n8933) );
  NAND2_X1 U11481 ( .A1(n13214), .A2(n8943), .ZN(n8932) );
  NAND2_X1 U11482 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U11483 ( .A1(n13696), .A2(n8946), .ZN(n8936) );
  NAND2_X1 U11484 ( .A1(n13213), .A2(n8943), .ZN(n8935) );
  NAND2_X1 U11485 ( .A1(n8936), .A2(n8935), .ZN(n8938) );
  AOI22_X1 U11486 ( .A1(n13696), .A2(n8943), .B1(n6565), .B2(n13213), .ZN(
        n8937) );
  NAND2_X1 U11487 ( .A1(n13361), .A2(n8943), .ZN(n8941) );
  NAND2_X1 U11488 ( .A1(n13212), .A2(n8946), .ZN(n8940) );
  AOI22_X1 U11489 ( .A1(n13361), .A2(n6565), .B1(n13212), .B2(n8943), .ZN(
        n8942) );
  AND2_X1 U11490 ( .A1(n13211), .A2(n8943), .ZN(n8944) );
  AOI21_X1 U11491 ( .B1(n13347), .B2(n6565), .A(n8944), .ZN(n8947) );
  INV_X1 U11492 ( .A(n8947), .ZN(n8945) );
  AOI22_X1 U11493 ( .A1(n13598), .A2(n6565), .B1(n13210), .B2(n8943), .ZN(
        n8956) );
  OAI22_X1 U11494 ( .A1(n7422), .A2(n8946), .B1(n13096), .B2(n8943), .ZN(n8955) );
  OAI22_X1 U11495 ( .A1(n13596), .A2(n8943), .B1(n9837), .B2(n6565), .ZN(n8985) );
  AOI22_X1 U11496 ( .A1(n13316), .A2(n8943), .B1(n8946), .B2(n13209), .ZN(
        n8986) );
  NOR2_X1 U11497 ( .A1(n8985), .A2(n8986), .ZN(n8954) );
  AOI21_X1 U11498 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8953) );
  OAI22_X1 U11499 ( .A1(n13689), .A2(n8946), .B1(n13189), .B2(n8943), .ZN(
        n8948) );
  INV_X1 U11500 ( .A(n8948), .ZN(n8949) );
  INV_X1 U11501 ( .A(n8951), .ZN(n8952) );
  INV_X1 U11502 ( .A(n8954), .ZN(n8959) );
  INV_X1 U11503 ( .A(n8955), .ZN(n8958) );
  INV_X1 U11504 ( .A(n8956), .ZN(n8957) );
  NAND3_X1 U11505 ( .A1(n8959), .A2(n8958), .A3(n8957), .ZN(n8975) );
  INV_X1 U11506 ( .A(SI_29_), .ZN(n13091) );
  NAND2_X1 U11507 ( .A1(n8962), .A2(n13091), .ZN(n8963) );
  MUX2_X1 U11508 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6568), .Z(n8965) );
  XNOR2_X1 U11509 ( .A(n8965), .B(SI_30_), .ZN(n8976) );
  NAND2_X1 U11510 ( .A1(n8965), .A2(SI_30_), .ZN(n8966) );
  MUX2_X1 U11511 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6551), .Z(n8967) );
  XNOR2_X1 U11512 ( .A(n8967), .B(SI_31_), .ZN(n8968) );
  INV_X1 U11513 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13589) );
  NOR2_X1 U11514 ( .A1(n6566), .A2(n13589), .ZN(n8974) );
  INV_X1 U11515 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8971) );
  NOR2_X1 U11516 ( .A1(n8182), .A2(n8971), .ZN(n8973) );
  INV_X1 U11517 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13678) );
  NOR2_X1 U11518 ( .A1(n7691), .A2(n13678), .ZN(n8972) );
  XNOR2_X1 U11519 ( .A(n13680), .B(n13302), .ZN(n9010) );
  MUX2_X1 U11520 ( .A(n8946), .B(n13302), .S(n13680), .Z(n8989) );
  NAND2_X1 U11521 ( .A1(n13302), .A2(n8946), .ZN(n8988) );
  INV_X1 U11522 ( .A(n8976), .ZN(n8977) );
  NAND2_X1 U11523 ( .A1(n12213), .A2(n7702), .ZN(n8981) );
  INV_X1 U11524 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12214) );
  OR2_X1 U11525 ( .A1(n8979), .A2(n12214), .ZN(n8980) );
  OAI211_X1 U11526 ( .C1(n11732), .C2(n9831), .A(n6564), .B(n9835), .ZN(n8982)
         );
  AOI21_X1 U11527 ( .B1(n13302), .B2(n8943), .A(n8982), .ZN(n8983) );
  OAI22_X1 U11528 ( .A1(n13684), .A2(n8943), .B1(n8984), .B2(n8983), .ZN(n8992) );
  INV_X1 U11529 ( .A(n8984), .ZN(n13208) );
  AOI22_X1 U11530 ( .A1(n8992), .A2(n8993), .B1(n8986), .B2(n8985), .ZN(n8987)
         );
  AOI21_X1 U11531 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(n8990) );
  INV_X1 U11532 ( .A(n13680), .ZN(n13299) );
  INV_X1 U11533 ( .A(n13302), .ZN(n8995) );
  NAND3_X1 U11534 ( .A1(n13299), .A2(n8995), .A3(n8943), .ZN(n8997) );
  NAND3_X1 U11535 ( .A1(n13680), .A2(n8822), .A3(n13302), .ZN(n8996) );
  INV_X1 U11536 ( .A(n9035), .ZN(n9001) );
  INV_X1 U11537 ( .A(n9835), .ZN(n9007) );
  NOR2_X1 U11538 ( .A1(n9009), .A2(n9694), .ZN(n8999) );
  OR2_X1 U11539 ( .A1(n9939), .A2(P2_U3088), .ZN(n11637) );
  INV_X1 U11540 ( .A(n11637), .ZN(n9006) );
  MUX2_X1 U11541 ( .A(n9009), .B(n6564), .S(n9831), .Z(n9003) );
  NAND2_X1 U11542 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  NAND4_X1 U11543 ( .A1(n14891), .A2(n9946), .A3(n9007), .A4(n13518), .ZN(
        n9008) );
  OAI211_X1 U11544 ( .C1(n9009), .C2(n11637), .A(n9008), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9037) );
  INV_X1 U11545 ( .A(n9010), .ZN(n9031) );
  XNOR2_X1 U11546 ( .A(n13361), .B(n9011), .ZN(n13356) );
  XOR2_X1 U11547 ( .A(n13218), .B(n13642), .Z(n13454) );
  XNOR2_X1 U11548 ( .A(n13647), .B(n13219), .ZN(n13468) );
  XNOR2_X1 U11549 ( .A(n13718), .B(n9012), .ZN(n13559) );
  NOR2_X1 U11550 ( .A1(n9014), .A2(n9013), .ZN(n11413) );
  AND2_X1 U11551 ( .A1(n9016), .A2(n9015), .ZN(n11131) );
  OAI21_X1 U11552 ( .B1(n7655), .B2(n11004), .A(n9698), .ZN(n11745) );
  NAND4_X1 U11553 ( .A1(n11006), .A2(n10183), .A3(n9831), .A4(n11745), .ZN(
        n9017) );
  XNOR2_X1 U11554 ( .A(n10989), .B(n13231), .ZN(n10991) );
  NAND4_X1 U11555 ( .A1(n10908), .A2(n11131), .A3(n9019), .A4(n10991), .ZN(
        n9020) );
  NOR3_X1 U11556 ( .A1(n9020), .A2(n11262), .A3(n11176), .ZN(n9021) );
  XNOR2_X1 U11557 ( .A(n13578), .B(n13224), .ZN(n11489) );
  NAND4_X1 U11558 ( .A1(n11413), .A2(n9021), .A3(n11489), .A4(n11345), .ZN(
        n9022) );
  NOR4_X1 U11559 ( .A1(n13512), .A2(n13545), .A3(n13559), .A4(n9022), .ZN(
        n9024) );
  NAND4_X1 U11560 ( .A1(n13468), .A2(n9024), .A3(n13491), .A4(n9023), .ZN(
        n9025) );
  NOR4_X1 U11561 ( .A1(n13416), .A2(n13454), .A3(n13447), .A4(n9025), .ZN(
        n9026) );
  NAND4_X1 U11562 ( .A1(n13372), .A2(n9026), .A3(n13382), .A4(n13401), .ZN(
        n9027) );
  NOR4_X1 U11563 ( .A1(n13330), .A2(n13341), .A3(n13356), .A4(n9027), .ZN(
        n9030) );
  XNOR2_X1 U11564 ( .A(n13311), .B(n13208), .ZN(n9029) );
  NAND4_X1 U11565 ( .A1(n9031), .A2(n9030), .A3(n9029), .A4(n9028), .ZN(n9032)
         );
  XNOR2_X1 U11566 ( .A(n9032), .B(n13292), .ZN(n9033) );
  NOR3_X1 U11567 ( .A1(n9033), .A2(n6564), .A3(n11637), .ZN(n9034) );
  OAI21_X1 U11568 ( .B1(n9035), .B2(n9831), .A(n9034), .ZN(n9036) );
  NAND3_X1 U11569 ( .A1(n9038), .A2(n9037), .A3(n9036), .ZN(P2_U3328) );
  NAND4_X1 U11570 ( .A1(n9041), .A2(n9040), .A3(n15206), .A4(n9254), .ZN(n9042) );
  INV_X1 U11571 ( .A(n9042), .ZN(n9046) );
  INV_X1 U11572 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9048) );
  INV_X1 U11573 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11574 ( .A1(n9058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9057) );
  MUX2_X1 U11575 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9057), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9060) );
  INV_X1 U11576 ( .A(n9135), .ZN(n9059) );
  NAND3_X1 U11577 ( .A1(n9383), .A2(n9062), .A3(n9061), .ZN(n9063) );
  NAND2_X1 U11578 ( .A1(n9063), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9065) );
  INV_X1 U11579 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11580 ( .A1(n12190), .A2(n10611), .ZN(n9066) );
  NAND2_X1 U11581 ( .A1(n12180), .A2(n9066), .ZN(n9068) );
  NAND2_X1 U11582 ( .A1(n6651), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11583 ( .A1(n9068), .A2(n10934), .ZN(n9070) );
  INV_X1 U11584 ( .A(n10611), .ZN(n9683) );
  OAI21_X1 U11585 ( .B1(n9683), .B2(n12014), .A(n12012), .ZN(n9069) );
  NAND2_X1 U11586 ( .A1(n9070), .A2(n9069), .ZN(n10626) );
  NAND2_X1 U11587 ( .A1(n6555), .A2(n10611), .ZN(n9684) );
  INV_X1 U11588 ( .A(n9684), .ZN(n12185) );
  NAND3_X1 U11589 ( .A1(n10626), .A2(n12185), .A3(n15098), .ZN(n9072) );
  NOR2_X1 U11590 ( .A1(n12012), .A2(n10611), .ZN(n9071) );
  NAND2_X1 U11591 ( .A1(n6555), .A2(n9071), .ZN(n9682) );
  AND2_X1 U11592 ( .A1(n9072), .A2(n9682), .ZN(n11591) );
  NAND2_X1 U11593 ( .A1(n12180), .A2(n10611), .ZN(n15123) );
  OR2_X1 U11594 ( .A1(n15123), .A2(n12190), .ZN(n12946) );
  AND2_X1 U11595 ( .A1(n11591), .A2(n12946), .ZN(n14611) );
  INV_X1 U11596 ( .A(n9191), .ZN(n9074) );
  NAND2_X1 U11597 ( .A1(n9917), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11598 ( .A1(n9910), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11599 ( .A1(n9869), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11600 ( .A1(n15396), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U11601 ( .A1(n9209), .A2(n9208), .ZN(n9079) );
  NAND2_X1 U11602 ( .A1(n9079), .A2(n15210), .ZN(n9221) );
  NAND2_X1 U11603 ( .A1(n9913), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11604 ( .A1(n9895), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11605 ( .A1(n9221), .A2(n9220), .ZN(n9082) );
  NAND2_X1 U11606 ( .A1(n9909), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11607 ( .A1(n9901), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11608 ( .A1(n9237), .A2(n9236), .ZN(n9085) );
  NAND2_X1 U11609 ( .A1(n9919), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11610 ( .A1(n9251), .A2(n9086), .ZN(n9088) );
  NAND2_X1 U11611 ( .A1(n9922), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11612 ( .A1(n9926), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11613 ( .A1(n9925), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9089) );
  INV_X1 U11614 ( .A(n9271), .ZN(n9090) );
  NAND2_X1 U11615 ( .A1(n9932), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U11616 ( .A1(n9936), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11617 ( .A1(n9935), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11618 ( .A1(n10091), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U11619 ( .A1(n10090), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U11620 ( .A1(n10130), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11621 ( .A1(n15303), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11622 ( .A1(n10135), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11623 ( .A1(n10137), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9099) );
  NAND2_X2 U11624 ( .A1(n9101), .A2(n10157), .ZN(n9103) );
  NAND2_X1 U11625 ( .A1(n10463), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9105) );
  INV_X1 U11626 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U11627 ( .A1(n10465), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U11628 ( .A1(n10672), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U11629 ( .A1(n10671), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11630 ( .A1(n10702), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11631 ( .A1(n10704), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11632 ( .A1(n10829), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11633 ( .A1(n10831), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11634 ( .A1(n11202), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11635 ( .A1(n11204), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U11636 ( .A1(n15248), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9115) );
  INV_X1 U11637 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U11638 ( .A1(n11299), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11639 ( .A1(n11408), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11640 ( .A1(n11407), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9119) );
  AND2_X1 U11641 ( .A1(n9120), .A2(n9119), .ZN(n9483) );
  XNOR2_X1 U11642 ( .A(n11734), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11643 ( .A1(n11734), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9121) );
  XNOR2_X1 U11644 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9509) );
  NAND2_X1 U11645 ( .A1(n11639), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9123) );
  XNOR2_X1 U11646 ( .A(n11676), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11647 ( .A1(n11676), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9127) );
  NOR2_X1 U11648 ( .A1(n14388), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11649 ( .A1(n14388), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9129) );
  AND2_X1 U11650 ( .A1(n14385), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U11651 ( .A1(n13734), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9131) );
  AND2_X1 U11652 ( .A1(n13731), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11653 ( .A1(n11726), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9133) );
  XNOR2_X1 U11654 ( .A(n14381), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n11991) );
  XNOR2_X1 U11655 ( .A(n11993), .B(n11991), .ZN(n13087) );
  INV_X1 U11656 ( .A(n9162), .ZN(n9140) );
  XNOR2_X2 U11657 ( .A(n9138), .B(n9161), .ZN(n9623) );
  NAND2_X1 U11658 ( .A1(n9635), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9139) );
  NAND2_X4 U11659 ( .A1(n9623), .A2(n12718), .ZN(n9179) );
  NAND2_X1 U11660 ( .A1(n13087), .A2(n12004), .ZN(n9143) );
  NAND2_X1 U11661 ( .A1(n9565), .A2(SI_29_), .ZN(n9142) );
  NAND2_X2 U11662 ( .A1(n9143), .A2(n9142), .ZN(n12385) );
  INV_X1 U11663 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U11664 ( .A1(n15304), .A2(n10820), .ZN(n9144) );
  INV_X1 U11665 ( .A(n9366), .ZN(n9148) );
  INV_X1 U11666 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9147) );
  INV_X1 U11667 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9150) );
  INV_X1 U11668 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15291) );
  INV_X1 U11669 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9154) );
  INV_X1 U11670 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9156) );
  INV_X1 U11671 ( .A(n9544), .ZN(n9158) );
  INV_X1 U11672 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12574) );
  INV_X1 U11673 ( .A(n9568), .ZN(n9160) );
  INV_X1 U11674 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11675 ( .A1(n9160), .A2(n9159), .ZN(n12381) );
  INV_X1 U11676 ( .A(n9167), .ZN(n9164) );
  INV_X1 U11677 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11678 ( .A1(n9164), .A2(n9163), .ZN(n13082) );
  NAND2_X2 U11679 ( .A1(n9170), .A2(n9169), .ZN(n9423) );
  INV_X2 U11680 ( .A(n9175), .ZN(n9478) );
  INV_X1 U11681 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U11682 ( .A1(n9555), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9172) );
  NAND2_X2 U11683 ( .A1(n12380), .A2(n13090), .ZN(n11984) );
  NAND2_X1 U11684 ( .A1(n9571), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9171) );
  OAI211_X1 U11685 ( .C1(n6553), .C2(n12382), .A(n9172), .B(n9171), .ZN(n9173)
         );
  INV_X1 U11686 ( .A(n9173), .ZN(n9174) );
  NAND2_X1 U11687 ( .A1(n11990), .A2(n9174), .ZN(n12750) );
  XNOR2_X1 U11688 ( .A(n12385), .B(n12750), .ZN(n12176) );
  INV_X1 U11689 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9176) );
  INV_X1 U11690 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10557) );
  INV_X1 U11691 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10330) );
  OR2_X1 U11692 ( .A1(n9275), .A2(n10330), .ZN(n9177) );
  INV_X1 U11693 ( .A(SI_1_), .ZN(n9874) );
  XNOR2_X1 U11694 ( .A(n9178), .B(n9191), .ZN(n9875) );
  INV_X1 U11695 ( .A(n10356), .ZN(n9180) );
  INV_X1 U11696 ( .A(n10568), .ZN(n10331) );
  NAND2_X1 U11697 ( .A1(n9460), .A2(n10331), .ZN(n9182) );
  NAND2_X1 U11698 ( .A1(n9555), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9188) );
  INV_X1 U11699 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n9183) );
  OR2_X1 U11700 ( .A1(n11984), .A2(n9183), .ZN(n9187) );
  INV_X1 U11701 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14947) );
  INV_X1 U11702 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n14942) );
  NAND2_X1 U11703 ( .A1(n9189), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U11704 ( .A1(n9191), .A2(n9190), .ZN(n9192) );
  MUX2_X1 U11705 ( .A(n9192), .B(SI_0_), .S(n6568), .Z(n13093) );
  MUX2_X1 U11706 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13093), .S(n9179), .Z(n11756)
         );
  INV_X1 U11707 ( .A(n11756), .ZN(n14934) );
  INV_X1 U11708 ( .A(n13014), .ZN(n9193) );
  NAND2_X1 U11709 ( .A1(n9555), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9198) );
  INV_X1 U11710 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15100) );
  OR2_X1 U11711 ( .A1(n9423), .A2(n15100), .ZN(n9197) );
  INV_X1 U11712 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15120) );
  OR2_X1 U11713 ( .A1(n9275), .A2(n15120), .ZN(n9196) );
  INV_X1 U11714 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9194) );
  OR2_X1 U11715 ( .A1(n11984), .A2(n9194), .ZN(n9195) );
  XNOR2_X1 U11716 ( .A(n9200), .B(n9199), .ZN(n9887) );
  OR2_X1 U11717 ( .A1(n9487), .A2(n9887), .ZN(n9202) );
  OR2_X1 U11718 ( .A1(n12005), .A2(SI_2_), .ZN(n9201) );
  NAND2_X1 U11719 ( .A1(n13008), .A2(n15099), .ZN(n12022) );
  NAND2_X1 U11720 ( .A1(n9571), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9207) );
  OR2_X1 U11721 ( .A1(n9423), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9206) );
  INV_X1 U11722 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10341) );
  OR2_X1 U11723 ( .A1(n9275), .A2(n10341), .ZN(n9205) );
  INV_X1 U11724 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10340) );
  OR2_X1 U11725 ( .A1(n6557), .A2(n10340), .ZN(n9204) );
  XNOR2_X1 U11726 ( .A(n9209), .B(n9208), .ZN(n9885) );
  OR2_X1 U11727 ( .A1(n9487), .A2(n9885), .ZN(n9211) );
  OR2_X1 U11728 ( .A1(n12005), .A2(SI_3_), .ZN(n9210) );
  OR2_X2 U11729 ( .A1(n9585), .A2(n11098), .ZN(n12026) );
  NAND2_X1 U11730 ( .A1(n9585), .A2(n11098), .ZN(n12025) );
  AND2_X2 U11731 ( .A1(n12026), .A2(n12025), .ZN(n12162) );
  NAND2_X1 U11732 ( .A1(n11087), .A2(n12162), .ZN(n9212) );
  NAND2_X1 U11733 ( .A1(n6559), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9217) );
  INV_X1 U11734 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10361) );
  OR2_X1 U11735 ( .A1(n6553), .A2(n10361), .ZN(n9216) );
  AND2_X1 U11736 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9213) );
  NOR2_X1 U11737 ( .A1(n9227), .A2(n9213), .ZN(n15091) );
  OR2_X1 U11738 ( .A1(n9478), .A2(n15091), .ZN(n9215) );
  INV_X1 U11739 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10372) );
  OR2_X1 U11740 ( .A1(n6558), .A2(n10372), .ZN(n9214) );
  NAND4_X1 U11741 ( .A1(n9217), .A2(n9216), .A3(n9215), .A4(n9214), .ZN(n12611) );
  NAND2_X1 U11742 ( .A1(n9218), .A2(n15206), .ZN(n9234) );
  NAND2_X1 U11743 ( .A1(n9234), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9219) );
  XNOR2_X1 U11744 ( .A(n9221), .B(n9220), .ZN(n9889) );
  OR2_X1 U11745 ( .A1(n9487), .A2(n9889), .ZN(n9223) );
  OR2_X1 U11746 ( .A1(n12005), .A2(SI_4_), .ZN(n9222) );
  OAI211_X1 U11747 ( .C1(n10373), .C2(n9179), .A(n9223), .B(n9222), .ZN(n15090) );
  NAND2_X1 U11748 ( .A1(n12611), .A2(n15090), .ZN(n12030) );
  NAND2_X1 U11749 ( .A1(n15083), .A2(n15082), .ZN(n9224) );
  NAND2_X1 U11750 ( .A1(n6559), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9233) );
  INV_X1 U11751 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9225) );
  OR2_X1 U11752 ( .A1(n6553), .A2(n9225), .ZN(n9232) );
  NOR2_X1 U11753 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  OR2_X1 U11754 ( .A1(n9241), .A2(n9228), .ZN(n10936) );
  INV_X1 U11755 ( .A(n10936), .ZN(n11246) );
  OR2_X1 U11756 ( .A1(n9478), .A2(n11246), .ZN(n9231) );
  INV_X1 U11757 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9229) );
  OR2_X1 U11758 ( .A1(n6558), .A2(n9229), .ZN(n9230) );
  NAND4_X1 U11759 ( .A1(n9233), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(n12610) );
  NAND2_X1 U11760 ( .A1(n9252), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9235) );
  XNOR2_X1 U11761 ( .A(n9235), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10383) );
  XNOR2_X1 U11762 ( .A(n9237), .B(n9236), .ZN(n9883) );
  OR2_X1 U11763 ( .A1(n9487), .A2(n9883), .ZN(n9239) );
  OR2_X1 U11764 ( .A1(n12005), .A2(SI_5_), .ZN(n9238) );
  OAI211_X1 U11765 ( .C1(n10383), .C2(n9179), .A(n9239), .B(n9238), .ZN(n11240) );
  XNOR2_X1 U11766 ( .A(n12610), .B(n11240), .ZN(n10921) );
  INV_X1 U11767 ( .A(n10921), .ZN(n12165) );
  NAND2_X1 U11768 ( .A1(n10919), .A2(n12165), .ZN(n9240) );
  OR2_X1 U11769 ( .A1(n12610), .A2(n11240), .ZN(n12009) );
  NOR2_X1 U11770 ( .A1(n9241), .A2(n15331), .ZN(n9242) );
  OR2_X1 U11771 ( .A1(n9263), .A2(n9242), .ZN(n15075) );
  NAND2_X1 U11772 ( .A1(n9175), .A2(n15075), .ZN(n9249) );
  INV_X1 U11773 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9243) );
  OR2_X1 U11774 ( .A1(n9369), .A2(n9243), .ZN(n9248) );
  INV_X1 U11775 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9244) );
  OR2_X1 U11776 ( .A1(n6558), .A2(n9244), .ZN(n9247) );
  INV_X1 U11777 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9245) );
  OR2_X1 U11778 ( .A1(n11984), .A2(n9245), .ZN(n9246) );
  NAND4_X1 U11779 ( .A1(n9249), .A2(n9248), .A3(n9247), .A4(n9246), .ZN(n12609) );
  INV_X1 U11780 ( .A(SI_6_), .ZN(n9879) );
  OR2_X1 U11781 ( .A1(n12005), .A2(n9879), .ZN(n9260) );
  XNOR2_X1 U11782 ( .A(n9922), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9250) );
  XNOR2_X1 U11783 ( .A(n9251), .B(n9250), .ZN(n9880) );
  OR2_X1 U11784 ( .A1(n9487), .A2(n9880), .ZN(n9259) );
  NOR2_X1 U11785 ( .A1(n9255), .A2(n9415), .ZN(n9253) );
  MUX2_X1 U11786 ( .A(n9415), .B(n9253), .S(P3_IR_REG_6__SCAN_IN), .Z(n9257)
         );
  NAND2_X1 U11787 ( .A1(n9255), .A2(n9254), .ZN(n9280) );
  INV_X1 U11788 ( .A(n9280), .ZN(n9256) );
  INV_X1 U11789 ( .A(n14962), .ZN(n10815) );
  NAND2_X1 U11790 ( .A1(n9460), .A2(n10815), .ZN(n9258) );
  NAND2_X1 U11791 ( .A1(n12609), .A2(n15078), .ZN(n12036) );
  NAND2_X1 U11792 ( .A1(n6559), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9269) );
  INV_X1 U11793 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9261) );
  OR2_X1 U11794 ( .A1(n6557), .A2(n9261), .ZN(n9268) );
  OR2_X1 U11795 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  AND2_X1 U11796 ( .A1(n9292), .A2(n9264), .ZN(n11476) );
  OR2_X1 U11797 ( .A1(n9478), .A2(n11476), .ZN(n9267) );
  INV_X1 U11798 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9265) );
  OR2_X1 U11799 ( .A1(n9369), .A2(n9265), .ZN(n9266) );
  NAND4_X1 U11800 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n12608) );
  NAND2_X1 U11801 ( .A1(n9280), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9270) );
  OR2_X1 U11802 ( .A1(n12005), .A2(SI_7_), .ZN(n9274) );
  XNOR2_X1 U11803 ( .A(n9272), .B(n9271), .ZN(n9892) );
  OR2_X1 U11804 ( .A1(n9487), .A2(n9892), .ZN(n9273) );
  OAI211_X1 U11805 ( .C1(n14982), .C2(n9179), .A(n9274), .B(n9273), .ZN(n11471) );
  OR2_X1 U11806 ( .A1(n12608), .A2(n11471), .ZN(n12042) );
  NAND2_X1 U11807 ( .A1(n12608), .A2(n11471), .ZN(n12041) );
  INV_X1 U11808 ( .A(n15056), .ZN(n11284) );
  NAND2_X1 U11809 ( .A1(n6559), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9279) );
  INV_X1 U11810 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10817) );
  OR2_X1 U11811 ( .A1(n9369), .A2(n10817), .ZN(n9278) );
  XNOR2_X1 U11812 ( .A(n9292), .B(n15304), .ZN(n15067) );
  OR2_X1 U11813 ( .A1(n9478), .A2(n15067), .ZN(n9277) );
  INV_X1 U11814 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10795) );
  OR2_X1 U11815 ( .A1(n6558), .A2(n10795), .ZN(n9276) );
  INV_X1 U11816 ( .A(n9315), .ZN(n9284) );
  NAND2_X1 U11817 ( .A1(n9281), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9282) );
  MUX2_X1 U11818 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9282), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n9283) );
  INV_X1 U11819 ( .A(SI_8_), .ZN(n9872) );
  OR2_X1 U11820 ( .A1(n12005), .A2(n9872), .ZN(n9290) );
  OR2_X1 U11821 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  NAND2_X1 U11822 ( .A1(n9288), .A2(n9287), .ZN(n9873) );
  OR2_X1 U11823 ( .A1(n9487), .A2(n9873), .ZN(n9289) );
  OAI211_X1 U11824 ( .C1(n9179), .C2(n14995), .A(n9290), .B(n9289), .ZN(n15066) );
  NAND2_X1 U11825 ( .A1(n15055), .A2(n15061), .ZN(n9291) );
  INV_X1 U11826 ( .A(n15066), .ZN(n12046) );
  OR2_X1 U11827 ( .A1(n15045), .A2(n12046), .ZN(n12048) );
  NAND2_X1 U11828 ( .A1(n6559), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9298) );
  OAI21_X1 U11829 ( .B1(n9292), .B2(P3_REG3_REG_8__SCAN_IN), .A(
        P3_REG3_REG_9__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11830 ( .A1(n9293), .A2(n9307), .ZN(n15049) );
  INV_X1 U11831 ( .A(n15049), .ZN(n9294) );
  OR2_X1 U11832 ( .A1(n9423), .A2(n9294), .ZN(n9297) );
  INV_X1 U11833 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15307) );
  OR2_X1 U11834 ( .A1(n6553), .A2(n15307), .ZN(n9296) );
  INV_X1 U11835 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15236) );
  OR2_X1 U11836 ( .A1(n6558), .A2(n15236), .ZN(n9295) );
  NAND4_X1 U11837 ( .A1(n9298), .A2(n9297), .A3(n9296), .A4(n9295), .ZN(n12607) );
  OR2_X1 U11838 ( .A1(n9315), .A2(n9415), .ZN(n9299) );
  XNOR2_X1 U11839 ( .A(n9299), .B(n9313), .ZN(n10868) );
  OR2_X1 U11840 ( .A1(n12005), .A2(SI_9_), .ZN(n9305) );
  OR2_X1 U11841 ( .A1(n9301), .A2(n9300), .ZN(n9302) );
  AND2_X1 U11842 ( .A1(n9303), .A2(n9302), .ZN(n9876) );
  OR2_X1 U11843 ( .A1(n9487), .A2(n9876), .ZN(n9304) );
  OAI211_X1 U11844 ( .C1(n10868), .C2(n9179), .A(n9305), .B(n9304), .ZN(n15052) );
  OR2_X1 U11845 ( .A1(n12607), .A2(n15052), .ZN(n12052) );
  INV_X1 U11846 ( .A(n12052), .ZN(n9306) );
  NAND2_X1 U11847 ( .A1(n12607), .A2(n15052), .ZN(n12051) );
  NAND2_X1 U11848 ( .A1(n6559), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9312) );
  INV_X1 U11849 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10858) );
  OR2_X1 U11850 ( .A1(n6557), .A2(n10858), .ZN(n9311) );
  NAND2_X1 U11851 ( .A1(n9307), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9308) );
  AND2_X1 U11852 ( .A1(n9340), .A2(n9308), .ZN(n15034) );
  OR2_X1 U11853 ( .A1(n9478), .A2(n15034), .ZN(n9310) );
  INV_X1 U11854 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10859) );
  OR2_X1 U11855 ( .A1(n6553), .A2(n10859), .ZN(n9309) );
  INV_X1 U11856 ( .A(n9313), .ZN(n9314) );
  NAND2_X1 U11857 ( .A1(n9315), .A2(n9314), .ZN(n9334) );
  NAND2_X1 U11858 ( .A1(n9334), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9317) );
  INV_X1 U11859 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9316) );
  OR2_X1 U11860 ( .A1(n12005), .A2(SI_10_), .ZN(n9323) );
  OR2_X1 U11861 ( .A1(n9319), .A2(n9318), .ZN(n9320) );
  AND2_X1 U11862 ( .A1(n9321), .A2(n9320), .ZN(n9881) );
  OR2_X1 U11863 ( .A1(n9487), .A2(n9881), .ZN(n9322) );
  OAI211_X1 U11864 ( .C1(n10871), .C2(n9179), .A(n9323), .B(n9322), .ZN(n15033) );
  OR2_X1 U11865 ( .A1(n15044), .A2(n15033), .ZN(n12056) );
  NAND2_X1 U11866 ( .A1(n15044), .A2(n15033), .ZN(n12055) );
  NAND2_X1 U11867 ( .A1(n12056), .A2(n12055), .ZN(n15027) );
  INV_X1 U11868 ( .A(n15027), .ZN(n12159) );
  NAND2_X1 U11869 ( .A1(n6559), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9329) );
  INV_X1 U11870 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9324) );
  OR2_X1 U11871 ( .A1(n6557), .A2(n9324), .ZN(n9328) );
  INV_X1 U11872 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11384) );
  XNOR2_X1 U11873 ( .A(n9340), .B(n11384), .ZN(n12553) );
  OR2_X1 U11874 ( .A1(n9423), .A2(n12553), .ZN(n9327) );
  INV_X1 U11875 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9325) );
  OR2_X1 U11876 ( .A1(n9369), .A2(n9325), .ZN(n9326) );
  NAND4_X1 U11877 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n12606) );
  OR2_X1 U11878 ( .A1(n6773), .A2(n9330), .ZN(n9332) );
  AND2_X1 U11879 ( .A1(n9333), .A2(n9332), .ZN(n9896) );
  OR2_X1 U11880 ( .A1(n9487), .A2(n9896), .ZN(n9338) );
  OR2_X1 U11881 ( .A1(n12005), .A2(SI_11_), .ZN(n9337) );
  OAI21_X1 U11882 ( .B1(n9334), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9335) );
  XNOR2_X1 U11883 ( .A(n9335), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11549) );
  INV_X1 U11884 ( .A(n11549), .ZN(n11389) );
  NAND2_X1 U11885 ( .A1(n9460), .A2(n11389), .ZN(n9336) );
  NAND2_X1 U11886 ( .A1(n12606), .A2(n14603), .ZN(n12060) );
  NAND2_X1 U11887 ( .A1(n12059), .A2(n12060), .ZN(n14598) );
  NAND2_X1 U11888 ( .A1(n6559), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9345) );
  OAI21_X1 U11889 ( .B1(n9340), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n9341) );
  AND2_X1 U11890 ( .A1(n9341), .A2(n9366), .ZN(n12485) );
  OR2_X1 U11891 ( .A1(n9423), .A2(n12485), .ZN(n9344) );
  INV_X1 U11892 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11598) );
  OR2_X1 U11893 ( .A1(n9369), .A2(n11598), .ZN(n9343) );
  INV_X1 U11894 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14615) );
  OR2_X1 U11895 ( .A1(n6558), .A2(n14615), .ZN(n9342) );
  NAND4_X1 U11896 ( .A1(n9345), .A2(n9344), .A3(n9343), .A4(n9342), .ZN(n12605) );
  OR2_X1 U11897 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U11898 ( .A1(n9349), .A2(n9348), .ZN(n9914) );
  OR2_X1 U11899 ( .A1(n9914), .A2(n9487), .ZN(n9356) );
  NAND2_X1 U11900 ( .A1(n9351), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9352) );
  MUX2_X1 U11901 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9352), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9353) );
  NAND2_X1 U11902 ( .A1(n9353), .A2(n9055), .ZN(n12619) );
  INV_X1 U11903 ( .A(n12619), .ZN(n12625) );
  NAND2_X1 U11904 ( .A1(n9460), .A2(n12625), .ZN(n9355) );
  NAND2_X1 U11905 ( .A1(n9565), .A2(SI_12_), .ZN(n9354) );
  AND2_X1 U11906 ( .A1(n12059), .A2(n12064), .ZN(n14581) );
  NAND2_X1 U11907 ( .A1(n9357), .A2(n10158), .ZN(n9358) );
  NAND2_X1 U11908 ( .A1(n9359), .A2(n9358), .ZN(n9933) );
  OR2_X1 U11909 ( .A1(n9933), .A2(n9487), .ZN(n9364) );
  NAND2_X1 U11910 ( .A1(n9055), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9360) );
  MUX2_X1 U11911 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9360), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9361) );
  INV_X1 U11912 ( .A(n9361), .ZN(n9362) );
  NOR2_X1 U11913 ( .A1(n9362), .A2(n9383), .ZN(n12620) );
  AOI22_X1 U11914 ( .A1(n9565), .A2(SI_13_), .B1(n9460), .B2(n12620), .ZN(
        n9363) );
  NAND2_X1 U11915 ( .A1(n9364), .A2(n9363), .ZN(n14592) );
  NAND2_X1 U11916 ( .A1(n6559), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9373) );
  INV_X1 U11917 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9365) );
  OR2_X1 U11918 ( .A1(n6558), .A2(n9365), .ZN(n9372) );
  NAND2_X1 U11919 ( .A1(n9366), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9367) );
  AND2_X1 U11920 ( .A1(n9389), .A2(n9367), .ZN(n12539) );
  OR2_X1 U11921 ( .A1(n9478), .A2(n12539), .ZN(n9371) );
  INV_X1 U11922 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n9368) );
  OR2_X1 U11923 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND4_X1 U11924 ( .A1(n9373), .A2(n9372), .A3(n9371), .A4(n9370), .ZN(n12604) );
  AND2_X1 U11925 ( .A1(n14592), .A2(n12439), .ZN(n9376) );
  INV_X1 U11926 ( .A(n9376), .ZN(n12070) );
  AND2_X1 U11927 ( .A1(n14581), .A2(n12070), .ZN(n9374) );
  OR2_X1 U11928 ( .A1(n14592), .A2(n12439), .ZN(n12075) );
  INV_X1 U11929 ( .A(n12075), .ZN(n9377) );
  INV_X1 U11930 ( .A(n12064), .ZN(n9375) );
  NAND2_X1 U11931 ( .A1(n12605), .A2(n14610), .ZN(n12063) );
  OR2_X1 U11932 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  NAND2_X1 U11933 ( .A1(n9382), .A2(n9381), .ZN(n10035) );
  OR2_X1 U11934 ( .A1(n10035), .A2(n9487), .ZN(n9388) );
  OR2_X1 U11935 ( .A1(n9383), .A2(n9415), .ZN(n9385) );
  XNOR2_X1 U11936 ( .A(n9385), .B(n9384), .ZN(n12634) );
  INV_X1 U11937 ( .A(n12634), .ZN(n9386) );
  AOI22_X1 U11938 ( .A1(n9565), .A2(SI_14_), .B1(n9460), .B2(n9386), .ZN(n9387) );
  NAND2_X1 U11939 ( .A1(n9388), .A2(n9387), .ZN(n13002) );
  NAND2_X1 U11940 ( .A1(n6559), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9395) );
  INV_X1 U11941 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11666) );
  OR2_X1 U11942 ( .A1(n9369), .A2(n11666), .ZN(n9394) );
  NAND2_X1 U11943 ( .A1(n9389), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9390) );
  AND2_X1 U11944 ( .A1(n9404), .A2(n9390), .ZN(n12442) );
  OR2_X1 U11945 ( .A1(n9478), .A2(n12442), .ZN(n9393) );
  INV_X1 U11946 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n9391) );
  OR2_X1 U11947 ( .A1(n6557), .A2(n9391), .ZN(n9392) );
  OR2_X1 U11948 ( .A1(n13002), .A2(n14591), .ZN(n12071) );
  NAND2_X1 U11949 ( .A1(n13002), .A2(n14591), .ZN(n12926) );
  NAND2_X1 U11950 ( .A1(n12071), .A2(n12926), .ZN(n12168) );
  OR2_X1 U11951 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  NAND2_X1 U11952 ( .A1(n9399), .A2(n9398), .ZN(n10094) );
  OR2_X1 U11953 ( .A1(n10094), .A2(n9487), .ZN(n9403) );
  OR2_X1 U11954 ( .A1(n9400), .A2(n9415), .ZN(n9401) );
  XNOR2_X1 U11955 ( .A(n9401), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U11956 ( .A1(n9565), .A2(SI_15_), .B1(n9460), .B2(n12660), .ZN(
        n9402) );
  NAND2_X1 U11957 ( .A1(n9403), .A2(n9402), .ZN(n12930) );
  INV_X1 U11958 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14573) );
  OR2_X1 U11959 ( .A1(n6558), .A2(n14573), .ZN(n9409) );
  INV_X1 U11960 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n15434) );
  OR2_X1 U11961 ( .A1(n11984), .A2(n15434), .ZN(n9408) );
  NAND2_X1 U11962 ( .A1(n9404), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9405) );
  AND2_X1 U11963 ( .A1(n9421), .A2(n9405), .ZN(n12931) );
  OR2_X1 U11964 ( .A1(n9478), .A2(n12931), .ZN(n9407) );
  INV_X1 U11965 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14565) );
  OR2_X1 U11966 ( .A1(n6553), .A2(n14565), .ZN(n9406) );
  NAND4_X1 U11967 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n12602) );
  NAND2_X1 U11968 ( .A1(n12930), .A2(n12912), .ZN(n12080) );
  AND2_X1 U11969 ( .A1(n12926), .A2(n12080), .ZN(n9410) );
  OR2_X1 U11970 ( .A1(n12930), .A2(n12912), .ZN(n12073) );
  OR2_X1 U11971 ( .A1(n9412), .A2(n9411), .ZN(n9413) );
  NAND2_X1 U11972 ( .A1(n9414), .A2(n9413), .ZN(n10128) );
  OR2_X1 U11973 ( .A1(n10128), .A2(n9487), .ZN(n9420) );
  OR2_X1 U11974 ( .A1(n9416), .A2(n9415), .ZN(n9418) );
  XNOR2_X1 U11975 ( .A(n9418), .B(n9417), .ZN(n12674) );
  INV_X1 U11976 ( .A(n12674), .ZN(n12653) );
  AOI22_X1 U11977 ( .A1(n9565), .A2(SI_16_), .B1(n9460), .B2(n12653), .ZN(
        n9419) );
  NAND2_X1 U11978 ( .A1(n9420), .A2(n9419), .ZN(n12405) );
  NAND2_X1 U11979 ( .A1(n6559), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9427) );
  INV_X1 U11980 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12996) );
  OR2_X1 U11981 ( .A1(n6558), .A2(n12996), .ZN(n9426) );
  NAND2_X1 U11982 ( .A1(n9421), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9422) );
  AND2_X1 U11983 ( .A1(n9436), .A2(n9422), .ZN(n12917) );
  OR2_X1 U11984 ( .A1(n9478), .A2(n12917), .ZN(n9425) );
  INV_X1 U11985 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12918) );
  OR2_X1 U11986 ( .A1(n9369), .A2(n12918), .ZN(n9424) );
  OR2_X1 U11987 ( .A1(n12405), .A2(n12925), .ZN(n12074) );
  NAND2_X1 U11988 ( .A1(n12405), .A2(n12925), .ZN(n12081) );
  NAND2_X1 U11989 ( .A1(n12916), .A2(n12915), .ZN(n12914) );
  OR2_X1 U11990 ( .A1(n9429), .A2(n9428), .ZN(n9430) );
  NAND2_X1 U11991 ( .A1(n9431), .A2(n9430), .ZN(n10133) );
  OR2_X1 U11992 ( .A1(n10133), .A2(n9487), .ZN(n9435) );
  NAND2_X1 U11993 ( .A1(n9432), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9433) );
  XNOR2_X1 U11994 ( .A(n9433), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U11995 ( .A1(n9565), .A2(SI_17_), .B1(n9460), .B2(n12705), .ZN(
        n9434) );
  NAND2_X1 U11996 ( .A1(n6559), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9441) );
  INV_X1 U11997 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12992) );
  OR2_X1 U11998 ( .A1(n6558), .A2(n12992), .ZN(n9440) );
  NAND2_X1 U11999 ( .A1(n9436), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9437) );
  AND2_X1 U12000 ( .A1(n9450), .A2(n9437), .ZN(n12904) );
  OR2_X1 U12001 ( .A1(n9478), .A2(n12904), .ZN(n9439) );
  INV_X1 U12002 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12905) );
  OR2_X1 U12003 ( .A1(n6553), .A2(n12905), .ZN(n9438) );
  OR2_X1 U12004 ( .A1(n12903), .A2(n12913), .ZN(n12090) );
  NAND2_X1 U12005 ( .A1(n12903), .A2(n12913), .ZN(n12087) );
  NAND2_X1 U12006 ( .A1(n12090), .A2(n12087), .ZN(n12896) );
  INV_X1 U12007 ( .A(n12896), .ZN(n12901) );
  OR2_X1 U12008 ( .A1(n6774), .A2(n9442), .ZN(n9444) );
  NAND2_X1 U12009 ( .A1(n9445), .A2(n9444), .ZN(n10179) );
  OR2_X1 U12010 ( .A1(n10179), .A2(n9487), .ZN(n9449) );
  NAND2_X1 U12011 ( .A1(n9446), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9447) );
  XNOR2_X1 U12012 ( .A(n9447), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U12013 ( .A1(n9565), .A2(SI_18_), .B1(n9460), .B2(n12716), .ZN(
        n9448) );
  NAND2_X1 U12014 ( .A1(n9555), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9455) );
  INV_X1 U12015 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n15365) );
  OR2_X1 U12016 ( .A1(n11984), .A2(n15365), .ZN(n9454) );
  NAND2_X1 U12017 ( .A1(n9450), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9451) );
  AND2_X1 U12018 ( .A1(n9463), .A2(n9451), .ZN(n12886) );
  OR2_X1 U12019 ( .A1(n9478), .A2(n12886), .ZN(n9453) );
  INV_X1 U12020 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12887) );
  OR2_X1 U12021 ( .A1(n6553), .A2(n12887), .ZN(n9452) );
  NAND2_X1 U12022 ( .A1(n12986), .A2(n12900), .ZN(n12088) );
  NAND2_X1 U12023 ( .A1(n12890), .A2(n12089), .ZN(n12876) );
  INV_X1 U12024 ( .A(n12876), .ZN(n9470) );
  OR2_X1 U12025 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U12026 ( .A1(n9459), .A2(n9458), .ZN(n10256) );
  NAND2_X1 U12027 ( .A1(n10256), .A2(n12004), .ZN(n9462) );
  AOI22_X1 U12028 ( .A1(n9565), .A2(n10255), .B1(n9460), .B2(n6555), .ZN(n9461) );
  NAND2_X1 U12029 ( .A1(n6559), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9468) );
  INV_X1 U12030 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12984) );
  OR2_X1 U12031 ( .A1(n6557), .A2(n12984), .ZN(n9467) );
  NAND2_X1 U12032 ( .A1(n9463), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9464) );
  AND2_X1 U12033 ( .A1(n9476), .A2(n9464), .ZN(n12877) );
  OR2_X1 U12034 ( .A1(n9478), .A2(n12877), .ZN(n9466) );
  INV_X1 U12035 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12878) );
  OR2_X1 U12036 ( .A1(n9369), .A2(n12878), .ZN(n9465) );
  NAND4_X1 U12037 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n12884) );
  NAND2_X1 U12038 ( .A1(n13062), .A2(n12884), .ZN(n12094) );
  INV_X1 U12039 ( .A(n12095), .ZN(n9469) );
  NAND2_X1 U12040 ( .A1(n9471), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U12041 ( .A1(n9473), .A2(n9472), .ZN(n10505) );
  OR2_X1 U12042 ( .A1(n12005), .A2(n10504), .ZN(n9474) );
  NAND2_X1 U12043 ( .A1(n9555), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9482) );
  INV_X1 U12044 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13056) );
  OR2_X1 U12045 ( .A1(n11984), .A2(n13056), .ZN(n9481) );
  NAND2_X1 U12046 ( .A1(n9476), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U12047 ( .A1(n9490), .A2(n9477), .ZN(n12533) );
  INV_X1 U12048 ( .A(n12533), .ZN(n12863) );
  OR2_X1 U12049 ( .A1(n9478), .A2(n12863), .ZN(n9480) );
  INV_X1 U12050 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12864) );
  OR2_X1 U12051 ( .A1(n6553), .A2(n12864), .ZN(n9479) );
  XNOR2_X1 U12052 ( .A(n12866), .B(n12872), .ZN(n12858) );
  INV_X1 U12053 ( .A(n12858), .ZN(n12855) );
  NAND2_X1 U12054 ( .A1(n12856), .A2(n12855), .ZN(n12854) );
  OR2_X1 U12055 ( .A1(n12866), .A2(n12872), .ZN(n12100) );
  NAND2_X1 U12056 ( .A1(n12854), .A2(n12100), .ZN(n12847) );
  OR2_X1 U12057 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  NAND2_X1 U12058 ( .A1(n9486), .A2(n9485), .ZN(n10675) );
  INV_X1 U12059 ( .A(SI_21_), .ZN(n10674) );
  OR2_X1 U12060 ( .A1(n12005), .A2(n10674), .ZN(n9488) );
  NAND2_X1 U12061 ( .A1(n9490), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U12062 ( .A1(n9502), .A2(n9491), .ZN(n12849) );
  NAND2_X1 U12063 ( .A1(n9570), .A2(n12849), .ZN(n9496) );
  INV_X1 U12064 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12974) );
  OR2_X1 U12065 ( .A1(n6557), .A2(n12974), .ZN(n9495) );
  INV_X1 U12066 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13052) );
  OR2_X1 U12067 ( .A1(n11984), .A2(n13052), .ZN(n9494) );
  INV_X1 U12068 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n9492) );
  OR2_X1 U12069 ( .A1(n9369), .A2(n9492), .ZN(n9493) );
  NAND4_X1 U12070 ( .A1(n9496), .A2(n9495), .A3(n9494), .A4(n9493), .ZN(n12860) );
  NOR2_X1 U12071 ( .A1(n12848), .A2(n12834), .ZN(n12106) );
  NAND2_X1 U12072 ( .A1(n12848), .A2(n12834), .ZN(n12105) );
  XNOR2_X1 U12073 ( .A(n9498), .B(n9497), .ZN(n10698) );
  NAND2_X1 U12074 ( .A1(n10698), .A2(n12004), .ZN(n9501) );
  OR2_X1 U12075 ( .A1(n12005), .A2(n9499), .ZN(n9500) );
  NAND2_X1 U12076 ( .A1(n9502), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U12077 ( .A1(n9515), .A2(n9503), .ZN(n12838) );
  NAND2_X1 U12078 ( .A1(n9570), .A2(n12838), .ZN(n9508) );
  NAND2_X1 U12079 ( .A1(n9555), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9507) );
  INV_X1 U12080 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13048) );
  OR2_X1 U12081 ( .A1(n11984), .A2(n13048), .ZN(n9506) );
  INV_X1 U12082 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9504) );
  OR2_X1 U12083 ( .A1(n9369), .A2(n9504), .ZN(n9505) );
  NAND4_X1 U12084 ( .A1(n9508), .A2(n9507), .A3(n9506), .A4(n9505), .ZN(n12818) );
  XNOR2_X1 U12085 ( .A(n9510), .B(n9509), .ZN(n10958) );
  NAND2_X1 U12086 ( .A1(n10958), .A2(n12004), .ZN(n9512) );
  OR2_X1 U12087 ( .A1(n12005), .A2(n10960), .ZN(n9511) );
  INV_X1 U12088 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U12089 ( .A1(n9555), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U12090 ( .A1(n9571), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9513) );
  AND2_X1 U12091 ( .A1(n9514), .A2(n9513), .ZN(n9518) );
  NAND2_X1 U12092 ( .A1(n9515), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U12093 ( .A1(n9524), .A2(n9516), .ZN(n12825) );
  NAND2_X1 U12094 ( .A1(n12825), .A2(n9570), .ZN(n9517) );
  XNOR2_X1 U12095 ( .A(n12824), .B(n12803), .ZN(n12822) );
  OR2_X1 U12096 ( .A1(n12824), .A2(n12833), .ZN(n12119) );
  INV_X1 U12097 ( .A(n12119), .ZN(n9520) );
  XNOR2_X1 U12098 ( .A(n9521), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U12099 ( .A1(n11317), .A2(n12004), .ZN(n9523) );
  INV_X1 U12100 ( .A(SI_24_), .ZN(n11318) );
  OR2_X1 U12101 ( .A1(n12005), .A2(n11318), .ZN(n9522) );
  NAND2_X1 U12102 ( .A1(n9524), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U12103 ( .A1(n9534), .A2(n9525), .ZN(n12811) );
  NAND2_X1 U12104 ( .A1(n12811), .A2(n9570), .ZN(n9528) );
  AOI22_X1 U12105 ( .A1(n9555), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n6559), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U12106 ( .A1(n9184), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9526) );
  OR2_X1 U12107 ( .A1(n12810), .A2(n12821), .ZN(n12120) );
  NAND2_X1 U12108 ( .A1(n12810), .A2(n12821), .ZN(n12121) );
  NAND2_X1 U12109 ( .A1(n12809), .A2(n9529), .ZN(n12808) );
  XNOR2_X1 U12110 ( .A(n9531), .B(n9530), .ZN(n11402) );
  NAND2_X1 U12111 ( .A1(n11402), .A2(n12004), .ZN(n9533) );
  OR2_X1 U12112 ( .A1(n12005), .A2(n15435), .ZN(n9532) );
  NAND2_X1 U12113 ( .A1(n9534), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U12114 ( .A1(n9544), .A2(n9535), .ZN(n12797) );
  NAND2_X1 U12115 ( .A1(n12797), .A2(n9570), .ZN(n9538) );
  AOI22_X1 U12116 ( .A1(n9555), .A2(P3_REG1_REG_25__SCAN_IN), .B1(n6559), .B2(
        P3_REG0_REG_25__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U12117 ( .A1(n9184), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U12118 ( .A1(n12499), .A2(n12806), .ZN(n9539) );
  INV_X1 U12119 ( .A(n9539), .ZN(n12126) );
  XNOR2_X1 U12120 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n9540) );
  XNOR2_X1 U12121 ( .A(n9541), .B(n9540), .ZN(n11501) );
  NAND2_X1 U12122 ( .A1(n11501), .A2(n12004), .ZN(n9543) );
  OR2_X1 U12123 ( .A1(n12005), .A2(n11502), .ZN(n9542) );
  NAND2_X1 U12124 ( .A1(n9544), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U12125 ( .A1(n9553), .A2(n9545), .ZN(n12783) );
  NAND2_X1 U12126 ( .A1(n12783), .A2(n9570), .ZN(n9550) );
  INV_X1 U12127 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U12128 ( .A1(n9184), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U12129 ( .A1(n9571), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9546) );
  OAI211_X1 U12130 ( .C1(n6558), .C2(n12953), .A(n9547), .B(n9546), .ZN(n9548)
         );
  INV_X1 U12131 ( .A(n9548), .ZN(n9549) );
  NOR2_X1 U12132 ( .A1(n12579), .A2(n12765), .ZN(n12127) );
  XOR2_X1 U12133 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .Z(n9551) );
  XNOR2_X1 U12134 ( .A(n9552), .B(n9551), .ZN(n11588) );
  AOI22_X2 U12135 ( .A1(n11588), .A2(n12004), .B1(SI_27_), .B2(n9565), .ZN(
        n13032) );
  NAND2_X1 U12136 ( .A1(n9553), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U12137 ( .A1(n9568), .A2(n9554), .ZN(n12770) );
  NAND2_X1 U12138 ( .A1(n12770), .A2(n9570), .ZN(n9560) );
  INV_X1 U12139 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n15289) );
  NAND2_X1 U12140 ( .A1(n9184), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U12141 ( .A1(n9555), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9556) );
  OAI211_X1 U12142 ( .C1(n11984), .C2(n15289), .A(n9557), .B(n9556), .ZN(n9558) );
  INV_X1 U12143 ( .A(n9558), .ZN(n9559) );
  NOR2_X1 U12144 ( .A1(n13032), .A2(n12777), .ZN(n9562) );
  INV_X1 U12145 ( .A(n13032), .ZN(n9561) );
  INV_X1 U12146 ( .A(n9562), .ZN(n12138) );
  XNOR2_X1 U12147 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n9563) );
  XNOR2_X1 U12148 ( .A(n9564), .B(n9563), .ZN(n11728) );
  NAND2_X1 U12149 ( .A1(n11728), .A2(n12004), .ZN(n9567) );
  NAND2_X1 U12150 ( .A1(n9565), .A2(SI_28_), .ZN(n9566) );
  INV_X1 U12151 ( .A(n13029), .ZN(n9577) );
  NAND2_X1 U12152 ( .A1(n9568), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U12153 ( .A1(n12381), .A2(n9569), .ZN(n12755) );
  NAND2_X1 U12154 ( .A1(n12755), .A2(n9570), .ZN(n9576) );
  INV_X1 U12155 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U12156 ( .A1(n6559), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9573) );
  NAND2_X1 U12157 ( .A1(n9184), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9572) );
  OAI211_X1 U12158 ( .C1(n6557), .C2(n12945), .A(n9573), .B(n9572), .ZN(n9574)
         );
  INV_X1 U12159 ( .A(n9574), .ZN(n9575) );
  NAND2_X1 U12160 ( .A1(n9576), .A2(n9575), .ZN(n12597) );
  NAND2_X1 U12161 ( .A1(n9577), .A2(n12766), .ZN(n12139) );
  INV_X1 U12162 ( .A(n12139), .ZN(n9578) );
  NAND2_X1 U12163 ( .A1(n13029), .A2(n12597), .ZN(n12146) );
  INV_X1 U12164 ( .A(n12146), .ZN(n9579) );
  NAND2_X1 U12165 ( .A1(n13009), .A2(n11756), .ZN(n13007) );
  NAND2_X1 U12166 ( .A1(n13006), .A2(n15108), .ZN(n9581) );
  NAND2_X1 U12167 ( .A1(n9581), .A2(n9580), .ZN(n15112) );
  INV_X1 U12168 ( .A(n15099), .ZN(n9582) );
  OR2_X1 U12169 ( .A1(n13008), .A2(n9582), .ZN(n11088) );
  INV_X1 U12170 ( .A(n11088), .ZN(n9583) );
  NAND2_X1 U12171 ( .A1(n15112), .A2(n9584), .ZN(n11093) );
  INV_X1 U12172 ( .A(n11098), .ZN(n9586) );
  NAND2_X1 U12173 ( .A1(n9585), .A2(n9586), .ZN(n9587) );
  INV_X1 U12174 ( .A(n15090), .ZN(n9588) );
  AND2_X1 U12175 ( .A1(n12611), .A2(n9588), .ZN(n9589) );
  INV_X1 U12176 ( .A(n11240), .ZN(n12008) );
  OR2_X1 U12177 ( .A1(n12610), .A2(n12008), .ZN(n9590) );
  INV_X1 U12178 ( .A(n15078), .ZN(n11505) );
  NAND2_X1 U12179 ( .A1(n12609), .A2(n11505), .ZN(n11283) );
  INV_X1 U12180 ( .A(n15061), .ZN(n12161) );
  INV_X1 U12181 ( .A(n11471), .ZN(n9592) );
  NAND2_X1 U12182 ( .A1(n12608), .A2(n9592), .ZN(n15058) );
  AND2_X1 U12183 ( .A1(n12161), .A2(n15058), .ZN(n9593) );
  AND2_X1 U12184 ( .A1(n11283), .A2(n9593), .ZN(n9598) );
  INV_X1 U12185 ( .A(n9593), .ZN(n9594) );
  OR2_X1 U12186 ( .A1(n9594), .A2(n15056), .ZN(n9596) );
  OR2_X1 U12187 ( .A1(n15045), .A2(n15066), .ZN(n9595) );
  NAND2_X1 U12188 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  NAND2_X1 U12189 ( .A1(n12052), .A2(n12051), .ZN(n15041) );
  NAND2_X1 U12190 ( .A1(n15042), .A2(n15041), .ZN(n15040) );
  INV_X1 U12191 ( .A(n15052), .ZN(n9599) );
  NAND2_X1 U12192 ( .A1(n12607), .A2(n9599), .ZN(n9600) );
  NAND2_X1 U12193 ( .A1(n15040), .A2(n9600), .ZN(n15028) );
  INV_X1 U12194 ( .A(n15033), .ZN(n9601) );
  NAND2_X1 U12195 ( .A1(n15044), .A2(n9601), .ZN(n9602) );
  OR2_X1 U12196 ( .A1(n11593), .A2(n6607), .ZN(n9603) );
  INV_X1 U12197 ( .A(n14610), .ZN(n12491) );
  NAND2_X1 U12198 ( .A1(n12605), .A2(n12491), .ZN(n14586) );
  OR2_X1 U12199 ( .A1(n6607), .A2(n14586), .ZN(n9605) );
  NAND2_X1 U12200 ( .A1(n14592), .A2(n12604), .ZN(n9604) );
  NAND2_X1 U12201 ( .A1(n13002), .A2(n12603), .ZN(n9606) );
  NAND2_X1 U12202 ( .A1(n9607), .A2(n9606), .ZN(n12923) );
  AND2_X1 U12203 ( .A1(n12930), .A2(n12602), .ZN(n9608) );
  NAND2_X1 U12204 ( .A1(n12405), .A2(n12601), .ZN(n9609) );
  NAND2_X1 U12205 ( .A1(n12903), .A2(n12883), .ZN(n9610) );
  NAND2_X2 U12206 ( .A1(n7597), .A2(n6571), .ZN(n12882) );
  INV_X1 U12207 ( .A(n12900), .ZN(n12600) );
  OR2_X1 U12208 ( .A1(n12986), .A2(n12600), .ZN(n9611) );
  INV_X1 U12209 ( .A(n12884), .ZN(n12531) );
  OR2_X1 U12210 ( .A1(n13062), .A2(n12531), .ZN(n9613) );
  NAND2_X1 U12211 ( .A1(n12866), .A2(n12599), .ZN(n9614) );
  OR2_X1 U12212 ( .A1(n12848), .A2(n12860), .ZN(n12104) );
  NAND2_X1 U12213 ( .A1(n12848), .A2(n12860), .ZN(n12103) );
  AND2_X1 U12214 ( .A1(n12837), .A2(n12818), .ZN(n9617) );
  OR2_X1 U12215 ( .A1(n12837), .A2(n12818), .ZN(n9616) );
  NAND2_X1 U12216 ( .A1(n12824), .A2(n12803), .ZN(n9619) );
  NAND2_X1 U12217 ( .A1(n12810), .A2(n12791), .ZN(n9620) );
  NAND2_X1 U12218 ( .A1(n12790), .A2(n12789), .ZN(n12788) );
  XNOR2_X1 U12219 ( .A(n9622), .B(n12176), .ZN(n9632) );
  NAND2_X1 U12220 ( .A1(n12180), .A2(n12190), .ZN(n9666) );
  NAND2_X1 U12221 ( .A1(n9683), .A2(n12014), .ZN(n12184) );
  INV_X1 U12222 ( .A(n9623), .ZN(n12187) );
  NAND2_X1 U12223 ( .A1(n12187), .A2(n10376), .ZN(n10355) );
  NAND2_X1 U12224 ( .A1(n9179), .A2(n10355), .ZN(n10641) );
  INV_X1 U12225 ( .A(n10641), .ZN(n9624) );
  INV_X1 U12226 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n9627) );
  NAND2_X1 U12227 ( .A1(n6559), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9626) );
  NAND2_X1 U12228 ( .A1(n9184), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9625) );
  OAI211_X1 U12229 ( .C1(n9627), .C2(n6557), .A(n9626), .B(n9625), .ZN(n9628)
         );
  INV_X1 U12230 ( .A(n9628), .ZN(n9629) );
  AND2_X1 U12231 ( .A1(n12187), .A2(P3_B_REG_SCAN_IN), .ZN(n9630) );
  OR2_X1 U12232 ( .A1(n15105), .A2(n9630), .ZN(n12742) );
  OAI22_X1 U12233 ( .A1(n12766), .A2(n15107), .B1(n12148), .B2(n12742), .ZN(
        n9631) );
  NAND2_X1 U12234 ( .A1(n9633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9634) );
  MUX2_X1 U12235 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9634), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9636) );
  INV_X1 U12236 ( .A(n9637), .ZN(n9643) );
  NAND2_X1 U12237 ( .A1(n9643), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9638) );
  MUX2_X1 U12238 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9638), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9639) );
  NAND2_X1 U12239 ( .A1(n9639), .A2(n9633), .ZN(n11404) );
  INV_X1 U12240 ( .A(n9640), .ZN(n9641) );
  NAND2_X1 U12241 ( .A1(n9641), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9642) );
  MUX2_X1 U12242 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9642), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9644) );
  NAND2_X1 U12243 ( .A1(n9644), .A2(n9643), .ZN(n11320) );
  XNOR2_X1 U12244 ( .A(n11320), .B(P3_B_REG_SCAN_IN), .ZN(n9645) );
  NAND2_X1 U12245 ( .A1(n11404), .A2(n9645), .ZN(n9646) );
  INV_X1 U12246 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U12247 ( .A1(n10008), .A2(n9647), .ZN(n9649) );
  NAND2_X1 U12248 ( .A1(n11504), .A2(n11320), .ZN(n9648) );
  INV_X1 U12249 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U12250 ( .A1(n10008), .A2(n9650), .ZN(n9652) );
  NAND2_X1 U12251 ( .A1(n11504), .A2(n11404), .ZN(n9651) );
  NAND2_X1 U12252 ( .A1(n13079), .A2(n13077), .ZN(n9681) );
  NOR2_X1 U12253 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .ZN(
        n9656) );
  NOR4_X1 U12254 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9655) );
  NOR4_X1 U12255 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n9654) );
  NOR4_X1 U12256 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n9653) );
  NAND4_X1 U12257 ( .A1(n9656), .A2(n9655), .A3(n9654), .A4(n9653), .ZN(n9662)
         );
  NOR4_X1 U12258 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9660) );
  NOR4_X1 U12259 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n9659) );
  NOR4_X1 U12260 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9658) );
  NOR4_X1 U12261 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9657) );
  NAND4_X1 U12262 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n9661)
         );
  OAI21_X1 U12263 ( .B1(n9662), .B2(n9661), .A(n10008), .ZN(n9678) );
  INV_X1 U12264 ( .A(n9678), .ZN(n9670) );
  NOR2_X1 U12265 ( .A1(n9681), .A2(n9670), .ZN(n10628) );
  NOR2_X1 U12266 ( .A1(n11404), .A2(n11320), .ZN(n9663) );
  NAND2_X1 U12267 ( .A1(n9059), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9665) );
  XNOR2_X1 U12268 ( .A(n9665), .B(n9134), .ZN(n10353) );
  NOR2_X1 U12269 ( .A1(n9684), .A2(n12143), .ZN(n10972) );
  NAND2_X1 U12270 ( .A1(n10624), .A2(n10972), .ZN(n10640) );
  OR2_X1 U12271 ( .A1(n10611), .A2(n12014), .ZN(n12183) );
  NOR2_X1 U12272 ( .A1(n9666), .A2(n12183), .ZN(n10629) );
  NAND2_X1 U12273 ( .A1(n10624), .A2(n10629), .ZN(n9667) );
  NAND2_X1 U12274 ( .A1(n10640), .A2(n9667), .ZN(n9668) );
  NAND2_X1 U12275 ( .A1(n10628), .A2(n9668), .ZN(n9672) );
  INV_X1 U12276 ( .A(n13079), .ZN(n9669) );
  NAND2_X1 U12277 ( .A1(n9669), .A2(n9686), .ZN(n9679) );
  NAND3_X1 U12278 ( .A1(n10643), .A2(n10624), .A3(n10626), .ZN(n9671) );
  INV_X1 U12279 ( .A(n12385), .ZN(n9674) );
  INV_X1 U12280 ( .A(n9675), .ZN(n9676) );
  AND2_X1 U12281 ( .A1(n9678), .A2(n10624), .ZN(n9680) );
  NAND2_X1 U12282 ( .A1(n9684), .A2(n12133), .ZN(n10632) );
  NAND2_X1 U12283 ( .A1(n9682), .A2(n12143), .ZN(n10926) );
  AND2_X1 U12284 ( .A1(n10632), .A2(n10926), .ZN(n10928) );
  OAI22_X1 U12285 ( .A1(n12180), .A2(n12012), .B1(n9683), .B2(n15098), .ZN(
        n9685) );
  AOI21_X1 U12286 ( .B1(n9685), .B2(n9684), .A(n12133), .ZN(n9687) );
  MUX2_X1 U12287 ( .A(n10928), .B(n9687), .S(n9686), .Z(n9688) );
  INV_X1 U12288 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12289 ( .A1(n15179), .A2(n9689), .ZN(n9690) );
  INV_X1 U12290 ( .A(n15098), .ZN(n15065) );
  AND2_X1 U12291 ( .A1(n15181), .A2(n15065), .ZN(n12938) );
  NAND2_X1 U12292 ( .A1(n9693), .A2(n9692), .ZN(P3_U3488) );
  NAND2_X1 U12293 ( .A1(n8764), .A2(n9714), .ZN(n9696) );
  INV_X1 U12294 ( .A(n9696), .ZN(n9695) );
  OAI22_X1 U12295 ( .A1(n9698), .A2(n13528), .B1(n11004), .B2(n6560), .ZN(
        n10163) );
  NAND2_X1 U12296 ( .A1(n10160), .A2(n9699), .ZN(n10221) );
  XNOR2_X1 U12297 ( .A(n9807), .B(n11071), .ZN(n9700) );
  NAND2_X1 U12298 ( .A1(n13234), .A2(n9714), .ZN(n9701) );
  NAND2_X1 U12299 ( .A1(n9700), .A2(n9701), .ZN(n9705) );
  INV_X1 U12300 ( .A(n9700), .ZN(n9703) );
  INV_X1 U12301 ( .A(n9701), .ZN(n9702) );
  NAND2_X1 U12302 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  AND2_X1 U12303 ( .A1(n9705), .A2(n9704), .ZN(n10222) );
  INV_X1 U12304 ( .A(n10323), .ZN(n9707) );
  XNOR2_X1 U12305 ( .A(n9807), .B(n10273), .ZN(n9709) );
  AND2_X1 U12306 ( .A1(n13233), .A2(n13564), .ZN(n9708) );
  XNOR2_X1 U12307 ( .A(n9709), .B(n9708), .ZN(n10322) );
  INV_X1 U12308 ( .A(n10322), .ZN(n9706) );
  XNOR2_X1 U12309 ( .A(n10393), .B(n9807), .ZN(n9711) );
  AND2_X1 U12310 ( .A1(n13232), .A2(n13564), .ZN(n9710) );
  OR2_X1 U12311 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  NAND2_X1 U12312 ( .A1(n9711), .A2(n9710), .ZN(n9712) );
  AND2_X1 U12313 ( .A1(n9713), .A2(n9712), .ZN(n10258) );
  XNOR2_X1 U12314 ( .A(n10989), .B(n9824), .ZN(n9715) );
  NAND2_X1 U12315 ( .A1(n13231), .A2(n13564), .ZN(n9716) );
  NAND2_X1 U12316 ( .A1(n9715), .A2(n9716), .ZN(n9720) );
  INV_X1 U12317 ( .A(n9715), .ZN(n9718) );
  INV_X1 U12318 ( .A(n9716), .ZN(n9717) );
  NAND2_X1 U12319 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  XNOR2_X1 U12320 ( .A(n14910), .B(n9824), .ZN(n9721) );
  NAND2_X1 U12321 ( .A1(n13230), .A2(n9813), .ZN(n9722) );
  XNOR2_X1 U12322 ( .A(n9721), .B(n9722), .ZN(n10570) );
  INV_X1 U12323 ( .A(n9721), .ZN(n9724) );
  INV_X1 U12324 ( .A(n9722), .ZN(n9723) );
  NAND2_X1 U12325 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  XNOR2_X1 U12326 ( .A(n14917), .B(n9807), .ZN(n9728) );
  NAND2_X1 U12327 ( .A1(n13229), .A2(n9813), .ZN(n9726) );
  XNOR2_X1 U12328 ( .A(n9728), .B(n9726), .ZN(n10649) );
  NAND2_X1 U12329 ( .A1(n10650), .A2(n10649), .ZN(n9730) );
  INV_X1 U12330 ( .A(n9726), .ZN(n9727) );
  NAND2_X1 U12331 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  XNOR2_X1 U12332 ( .A(n10913), .B(n9824), .ZN(n9731) );
  NAND2_X1 U12333 ( .A1(n13228), .A2(n9813), .ZN(n9732) );
  NAND2_X1 U12334 ( .A1(n9731), .A2(n9732), .ZN(n10734) );
  INV_X1 U12335 ( .A(n9731), .ZN(n9734) );
  INV_X1 U12336 ( .A(n9732), .ZN(n9733) );
  NAND2_X1 U12337 ( .A1(n9734), .A2(n9733), .ZN(n10733) );
  XNOR2_X1 U12338 ( .A(n11250), .B(n9824), .ZN(n9738) );
  NAND2_X1 U12339 ( .A1(n13227), .A2(n9813), .ZN(n9737) );
  XNOR2_X1 U12340 ( .A(n9738), .B(n9737), .ZN(n10964) );
  NAND2_X1 U12341 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  XNOR2_X1 U12342 ( .A(n11277), .B(n9807), .ZN(n9740) );
  AND2_X1 U12343 ( .A1(n13226), .A2(n13564), .ZN(n9741) );
  NAND2_X1 U12344 ( .A1(n9740), .A2(n9741), .ZN(n9745) );
  INV_X1 U12345 ( .A(n9740), .ZN(n9743) );
  INV_X1 U12346 ( .A(n9741), .ZN(n9742) );
  NAND2_X1 U12347 ( .A1(n9743), .A2(n9742), .ZN(n9744) );
  AND2_X1 U12348 ( .A1(n9745), .A2(n9744), .ZN(n11193) );
  XNOR2_X1 U12349 ( .A(n11479), .B(n9807), .ZN(n9746) );
  NAND2_X1 U12350 ( .A1(n13225), .A2(n9813), .ZN(n9747) );
  XNOR2_X1 U12351 ( .A(n9746), .B(n9747), .ZN(n11333) );
  INV_X1 U12352 ( .A(n9746), .ZN(n9748) );
  NAND2_X1 U12353 ( .A1(n9748), .A2(n9747), .ZN(n11430) );
  XNOR2_X1 U12354 ( .A(n13578), .B(n9807), .ZN(n9749) );
  NAND2_X1 U12355 ( .A1(n13224), .A2(n9813), .ZN(n9750) );
  XNOR2_X1 U12356 ( .A(n9749), .B(n9750), .ZN(n11431) );
  INV_X1 U12357 ( .A(n9749), .ZN(n9751) );
  NAND2_X1 U12358 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U12359 ( .A1(n11434), .A2(n9752), .ZN(n11560) );
  XNOR2_X1 U12360 ( .A(n11575), .B(n9807), .ZN(n9753) );
  AND2_X1 U12361 ( .A1(n13223), .A2(n13564), .ZN(n9754) );
  NAND2_X1 U12362 ( .A1(n9753), .A2(n9754), .ZN(n9760) );
  INV_X1 U12363 ( .A(n9753), .ZN(n9756) );
  INV_X1 U12364 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U12365 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NAND2_X1 U12366 ( .A1(n9760), .A2(n9757), .ZN(n11559) );
  INV_X1 U12367 ( .A(n11559), .ZN(n9758) );
  XNOR2_X1 U12368 ( .A(n13718), .B(n9807), .ZN(n9761) );
  NAND2_X1 U12369 ( .A1(n13222), .A2(n9813), .ZN(n9762) );
  XNOR2_X1 U12370 ( .A(n9761), .B(n9762), .ZN(n11657) );
  XNOR2_X1 U12371 ( .A(n13715), .B(n9824), .ZN(n14626) );
  NAND2_X1 U12372 ( .A1(n13519), .A2(n9813), .ZN(n13203) );
  INV_X1 U12373 ( .A(n9761), .ZN(n9763) );
  AND2_X1 U12374 ( .A1(n9763), .A2(n9762), .ZN(n13199) );
  AOI21_X1 U12375 ( .B1(n14626), .B2(n13203), .A(n13199), .ZN(n9764) );
  XNOR2_X1 U12376 ( .A(n14637), .B(n9807), .ZN(n9768) );
  NAND2_X1 U12377 ( .A1(n13221), .A2(n9813), .ZN(n9769) );
  XNOR2_X1 U12378 ( .A(n9768), .B(n9769), .ZN(n14631) );
  NAND2_X1 U12379 ( .A1(n9767), .A2(n9766), .ZN(n14630) );
  INV_X1 U12380 ( .A(n9768), .ZN(n9770) );
  NAND2_X1 U12381 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  XNOR2_X1 U12382 ( .A(n13656), .B(n9807), .ZN(n9772) );
  NAND2_X1 U12383 ( .A1(n13517), .A2(n9813), .ZN(n9773) );
  XNOR2_X1 U12384 ( .A(n9772), .B(n9773), .ZN(n13137) );
  NAND2_X2 U12385 ( .A1(n13136), .A2(n13137), .ZN(n13135) );
  INV_X1 U12386 ( .A(n9772), .ZN(n9774) );
  NAND2_X1 U12387 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  XNOR2_X1 U12388 ( .A(n13651), .B(n9807), .ZN(n9776) );
  AND2_X1 U12389 ( .A1(n13220), .A2(n13564), .ZN(n9777) );
  NAND2_X1 U12390 ( .A1(n9776), .A2(n9777), .ZN(n9782) );
  INV_X1 U12391 ( .A(n9776), .ZN(n9779) );
  INV_X1 U12392 ( .A(n9777), .ZN(n9778) );
  NAND2_X1 U12393 ( .A1(n9779), .A2(n9778), .ZN(n9780) );
  NAND2_X1 U12394 ( .A1(n9782), .A2(n9780), .ZN(n13172) );
  XNOR2_X1 U12395 ( .A(n13647), .B(n9807), .ZN(n9783) );
  NAND2_X1 U12396 ( .A1(n13219), .A2(n9813), .ZN(n9784) );
  XNOR2_X1 U12397 ( .A(n9783), .B(n9784), .ZN(n13112) );
  NAND2_X2 U12398 ( .A1(n13113), .A2(n13112), .ZN(n13111) );
  INV_X1 U12399 ( .A(n9783), .ZN(n9785) );
  NAND2_X1 U12400 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  XNOR2_X1 U12401 ( .A(n13642), .B(n9824), .ZN(n9787) );
  NAND2_X1 U12402 ( .A1(n13218), .A2(n9813), .ZN(n9788) );
  AND2_X1 U12403 ( .A1(n9787), .A2(n9788), .ZN(n13154) );
  INV_X1 U12404 ( .A(n9787), .ZN(n9790) );
  INV_X1 U12405 ( .A(n9788), .ZN(n9789) );
  NAND2_X1 U12406 ( .A1(n9790), .A2(n9789), .ZN(n13155) );
  XNOR2_X1 U12407 ( .A(n13636), .B(n9807), .ZN(n9793) );
  NAND2_X1 U12408 ( .A1(n13217), .A2(n9813), .ZN(n9791) );
  XNOR2_X1 U12409 ( .A(n9793), .B(n9791), .ZN(n13119) );
  INV_X1 U12410 ( .A(n9791), .ZN(n9792) );
  XNOR2_X1 U12411 ( .A(n13705), .B(n9824), .ZN(n9794) );
  AND2_X1 U12412 ( .A1(n13216), .A2(n13564), .ZN(n13164) );
  NAND2_X1 U12413 ( .A1(n13165), .A2(n13164), .ZN(n9798) );
  INV_X1 U12414 ( .A(n9794), .ZN(n9795) );
  NAND2_X1 U12415 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  XNOR2_X1 U12416 ( .A(n13408), .B(n9824), .ZN(n9799) );
  AND2_X1 U12417 ( .A1(n13215), .A2(n13564), .ZN(n13103) );
  INV_X1 U12418 ( .A(n9799), .ZN(n9800) );
  NAND2_X1 U12419 ( .A1(n9801), .A2(n9800), .ZN(n9802) );
  XNOR2_X1 U12420 ( .A(n13620), .B(n9807), .ZN(n9805) );
  NAND2_X1 U12421 ( .A1(n13214), .A2(n9813), .ZN(n9803) );
  XNOR2_X1 U12422 ( .A(n9805), .B(n9803), .ZN(n13147) );
  INV_X1 U12423 ( .A(n9803), .ZN(n9804) );
  NAND2_X1 U12424 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  XNOR2_X1 U12425 ( .A(n13696), .B(n9807), .ZN(n9810) );
  NAND2_X1 U12426 ( .A1(n13213), .A2(n9813), .ZN(n9808) );
  XNOR2_X1 U12427 ( .A(n9810), .B(n9808), .ZN(n13127) );
  INV_X1 U12428 ( .A(n9808), .ZN(n9809) );
  NAND2_X1 U12429 ( .A1(n9810), .A2(n9809), .ZN(n9811) );
  XNOR2_X1 U12430 ( .A(n13361), .B(n9824), .ZN(n9814) );
  NAND2_X1 U12431 ( .A1(n13212), .A2(n9813), .ZN(n9815) );
  NAND2_X1 U12432 ( .A1(n9814), .A2(n9815), .ZN(n9819) );
  INV_X1 U12433 ( .A(n9814), .ZN(n9817) );
  INV_X1 U12434 ( .A(n9815), .ZN(n9816) );
  NAND2_X1 U12435 ( .A1(n9817), .A2(n9816), .ZN(n9818) );
  NAND2_X1 U12436 ( .A1(n9819), .A2(n9818), .ZN(n13186) );
  XNOR2_X1 U12437 ( .A(n13689), .B(n9824), .ZN(n9820) );
  NOR2_X1 U12438 ( .A1(n13189), .A2(n13528), .ZN(n9821) );
  XNOR2_X1 U12439 ( .A(n9820), .B(n9821), .ZN(n13095) );
  INV_X1 U12440 ( .A(n9820), .ZN(n9823) );
  INV_X1 U12441 ( .A(n9821), .ZN(n9822) );
  OR2_X1 U12442 ( .A1(n13096), .A2(n13528), .ZN(n9825) );
  XNOR2_X1 U12443 ( .A(n9825), .B(n9824), .ZN(n9826) );
  XNOR2_X1 U12444 ( .A(n9827), .B(n9826), .ZN(n9834) );
  NAND2_X1 U12445 ( .A1(n10980), .A2(n10978), .ZN(n9828) );
  OR2_X1 U12446 ( .A1(n9828), .A2(n14890), .ZN(n9841) );
  OR2_X1 U12447 ( .A1(n9841), .A2(n14893), .ZN(n9836) );
  INV_X1 U12448 ( .A(n9938), .ZN(n9829) );
  NAND2_X1 U12449 ( .A1(n14902), .A2(n9829), .ZN(n9830) );
  NAND2_X1 U12450 ( .A1(n11744), .A2(n9831), .ZN(n10985) );
  OR2_X1 U12451 ( .A1(n9837), .A2(n13188), .ZN(n9839) );
  OR2_X1 U12452 ( .A1(n13189), .A2(n13190), .ZN(n9838) );
  NAND2_X1 U12453 ( .A1(n9839), .A2(n9838), .ZN(n13324) );
  AOI22_X1 U12454 ( .A1(n14635), .A2(n13324), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9848) );
  NAND2_X1 U12455 ( .A1(n9841), .A2(n9840), .ZN(n9844) );
  AND2_X1 U12456 ( .A1(n9842), .A2(n10977), .ZN(n9843) );
  NAND2_X1 U12457 ( .A1(n9844), .A2(n9843), .ZN(n10164) );
  NAND2_X1 U12458 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  INV_X1 U12459 ( .A(n9939), .ZN(n9849) );
  OR2_X2 U12460 ( .A1(n10080), .A2(n10297), .ZN(n13959) );
  INV_X2 U12461 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U12462 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9857) );
  INV_X1 U12463 ( .A(n9852), .ZN(n9856) );
  OR2_X1 U12464 ( .A1(n10296), .A2(P1_U3086), .ZN(n11982) );
  NAND2_X1 U12465 ( .A1(n10291), .A2(n11982), .ZN(n9862) );
  NAND2_X1 U12466 ( .A1(n11928), .A2(n10296), .ZN(n9854) );
  NAND2_X1 U12467 ( .A1(n9854), .A2(n9853), .ZN(n9861) );
  INV_X1 U12468 ( .A(n9861), .ZN(n9855) );
  AND2_X1 U12469 ( .A1(n9862), .A2(n9855), .ZN(n10051) );
  AOI211_X1 U12470 ( .C1(n9857), .C2(n9856), .A(n10189), .B(n14715), .ZN(n9867) );
  NAND2_X1 U12471 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10476) );
  NOR2_X1 U12472 ( .A1(n9859), .A2(n10476), .ZN(n10200) );
  INV_X1 U12473 ( .A(n10051), .ZN(n9860) );
  AOI211_X1 U12474 ( .C1(n9859), .C2(n10476), .A(n10200), .B(n14719), .ZN(
        n9866) );
  NOR2_X1 U12475 ( .A1(n14757), .A2(n9870), .ZN(n9865) );
  INV_X1 U12476 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9863) );
  OAI22_X1 U12477 ( .A1(n14761), .A2(n9863), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8320), .ZN(n9864) );
  OR4_X1 U12478 ( .A1(n9867), .A2(n9866), .A3(n9865), .A4(n9864), .ZN(P1_U3244) );
  AND2_X1 U12479 ( .A1(n6568), .A2(P1_U3086), .ZN(n14375) );
  INV_X2 U12480 ( .A(n14375), .ZN(n14384) );
  AND2_X1 U12481 ( .A1(n9902), .A2(P1_U3086), .ZN(n11633) );
  INV_X2 U12482 ( .A(n11633), .ZN(n14390) );
  OAI222_X1 U12483 ( .A1(n14384), .A2(n9869), .B1(n14390), .B2(n6656), .C1(
        n6548), .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U12484 ( .A1(n14384), .A2(n9871), .B1(n14390), .B2(n9916), .C1(
        P1_U3086), .C2(n9870), .ZN(P1_U3354) );
  NOR2_X1 U12485 ( .A1(n6568), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13084) );
  INV_X1 U12486 ( .A(n13084), .ZN(n13089) );
  OAI222_X1 U12487 ( .A1(n13089), .A2(n9873), .B1(n13092), .B2(n9872), .C1(
        P3_U3151), .C2(n14995), .ZN(P3_U3287) );
  OAI222_X1 U12488 ( .A1(n13089), .A2(n9875), .B1(n13092), .B2(n9874), .C1(
        P3_U3151), .C2(n10568), .ZN(P3_U3294) );
  INV_X1 U12489 ( .A(SI_9_), .ZN(n9878) );
  INV_X1 U12490 ( .A(n9876), .ZN(n9877) );
  OAI222_X1 U12491 ( .A1(P3_U3151), .A2(n6776), .B1(n13092), .B2(n9878), .C1(
        n13089), .C2(n9877), .ZN(P3_U3286) );
  OAI222_X1 U12492 ( .A1(n14384), .A2(n15396), .B1(n14390), .B2(n9905), .C1(
        n10204), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U12493 ( .A1(P3_U3151), .A2(n14962), .B1(n13089), .B2(n9880), .C1(
        n9879), .C2(n13092), .ZN(P3_U3289) );
  INV_X1 U12494 ( .A(n9881), .ZN(n9882) );
  OAI222_X1 U12495 ( .A1(P3_U3151), .A2(n11396), .B1(n13092), .B2(n15445), 
        .C1(n13089), .C2(n9882), .ZN(P3_U3285) );
  INV_X1 U12496 ( .A(n13092), .ZN(n9891) );
  AOI222_X1 U12497 ( .A1(n9883), .A2(n13084), .B1(SI_5_), .B2(n9891), .C1(
        n10383), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9884) );
  INV_X1 U12498 ( .A(n9884), .ZN(P3_U3290) );
  AOI222_X1 U12499 ( .A1(n9885), .A2(n13084), .B1(n10519), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n9891), .C2(SI_3_), .ZN(n9886) );
  INV_X1 U12500 ( .A(n9886), .ZN(P3_U3292) );
  AOI222_X1 U12501 ( .A1(n10548), .A2(P3_STATE_REG_SCAN_IN), .B1(n9887), .B2(
        n13084), .C1(n9891), .C2(SI_2_), .ZN(n9888) );
  INV_X1 U12502 ( .A(n9888), .ZN(P3_U3293) );
  AOI222_X1 U12503 ( .A1(n9889), .A2(n13084), .B1(n10373), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n9891), .ZN(n9890) );
  INV_X1 U12504 ( .A(n9890), .ZN(P3_U3291) );
  AOI222_X1 U12505 ( .A1(n9892), .A2(n13084), .B1(SI_7_), .B2(n9891), .C1(
        n14982), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9893) );
  INV_X1 U12506 ( .A(n9893), .ZN(P3_U3288) );
  INV_X1 U12507 ( .A(n9894), .ZN(n9912) );
  OAI222_X1 U12508 ( .A1(n14384), .A2(n9895), .B1(n14390), .B2(n9912), .C1(
        n10488), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12509 ( .A(n9896), .ZN(n9897) );
  OAI222_X1 U12510 ( .A1(P3_U3151), .A2(n11389), .B1(n13092), .B2(n9898), .C1(
        n13089), .C2(n9897), .ZN(P3_U3284) );
  INV_X1 U12511 ( .A(n9899), .ZN(n9908) );
  INV_X1 U12512 ( .A(n10246), .ZN(n9900) );
  OAI222_X1 U12513 ( .A1(n14384), .A2(n9901), .B1(n14390), .B2(n9908), .C1(
        n9900), .C2(P1_U3086), .ZN(P1_U3350) );
  AND2_X1 U12514 ( .A1(n6568), .A2(P2_U3088), .ZN(n13727) );
  INV_X1 U12515 ( .A(n10120), .ZN(n9904) );
  OAI222_X1 U12516 ( .A1(n13736), .A2(n9906), .B1(n11298), .B2(n9905), .C1(
        P2_U3088), .C2(n9904), .ZN(P2_U3324) );
  INV_X1 U12517 ( .A(n9986), .ZN(n9907) );
  OAI222_X1 U12518 ( .A1(n13736), .A2(n9909), .B1(n11298), .B2(n9908), .C1(
        P2_U3088), .C2(n9907), .ZN(P2_U3322) );
  INV_X2 U12519 ( .A(n13727), .ZN(n11298) );
  OAI222_X1 U12520 ( .A1(n13736), .A2(n9910), .B1(n11298), .B2(n6656), .C1(
        P2_U3088), .C2(n9962), .ZN(P2_U3325) );
  INV_X1 U12521 ( .A(n10001), .ZN(n9911) );
  OAI222_X1 U12522 ( .A1(n13736), .A2(n9913), .B1(n11298), .B2(n9912), .C1(
        P2_U3088), .C2(n9911), .ZN(P2_U3323) );
  OAI222_X1 U12523 ( .A1(n13092), .A2(n9915), .B1(n13089), .B2(n9914), .C1(
        n12619), .C2(P3_U3151), .ZN(P3_U3283) );
  OAI222_X1 U12524 ( .A1(P2_U3088), .A2(n10036), .B1(n13736), .B2(n9917), .C1(
        n11298), .C2(n9916), .ZN(P2_U3326) );
  INV_X1 U12525 ( .A(n10421), .ZN(n9920) );
  INV_X1 U12526 ( .A(n9918), .ZN(n9921) );
  OAI222_X1 U12527 ( .A1(n9920), .A2(P1_U3086), .B1(n14390), .B2(n9921), .C1(
        n9919), .C2(n14384), .ZN(P1_U3349) );
  OAI222_X1 U12528 ( .A1(n13736), .A2(n9922), .B1(n11298), .B2(n9921), .C1(
        P2_U3088), .C2(n9989), .ZN(P2_U3321) );
  INV_X1 U12529 ( .A(n9923), .ZN(n9927) );
  INV_X1 U12530 ( .A(n13240), .ZN(n9924) );
  OAI222_X1 U12531 ( .A1(n13736), .A2(n9925), .B1(n11298), .B2(n9927), .C1(
        P2_U3088), .C2(n9924), .ZN(P2_U3320) );
  INV_X1 U12532 ( .A(n10433), .ZN(n9928) );
  OAI222_X1 U12533 ( .A1(n9928), .A2(P1_U3086), .B1(n14390), .B2(n9927), .C1(
        n9926), .C2(n14384), .ZN(P1_U3348) );
  INV_X1 U12534 ( .A(n10315), .ZN(n9929) );
  OAI222_X1 U12535 ( .A1(P1_U3086), .A2(n9929), .B1(n14390), .B2(n9931), .C1(
        n15351), .C2(n14384), .ZN(P1_U3347) );
  INV_X1 U12536 ( .A(n13258), .ZN(n9930) );
  OAI222_X1 U12537 ( .A1(n13736), .A2(n9932), .B1(n11298), .B2(n9931), .C1(
        n9930), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U12538 ( .A(n12620), .ZN(n15006) );
  INV_X1 U12539 ( .A(SI_13_), .ZN(n9934) );
  OAI222_X1 U12540 ( .A1(P3_U3151), .A2(n15006), .B1(n13092), .B2(n9934), .C1(
        n13089), .C2(n9933), .ZN(P3_U3282) );
  INV_X1 U12541 ( .A(n10067), .ZN(n10105) );
  OAI222_X1 U12542 ( .A1(n13736), .A2(n9935), .B1(n11298), .B2(n9937), .C1(
        n10105), .C2(P2_U3088), .ZN(P2_U3318) );
  OAI222_X1 U12543 ( .A1(P1_U3086), .A2(n10308), .B1(n14390), .B2(n9937), .C1(
        n9936), .C2(n14384), .ZN(P1_U3346) );
  INV_X1 U12544 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U12545 ( .A1(n9939), .A2(n9938), .ZN(n9941) );
  NAND2_X1 U12546 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NAND2_X1 U12547 ( .A1(n9943), .A2(n9942), .ZN(n9961) );
  NOR2_X2 U12548 ( .A1(n9961), .A2(P2_U3088), .ZN(n14855) );
  AND2_X1 U12549 ( .A1(n9945), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9944) );
  NAND2_X1 U12550 ( .A1(n9961), .A2(n9944), .ZN(n14862) );
  NAND2_X1 U12551 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10444) );
  INV_X1 U12552 ( .A(n10444), .ZN(n9959) );
  OR2_X1 U12553 ( .A1(n9945), .A2(P2_U3088), .ZN(n13729) );
  NOR2_X1 U12554 ( .A1(n13729), .A2(n9946), .ZN(n9947) );
  NAND2_X1 U12555 ( .A1(n9961), .A2(n9947), .ZN(n14850) );
  XNOR2_X1 U12556 ( .A(n9986), .B(n9948), .ZN(n9956) );
  INV_X1 U12557 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9949) );
  XNOR2_X1 U12558 ( .A(n10120), .B(n9949), .ZN(n10116) );
  XNOR2_X1 U12559 ( .A(n10036), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n10044) );
  AND2_X1 U12560 ( .A1(n6810), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U12561 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U12562 ( .A1(n6946), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12563 ( .A1(n10042), .A2(n9950), .ZN(n14805) );
  XNOR2_X1 U12564 ( .A(n9962), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14806) );
  NAND2_X1 U12565 ( .A1(n14805), .A2(n14806), .ZN(n14804) );
  INV_X1 U12566 ( .A(n9962), .ZN(n14807) );
  NAND2_X1 U12567 ( .A1(n14807), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U12568 ( .A1(n14804), .A2(n9951), .ZN(n10115) );
  NAND2_X1 U12569 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  NAND2_X1 U12570 ( .A1(n10120), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12571 ( .A1(n10114), .A2(n9952), .ZN(n9997) );
  INV_X1 U12572 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9953) );
  XNOR2_X1 U12573 ( .A(n10001), .B(n9953), .ZN(n9998) );
  NAND2_X1 U12574 ( .A1(n9997), .A2(n9998), .ZN(n9996) );
  NAND2_X1 U12575 ( .A1(n10001), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9954) );
  NAND2_X1 U12576 ( .A1(n9996), .A2(n9954), .ZN(n9955) );
  NAND2_X1 U12577 ( .A1(n9955), .A2(n9956), .ZN(n9981) );
  OAI21_X1 U12578 ( .B1(n9956), .B2(n9955), .A(n9981), .ZN(n9957) );
  NOR2_X1 U12579 ( .A1(n14850), .A2(n9957), .ZN(n9958) );
  AOI211_X1 U12580 ( .C1(n14838), .C2(n9986), .A(n9959), .B(n9958), .ZN(n9978)
         );
  NOR2_X1 U12581 ( .A1(n13729), .A2(n13733), .ZN(n9960) );
  AND2_X1 U12582 ( .A1(n9961), .A2(n9960), .ZN(n14857) );
  MUX2_X1 U12583 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11083), .S(n10120), .Z(
        n9968) );
  INV_X1 U12584 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11075) );
  MUX2_X1 U12585 ( .A(n11075), .B(P2_REG2_REG_2__SCAN_IN), .S(n9962), .Z(
        n14814) );
  MUX2_X1 U12586 ( .A(n9963), .B(P2_REG2_REG_1__SCAN_IN), .S(n10036), .Z(n9965) );
  AND2_X1 U12587 ( .A1(n6810), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12588 ( .A1(n9965), .A2(n9964), .ZN(n10039) );
  NAND2_X1 U12589 ( .A1(n6946), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12590 ( .A1(n10039), .A2(n9966), .ZN(n14815) );
  NAND2_X1 U12591 ( .A1(n14814), .A2(n14815), .ZN(n14813) );
  NAND2_X1 U12592 ( .A1(n14807), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12593 ( .A1(n14813), .A2(n10121), .ZN(n9967) );
  NAND2_X1 U12594 ( .A1(n9968), .A2(n9967), .ZN(n10124) );
  NAND2_X1 U12595 ( .A1(n10120), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U12596 ( .A1(n10124), .A2(n10003), .ZN(n9970) );
  MUX2_X1 U12597 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11066), .S(n10001), .Z(
        n9969) );
  NAND2_X1 U12598 ( .A1(n9970), .A2(n9969), .ZN(n10005) );
  NAND2_X1 U12599 ( .A1(n10001), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U12600 ( .A1(n10005), .A2(n9974), .ZN(n9973) );
  MUX2_X1 U12601 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9971), .S(n9986), .Z(n9972)
         );
  NAND2_X1 U12602 ( .A1(n9973), .A2(n9972), .ZN(n9992) );
  MUX2_X1 U12603 ( .A(n9971), .B(P2_REG2_REG_5__SCAN_IN), .S(n9986), .Z(n9975)
         );
  NAND3_X1 U12604 ( .A1(n10005), .A2(n9975), .A3(n9974), .ZN(n9976) );
  NAND3_X1 U12605 ( .A1(n14857), .A2(n9992), .A3(n9976), .ZN(n9977) );
  OAI211_X1 U12606 ( .C1(n9979), .C2(n14848), .A(n9978), .B(n9977), .ZN(
        P2_U3219) );
  AND2_X1 U12607 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10575) );
  MUX2_X1 U12608 ( .A(n7749), .B(P2_REG1_REG_6__SCAN_IN), .S(n9989), .Z(n9983)
         );
  NAND2_X1 U12609 ( .A1(n9986), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U12610 ( .A1(n9981), .A2(n9980), .ZN(n9982) );
  NAND2_X1 U12611 ( .A1(n9982), .A2(n9983), .ZN(n10055) );
  OAI21_X1 U12612 ( .B1(n9983), .B2(n9982), .A(n10055), .ZN(n9984) );
  NOR2_X1 U12613 ( .A1(n14850), .A2(n9984), .ZN(n9985) );
  AOI211_X1 U12614 ( .C1(n14838), .C2(n10061), .A(n10575), .B(n9985), .ZN(
        n9995) );
  NAND2_X1 U12615 ( .A1(n9986), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U12616 ( .A1(n9992), .A2(n9990), .ZN(n9988) );
  MUX2_X1 U12617 ( .A(n11123), .B(P2_REG2_REG_6__SCAN_IN), .S(n9989), .Z(n9987) );
  NAND2_X1 U12618 ( .A1(n9988), .A2(n9987), .ZN(n13243) );
  MUX2_X1 U12619 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11123), .S(n9989), .Z(n9991) );
  NAND3_X1 U12620 ( .A1(n9992), .A2(n9991), .A3(n9990), .ZN(n9993) );
  NAND3_X1 U12621 ( .A1(n14857), .A2(n13243), .A3(n9993), .ZN(n9994) );
  OAI211_X1 U12622 ( .C1(n7276), .C2(n14848), .A(n9995), .B(n9994), .ZN(
        P2_U3220) );
  AND2_X1 U12623 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10262) );
  OAI21_X1 U12624 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n9999) );
  NOR2_X1 U12625 ( .A1(n14850), .A2(n9999), .ZN(n10000) );
  AOI211_X1 U12626 ( .C1(n14838), .C2(n10001), .A(n10262), .B(n10000), .ZN(
        n10007) );
  MUX2_X1 U12627 ( .A(n11066), .B(P2_REG2_REG_4__SCAN_IN), .S(n10001), .Z(
        n10002) );
  NAND3_X1 U12628 ( .A1(n10124), .A2(n10003), .A3(n10002), .ZN(n10004) );
  NAND3_X1 U12629 ( .A1(n14857), .A2(n10005), .A3(n10004), .ZN(n10006) );
  OAI211_X1 U12630 ( .C1(n6791), .C2(n14848), .A(n10007), .B(n10006), .ZN(
        P2_U3218) );
  INV_X1 U12631 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15378) );
  NOR2_X1 U12632 ( .A1(n10034), .A2(n15378), .ZN(P3_U3251) );
  INV_X1 U12633 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U12634 ( .A1(n10034), .A2(n10009), .ZN(P3_U3263) );
  INV_X1 U12635 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n15452) );
  NOR2_X1 U12636 ( .A1(n10034), .A2(n15452), .ZN(P3_U3258) );
  INV_X1 U12637 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10010) );
  NOR2_X1 U12638 ( .A1(n10034), .A2(n10010), .ZN(P3_U3262) );
  INV_X1 U12639 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U12640 ( .A1(n10034), .A2(n10011), .ZN(P3_U3256) );
  INV_X1 U12641 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10012) );
  NOR2_X1 U12642 ( .A1(n10034), .A2(n10012), .ZN(P3_U3253) );
  INV_X1 U12643 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U12644 ( .A1(n10034), .A2(n10013), .ZN(P3_U3252) );
  INV_X1 U12645 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U12646 ( .A1(n10034), .A2(n10014), .ZN(P3_U3244) );
  INV_X1 U12647 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U12648 ( .A1(n10034), .A2(n10015), .ZN(P3_U3247) );
  INV_X1 U12649 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15232) );
  NOR2_X1 U12650 ( .A1(n10034), .A2(n15232), .ZN(P3_U3254) );
  INV_X1 U12651 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U12652 ( .A1(n10034), .A2(n10016), .ZN(P3_U3259) );
  INV_X1 U12653 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U12654 ( .A1(n10034), .A2(n10017), .ZN(P3_U3241) );
  INV_X1 U12655 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U12656 ( .A1(n10034), .A2(n10018), .ZN(P3_U3257) );
  INV_X1 U12657 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U12658 ( .A1(n10034), .A2(n10019), .ZN(P3_U3240) );
  INV_X1 U12659 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U12660 ( .A1(n10034), .A2(n15246), .ZN(P3_U3255) );
  INV_X1 U12661 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10020) );
  NOR2_X1 U12662 ( .A1(n10034), .A2(n10020), .ZN(P3_U3250) );
  INV_X1 U12663 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10021) );
  NOR2_X1 U12664 ( .A1(n10034), .A2(n10021), .ZN(P3_U3249) );
  INV_X1 U12665 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U12666 ( .A1(n10034), .A2(n10022), .ZN(P3_U3248) );
  INV_X1 U12667 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10023) );
  NOR2_X1 U12668 ( .A1(n10034), .A2(n10023), .ZN(P3_U3238) );
  INV_X1 U12669 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U12670 ( .A1(n10034), .A2(n10024), .ZN(P3_U3246) );
  INV_X1 U12671 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10025) );
  NOR2_X1 U12672 ( .A1(n10034), .A2(n10025), .ZN(P3_U3245) );
  INV_X1 U12673 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U12674 ( .A1(n10034), .A2(n10026), .ZN(P3_U3235) );
  INV_X1 U12675 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U12676 ( .A1(n10034), .A2(n10027), .ZN(P3_U3236) );
  INV_X1 U12677 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U12678 ( .A1(n10034), .A2(n10028), .ZN(P3_U3243) );
  INV_X1 U12679 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U12680 ( .A1(n10034), .A2(n10029), .ZN(P3_U3260) );
  INV_X1 U12681 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U12682 ( .A1(n10034), .A2(n10030), .ZN(P3_U3234) );
  INV_X1 U12683 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U12684 ( .A1(n10034), .A2(n10031), .ZN(P3_U3237) );
  INV_X1 U12685 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U12686 ( .A1(n10034), .A2(n10032), .ZN(P3_U3242) );
  INV_X1 U12687 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10033) );
  NOR2_X1 U12688 ( .A1(n10034), .A2(n10033), .ZN(P3_U3239) );
  INV_X1 U12689 ( .A(SI_14_), .ZN(n15394) );
  OAI222_X1 U12690 ( .A1(P3_U3151), .A2(n12634), .B1(n13092), .B2(n15394), 
        .C1(n13089), .C2(n10035), .ZN(P3_U3281) );
  MUX2_X1 U12691 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9963), .S(n10036), .Z(
        n10037) );
  OAI21_X1 U12692 ( .B1(n11737), .B2(n7656), .A(n10037), .ZN(n10038) );
  NAND3_X1 U12693 ( .A1(n14857), .A2(n10039), .A3(n10038), .ZN(n10040) );
  OAI21_X1 U12694 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n11007), .A(n10040), .ZN(
        n10041) );
  AOI21_X1 U12695 ( .B1(n6946), .B2(n14838), .A(n10041), .ZN(n10046) );
  OAI211_X1 U12696 ( .C1(n10044), .C2(n10043), .A(n14833), .B(n10042), .ZN(
        n10045) );
  OAI211_X1 U12697 ( .C1(n6742), .C2(n14848), .A(n10046), .B(n10045), .ZN(
        P2_U3215) );
  INV_X1 U12698 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10053) );
  INV_X1 U12699 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10048) );
  OAI21_X1 U12700 ( .B1(n6705), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10047), .ZN(
        n10479) );
  AOI21_X1 U12701 ( .B1(n6705), .B2(n10048), .A(n10479), .ZN(n10049) );
  INV_X1 U12702 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10480) );
  XNOR2_X1 U12703 ( .A(n10049), .B(n10480), .ZN(n10050) );
  AOI22_X1 U12704 ( .A1(n10051), .A2(n10050), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10052) );
  OAI21_X1 U12705 ( .B1(n14761), .B2(n10053), .A(n10052), .ZN(P1_U3243) );
  MUX2_X1 U12706 ( .A(n10104), .B(P2_REG1_REG_9__SCAN_IN), .S(n10067), .Z(
        n10060) );
  NAND2_X1 U12707 ( .A1(n10061), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10054) );
  NAND2_X1 U12708 ( .A1(n10055), .A2(n10054), .ZN(n13238) );
  MUX2_X1 U12709 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7770), .S(n13240), .Z(
        n13239) );
  NAND2_X1 U12710 ( .A1(n13238), .A2(n13239), .ZN(n13237) );
  NAND2_X1 U12711 ( .A1(n13240), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U12712 ( .A1(n13237), .A2(n10056), .ZN(n13251) );
  INV_X1 U12713 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10918) );
  MUX2_X1 U12714 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10918), .S(n13258), .Z(
        n13252) );
  NAND2_X1 U12715 ( .A1(n13251), .A2(n13252), .ZN(n13250) );
  NAND2_X1 U12716 ( .A1(n13258), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10057) );
  NAND2_X1 U12717 ( .A1(n13250), .A2(n10057), .ZN(n10059) );
  OR2_X1 U12718 ( .A1(n10059), .A2(n10060), .ZN(n10107) );
  INV_X1 U12719 ( .A(n10107), .ZN(n10058) );
  AOI21_X1 U12720 ( .B1(n10060), .B2(n10059), .A(n10058), .ZN(n10077) );
  NAND2_X1 U12721 ( .A1(n10061), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13242) );
  NAND2_X1 U12722 ( .A1(n13243), .A2(n13242), .ZN(n10063) );
  MUX2_X1 U12723 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11136), .S(n13240), .Z(
        n10062) );
  NAND2_X1 U12724 ( .A1(n10063), .A2(n10062), .ZN(n13255) );
  NAND2_X1 U12725 ( .A1(n13240), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U12726 ( .A1(n13255), .A2(n13254), .ZN(n10065) );
  MUX2_X1 U12727 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11105), .S(n13258), .Z(
        n10064) );
  NAND2_X1 U12728 ( .A1(n10065), .A2(n10064), .ZN(n13257) );
  NAND2_X1 U12729 ( .A1(n13258), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U12730 ( .A1(n13257), .A2(n10066), .ZN(n10069) );
  INV_X1 U12731 ( .A(n10069), .ZN(n10071) );
  MUX2_X1 U12732 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11248), .S(n10067), .Z(
        n10070) );
  MUX2_X1 U12733 ( .A(n11248), .B(P2_REG2_REG_9__SCAN_IN), .S(n10067), .Z(
        n10068) );
  OR2_X1 U12734 ( .A1(n10069), .A2(n10068), .ZN(n10096) );
  OAI21_X1 U12735 ( .B1(n10071), .B2(n10070), .A(n10096), .ZN(n10075) );
  NOR2_X1 U12736 ( .A1(n10072), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10967) );
  AOI21_X1 U12737 ( .B1(n14855), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10967), .ZN(
        n10073) );
  OAI21_X1 U12738 ( .B1(n10105), .B2(n14862), .A(n10073), .ZN(n10074) );
  AOI21_X1 U12739 ( .B1(n14857), .B2(n10075), .A(n10074), .ZN(n10076) );
  OAI21_X1 U12740 ( .B1(n10077), .B2(n14850), .A(n10076), .ZN(P2_U3223) );
  INV_X1 U12741 ( .A(n10291), .ZN(n11979) );
  INV_X1 U12742 ( .A(n10078), .ZN(n10079) );
  INV_X1 U12743 ( .A(n10080), .ZN(n10086) );
  INV_X1 U12744 ( .A(n10081), .ZN(n10082) );
  AOI22_X1 U12745 ( .A1(n14764), .A2(n10083), .B1(n10086), .B2(n10082), .ZN(
        P1_U3445) );
  INV_X1 U12746 ( .A(n10084), .ZN(n10085) );
  AOI22_X1 U12747 ( .A1(n14764), .A2(n10087), .B1(n10086), .B2(n10085), .ZN(
        P1_U3446) );
  INV_X1 U12748 ( .A(n14761), .ZN(n10945) );
  NOR2_X1 U12749 ( .A1(n10945), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12750 ( .A(n10088), .ZN(n10092) );
  INV_X1 U12751 ( .A(n14824), .ZN(n10089) );
  OAI222_X1 U12752 ( .A1(n13736), .A2(n10090), .B1(n11298), .B2(n10092), .C1(
        P2_U3088), .C2(n10089), .ZN(P2_U3317) );
  INV_X1 U12753 ( .A(n10760), .ZN(n10093) );
  OAI222_X1 U12754 ( .A1(n10093), .A2(P1_U3086), .B1(n14390), .B2(n10092), 
        .C1(n10091), .C2(n14384), .ZN(P1_U3345) );
  INV_X1 U12755 ( .A(n12660), .ZN(n14566) );
  OAI222_X1 U12756 ( .A1(P3_U3151), .A2(n14566), .B1(n13092), .B2(n15383), 
        .C1(n13089), .C2(n10094), .ZN(P3_U3280) );
  NAND2_X1 U12757 ( .A1(n10105), .A2(n11248), .ZN(n10095) );
  NAND2_X1 U12758 ( .A1(n10096), .A2(n10095), .ZN(n14826) );
  MUX2_X1 U12759 ( .A(n11267), .B(P2_REG2_REG_10__SCAN_IN), .S(n14824), .Z(
        n14827) );
  OR2_X1 U12760 ( .A1(n14826), .A2(n14827), .ZN(n14828) );
  NAND2_X1 U12761 ( .A1(n14824), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10097) );
  AND2_X1 U12762 ( .A1(n14828), .A2(n10097), .ZN(n10099) );
  MUX2_X1 U12763 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11347), .S(n10138), .Z(
        n10098) );
  NAND2_X1 U12764 ( .A1(n10099), .A2(n10098), .ZN(n10147) );
  OAI21_X1 U12765 ( .B1(n10099), .B2(n10098), .A(n10147), .ZN(n10103) );
  INV_X1 U12766 ( .A(n10138), .ZN(n10143) );
  NOR2_X1 U12767 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15348), .ZN(n10100) );
  AOI21_X1 U12768 ( .B1(n14855), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10100), 
        .ZN(n10101) );
  OAI21_X1 U12769 ( .B1(n10143), .B2(n14862), .A(n10101), .ZN(n10102) );
  AOI21_X1 U12770 ( .B1(n10103), .B2(n14857), .A(n10102), .ZN(n10113) );
  NAND2_X1 U12771 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  NAND2_X1 U12772 ( .A1(n10107), .A2(n10106), .ZN(n14820) );
  INV_X1 U12773 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10108) );
  MUX2_X1 U12774 ( .A(n10108), .B(P2_REG1_REG_10__SCAN_IN), .S(n14824), .Z(
        n14821) );
  OR2_X1 U12775 ( .A1(n14820), .A2(n14821), .ZN(n14818) );
  NAND2_X1 U12776 ( .A1(n14824), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12777 ( .A1(n14818), .A2(n10109), .ZN(n10111) );
  INV_X1 U12778 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11500) );
  MUX2_X1 U12779 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11500), .S(n10138), .Z(
        n10110) );
  NAND2_X1 U12780 ( .A1(n10111), .A2(n10110), .ZN(n10140) );
  OAI211_X1 U12781 ( .C1(n10111), .C2(n10110), .A(n10140), .B(n14833), .ZN(
        n10112) );
  NAND2_X1 U12782 ( .A1(n10113), .A2(n10112), .ZN(P2_U3225) );
  INV_X1 U12783 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10127) );
  INV_X1 U12784 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U12785 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10327), .ZN(n10119) );
  OAI211_X1 U12786 ( .C1(n10116), .C2(n10115), .A(n14833), .B(n10114), .ZN(
        n10117) );
  INV_X1 U12787 ( .A(n10117), .ZN(n10118) );
  AOI211_X1 U12788 ( .C1(n14838), .C2(n10120), .A(n10119), .B(n10118), .ZN(
        n10126) );
  MUX2_X1 U12789 ( .A(n11083), .B(P2_REG2_REG_3__SCAN_IN), .S(n10120), .Z(
        n10122) );
  NAND3_X1 U12790 ( .A1(n10122), .A2(n14813), .A3(n10121), .ZN(n10123) );
  NAND3_X1 U12791 ( .A1(n14857), .A2(n10124), .A3(n10123), .ZN(n10125) );
  OAI211_X1 U12792 ( .C1(n10127), .C2(n14848), .A(n10126), .B(n10125), .ZN(
        P2_U3217) );
  OAI222_X1 U12793 ( .A1(P3_U3151), .A2(n12674), .B1(n13092), .B2(n15337), 
        .C1(n13089), .C2(n10128), .ZN(P3_U3279) );
  INV_X1 U12794 ( .A(n10952), .ZN(n10131) );
  INV_X1 U12795 ( .A(n10129), .ZN(n10132) );
  OAI222_X1 U12796 ( .A1(P1_U3086), .A2(n10131), .B1(n14390), .B2(n10132), 
        .C1(n10130), .C2(n14384), .ZN(P1_U3344) );
  OAI222_X1 U12797 ( .A1(n13736), .A2(n15303), .B1(n11298), .B2(n10132), .C1(
        n10143), .C2(P2_U3088), .ZN(P2_U3316) );
  INV_X1 U12798 ( .A(n12705), .ZN(n12695) );
  OAI222_X1 U12799 ( .A1(P3_U3151), .A2(n12695), .B1(n13092), .B2(n15251), 
        .C1(n13089), .C2(n10133), .ZN(P3_U3278) );
  INV_X1 U12800 ( .A(n13978), .ZN(n10947) );
  INV_X1 U12801 ( .A(n10134), .ZN(n10136) );
  OAI222_X1 U12802 ( .A1(P1_U3086), .A2(n10947), .B1(n14390), .B2(n10136), 
        .C1(n10135), .C2(n14384), .ZN(P1_U3343) );
  INV_X1 U12803 ( .A(n10144), .ZN(n10234) );
  OAI222_X1 U12804 ( .A1(n13736), .A2(n10137), .B1(n11298), .B2(n10136), .C1(
        n10234), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U12805 ( .A1(n10138), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10139) );
  AND2_X1 U12806 ( .A1(n10140), .A2(n10139), .ZN(n10142) );
  MUX2_X1 U12807 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10227), .S(n10144), .Z(
        n10141) );
  NAND2_X1 U12808 ( .A1(n10142), .A2(n10141), .ZN(n10229) );
  OAI21_X1 U12809 ( .B1(n10142), .B2(n10141), .A(n10229), .ZN(n10153) );
  NAND2_X1 U12810 ( .A1(n10143), .A2(n11347), .ZN(n10145) );
  MUX2_X1 U12811 ( .A(n13575), .B(P2_REG2_REG_12__SCAN_IN), .S(n10144), .Z(
        n10146) );
  AOI21_X1 U12812 ( .B1(n10147), .B2(n10145), .A(n10146), .ZN(n10233) );
  AND3_X1 U12813 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10148) );
  OAI21_X1 U12814 ( .B1(n10233), .B2(n10148), .A(n14857), .ZN(n10151) );
  NOR2_X1 U12815 ( .A1(n10149), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11440) );
  AOI21_X1 U12816 ( .B1(n14855), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n11440), 
        .ZN(n10150) );
  OAI211_X1 U12817 ( .C1(n14862), .C2(n10234), .A(n10151), .B(n10150), .ZN(
        n10152) );
  AOI21_X1 U12818 ( .B1(n14833), .B2(n10153), .A(n10152), .ZN(n10154) );
  INV_X1 U12819 ( .A(n10154), .ZN(P2_U3226) );
  INV_X1 U12820 ( .A(n10155), .ZN(n10159) );
  INV_X1 U12821 ( .A(n14681), .ZN(n10156) );
  OAI222_X1 U12822 ( .A1(n14384), .A2(n10157), .B1(n14390), .B2(n10159), .C1(
        P1_U3086), .C2(n10156), .ZN(P1_U3342) );
  INV_X1 U12823 ( .A(n10880), .ZN(n10889) );
  OAI222_X1 U12824 ( .A1(P2_U3088), .A2(n10889), .B1(n11298), .B2(n10159), 
        .C1(n10158), .C2(n13736), .ZN(P2_U3314) );
  INV_X1 U12825 ( .A(n10160), .ZN(n10161) );
  AOI21_X1 U12826 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(n10168) );
  OR2_X1 U12827 ( .A1(n10164), .A2(P2_U3088), .ZN(n10218) );
  AOI22_X1 U12828 ( .A1(n6562), .A2(n14638), .B1(n10218), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10167) );
  INV_X1 U12829 ( .A(n7655), .ZN(n10165) );
  OAI22_X1 U12830 ( .A1(n10165), .A2(n13190), .B1(n10277), .B2(n13188), .ZN(
        n11000) );
  NAND2_X1 U12831 ( .A1(n14635), .A2(n11000), .ZN(n10166) );
  OAI211_X1 U12832 ( .C1(n10168), .C2(n13202), .A(n10167), .B(n10166), .ZN(
        P2_U3194) );
  NAND2_X1 U12833 ( .A1(n8764), .A2(n13516), .ZN(n10467) );
  AOI22_X1 U12834 ( .A1(n11004), .A2(n14638), .B1(n10218), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10172) );
  AOI21_X1 U12835 ( .B1(n7655), .B2(n9813), .A(n11004), .ZN(n10169) );
  OAI22_X1 U12836 ( .A1(n11005), .A2(n10169), .B1(n9813), .B2(n11752), .ZN(
        n10170) );
  NAND2_X1 U12837 ( .A1(n14633), .A2(n10170), .ZN(n10171) );
  OAI211_X1 U12838 ( .C1(n10467), .C2(n13178), .A(n10172), .B(n10171), .ZN(
        P2_U3204) );
  INV_X1 U12839 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10178) );
  INV_X1 U12840 ( .A(n10300), .ZN(n10176) );
  INV_X1 U12841 ( .A(n12209), .ZN(n10175) );
  NAND2_X1 U12842 ( .A1(n8672), .A2(n10175), .ZN(n10173) );
  AND2_X1 U12843 ( .A1(n10173), .A2(n10454), .ZN(n11935) );
  OAI21_X1 U12844 ( .B1(n14793), .B2(n14522), .A(n11935), .ZN(n10174) );
  OR2_X1 U12845 ( .A1(n12212), .A2(n14210), .ZN(n10748) );
  OAI211_X1 U12846 ( .C1(n10176), .C2(n10175), .A(n10174), .B(n10748), .ZN(
        n14336) );
  NAND2_X1 U12847 ( .A1(n14336), .A2(n14796), .ZN(n10177) );
  OAI21_X1 U12848 ( .B1(n14796), .B2(n10178), .A(n10177), .ZN(P1_U3459) );
  INV_X1 U12849 ( .A(n12716), .ZN(n10180) );
  OAI222_X1 U12850 ( .A1(P3_U3151), .A2(n10180), .B1(n13092), .B2(n15448), 
        .C1(n13089), .C2(n10179), .ZN(P3_U3277) );
  XNOR2_X1 U12851 ( .A(n10181), .B(n10183), .ZN(n11078) );
  INV_X1 U12852 ( .A(n10268), .ZN(n10182) );
  AOI211_X1 U12853 ( .C1(n7671), .C2(n11002), .A(n9813), .B(n10182), .ZN(
        n11073) );
  AOI21_X1 U12854 ( .B1(n14918), .B2(n7671), .A(n11073), .ZN(n10187) );
  XNOR2_X1 U12855 ( .A(n10184), .B(n10183), .ZN(n10186) );
  OAI22_X1 U12856 ( .A1(n10185), .A2(n13190), .B1(n7221), .B2(n13188), .ZN(
        n10219) );
  AOI21_X1 U12857 ( .B1(n10186), .B2(n13540), .A(n10219), .ZN(n11074) );
  OAI211_X1 U12858 ( .C1(n14921), .C2(n11078), .A(n10187), .B(n11074), .ZN(
        n10388) );
  NAND2_X1 U12859 ( .A1(n14908), .A2(n10388), .ZN(n10188) );
  OAI21_X1 U12860 ( .B1(n14908), .B2(n7658), .A(n10188), .ZN(P2_U3436) );
  INV_X1 U12861 ( .A(n10488), .ZN(n10209) );
  INV_X1 U12862 ( .A(n10204), .ZN(n10406) );
  INV_X1 U12863 ( .A(n6548), .ZN(n10203) );
  INV_X1 U12864 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U12865 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10190), .S(n6548), .Z(
        n10496) );
  NOR2_X1 U12866 ( .A1(n10497), .A2(n10496), .ZN(n10495) );
  INV_X1 U12867 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U12868 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10191), .S(n10204), .Z(
        n10401) );
  NOR2_X1 U12869 ( .A1(n10402), .A2(n10401), .ZN(n10400) );
  INV_X1 U12870 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10192) );
  MUX2_X1 U12871 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10192), .S(n10488), .Z(
        n10482) );
  NOR2_X1 U12872 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  XOR2_X1 U12873 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10246), .Z(n10245) );
  NAND2_X1 U12874 ( .A1(n10244), .A2(n10245), .ZN(n10243) );
  INV_X1 U12875 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10193) );
  MUX2_X1 U12876 ( .A(n10193), .B(P1_REG1_REG_6__SCAN_IN), .S(n10421), .Z(
        n10420) );
  NOR2_X1 U12877 ( .A1(n10419), .A2(n10420), .ZN(n10418) );
  INV_X1 U12878 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U12879 ( .A(n10194), .B(P1_REG1_REG_7__SCAN_IN), .S(n10433), .Z(
        n10431) );
  NOR2_X1 U12880 ( .A1(n10432), .A2(n10431), .ZN(n10430) );
  INV_X1 U12881 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10195) );
  MUX2_X1 U12882 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10195), .S(n10315), .Z(
        n10196) );
  NAND2_X1 U12883 ( .A1(n10197), .A2(n10196), .ZN(n10310) );
  OAI21_X1 U12884 ( .B1(n10197), .B2(n10196), .A(n10310), .ZN(n10216) );
  INV_X1 U12885 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12886 ( .A1(n14726), .A2(n10315), .ZN(n10198) );
  NAND2_X1 U12887 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11626) );
  OAI211_X1 U12888 ( .C1(n10199), .C2(n14761), .A(n10198), .B(n11626), .ZN(
        n10215) );
  AOI21_X1 U12889 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10201), .A(n10200), .ZN(
        n10494) );
  INV_X1 U12890 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10202) );
  MUX2_X1 U12891 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10202), .S(n6548), .Z(
        n10493) );
  NOR2_X1 U12892 ( .A1(n10494), .A2(n10493), .ZN(n10492) );
  AOI21_X1 U12893 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n10203), .A(n10492), .ZN(
        n10405) );
  INV_X1 U12894 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10205) );
  MUX2_X1 U12895 ( .A(n10205), .B(P1_REG2_REG_3__SCAN_IN), .S(n10204), .Z(
        n10206) );
  INV_X1 U12896 ( .A(n10206), .ZN(n10404) );
  NOR2_X1 U12897 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  AOI21_X1 U12898 ( .B1(n10406), .B2(P1_REG2_REG_3__SCAN_IN), .A(n10403), .ZN(
        n10486) );
  INV_X1 U12899 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U12900 ( .A(n10207), .B(P1_REG2_REG_4__SCAN_IN), .S(n10488), .Z(
        n10208) );
  INV_X1 U12901 ( .A(n10208), .ZN(n10485) );
  NOR2_X1 U12902 ( .A1(n10486), .A2(n10485), .ZN(n10484) );
  XNOR2_X1 U12903 ( .A(n10246), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n10249) );
  XNOR2_X1 U12904 ( .A(n10421), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n10416) );
  AOI21_X1 U12905 ( .B1(n10421), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6618), .ZN(
        n10429) );
  XNOR2_X1 U12906 ( .A(n10433), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n10428) );
  INV_X1 U12907 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10210) );
  MUX2_X1 U12908 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10210), .S(n10315), .Z(
        n10211) );
  INV_X1 U12909 ( .A(n10211), .ZN(n10212) );
  AOI211_X1 U12910 ( .C1(n10213), .C2(n10212), .A(n14719), .B(n10314), .ZN(
        n10214) );
  AOI211_X1 U12911 ( .C1(n14753), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n10217) );
  INV_X1 U12912 ( .A(n10217), .ZN(P1_U3251) );
  AOI22_X1 U12913 ( .A1(n14635), .A2(n10219), .B1(n10218), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10225) );
  OAI21_X1 U12914 ( .B1(n10222), .B2(n10221), .A(n10220), .ZN(n10223) );
  NAND2_X1 U12915 ( .A1(n14633), .A2(n10223), .ZN(n10224) );
  OAI211_X1 U12916 ( .C1(n11071), .C2(n13183), .A(n10225), .B(n10224), .ZN(
        P2_U3209) );
  INV_X1 U12917 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U12918 ( .A(n10226), .B(P2_REG1_REG_13__SCAN_IN), .S(n10880), .Z(
        n10232) );
  NAND2_X1 U12919 ( .A1(n10234), .A2(n10227), .ZN(n10228) );
  NAND2_X1 U12920 ( .A1(n10229), .A2(n10228), .ZN(n10231) );
  INV_X1 U12921 ( .A(n10882), .ZN(n10230) );
  AOI211_X1 U12922 ( .C1(n10232), .C2(n10231), .A(n14850), .B(n10230), .ZN(
        n10242) );
  AOI21_X1 U12923 ( .B1(n13575), .B2(n10234), .A(n10233), .ZN(n10237) );
  MUX2_X1 U12924 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10235), .S(n10880), .Z(
        n10236) );
  NAND2_X1 U12925 ( .A1(n10237), .A2(n10236), .ZN(n10888) );
  OAI211_X1 U12926 ( .C1(n10237), .C2(n10236), .A(n10888), .B(n14857), .ZN(
        n10240) );
  NOR2_X1 U12927 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11563), .ZN(n10238) );
  AOI21_X1 U12928 ( .B1(n14855), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10238), 
        .ZN(n10239) );
  OAI211_X1 U12929 ( .C1(n14862), .C2(n10889), .A(n10240), .B(n10239), .ZN(
        n10241) );
  OR2_X1 U12930 ( .A1(n10242), .A2(n10241), .ZN(P2_U3227) );
  OAI21_X1 U12931 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(n10253) );
  INV_X1 U12932 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14446) );
  NAND2_X1 U12933 ( .A1(n14726), .A2(n10246), .ZN(n10247) );
  NAND2_X1 U12934 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11220) );
  OAI211_X1 U12935 ( .C1(n14446), .C2(n14761), .A(n10247), .B(n11220), .ZN(
        n10252) );
  AOI211_X1 U12936 ( .C1(n10250), .C2(n10249), .A(n14719), .B(n10248), .ZN(
        n10251) );
  AOI211_X1 U12937 ( .C1(n14753), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        n10254) );
  INV_X1 U12938 ( .A(n10254), .ZN(P1_U3248) );
  OAI222_X1 U12939 ( .A1(n13089), .A2(n10256), .B1(n13092), .B2(n10255), .C1(
        P3_U3151), .C2(n6555), .ZN(P3_U3276) );
  OAI21_X1 U12940 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10266) );
  NAND2_X1 U12941 ( .A1(n13233), .A2(n13518), .ZN(n10261) );
  NAND2_X1 U12942 ( .A1(n13231), .A2(n13516), .ZN(n10260) );
  NAND2_X1 U12943 ( .A1(n10261), .A2(n10260), .ZN(n10396) );
  AOI21_X1 U12944 ( .B1(n14635), .B2(n10396), .A(n10262), .ZN(n10264) );
  NAND2_X1 U12945 ( .A1(n14638), .A2(n10393), .ZN(n10263) );
  OAI211_X1 U12946 ( .C1(n14643), .C2(n11061), .A(n10264), .B(n10263), .ZN(
        n10265) );
  AOI21_X1 U12947 ( .B1(n14633), .B2(n10266), .A(n10265), .ZN(n10267) );
  INV_X1 U12948 ( .A(n10267), .ZN(P2_U3202) );
  NAND2_X1 U12949 ( .A1(n10268), .A2(n10273), .ZN(n10269) );
  NAND2_X1 U12950 ( .A1(n10269), .A2(n13528), .ZN(n10270) );
  NOR2_X1 U12951 ( .A1(n10391), .A2(n10270), .ZN(n11081) );
  XNOR2_X1 U12952 ( .A(n10271), .B(n10274), .ZN(n11086) );
  NOR2_X1 U12953 ( .A1(n11086), .A2(n14921), .ZN(n10272) );
  AOI211_X1 U12954 ( .C1(n14918), .C2(n10273), .A(n11081), .B(n10272), .ZN(
        n10279) );
  XNOR2_X1 U12955 ( .A(n10275), .B(n10274), .ZN(n10278) );
  OAI22_X1 U12956 ( .A1(n10277), .A2(n13190), .B1(n10276), .B2(n13188), .ZN(
        n10324) );
  AOI21_X1 U12957 ( .B1(n10278), .B2(n13540), .A(n10324), .ZN(n11082) );
  NAND2_X1 U12958 ( .A1(n10279), .A2(n11082), .ZN(n10412) );
  NAND2_X1 U12959 ( .A1(n10412), .A2(n14908), .ZN(n10280) );
  OAI21_X1 U12960 ( .B1(n14908), .B2(n7674), .A(n10280), .ZN(P2_U3439) );
  XNOR2_X1 U12961 ( .A(n10283), .B(n12364), .ZN(n10523) );
  XOR2_X1 U12962 ( .A(n10526), .B(n10523), .Z(n10288) );
  OR2_X1 U12963 ( .A1(n8672), .A2(n12345), .ZN(n10285) );
  AOI22_X1 U12964 ( .A1(n12362), .A2(n12209), .B1(n10286), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U12965 ( .A1(n10285), .A2(n10284), .ZN(n10475) );
  AOI222_X1 U12966 ( .A1(n13961), .A2(n12362), .B1(n12209), .B2(n11448), .C1(
        n10286), .C2(P1_REG1_REG_0__SCAN_IN), .ZN(n10474) );
  MUX2_X1 U12967 ( .A(n10475), .B(n12343), .S(n10474), .Z(n10287) );
  AOI21_X1 U12968 ( .B1(n10288), .B2(n10287), .A(n10524), .ZN(n10307) );
  INV_X1 U12969 ( .A(n10716), .ZN(n10290) );
  NAND3_X1 U12970 ( .A1(n10717), .A2(n10290), .A3(n10289), .ZN(n10295) );
  NOR2_X1 U12971 ( .A1(n10295), .A2(n10291), .ZN(n10294) );
  INV_X1 U12972 ( .A(n10294), .ZN(n10304) );
  INV_X1 U12973 ( .A(n11928), .ZN(n10292) );
  NAND2_X1 U12974 ( .A1(n14788), .A2(n10292), .ZN(n10293) );
  AND2_X1 U12975 ( .A1(n10294), .A2(n11978), .ZN(n13795) );
  NOR2_X1 U12976 ( .A1(n8675), .A2(n14210), .ZN(n10452) );
  NAND2_X1 U12977 ( .A1(n10295), .A2(n10301), .ZN(n10299) );
  AND3_X1 U12978 ( .A1(n11978), .A2(n10297), .A3(n10296), .ZN(n10298) );
  NAND2_X1 U12979 ( .A1(n10299), .A2(n10298), .ZN(n10665) );
  OR2_X1 U12980 ( .A1(n10665), .A2(P1_U3086), .ZN(n12208) );
  AOI22_X1 U12981 ( .A1(n13795), .A2(n10452), .B1(n12208), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12982 ( .A1(n13795), .A2(n14174), .ZN(n13904) );
  INV_X1 U12983 ( .A(n13904), .ZN(n13883) );
  AND2_X1 U12984 ( .A1(n10300), .A2(n11929), .ZN(n10720) );
  INV_X1 U12985 ( .A(n10720), .ZN(n10303) );
  INV_X1 U12986 ( .A(n10301), .ZN(n10302) );
  OAI21_X2 U12987 ( .B1(n10304), .B2(n10303), .A(n14526), .ZN(n13936) );
  AOI22_X1 U12988 ( .A1(n13883), .A2(n13961), .B1(n8662), .B2(n13936), .ZN(
        n10305) );
  OAI211_X1 U12989 ( .C1(n10307), .C2(n13938), .A(n10306), .B(n10305), .ZN(
        P1_U3222) );
  INV_X1 U12990 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U12991 ( .A(n10309), .B(P1_REG1_REG_9__SCAN_IN), .S(n10308), .Z(
        n10312) );
  OAI21_X1 U12992 ( .B1(n10312), .B2(n10311), .A(n10581), .ZN(n10320) );
  INV_X1 U12993 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14395) );
  NAND2_X1 U12994 ( .A1(n14726), .A2(n10582), .ZN(n10313) );
  NAND2_X1 U12995 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11718) );
  OAI211_X1 U12996 ( .C1(n14395), .C2(n14761), .A(n10313), .B(n11718), .ZN(
        n10319) );
  XNOR2_X1 U12997 ( .A(n10582), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U12998 ( .A1(n10317), .A2(n10316), .ZN(n10578) );
  AOI211_X1 U12999 ( .C1(n10317), .C2(n10316), .A(n14719), .B(n10578), .ZN(
        n10318) );
  AOI211_X1 U13000 ( .C1(n14753), .C2(n10320), .A(n10319), .B(n10318), .ZN(
        n10321) );
  INV_X1 U13001 ( .A(n10321), .ZN(P1_U3252) );
  XNOR2_X1 U13002 ( .A(n10323), .B(n10322), .ZN(n10329) );
  AOI22_X1 U13003 ( .A1(n14635), .A2(n10324), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10325) );
  OAI21_X1 U13004 ( .B1(n11079), .B2(n13183), .A(n10325), .ZN(n10326) );
  AOI21_X1 U13005 ( .B1(n9845), .B2(n10327), .A(n10326), .ZN(n10328) );
  OAI21_X1 U13006 ( .B1(n10329), .B2(n13202), .A(n10328), .ZN(P2_U3190) );
  MUX2_X1 U13007 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n14941), .Z(n10348) );
  INV_X1 U13008 ( .A(n10373), .ZN(n10609) );
  MUX2_X1 U13009 ( .A(n10330), .B(n10557), .S(n12718), .Z(n10332) );
  NAND2_X1 U13010 ( .A1(n10332), .A2(n10331), .ZN(n10543) );
  INV_X1 U13011 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U13012 ( .A1(n10333), .A2(n10568), .ZN(n10334) );
  NAND2_X1 U13013 ( .A1(n10543), .A2(n10334), .ZN(n10554) );
  INV_X1 U13014 ( .A(n10554), .ZN(n10336) );
  MUX2_X1 U13015 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n6550), .Z(n10335) );
  INV_X1 U13016 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n14948) );
  NOR2_X1 U13017 ( .A1(n10335), .A2(n14948), .ZN(n10553) );
  NAND2_X1 U13018 ( .A1(n10336), .A2(n10553), .ZN(n10556) );
  INV_X1 U13019 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10368) );
  MUX2_X1 U13020 ( .A(n15120), .B(n10368), .S(n6550), .Z(n10337) );
  NAND2_X1 U13021 ( .A1(n10337), .A2(n10548), .ZN(n10508) );
  INV_X1 U13022 ( .A(n10337), .ZN(n10338) );
  NAND2_X1 U13023 ( .A1(n10338), .A2(n6714), .ZN(n10339) );
  NAND2_X1 U13024 ( .A1(n10508), .A2(n10339), .ZN(n10542) );
  AOI21_X1 U13025 ( .B1(n10556), .B2(n10543), .A(n10542), .ZN(n10506) );
  INV_X1 U13026 ( .A(n10508), .ZN(n10346) );
  MUX2_X1 U13027 ( .A(n10341), .B(n10340), .S(n14941), .Z(n10342) );
  NAND2_X1 U13028 ( .A1(n10342), .A2(n10519), .ZN(n10347) );
  INV_X1 U13029 ( .A(n10342), .ZN(n10343) );
  NAND2_X1 U13030 ( .A1(n10343), .A2(n10370), .ZN(n10344) );
  NAND2_X1 U13031 ( .A1(n10347), .A2(n10344), .ZN(n10507) );
  INV_X1 U13032 ( .A(n10507), .ZN(n10345) );
  OAI21_X1 U13033 ( .B1(n10506), .B2(n10346), .A(n10345), .ZN(n10510) );
  NAND2_X1 U13034 ( .A1(n10510), .A2(n10347), .ZN(n10591) );
  XNOR2_X1 U13035 ( .A(n10348), .B(n10373), .ZN(n10590) );
  NAND2_X1 U13036 ( .A1(n10591), .A2(n10590), .ZN(n10589) );
  OAI21_X1 U13037 ( .B1(n10348), .B2(n10609), .A(n10589), .ZN(n10800) );
  MUX2_X1 U13038 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n14941), .Z(n10349) );
  NOR2_X1 U13039 ( .A1(n10349), .A2(n10814), .ZN(n10798) );
  INV_X1 U13040 ( .A(n10798), .ZN(n10350) );
  NAND2_X1 U13041 ( .A1(n10349), .A2(n10814), .ZN(n10799) );
  NAND2_X1 U13042 ( .A1(n10350), .A2(n10799), .ZN(n10351) );
  XNOR2_X1 U13043 ( .A(n10800), .B(n10351), .ZN(n10385) );
  INV_X1 U13044 ( .A(n12598), .ZN(n12612) );
  NAND2_X1 U13045 ( .A1(n12612), .A2(n9623), .ZN(n15017) );
  NAND2_X1 U13046 ( .A1(n12133), .A2(n10353), .ZN(n10352) );
  NAND2_X1 U13047 ( .A1(n9179), .A2(n10352), .ZN(n10364) );
  OR2_X1 U13048 ( .A1(n10353), .A2(P3_U3151), .ZN(n12192) );
  INV_X1 U13049 ( .A(n12192), .ZN(n10354) );
  NOR2_X1 U13050 ( .A1(n10624), .A2(n10354), .ZN(n10363) );
  MUX2_X1 U13051 ( .A(n10377), .B(n12598), .S(n12187), .Z(n15007) );
  NOR2_X1 U13052 ( .A1(n10377), .A2(n10355), .ZN(n12732) );
  XNOR2_X1 U13053 ( .A(n10548), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10533) );
  NOR2_X1 U13054 ( .A1(n14942), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U13055 ( .A1(n10356), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10358) );
  OAI21_X1 U13056 ( .B1(n10568), .B2(n10357), .A(n10358), .ZN(n10550) );
  NAND2_X1 U13057 ( .A1(n10552), .A2(n10358), .ZN(n10532) );
  NAND2_X1 U13058 ( .A1(n10533), .A2(n10532), .ZN(n10531) );
  NAND2_X1 U13059 ( .A1(n10359), .A2(n10370), .ZN(n10360) );
  INV_X1 U13060 ( .A(n10360), .ZN(n10593) );
  MUX2_X1 U13061 ( .A(n10361), .B(P3_REG2_REG_4__SCAN_IN), .S(n10373), .Z(
        n10594) );
  AOI21_X1 U13062 ( .B1(n9225), .B2(n10362), .A(n10812), .ZN(n10381) );
  INV_X1 U13063 ( .A(n10363), .ZN(n10365) );
  AND2_X1 U13064 ( .A1(n10365), .A2(n10364), .ZN(n14978) );
  NOR2_X1 U13065 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9226), .ZN(n11243) );
  AOI21_X1 U13066 ( .B1(n14978), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11243), .ZN(
        n10380) );
  INV_X1 U13067 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10366) );
  NOR2_X1 U13068 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10366), .ZN(n10367) );
  OAI21_X1 U13069 ( .B1(n10568), .B2(n10367), .A(n6591), .ZN(n10558) );
  OR2_X1 U13070 ( .A1(n10558), .A2(n10557), .ZN(n10560) );
  OR2_X1 U13071 ( .A1(n10548), .A2(n10368), .ZN(n10369) );
  NAND2_X1 U13072 ( .A1(n10601), .A2(n10599), .ZN(n10371) );
  MUX2_X1 U13073 ( .A(n10372), .B(P3_REG1_REG_4__SCAN_IN), .S(n10373), .Z(
        n10598) );
  OR2_X1 U13074 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  NOR2_X1 U13075 ( .A1(n10375), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U13076 ( .A1(n10377), .A2(n10376), .ZN(n12737) );
  OAI21_X1 U13077 ( .B1(n10793), .B2(n10378), .A(n12737), .ZN(n10379) );
  OAI211_X1 U13078 ( .C1(n15023), .C2(n10381), .A(n10380), .B(n10379), .ZN(
        n10382) );
  AOI21_X1 U13079 ( .B1(n10383), .B2(n14981), .A(n10382), .ZN(n10384) );
  OAI21_X1 U13080 ( .B1(n10385), .B2(n15017), .A(n10384), .ZN(P3_U3187) );
  INV_X1 U13081 ( .A(n14890), .ZN(n10386) );
  NAND2_X1 U13082 ( .A1(n14931), .A2(n10388), .ZN(n10389) );
  OAI21_X1 U13083 ( .B1(n14931), .B2(n7659), .A(n10389), .ZN(P2_U3501) );
  XNOR2_X1 U13084 ( .A(n10390), .B(n10394), .ZN(n11069) );
  INV_X1 U13085 ( .A(n10391), .ZN(n10392) );
  AOI211_X1 U13086 ( .C1(n10393), .C2(n10392), .A(n9813), .B(n6697), .ZN(
        n11064) );
  AOI21_X1 U13087 ( .B1(n14918), .B2(n10393), .A(n11064), .ZN(n10398) );
  XNOR2_X1 U13088 ( .A(n10395), .B(n10394), .ZN(n10397) );
  AOI21_X1 U13089 ( .B1(n10397), .B2(n13540), .A(n10396), .ZN(n11065) );
  OAI211_X1 U13090 ( .C1(n14921), .C2(n11069), .A(n10398), .B(n11065), .ZN(
        n10414) );
  NAND2_X1 U13091 ( .A1(n10414), .A2(n14908), .ZN(n10399) );
  OAI21_X1 U13092 ( .B1(n14908), .B2(n7692), .A(n10399), .ZN(P2_U3442) );
  AOI211_X1 U13093 ( .C1(n10402), .C2(n10401), .A(n10400), .B(n14715), .ZN(
        n10411) );
  AOI211_X1 U13094 ( .C1(n10405), .C2(n10404), .A(n10403), .B(n14719), .ZN(
        n10410) );
  INV_X1 U13095 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14442) );
  NAND2_X1 U13096 ( .A1(n14726), .A2(n10406), .ZN(n10408) );
  NAND2_X1 U13097 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n10407) );
  OAI211_X1 U13098 ( .C1(n14442), .C2(n14761), .A(n10408), .B(n10407), .ZN(
        n10409) );
  OR3_X1 U13099 ( .A1(n10411), .A2(n10410), .A3(n10409), .ZN(P1_U3246) );
  NAND2_X1 U13100 ( .A1(n10412), .A2(n14931), .ZN(n10413) );
  OAI21_X1 U13101 ( .B1(n14931), .B2(n9949), .A(n10413), .ZN(P2_U3502) );
  NAND2_X1 U13102 ( .A1(n10414), .A2(n14931), .ZN(n10415) );
  OAI21_X1 U13103 ( .B1(n14931), .B2(n9953), .A(n10415), .ZN(P2_U3503) );
  AOI211_X1 U13104 ( .C1(n10417), .C2(n10416), .A(n14719), .B(n6618), .ZN(
        n10426) );
  AOI211_X1 U13105 ( .C1(n10420), .C2(n10419), .A(n14715), .B(n10418), .ZN(
        n10425) );
  NAND2_X1 U13106 ( .A1(n14726), .A2(n10421), .ZN(n10423) );
  NAND2_X1 U13107 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10422) );
  OAI211_X1 U13108 ( .C1(n15395), .C2(n14761), .A(n10423), .B(n10422), .ZN(
        n10424) );
  OR3_X1 U13109 ( .A1(n10426), .A2(n10425), .A3(n10424), .ZN(P1_U3249) );
  AOI211_X1 U13110 ( .C1(n10429), .C2(n10428), .A(n14719), .B(n10427), .ZN(
        n10437) );
  AOI211_X1 U13111 ( .C1(n10432), .C2(n10431), .A(n14715), .B(n10430), .ZN(
        n10436) );
  INV_X1 U13112 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14457) );
  NAND2_X1 U13113 ( .A1(n14726), .A2(n10433), .ZN(n10434) );
  NAND2_X1 U13114 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11454) );
  OAI211_X1 U13115 ( .C1(n14457), .C2(n14761), .A(n10434), .B(n11454), .ZN(
        n10435) );
  OR3_X1 U13116 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(P1_U3250) );
  OAI21_X1 U13117 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n10441) );
  NAND2_X1 U13118 ( .A1(n10441), .A2(n14633), .ZN(n10447) );
  NAND2_X1 U13119 ( .A1(n13232), .A2(n13518), .ZN(n10443) );
  NAND2_X1 U13120 ( .A1(n13230), .A2(n13516), .ZN(n10442) );
  AND2_X1 U13121 ( .A1(n10443), .A2(n10442), .ZN(n10994) );
  OAI21_X1 U13122 ( .B1(n13178), .B2(n10994), .A(n10444), .ZN(n10445) );
  AOI21_X1 U13123 ( .B1(n10989), .B2(n14638), .A(n10445), .ZN(n10446) );
  OAI211_X1 U13124 ( .C1(n14643), .C2(n10987), .A(n10447), .B(n10446), .ZN(
        P2_U3199) );
  NAND2_X1 U13125 ( .A1(n8662), .A2(n12209), .ZN(n10448) );
  NAND2_X1 U13126 ( .A1(n10723), .A2(n10448), .ZN(n11019) );
  OAI21_X1 U13127 ( .B1(n11759), .B2(n8672), .A(n14522), .ZN(n10451) );
  XNOR2_X1 U13128 ( .A(n13960), .B(n11019), .ZN(n10449) );
  AOI21_X1 U13129 ( .B1(n10449), .B2(n14522), .A(n13961), .ZN(n10450) );
  AOI21_X1 U13130 ( .B1(n14212), .B2(n10451), .A(n10450), .ZN(n10453) );
  NOR2_X1 U13131 ( .A1(n10453), .A2(n10452), .ZN(n11027) );
  XNOR2_X1 U13132 ( .A(n11759), .B(n10454), .ZN(n11025) );
  NAND2_X1 U13133 ( .A1(n11025), .A2(n14793), .ZN(n10455) );
  OAI211_X1 U13134 ( .C1(n11019), .C2(n14252), .A(n11027), .B(n10455), .ZN(
        n10458) );
  NAND2_X1 U13135 ( .A1(n10458), .A2(n14803), .ZN(n10457) );
  NAND2_X1 U13136 ( .A1(n14235), .A2(n8662), .ZN(n10456) );
  OAI211_X1 U13137 ( .C1(n14803), .C2(n6826), .A(n10457), .B(n10456), .ZN(
        P1_U3529) );
  INV_X1 U13138 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U13139 ( .A1(n10458), .A2(n14796), .ZN(n10460) );
  NAND2_X1 U13140 ( .A1(n11173), .A2(n8662), .ZN(n10459) );
  OAI211_X1 U13141 ( .C1(n14796), .C2(n10461), .A(n10460), .B(n10459), .ZN(
        P1_U3462) );
  INV_X1 U13142 ( .A(n13980), .ZN(n14695) );
  INV_X1 U13143 ( .A(n10462), .ZN(n10464) );
  OAI222_X1 U13144 ( .A1(P1_U3086), .A2(n14695), .B1(n14390), .B2(n10464), 
        .C1(n10463), .C2(n14384), .ZN(P1_U3341) );
  INV_X1 U13145 ( .A(n14837), .ZN(n10890) );
  OAI222_X1 U13146 ( .A1(n13736), .A2(n10465), .B1(n11298), .B2(n10464), .C1(
        n10890), .C2(P2_U3088), .ZN(P2_U3313) );
  NOR2_X1 U13147 ( .A1(n11745), .A2(n8756), .ZN(n10469) );
  AND2_X1 U13148 ( .A1(n13562), .A2(n6794), .ZN(n10466) );
  OR2_X1 U13149 ( .A1(n11745), .A2(n10466), .ZN(n10468) );
  NAND2_X1 U13150 ( .A1(n10468), .A2(n10467), .ZN(n11746) );
  AOI211_X1 U13151 ( .C1(n11004), .C2(n11744), .A(n10469), .B(n11746), .ZN(
        n10473) );
  NAND2_X1 U13152 ( .A1(n14929), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10470) );
  OAI21_X1 U13153 ( .B1(n14929), .B2(n10473), .A(n10470), .ZN(P2_U3499) );
  INV_X1 U13154 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10471) );
  OR2_X1 U13155 ( .A1(n14908), .A2(n10471), .ZN(n10472) );
  OAI21_X1 U13156 ( .B1(n14924), .B2(n10473), .A(n10472), .ZN(P2_U3430) );
  XNOR2_X1 U13157 ( .A(n10474), .B(n10475), .ZN(n12207) );
  MUX2_X1 U13158 ( .A(n10476), .B(n12207), .S(n6705), .Z(n10477) );
  AOI211_X1 U13159 ( .C1(n10480), .C2(n10479), .A(n13959), .B(n10478), .ZN(
        n10503) );
  AOI211_X1 U13160 ( .C1(n10483), .C2(n10482), .A(n10481), .B(n14715), .ZN(
        n10491) );
  AOI211_X1 U13161 ( .C1(n10486), .C2(n10485), .A(n10484), .B(n14719), .ZN(
        n10490) );
  NAND2_X1 U13162 ( .A1(n10945), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U13163 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n11230) );
  OAI211_X1 U13164 ( .C1(n14757), .C2(n10488), .A(n10487), .B(n11230), .ZN(
        n10489) );
  OR4_X1 U13165 ( .A1(n10503), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        P1_U3247) );
  AOI211_X1 U13166 ( .C1(n10494), .C2(n10493), .A(n10492), .B(n14719), .ZN(
        n10502) );
  AOI211_X1 U13167 ( .C1(n10497), .C2(n10496), .A(n10495), .B(n14715), .ZN(
        n10501) );
  AOI22_X1 U13168 ( .A1(n10945), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10498) );
  OAI21_X1 U13169 ( .B1(n6548), .B2(n14757), .A(n10498), .ZN(n10500) );
  OR4_X1 U13170 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        P1_U3245) );
  OAI222_X1 U13171 ( .A1(n13089), .A2(n10505), .B1(n13092), .B2(n10504), .C1(
        P3_U3151), .C2(n10611), .ZN(P3_U3275) );
  INV_X1 U13172 ( .A(n10506), .ZN(n10545) );
  NAND3_X1 U13173 ( .A1(n10545), .A2(n10508), .A3(n10507), .ZN(n10509) );
  AOI21_X1 U13174 ( .B1(n10510), .B2(n10509), .A(n15017), .ZN(n10518) );
  AOI21_X1 U13175 ( .B1(n10341), .B2(n10511), .A(n10595), .ZN(n10516) );
  INV_X1 U13176 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11099) );
  NOR2_X1 U13177 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11099), .ZN(n10790) );
  NAND2_X1 U13178 ( .A1(n10512), .A2(n10340), .ZN(n10513) );
  AOI21_X1 U13179 ( .B1(n10601), .B2(n10513), .A(n15015), .ZN(n10514) );
  AOI211_X1 U13180 ( .C1(n14978), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10790), .B(
        n10514), .ZN(n10515) );
  OAI21_X1 U13181 ( .B1(n10516), .B2(n15023), .A(n10515), .ZN(n10517) );
  AOI211_X1 U13182 ( .C1(n14981), .C2(n10519), .A(n10518), .B(n10517), .ZN(
        n10520) );
  INV_X1 U13183 ( .A(n10520), .ZN(P3_U3185) );
  AOI22_X1 U13184 ( .A1(n13958), .A2(n10521), .B1(n12362), .B2(n6552), .ZN(
        n10658) );
  INV_X1 U13185 ( .A(n10523), .ZN(n10525) );
  XOR2_X1 U13186 ( .A(n10661), .B(n10662), .Z(n10530) );
  NOR2_X1 U13187 ( .A1(n13921), .A2(n14766), .ZN(n10528) );
  NAND2_X1 U13188 ( .A1(n13795), .A2(n14172), .ZN(n13903) );
  OAI22_X1 U13189 ( .A1(n11232), .A2(n13903), .B1(n13904), .B2(n12212), .ZN(
        n10527) );
  AOI211_X1 U13190 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n12208), .A(n10528), .B(
        n10527), .ZN(n10529) );
  OAI21_X1 U13191 ( .B1(n10530), .B2(n13938), .A(n10529), .ZN(P1_U3237) );
  AOI22_X1 U13192 ( .A1(n14978), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10541) );
  OAI21_X1 U13193 ( .B1(n10533), .B2(n10532), .A(n10531), .ZN(n10534) );
  NAND2_X1 U13194 ( .A1(n12732), .A2(n10534), .ZN(n10540) );
  OAI21_X1 U13195 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(n10538) );
  NAND2_X1 U13196 ( .A1(n12737), .A2(n10538), .ZN(n10539) );
  NAND3_X1 U13197 ( .A1(n10541), .A2(n10540), .A3(n10539), .ZN(n10547) );
  NAND3_X1 U13198 ( .A1(n10556), .A2(n10543), .A3(n10542), .ZN(n10544) );
  AOI21_X1 U13199 ( .B1(n10545), .B2(n10544), .A(n15017), .ZN(n10546) );
  AOI211_X1 U13200 ( .C1(n14981), .C2(n10548), .A(n10547), .B(n10546), .ZN(
        n10549) );
  INV_X1 U13201 ( .A(n10549), .ZN(P3_U3184) );
  NAND2_X1 U13202 ( .A1(n10550), .A2(n10330), .ZN(n10551) );
  NAND2_X1 U13203 ( .A1(n10552), .A2(n10551), .ZN(n10566) );
  INV_X1 U13204 ( .A(n10553), .ZN(n14943) );
  NAND2_X1 U13205 ( .A1(n14943), .A2(n10554), .ZN(n10555) );
  AOI21_X1 U13206 ( .B1(n10556), .B2(n10555), .A(n15017), .ZN(n10565) );
  NAND2_X1 U13207 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  NAND2_X1 U13208 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  NAND2_X1 U13209 ( .A1(n12737), .A2(n10561), .ZN(n10563) );
  NAND2_X1 U13210 ( .A1(n14978), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10562) );
  OAI211_X1 U13211 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n6736), .A(n10563), .B(
        n10562), .ZN(n10564) );
  AOI211_X1 U13212 ( .C1(n12732), .C2(n10566), .A(n10565), .B(n10564), .ZN(
        n10567) );
  OAI21_X1 U13213 ( .B1(n10568), .B2(n15007), .A(n10567), .ZN(P3_U3183) );
  XOR2_X1 U13214 ( .A(n10570), .B(n10569), .Z(n10571) );
  NAND2_X1 U13215 ( .A1(n10571), .A2(n14633), .ZN(n10577) );
  OAI22_X1 U13216 ( .A1(n10573), .A2(n13190), .B1(n10572), .B2(n13188), .ZN(
        n11119) );
  NOR2_X1 U13217 ( .A1(n13183), .A2(n6936), .ZN(n10574) );
  AOI211_X1 U13218 ( .C1(n14635), .C2(n11119), .A(n10575), .B(n10574), .ZN(
        n10576) );
  OAI211_X1 U13219 ( .C1(n14643), .C2(n11126), .A(n10577), .B(n10576), .ZN(
        P2_U3211) );
  AOI21_X1 U13220 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n10582), .A(n10578), .ZN(
        n10580) );
  XNOR2_X1 U13221 ( .A(n10760), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n10579) );
  NOR2_X1 U13222 ( .A1(n10580), .A2(n10579), .ZN(n10759) );
  AOI211_X1 U13223 ( .C1(n10580), .C2(n10579), .A(n14719), .B(n10759), .ZN(
        n10588) );
  MUX2_X1 U13224 ( .A(n14801), .B(P1_REG1_REG_10__SCAN_IN), .S(n10760), .Z(
        n10584) );
  NOR2_X1 U13225 ( .A1(n10583), .A2(n10584), .ZN(n10754) );
  AOI211_X1 U13226 ( .C1(n10584), .C2(n10583), .A(n14715), .B(n10754), .ZN(
        n10587) );
  INV_X1 U13227 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14412) );
  NAND2_X1 U13228 ( .A1(n14726), .A2(n10760), .ZN(n10585) );
  NAND2_X1 U13229 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n13773)
         );
  OAI211_X1 U13230 ( .C1(n14412), .C2(n14761), .A(n10585), .B(n13773), .ZN(
        n10586) );
  OR3_X1 U13231 ( .A1(n10588), .A2(n10587), .A3(n10586), .ZN(P1_U3253) );
  OAI21_X1 U13232 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10592) );
  NAND2_X1 U13233 ( .A1(n10592), .A2(n14999), .ZN(n10608) );
  OR3_X1 U13234 ( .A1(n10595), .A2(n10594), .A3(n10593), .ZN(n10596) );
  AOI21_X1 U13235 ( .B1(n10597), .B2(n10596), .A(n15023), .ZN(n10606) );
  INV_X1 U13236 ( .A(n10598), .ZN(n10600) );
  NAND3_X1 U13237 ( .A1(n10601), .A2(n10600), .A3(n10599), .ZN(n10602) );
  AOI21_X1 U13238 ( .B1(n10603), .B2(n10602), .A(n15015), .ZN(n10605) );
  NAND2_X1 U13239 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n11151) );
  OAI21_X1 U13240 ( .B1(n15008), .B2(n14399), .A(n11151), .ZN(n10604) );
  NOR3_X1 U13241 ( .A1(n10606), .A2(n10605), .A3(n10604), .ZN(n10607) );
  OAI211_X1 U13242 ( .C1(n15007), .C2(n10609), .A(n10608), .B(n10607), .ZN(
        P3_U3186) );
  INV_X1 U13243 ( .A(n12183), .ZN(n10610) );
  NAND2_X1 U13244 ( .A1(n13079), .A2(n10610), .ZN(n10613) );
  NAND3_X1 U13245 ( .A1(n15104), .A2(n12421), .A3(n10614), .ZN(n10615) );
  NAND2_X1 U13246 ( .A1(n13007), .A2(n12421), .ZN(n10616) );
  NAND2_X1 U13247 ( .A1(n10617), .A2(n10616), .ZN(n10618) );
  NAND3_X1 U13248 ( .A1(n13015), .A2(n13014), .A3(n12462), .ZN(n10619) );
  OAI211_X1 U13249 ( .C1(n10620), .C2(n13007), .A(n10690), .B(n10619), .ZN(
        n10647) );
  NAND3_X1 U13250 ( .A1(n10628), .A2(n10626), .A3(n15098), .ZN(n10622) );
  NAND2_X1 U13251 ( .A1(n10643), .A2(n10629), .ZN(n10621) );
  NAND2_X1 U13252 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  OR2_X1 U13253 ( .A1(n10628), .A2(n15102), .ZN(n10625) );
  INV_X1 U13254 ( .A(n10626), .ZN(n10627) );
  OR2_X1 U13255 ( .A1(n10628), .A2(n10627), .ZN(n10634) );
  INV_X1 U13256 ( .A(n10629), .ZN(n10630) );
  OR2_X1 U13257 ( .A1(n10643), .A2(n10630), .ZN(n10631) );
  NAND4_X1 U13258 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10635) );
  NAND2_X1 U13259 ( .A1(n10635), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10638) );
  OAI21_X1 U13260 ( .B1(n10643), .B2(n10640), .A(n12192), .ZN(n10636) );
  INV_X1 U13261 ( .A(n10636), .ZN(n10637) );
  NOR2_X1 U13262 ( .A1(n12578), .A2(P3_U3151), .ZN(n14940) );
  OR2_X1 U13263 ( .A1(n14940), .A2(n6736), .ZN(n10645) );
  INV_X1 U13264 ( .A(n10640), .ZN(n12188) );
  AND2_X1 U13265 ( .A1(n12188), .A2(n10641), .ZN(n10639) );
  NAND2_X1 U13266 ( .A1(n10643), .A2(n10639), .ZN(n12575) );
  INV_X1 U13267 ( .A(n12575), .ZN(n14932) );
  NOR2_X1 U13268 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  AOI22_X1 U13269 ( .A1(n14932), .A2(n13008), .B1(n13009), .B2(n12555), .ZN(
        n10644) );
  OAI211_X1 U13270 ( .C1(n13018), .C2(n14935), .A(n10645), .B(n10644), .ZN(
        n10646) );
  AOI21_X1 U13271 ( .B1(n10647), .B2(n14938), .A(n10646), .ZN(n10648) );
  INV_X1 U13272 ( .A(n10648), .ZN(P3_U3162) );
  XNOR2_X1 U13273 ( .A(n10650), .B(n10649), .ZN(n10656) );
  NAND2_X1 U13274 ( .A1(n13230), .A2(n13518), .ZN(n10652) );
  NAND2_X1 U13275 ( .A1(n13228), .A2(n13516), .ZN(n10651) );
  AND2_X1 U13276 ( .A1(n10652), .A2(n10651), .ZN(n11133) );
  NAND2_X1 U13277 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n13235) );
  OAI21_X1 U13278 ( .B1(n13178), .B2(n11133), .A(n13235), .ZN(n10654) );
  NOR2_X1 U13279 ( .A1(n14643), .A2(n11139), .ZN(n10653) );
  AOI211_X1 U13280 ( .C1(n14917), .C2(n14638), .A(n10654), .B(n10653), .ZN(
        n10655) );
  OAI21_X1 U13281 ( .B1(n10656), .B2(n13202), .A(n10655), .ZN(P2_U3185) );
  AOI22_X1 U13282 ( .A1(n13957), .A2(n10521), .B1(n12362), .B2(n10685), .ZN(
        n11205) );
  OAI22_X1 U13283 ( .A1(n11232), .A2(n6589), .B1(n10846), .B2(n10522), .ZN(
        n10657) );
  XNOR2_X1 U13284 ( .A(n10657), .B(n12364), .ZN(n11206) );
  XOR2_X1 U13285 ( .A(n11205), .B(n11206), .Z(n10664) );
  INV_X1 U13286 ( .A(n10658), .ZN(n10659) );
  AOI211_X1 U13287 ( .C1(n10664), .C2(n10663), .A(n13938), .B(n11208), .ZN(
        n10669) );
  INV_X1 U13288 ( .A(n13903), .ZN(n13884) );
  AOI22_X1 U13289 ( .A1(n13884), .A2(n13956), .B1(n10685), .B2(n13936), .ZN(
        n10667) );
  MUX2_X1 U13290 ( .A(n13887), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n10666) );
  OAI211_X1 U13291 ( .C1(n8675), .C2(n13904), .A(n10667), .B(n10666), .ZN(
        n10668) );
  OR2_X1 U13292 ( .A1(n10669), .A2(n10668), .ZN(P1_U3218) );
  INV_X1 U13293 ( .A(n10670), .ZN(n10673) );
  INV_X1 U13294 ( .A(n10893), .ZN(n14861) );
  OAI222_X1 U13295 ( .A1(n13736), .A2(n10671), .B1(n11298), .B2(n10673), .C1(
        n14861), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13296 ( .A1(P1_U3086), .A2(n14710), .B1(n14390), .B2(n10673), 
        .C1(n10672), .C2(n14384), .ZN(P1_U3340) );
  OAI222_X1 U13297 ( .A1(n13089), .A2(n10675), .B1(n13092), .B2(n10674), .C1(
        P3_U3151), .C2(n10934), .ZN(P3_U3274) );
  OAI21_X1 U13298 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10851) );
  OAI21_X1 U13299 ( .B1(n11937), .B2(n10680), .A(n10679), .ZN(n10681) );
  AOI222_X1 U13300 ( .A1(n14522), .A2(n10681), .B1(n13956), .B2(n14172), .C1(
        n13958), .C2(n14174), .ZN(n10847) );
  OAI21_X1 U13301 ( .B1(n10722), .B2(n10846), .A(n14512), .ZN(n10682) );
  OR2_X1 U13302 ( .A1(n10838), .A2(n10682), .ZN(n10845) );
  NAND2_X1 U13303 ( .A1(n10847), .A2(n10845), .ZN(n10683) );
  AOI21_X1 U13304 ( .B1(n14793), .B2(n10851), .A(n10683), .ZN(n10687) );
  AOI22_X1 U13305 ( .A1(n11173), .A2(n10685), .B1(n14794), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n10684) );
  OAI21_X1 U13306 ( .B1(n10687), .B2(n14794), .A(n10684), .ZN(P1_U3468) );
  AOI22_X1 U13307 ( .A1(n14235), .A2(n10685), .B1(n14800), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n10686) );
  OAI21_X1 U13308 ( .B1(n10687), .B2(n14800), .A(n10686), .ZN(P1_U3531) );
  INV_X1 U13309 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U13310 ( .A1(n12777), .A2(n12612), .ZN(n10688) );
  OAI21_X1 U13311 ( .B1(n12612), .B2(n15260), .A(n10688), .ZN(P3_U3518) );
  XNOR2_X1 U13312 ( .A(n15099), .B(n12421), .ZN(n10783) );
  XNOR2_X1 U13313 ( .A(n10783), .B(n13008), .ZN(n10692) );
  NAND2_X1 U13314 ( .A1(n10690), .A2(n10689), .ZN(n10691) );
  NAND2_X1 U13315 ( .A1(n10691), .A2(n10692), .ZN(n10785) );
  OAI21_X1 U13316 ( .B1(n10692), .B2(n10691), .A(n10785), .ZN(n10696) );
  OR2_X1 U13317 ( .A1(n14940), .A2(n15100), .ZN(n10694) );
  AOI22_X1 U13318 ( .A1(n14932), .A2(n9585), .B1(n15104), .B2(n12555), .ZN(
        n10693) );
  OAI211_X1 U13319 ( .C1(n14935), .C2(n15099), .A(n10694), .B(n10693), .ZN(
        n10695) );
  AOI21_X1 U13320 ( .B1(n10696), .B2(n14938), .A(n10695), .ZN(n10697) );
  INV_X1 U13321 ( .A(n10697), .ZN(P3_U3177) );
  INV_X1 U13322 ( .A(n10698), .ZN(n10700) );
  OAI22_X1 U13323 ( .A1(n12190), .A2(P3_U3151), .B1(SI_22_), .B2(n13092), .ZN(
        n10699) );
  AOI21_X1 U13324 ( .B1(n10700), .B2(n13084), .A(n10699), .ZN(P3_U3273) );
  INV_X1 U13325 ( .A(n14725), .ZN(n10703) );
  INV_X1 U13326 ( .A(n10701), .ZN(n10705) );
  OAI222_X1 U13327 ( .A1(P1_U3086), .A2(n10703), .B1(n14390), .B2(n10705), 
        .C1(n10702), .C2(n14384), .ZN(P1_U3339) );
  OAI222_X1 U13328 ( .A1(P2_U3088), .A2(n11357), .B1(n11298), .B2(n10705), 
        .C1(n10704), .C2(n13736), .ZN(P2_U3311) );
  OR2_X1 U13329 ( .A1(n10706), .A2(n11934), .ZN(n10707) );
  NAND2_X1 U13330 ( .A1(n10708), .A2(n10707), .ZN(n14768) );
  INV_X1 U13331 ( .A(n14524), .ZN(n14076) );
  NAND2_X1 U13332 ( .A1(n14768), .A2(n14076), .ZN(n10715) );
  NAND2_X1 U13333 ( .A1(n10709), .A2(n11934), .ZN(n10710) );
  NAND2_X1 U13334 ( .A1(n10711), .A2(n10710), .ZN(n10713) );
  OAI22_X1 U13335 ( .A1(n12212), .A2(n14212), .B1(n11232), .B2(n14210), .ZN(
        n10712) );
  AOI21_X1 U13336 ( .B1(n10713), .B2(n14522), .A(n10712), .ZN(n10714) );
  AND2_X1 U13337 ( .A1(n10715), .A2(n10714), .ZN(n14770) );
  NOR2_X1 U13338 ( .A1(n10717), .A2(n10716), .ZN(n10718) );
  NAND2_X1 U13339 ( .A1(n10719), .A2(n10718), .ZN(n12199) );
  INV_X1 U13340 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10721) );
  OAI22_X1 U13341 ( .A1(n14529), .A2(n10202), .B1(n10721), .B2(n14526), .ZN(
        n10727) );
  INV_X1 U13342 ( .A(n10722), .ZN(n10725) );
  AOI21_X1 U13343 ( .B1(n6552), .B2(n10723), .A(n14252), .ZN(n10724) );
  NAND2_X1 U13344 ( .A1(n10725), .A2(n10724), .ZN(n14765) );
  NOR2_X1 U13345 ( .A1(n14516), .A2(n14765), .ZN(n10726) );
  AOI211_X1 U13346 ( .C1(n14225), .C2(n6552), .A(n10727), .B(n10726), .ZN(
        n10732) );
  INV_X1 U13347 ( .A(n10282), .ZN(n10729) );
  NAND2_X1 U13348 ( .A1(n10729), .A2(n11760), .ZN(n11926) );
  INV_X1 U13349 ( .A(n11926), .ZN(n10730) );
  NAND2_X1 U13350 ( .A1(n14529), .A2(n10730), .ZN(n14517) );
  INV_X1 U13351 ( .A(n14517), .ZN(n14087) );
  NAND2_X1 U13352 ( .A1(n14768), .A2(n14087), .ZN(n10731) );
  OAI211_X1 U13353 ( .C1(n14770), .C2(n14224), .A(n10732), .B(n10731), .ZN(
        P1_U3291) );
  NAND2_X1 U13354 ( .A1(n10734), .A2(n10733), .ZN(n10736) );
  XOR2_X1 U13355 ( .A(n10736), .B(n10735), .Z(n10744) );
  NAND2_X1 U13356 ( .A1(n13229), .A2(n13518), .ZN(n10738) );
  NAND2_X1 U13357 ( .A1(n13227), .A2(n13516), .ZN(n10737) );
  NAND2_X1 U13358 ( .A1(n10738), .A2(n10737), .ZN(n10910) );
  INV_X1 U13359 ( .A(n10910), .ZN(n10740) );
  OAI22_X1 U13360 ( .A1(n13178), .A2(n10740), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10739), .ZN(n10742) );
  NOR2_X1 U13361 ( .A1(n14643), .A2(n11106), .ZN(n10741) );
  AOI211_X1 U13362 ( .C1(n10913), .C2(n14638), .A(n10742), .B(n10741), .ZN(
        n10743) );
  OAI21_X1 U13363 ( .B1(n10744), .B2(n13202), .A(n10743), .ZN(P2_U3193) );
  NAND2_X1 U13364 ( .A1(n12598), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10745) );
  OAI21_X1 U13365 ( .B1(n12148), .B2(n12598), .A(n10745), .ZN(P3_U3521) );
  NAND2_X1 U13366 ( .A1(n14529), .A2(n14076), .ZN(n10746) );
  AOI21_X1 U13367 ( .B1(n14522), .B2(n14529), .A(n14233), .ZN(n10753) );
  INV_X1 U13368 ( .A(n11935), .ZN(n10752) );
  INV_X1 U13369 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10747) );
  OAI22_X1 U13370 ( .A1(n14224), .A2(n10748), .B1(n10747), .B2(n14526), .ZN(
        n10749) );
  AOI21_X1 U13371 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14224), .A(n10749), .ZN(
        n10751) );
  NOR2_X1 U13372 ( .A1(n14516), .A2(n14252), .ZN(n14168) );
  OAI21_X1 U13373 ( .B1(n14168), .B2(n14225), .A(n12209), .ZN(n10750) );
  OAI211_X1 U13374 ( .C1(n10753), .C2(n10752), .A(n10751), .B(n10750), .ZN(
        P1_U3293) );
  INV_X1 U13375 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10755) );
  MUX2_X1 U13376 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10755), .S(n10952), .Z(
        n10756) );
  NAND2_X1 U13377 ( .A1(n10757), .A2(n10756), .ZN(n10951) );
  OAI21_X1 U13378 ( .B1(n10757), .B2(n10756), .A(n10951), .ZN(n10766) );
  INV_X1 U13379 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14416) );
  NAND2_X1 U13380 ( .A1(n14726), .A2(n10952), .ZN(n10758) );
  NAND2_X1 U13381 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13885)
         );
  OAI211_X1 U13382 ( .C1(n14416), .C2(n14761), .A(n10758), .B(n13885), .ZN(
        n10765) );
  INV_X1 U13383 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10761) );
  MUX2_X1 U13384 ( .A(n10761), .B(P1_REG2_REG_11__SCAN_IN), .S(n10952), .Z(
        n10762) );
  AOI211_X1 U13385 ( .C1(n10763), .C2(n10762), .A(n14719), .B(n10942), .ZN(
        n10764) );
  AOI211_X1 U13386 ( .C1(n14753), .C2(n10766), .A(n10765), .B(n10764), .ZN(
        n10767) );
  INV_X1 U13387 ( .A(n10767), .ZN(P1_U3254) );
  INV_X1 U13388 ( .A(n10768), .ZN(n14781) );
  OAI21_X1 U13389 ( .B1(n10770), .B2(n11940), .A(n10769), .ZN(n10779) );
  INV_X1 U13390 ( .A(n10840), .ZN(n10772) );
  INV_X1 U13391 ( .A(n11039), .ZN(n10771) );
  AOI211_X1 U13392 ( .C1(n11789), .C2(n10772), .A(n14252), .B(n10771), .ZN(
        n11015) );
  INV_X1 U13393 ( .A(n10779), .ZN(n11018) );
  OAI21_X1 U13394 ( .B1(n10775), .B2(n10774), .A(n10773), .ZN(n10777) );
  OAI22_X1 U13395 ( .A1(n11456), .A2(n14210), .B1(n11782), .B2(n14212), .ZN(
        n10776) );
  AOI21_X1 U13396 ( .B1(n10777), .B2(n14522), .A(n10776), .ZN(n10778) );
  OAI21_X1 U13397 ( .B1(n11018), .B2(n14524), .A(n10778), .ZN(n11012) );
  AOI211_X1 U13398 ( .C1(n14781), .C2(n10779), .A(n11015), .B(n11012), .ZN(
        n10782) );
  AOI22_X1 U13399 ( .A1(n14235), .A2(n11789), .B1(n14800), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n10780) );
  OAI21_X1 U13400 ( .B1(n10782), .B2(n14800), .A(n10780), .ZN(P1_U3533) );
  AOI22_X1 U13401 ( .A1(n11173), .A2(n11789), .B1(n14794), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n10781) );
  OAI21_X1 U13402 ( .B1(n10782), .B2(n14794), .A(n10781), .ZN(P1_U3474) );
  INV_X1 U13403 ( .A(n13008), .ZN(n10788) );
  NAND2_X1 U13404 ( .A1(n10788), .A2(n10783), .ZN(n10784) );
  XNOR2_X1 U13405 ( .A(n11098), .B(n12421), .ZN(n11144) );
  XNOR2_X1 U13406 ( .A(n11144), .B(n9585), .ZN(n10786) );
  OAI211_X1 U13407 ( .C1(n10787), .C2(n10786), .A(n11147), .B(n14938), .ZN(
        n10792) );
  OAI22_X1 U13408 ( .A1(n10788), .A2(n12587), .B1(n14935), .B2(n11098), .ZN(
        n10789) );
  AOI211_X1 U13409 ( .C1(n14932), .C2(n12611), .A(n10790), .B(n10789), .ZN(
        n10791) );
  OAI211_X1 U13410 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12590), .A(n10792), .B(
        n10791), .ZN(P3_U3158) );
  AOI22_X1 U13411 ( .A1(n10815), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n9244), .B2(
        n14962), .ZN(n14960) );
  MUX2_X1 U13412 ( .A(n10795), .B(P3_REG1_REG_8__SCAN_IN), .S(n14995), .Z(
        n14988) );
  NAND2_X1 U13413 ( .A1(n14995), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10796) );
  AOI21_X1 U13414 ( .B1(n15236), .B2(n10797), .A(n10854), .ZN(n10827) );
  AOI21_X1 U13415 ( .B1(n10800), .B2(n10799), .A(n10798), .ZN(n14954) );
  MUX2_X1 U13416 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n14941), .Z(n10801) );
  XNOR2_X1 U13417 ( .A(n10801), .B(n14962), .ZN(n14953) );
  OAI22_X1 U13418 ( .A1(n14954), .A2(n14953), .B1(n10801), .B2(n14962), .ZN(
        n14980) );
  MUX2_X1 U13419 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n14941), .Z(n10802) );
  XNOR2_X1 U13420 ( .A(n10802), .B(n14982), .ZN(n14979) );
  INV_X1 U13421 ( .A(n10802), .ZN(n10803) );
  AOI22_X1 U13422 ( .A1(n14980), .A2(n14979), .B1(n14982), .B2(n10803), .ZN(
        n14987) );
  MUX2_X1 U13423 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n14941), .Z(n10804) );
  XNOR2_X1 U13424 ( .A(n10804), .B(n14995), .ZN(n14986) );
  OAI22_X1 U13425 ( .A1(n14987), .A2(n14986), .B1(n10804), .B2(n14995), .ZN(
        n10808) );
  MUX2_X1 U13426 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n14941), .Z(n10805) );
  NAND2_X1 U13427 ( .A1(n10805), .A2(n6776), .ZN(n10809) );
  NAND2_X1 U13428 ( .A1(n10808), .A2(n10809), .ZN(n10865) );
  INV_X1 U13429 ( .A(n10805), .ZN(n10806) );
  NAND2_X1 U13430 ( .A1(n10806), .A2(n10868), .ZN(n10864) );
  INV_X1 U13431 ( .A(n10864), .ZN(n10807) );
  NOR2_X1 U13432 ( .A1(n10865), .A2(n10807), .ZN(n10811) );
  AOI21_X1 U13433 ( .B1(n10809), .B2(n10864), .A(n10808), .ZN(n10810) );
  OAI21_X1 U13434 ( .B1(n10811), .B2(n10810), .A(n14999), .ZN(n10826) );
  AOI22_X1 U13435 ( .A1(n10815), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n9243), .B2(
        n14962), .ZN(n14956) );
  MUX2_X1 U13436 ( .A(n10817), .B(P3_REG2_REG_8__SCAN_IN), .S(n14995), .Z(
        n14994) );
  NAND2_X1 U13437 ( .A1(n14995), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10818) );
  AOI21_X1 U13438 ( .B1(n15307), .B2(n10819), .A(n10869), .ZN(n10823) );
  NOR2_X1 U13439 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10820), .ZN(n11686) );
  NOR2_X1 U13440 ( .A1(n15007), .A2(n6776), .ZN(n10821) );
  AOI211_X1 U13441 ( .C1(n14978), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n11686), .B(
        n10821), .ZN(n10822) );
  OAI21_X1 U13442 ( .B1(n10823), .B2(n15023), .A(n10822), .ZN(n10824) );
  INV_X1 U13443 ( .A(n10824), .ZN(n10825) );
  OAI211_X1 U13444 ( .C1(n10827), .C2(n15015), .A(n10826), .B(n10825), .ZN(
        P3_U3191) );
  INV_X1 U13445 ( .A(n13984), .ZN(n14740) );
  INV_X1 U13446 ( .A(n10828), .ZN(n10830) );
  OAI222_X1 U13447 ( .A1(P1_U3086), .A2(n14740), .B1(n14390), .B2(n10830), 
        .C1(n10829), .C2(n14384), .ZN(P1_U3338) );
  INV_X1 U13448 ( .A(n13270), .ZN(n13267) );
  OAI222_X1 U13449 ( .A1(n13736), .A2(n10831), .B1(n11298), .B2(n10830), .C1(
        n13267), .C2(P2_U3088), .ZN(P2_U3310) );
  OAI21_X1 U13450 ( .B1(n11936), .B2(n10833), .A(n10832), .ZN(n10834) );
  AOI222_X1 U13451 ( .A1(n14522), .A2(n10834), .B1(n13955), .B2(n14172), .C1(
        n13957), .C2(n14174), .ZN(n14773) );
  MUX2_X1 U13452 ( .A(n10207), .B(n14773), .S(n14529), .Z(n10844) );
  OAI21_X1 U13453 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(n14776) );
  OAI21_X1 U13454 ( .B1(n10838), .B2(n14774), .A(n14512), .ZN(n10839) );
  OR2_X1 U13455 ( .A1(n10840), .A2(n10839), .ZN(n14772) );
  INV_X1 U13456 ( .A(n14526), .ZN(n14222) );
  AOI22_X1 U13457 ( .A1(n14225), .A2(n11783), .B1(n14222), .B2(n11229), .ZN(
        n10841) );
  OAI21_X1 U13458 ( .B1(n14516), .B2(n14772), .A(n10841), .ZN(n10842) );
  AOI21_X1 U13459 ( .B1(n14776), .B2(n14233), .A(n10842), .ZN(n10843) );
  NAND2_X1 U13460 ( .A1(n10844), .A2(n10843), .ZN(P1_U3289) );
  OAI22_X1 U13461 ( .A1(n10846), .A2(n14525), .B1(n10845), .B2(n14516), .ZN(
        n10850) );
  OAI21_X1 U13462 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n14526), .A(n10847), .ZN(
        n10848) );
  MUX2_X1 U13463 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10848), .S(n14529), .Z(
        n10849) );
  AOI211_X1 U13464 ( .C1(n14233), .C2(n10851), .A(n10850), .B(n10849), .ZN(
        n10852) );
  INV_X1 U13465 ( .A(n10852), .ZN(P1_U3290) );
  NOR2_X1 U13466 ( .A1(n10868), .A2(n10853), .ZN(n10855) );
  AOI22_X1 U13467 ( .A1(n10871), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n10858), 
        .B2(n11396), .ZN(n10856) );
  AOI21_X1 U13468 ( .B1(n10857), .B2(n10856), .A(n11382), .ZN(n10879) );
  MUX2_X1 U13469 ( .A(n10859), .B(n10858), .S(n14941), .Z(n10860) );
  NAND2_X1 U13470 ( .A1(n10860), .A2(n10871), .ZN(n11386) );
  INV_X1 U13471 ( .A(n10860), .ZN(n10861) );
  NAND2_X1 U13472 ( .A1(n10861), .A2(n11396), .ZN(n10862) );
  NAND2_X1 U13473 ( .A1(n11386), .A2(n10862), .ZN(n10863) );
  AOI21_X1 U13474 ( .B1(n10865), .B2(n10864), .A(n10863), .ZN(n11388) );
  AND3_X1 U13475 ( .A1(n10865), .A2(n10864), .A3(n10863), .ZN(n10866) );
  OAI21_X1 U13476 ( .B1(n11388), .B2(n10866), .A(n14999), .ZN(n10878) );
  NOR2_X1 U13477 ( .A1(n10868), .A2(n10867), .ZN(n10870) );
  AOI22_X1 U13478 ( .A1(n10871), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n10859), 
        .B2(n11396), .ZN(n10872) );
  OAI221_X1 U13479 ( .B1(n11395), .B2(n10873), .C1(n11395), .C2(n10872), .A(
        n12732), .ZN(n10875) );
  AND2_X1 U13480 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n11707) );
  AOI21_X1 U13481 ( .B1(n14978), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11707), 
        .ZN(n10874) );
  OAI211_X1 U13482 ( .C1(n11396), .C2(n15007), .A(n10875), .B(n10874), .ZN(
        n10876) );
  INV_X1 U13483 ( .A(n10876), .ZN(n10877) );
  OAI211_X1 U13484 ( .C1(n10879), .C2(n15015), .A(n10878), .B(n10877), .ZN(
        P3_U3192) );
  NAND2_X1 U13485 ( .A1(n10880), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U13486 ( .A1(n10882), .A2(n10881), .ZN(n14835) );
  XNOR2_X1 U13487 ( .A(n14837), .B(n10883), .ZN(n14834) );
  AOI21_X1 U13488 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14837), .A(n14840), 
        .ZN(n10884) );
  NOR2_X1 U13489 ( .A1(n10884), .A2(n14861), .ZN(n10885) );
  XNOR2_X1 U13490 ( .A(n14861), .B(n10884), .ZN(n14852) );
  NOR2_X1 U13491 ( .A1(n15235), .A2(n14852), .ZN(n14851) );
  NOR2_X1 U13492 ( .A1(n10885), .A2(n14851), .ZN(n10887) );
  XNOR2_X1 U13493 ( .A(n11359), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n10886) );
  NOR2_X1 U13494 ( .A1(n10887), .A2(n10886), .ZN(n11358) );
  AOI211_X1 U13495 ( .C1(n10887), .C2(n10886), .A(n14850), .B(n11358), .ZN(
        n10903) );
  OAI21_X1 U13496 ( .B1(n10235), .B2(n10889), .A(n10888), .ZN(n10891) );
  NAND2_X1 U13497 ( .A1(n14837), .A2(n10891), .ZN(n10892) );
  XNOR2_X1 U13498 ( .A(n10891), .B(n10890), .ZN(n14844) );
  NAND2_X1 U13499 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14844), .ZN(n14843) );
  NAND2_X1 U13500 ( .A1(n10892), .A2(n14843), .ZN(n10894) );
  NAND2_X1 U13501 ( .A1(n10893), .A2(n10894), .ZN(n10895) );
  XNOR2_X1 U13502 ( .A(n10894), .B(n14861), .ZN(n14858) );
  NAND2_X1 U13503 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14858), .ZN(n14856) );
  NAND2_X1 U13504 ( .A1(n10895), .A2(n14856), .ZN(n10899) );
  NAND2_X1 U13505 ( .A1(n11357), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n10896) );
  OAI21_X1 U13506 ( .B1(n11357), .B2(P2_REG2_REG_16__SCAN_IN), .A(n10896), 
        .ZN(n10898) );
  INV_X1 U13507 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13532) );
  NAND2_X1 U13508 ( .A1(n11357), .A2(n13532), .ZN(n10897) );
  OAI211_X1 U13509 ( .C1(n11357), .C2(n13532), .A(n10899), .B(n10897), .ZN(
        n11356) );
  OAI211_X1 U13510 ( .C1(n10899), .C2(n10898), .A(n11356), .B(n14857), .ZN(
        n10901) );
  NOR2_X1 U13511 ( .A1(n7947), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14639) );
  AOI21_X1 U13512 ( .B1(n14855), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14639), 
        .ZN(n10900) );
  OAI211_X1 U13513 ( .C1(n14862), .C2(n11357), .A(n10901), .B(n10900), .ZN(
        n10902) );
  OR2_X1 U13514 ( .A1(n10903), .A2(n10902), .ZN(P2_U3230) );
  INV_X1 U13515 ( .A(n10904), .ZN(n10907) );
  INV_X1 U13516 ( .A(n10908), .ZN(n10906) );
  OAI21_X1 U13517 ( .B1(n10907), .B2(n10906), .A(n10905), .ZN(n11112) );
  XNOR2_X1 U13518 ( .A(n10909), .B(n10908), .ZN(n10911) );
  AOI21_X1 U13519 ( .B1(n10911), .B2(n13540), .A(n10910), .ZN(n11104) );
  INV_X1 U13520 ( .A(n11137), .ZN(n10912) );
  AOI211_X1 U13521 ( .C1(n10913), .C2(n10912), .A(n9813), .B(n11185), .ZN(
        n11109) );
  AOI21_X1 U13522 ( .B1(n14918), .B2(n10913), .A(n11109), .ZN(n10914) );
  OAI211_X1 U13523 ( .C1(n11112), .C2(n14921), .A(n11104), .B(n10914), .ZN(
        n10916) );
  NAND2_X1 U13524 ( .A1(n10916), .A2(n14908), .ZN(n10915) );
  OAI21_X1 U13525 ( .B1(n14908), .B2(n7793), .A(n10915), .ZN(P2_U3454) );
  NAND2_X1 U13526 ( .A1(n10916), .A2(n14931), .ZN(n10917) );
  OAI21_X1 U13527 ( .B1(n14931), .B2(n10918), .A(n10917), .ZN(P2_U3507) );
  XNOR2_X1 U13528 ( .A(n10919), .B(n10921), .ZN(n10933) );
  OAI21_X1 U13529 ( .B1(n10922), .B2(n10921), .A(n10920), .ZN(n10924) );
  INV_X1 U13530 ( .A(n12611), .ZN(n11241) );
  INV_X1 U13531 ( .A(n12609), .ZN(n11472) );
  OAI22_X1 U13532 ( .A1(n11241), .A2(n15107), .B1(n11472), .B2(n15105), .ZN(
        n10923) );
  AOI21_X1 U13533 ( .B1(n10924), .B2(n15039), .A(n10923), .ZN(n10925) );
  OAI21_X1 U13534 ( .B1(n11591), .B2(n10933), .A(n10925), .ZN(n15143) );
  INV_X1 U13535 ( .A(n15143), .ZN(n10940) );
  NAND2_X1 U13536 ( .A1(n13077), .A2(n10926), .ZN(n10927) );
  OAI21_X1 U13537 ( .B1(n13077), .B2(n10928), .A(n10927), .ZN(n10929) );
  INV_X1 U13538 ( .A(n10929), .ZN(n10930) );
  NAND2_X1 U13539 ( .A1(n10931), .A2(n10930), .ZN(n10935) );
  INV_X1 U13540 ( .A(n10933), .ZN(n15145) );
  OR2_X1 U13541 ( .A1(n15123), .A2(n10934), .ZN(n15025) );
  NOR2_X1 U13542 ( .A1(n15038), .A2(n15025), .ZN(n15126) );
  OR2_X1 U13543 ( .A1(n10935), .A2(n15102), .ZN(n10974) );
  INV_X1 U13544 ( .A(n10974), .ZN(n15093) );
  NOR2_X1 U13545 ( .A1(n11240), .A2(n15098), .ZN(n15144) );
  AOI22_X1 U13546 ( .A1(n15093), .A2(n15144), .B1(n15125), .B2(n10936), .ZN(
        n10937) );
  OAI21_X1 U13547 ( .B1(n9225), .B2(n15129), .A(n10937), .ZN(n10938) );
  AOI21_X1 U13548 ( .B1(n15145), .B2(n15126), .A(n10938), .ZN(n10939) );
  OAI21_X1 U13549 ( .B1(n10940), .B2(n15038), .A(n10939), .ZN(P3_U3228) );
  NOR2_X1 U13550 ( .A1(n13978), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10941) );
  AOI21_X1 U13551 ( .B1(n13978), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10941), 
        .ZN(n10944) );
  OAI21_X1 U13552 ( .B1(n10944), .B2(n10943), .A(n13965), .ZN(n10949) );
  NAND2_X1 U13553 ( .A1(n10945), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10946) );
  NAND2_X1 U13554 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13807)
         );
  OAI211_X1 U13555 ( .C1(n14757), .C2(n10947), .A(n10946), .B(n13807), .ZN(
        n10948) );
  AOI21_X1 U13556 ( .B1(n10949), .B2(n14749), .A(n10948), .ZN(n10957) );
  INV_X1 U13557 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10950) );
  MUX2_X1 U13558 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10950), .S(n13978), .Z(
        n10954) );
  OAI21_X1 U13559 ( .B1(n10954), .B2(n10953), .A(n13977), .ZN(n10955) );
  NAND2_X1 U13560 ( .A1(n10955), .A2(n14753), .ZN(n10956) );
  NAND2_X1 U13561 ( .A1(n10957), .A2(n10956), .ZN(P1_U3255) );
  NAND2_X1 U13562 ( .A1(n10958), .A2(n13084), .ZN(n10959) );
  OAI211_X1 U13563 ( .C1(n10960), .C2(n13092), .A(n10959), .B(n12192), .ZN(
        P3_U3272) );
  INV_X1 U13564 ( .A(n10961), .ZN(n10962) );
  AOI21_X1 U13565 ( .B1(n10964), .B2(n10963), .A(n10962), .ZN(n10971) );
  OAI22_X1 U13566 ( .A1(n10966), .A2(n13190), .B1(n10965), .B2(n13188), .ZN(
        n11182) );
  AOI21_X1 U13567 ( .B1(n14635), .B2(n11182), .A(n10967), .ZN(n10968) );
  OAI21_X1 U13568 ( .B1(n11247), .B2(n14643), .A(n10968), .ZN(n10969) );
  AOI21_X1 U13569 ( .B1(n11250), .B2(n14638), .A(n10969), .ZN(n10970) );
  OAI21_X1 U13570 ( .B1(n10971), .B2(n13202), .A(n10970), .ZN(P2_U3203) );
  NAND2_X1 U13571 ( .A1(n13009), .A2(n14934), .ZN(n12011) );
  NAND2_X1 U13572 ( .A1(n13014), .A2(n12011), .ZN(n14937) );
  NOR2_X1 U13573 ( .A1(n10972), .A2(n15065), .ZN(n10973) );
  AOI22_X1 U13574 ( .A1(n14937), .A2(n10973), .B1(n15043), .B2(n15104), .ZN(
        n11758) );
  MUX2_X1 U13575 ( .A(n11758), .B(n14942), .S(n15038), .Z(n10976) );
  AOI22_X1 U13576 ( .A1(n12889), .A2(n11756), .B1(n15125), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U13577 ( .A1(n10976), .A2(n10975), .ZN(P3_U3233) );
  AND2_X1 U13578 ( .A1(n14891), .A2(n10977), .ZN(n10979) );
  NAND4_X1 U13579 ( .A1(n10980), .A2(n10979), .A3(n14890), .A4(n10978), .ZN(
        n10981) );
  INV_X1 U13580 ( .A(n11114), .ZN(n10982) );
  NAND2_X1 U13581 ( .A1(n6794), .A2(n10982), .ZN(n10983) );
  XOR2_X1 U13582 ( .A(n10991), .B(n10984), .Z(n14906) );
  INV_X2 U13583 ( .A(n13552), .ZN(n13557) );
  NAND2_X1 U13584 ( .A1(n13557), .A2(n13292), .ZN(n13549) );
  OAI211_X1 U13585 ( .C1(n6697), .C2(n6938), .A(n13528), .B(n11125), .ZN(
        n14901) );
  INV_X1 U13586 ( .A(n10985), .ZN(n10986) );
  INV_X1 U13587 ( .A(n13573), .ZN(n13544) );
  INV_X1 U13588 ( .A(n10987), .ZN(n10988) );
  AOI22_X1 U13589 ( .A1(n13577), .A2(n10989), .B1(n13544), .B2(n10988), .ZN(
        n10990) );
  OAI21_X1 U13590 ( .B1(n13549), .B2(n14901), .A(n10990), .ZN(n10997) );
  XNOR2_X1 U13591 ( .A(n10992), .B(n10991), .ZN(n10993) );
  NAND2_X1 U13592 ( .A1(n10993), .A2(n13540), .ZN(n10995) );
  NAND2_X1 U13593 ( .A1(n10995), .A2(n10994), .ZN(n14903) );
  MUX2_X1 U13594 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14903), .S(n13557), .Z(
        n10996) );
  AOI211_X1 U13595 ( .C1(n13579), .C2(n14906), .A(n10997), .B(n10996), .ZN(
        n10998) );
  INV_X1 U13596 ( .A(n10998), .ZN(P2_U3260) );
  XNOR2_X1 U13597 ( .A(n11006), .B(n10999), .ZN(n11001) );
  AOI21_X1 U13598 ( .B1(n11001), .B2(n13540), .A(n11000), .ZN(n14896) );
  INV_X1 U13599 ( .A(n11002), .ZN(n11003) );
  AOI211_X1 U13600 ( .C1(n11004), .C2(n6562), .A(n9813), .B(n11003), .ZN(
        n14894) );
  XNOR2_X1 U13601 ( .A(n11006), .B(n11005), .ZN(n14899) );
  AOI22_X1 U13602 ( .A1(n13581), .A2(n14894), .B1(n13579), .B2(n14899), .ZN(
        n11011) );
  OAI22_X1 U13603 ( .A1(n13557), .A2(n9963), .B1(n11007), .B2(n13573), .ZN(
        n11008) );
  AOI21_X1 U13604 ( .B1(n13577), .B2(n6562), .A(n11008), .ZN(n11010) );
  OAI211_X1 U13605 ( .C1(n13552), .C2(n14896), .A(n11011), .B(n11010), .ZN(
        P2_U3264) );
  NAND2_X1 U13606 ( .A1(n11012), .A2(n14529), .ZN(n11017) );
  AOI22_X1 U13607 ( .A1(n14224), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n11219), 
        .B2(n14222), .ZN(n11013) );
  OAI21_X1 U13608 ( .B1(n11788), .B2(n14525), .A(n11013), .ZN(n11014) );
  AOI21_X1 U13609 ( .B1(n11015), .B2(n14194), .A(n11014), .ZN(n11016) );
  OAI211_X1 U13610 ( .C1(n11018), .C2(n14517), .A(n11017), .B(n11016), .ZN(
        P1_U3288) );
  INV_X1 U13611 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U13612 ( .A1(n14168), .A2(n11020), .ZN(n11022) );
  AOI22_X1 U13613 ( .A1(n14224), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14222), .ZN(n11021) );
  OAI211_X1 U13614 ( .C1(n11023), .C2(n14525), .A(n11022), .B(n11021), .ZN(
        n11024) );
  AOI21_X1 U13615 ( .B1(n14233), .B2(n11025), .A(n11024), .ZN(n11026) );
  OAI21_X1 U13616 ( .B1(n11027), .B2(n14224), .A(n11026), .ZN(P1_U3292) );
  OR2_X1 U13617 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  NAND2_X1 U13618 ( .A1(n11031), .A2(n11030), .ZN(n14782) );
  NAND2_X1 U13619 ( .A1(n14782), .A2(n14076), .ZN(n11038) );
  OAI21_X1 U13620 ( .B1(n11944), .B2(n11033), .A(n11032), .ZN(n11036) );
  NAND2_X1 U13621 ( .A1(n13953), .A2(n14172), .ZN(n11034) );
  OAI21_X1 U13622 ( .B1(n11787), .B2(n14212), .A(n11034), .ZN(n11035) );
  AOI21_X1 U13623 ( .B1(n11036), .B2(n14522), .A(n11035), .ZN(n11037) );
  AND2_X1 U13624 ( .A1(n11038), .A2(n11037), .ZN(n14784) );
  AOI21_X1 U13625 ( .B1(n11039), .B2(n11795), .A(n14252), .ZN(n11040) );
  NAND2_X1 U13626 ( .A1(n11040), .A2(n11054), .ZN(n14778) );
  AOI22_X1 U13627 ( .A1(n14224), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n11041), 
        .B2(n14222), .ZN(n11043) );
  NAND2_X1 U13628 ( .A1(n14225), .A2(n11795), .ZN(n11042) );
  OAI211_X1 U13629 ( .C1(n14778), .C2(n14516), .A(n11043), .B(n11042), .ZN(
        n11044) );
  AOI21_X1 U13630 ( .B1(n14782), .B2(n14087), .A(n11044), .ZN(n11045) );
  OAI21_X1 U13631 ( .B1(n14784), .B2(n14224), .A(n11045), .ZN(P1_U3287) );
  OAI21_X1 U13632 ( .B1(n11048), .B2(n11047), .A(n11046), .ZN(n11171) );
  INV_X1 U13633 ( .A(n11171), .ZN(n11060) );
  OAI21_X1 U13634 ( .B1(n11050), .B2(n11942), .A(n11049), .ZN(n11052) );
  OAI22_X1 U13635 ( .A1(n11456), .A2(n14212), .B1(n11719), .B2(n14210), .ZN(
        n11051) );
  AOI21_X1 U13636 ( .B1(n11052), .B2(n14522), .A(n11051), .ZN(n11053) );
  OAI21_X1 U13637 ( .B1(n11060), .B2(n14524), .A(n11053), .ZN(n11169) );
  NAND2_X1 U13638 ( .A1(n11169), .A2(n14529), .ZN(n11059) );
  XNOR2_X1 U13639 ( .A(n11054), .B(n11799), .ZN(n11055) );
  NOR2_X1 U13640 ( .A1(n11055), .A2(n14252), .ZN(n11170) );
  AOI22_X1 U13641 ( .A1(n14224), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n11453), 
        .B2(n14222), .ZN(n11056) );
  OAI21_X1 U13642 ( .B1(n6869), .B2(n14525), .A(n11056), .ZN(n11057) );
  AOI21_X1 U13643 ( .B1(n11170), .B2(n14194), .A(n11057), .ZN(n11058) );
  OAI211_X1 U13644 ( .C1(n11060), .C2(n14517), .A(n11059), .B(n11058), .ZN(
        P1_U3286) );
  OAI22_X1 U13645 ( .A1(n13486), .A2(n11062), .B1(n13573), .B2(n11061), .ZN(
        n11063) );
  AOI21_X1 U13646 ( .B1(n13581), .B2(n11064), .A(n11063), .ZN(n11068) );
  MUX2_X1 U13647 ( .A(n11066), .B(n11065), .S(n13557), .Z(n11067) );
  OAI211_X1 U13648 ( .C1(n13509), .C2(n11069), .A(n11068), .B(n11067), .ZN(
        P2_U3261) );
  OAI22_X1 U13649 ( .A1(n13486), .A2(n11071), .B1(n13573), .B2(n11070), .ZN(
        n11072) );
  AOI21_X1 U13650 ( .B1(n13581), .B2(n11073), .A(n11072), .ZN(n11077) );
  MUX2_X1 U13651 ( .A(n11075), .B(n11074), .S(n13557), .Z(n11076) );
  OAI211_X1 U13652 ( .C1(n13509), .C2(n11078), .A(n11077), .B(n11076), .ZN(
        P2_U3263) );
  OAI22_X1 U13653 ( .A1(n13486), .A2(n11079), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13573), .ZN(n11080) );
  AOI21_X1 U13654 ( .B1(n13581), .B2(n11081), .A(n11080), .ZN(n11085) );
  MUX2_X1 U13655 ( .A(n11083), .B(n11082), .S(n13557), .Z(n11084) );
  OAI211_X1 U13656 ( .C1(n13509), .C2(n11086), .A(n11085), .B(n11084), .ZN(
        P2_U3262) );
  XNOR2_X1 U13657 ( .A(n12162), .B(n11087), .ZN(n15137) );
  INV_X1 U13658 ( .A(n15137), .ZN(n11103) );
  INV_X1 U13659 ( .A(n15126), .ZN(n11102) );
  NAND2_X1 U13660 ( .A1(n15137), .A2(n15115), .ZN(n11096) );
  NAND2_X1 U13661 ( .A1(n15112), .A2(n11088), .ZN(n11089) );
  AOI21_X1 U13662 ( .B1(n11089), .B2(n12162), .A(n15110), .ZN(n11094) );
  NAND2_X1 U13663 ( .A1(n12611), .A2(n15043), .ZN(n11091) );
  NAND2_X1 U13664 ( .A1(n13008), .A2(n15046), .ZN(n11090) );
  NAND2_X1 U13665 ( .A1(n11091), .A2(n11090), .ZN(n11092) );
  AOI21_X1 U13666 ( .B1(n11094), .B2(n11093), .A(n11092), .ZN(n11095) );
  NAND2_X1 U13667 ( .A1(n11096), .A2(n11095), .ZN(n15135) );
  MUX2_X1 U13668 ( .A(n15135), .B(P3_REG2_REG_3__SCAN_IN), .S(n15038), .Z(
        n11097) );
  INV_X1 U13669 ( .A(n11097), .ZN(n11101) );
  NOR2_X1 U13670 ( .A1(n11098), .A2(n15098), .ZN(n15136) );
  AOI22_X1 U13671 ( .A1(n15093), .A2(n15136), .B1(n15125), .B2(n11099), .ZN(
        n11100) );
  OAI211_X1 U13672 ( .C1(n11103), .C2(n11102), .A(n11101), .B(n11100), .ZN(
        P3_U3230) );
  MUX2_X1 U13673 ( .A(n11105), .B(n11104), .S(n13557), .Z(n11111) );
  OAI22_X1 U13674 ( .A1(n13486), .A2(n11107), .B1(n13573), .B2(n11106), .ZN(
        n11108) );
  AOI21_X1 U13675 ( .B1(n11109), .B2(n13581), .A(n11108), .ZN(n11110) );
  OAI211_X1 U13676 ( .C1(n13509), .C2(n11112), .A(n11111), .B(n11110), .ZN(
        P2_U3257) );
  XOR2_X1 U13677 ( .A(n11115), .B(n11113), .Z(n11122) );
  INV_X1 U13678 ( .A(n11122), .ZN(n14913) );
  NAND2_X1 U13679 ( .A1(n13557), .A2(n11114), .ZN(n13395) );
  INV_X1 U13680 ( .A(n6794), .ZN(n11121) );
  NAND2_X1 U13681 ( .A1(n11116), .A2(n11115), .ZN(n11117) );
  AOI21_X1 U13682 ( .B1(n11118), .B2(n11117), .A(n13562), .ZN(n11120) );
  AOI211_X1 U13683 ( .C1(n11122), .C2(n11121), .A(n11120), .B(n11119), .ZN(
        n14912) );
  MUX2_X1 U13684 ( .A(n11123), .B(n14912), .S(n13557), .Z(n11129) );
  INV_X1 U13685 ( .A(n11138), .ZN(n11124) );
  AOI211_X1 U13686 ( .C1(n14910), .C2(n11125), .A(n9813), .B(n11124), .ZN(
        n14909) );
  OAI22_X1 U13687 ( .A1(n13486), .A2(n6936), .B1(n13573), .B2(n11126), .ZN(
        n11127) );
  AOI21_X1 U13688 ( .B1(n14909), .B2(n13581), .A(n11127), .ZN(n11128) );
  OAI211_X1 U13689 ( .C1(n14913), .C2(n13395), .A(n11129), .B(n11128), .ZN(
        P2_U3259) );
  XOR2_X1 U13690 ( .A(n11130), .B(n11131), .Z(n14922) );
  XNOR2_X1 U13691 ( .A(n11132), .B(n11131), .ZN(n11135) );
  INV_X1 U13692 ( .A(n11133), .ZN(n11134) );
  AOI21_X1 U13693 ( .B1(n11135), .B2(n13540), .A(n11134), .ZN(n14920) );
  MUX2_X1 U13694 ( .A(n14920), .B(n11136), .S(n13552), .Z(n11143) );
  AOI211_X1 U13695 ( .C1(n14917), .C2(n11138), .A(n9813), .B(n11137), .ZN(
        n14916) );
  INV_X1 U13696 ( .A(n14917), .ZN(n11140) );
  OAI22_X1 U13697 ( .A1(n13486), .A2(n11140), .B1(n13573), .B2(n11139), .ZN(
        n11141) );
  AOI21_X1 U13698 ( .B1(n14916), .B2(n13581), .A(n11141), .ZN(n11142) );
  OAI211_X1 U13699 ( .C1(n13509), .C2(n14922), .A(n11143), .B(n11142), .ZN(
        P2_U3258) );
  XNOR2_X1 U13700 ( .A(n15090), .B(n12421), .ZN(n11236) );
  XNOR2_X1 U13701 ( .A(n11236), .B(n12611), .ZN(n11149) );
  INV_X1 U13702 ( .A(n11144), .ZN(n11145) );
  NAND2_X1 U13703 ( .A1(n11145), .A2(n9585), .ZN(n11146) );
  OAI21_X1 U13704 ( .B1(n11149), .B2(n11148), .A(n11238), .ZN(n11150) );
  NAND2_X1 U13705 ( .A1(n11150), .A2(n14938), .ZN(n11155) );
  INV_X1 U13706 ( .A(n11151), .ZN(n11153) );
  INV_X1 U13707 ( .A(n9585), .ZN(n15106) );
  OAI22_X1 U13708 ( .A1(n15106), .A2(n12587), .B1(n14935), .B2(n15090), .ZN(
        n11152) );
  AOI211_X1 U13709 ( .C1(n14932), .C2(n12610), .A(n11153), .B(n11152), .ZN(
        n11154) );
  OAI211_X1 U13710 ( .C1(n15091), .C2(n12590), .A(n11155), .B(n11154), .ZN(
        P3_U3170) );
  OAI21_X1 U13711 ( .B1(n11157), .B2(n11158), .A(n11156), .ZN(n11330) );
  OAI211_X1 U13712 ( .C1(n11160), .C2(n8411), .A(n14522), .B(n11159), .ZN(
        n11325) );
  AOI22_X1 U13713 ( .A1(n13951), .A2(n14172), .B1(n14174), .B2(n13953), .ZN(
        n11627) );
  INV_X1 U13714 ( .A(n11161), .ZN(n11311) );
  OAI211_X1 U13715 ( .C1(n11632), .C2(n11162), .A(n11311), .B(n14512), .ZN(
        n11326) );
  NAND3_X1 U13716 ( .A1(n11325), .A2(n11627), .A3(n11326), .ZN(n11163) );
  AOI21_X1 U13717 ( .B1(n14793), .B2(n11330), .A(n11163), .ZN(n11168) );
  AOI22_X1 U13718 ( .A1(n14235), .A2(n11806), .B1(n14800), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n11164) );
  OAI21_X1 U13719 ( .B1(n11168), .B2(n14800), .A(n11164), .ZN(P1_U3536) );
  INV_X1 U13720 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11165) );
  OAI22_X1 U13721 ( .A1(n8752), .A2(n11632), .B1(n14796), .B2(n11165), .ZN(
        n11166) );
  INV_X1 U13722 ( .A(n11166), .ZN(n11167) );
  OAI21_X1 U13723 ( .B1(n11168), .B2(n14794), .A(n11167), .ZN(P1_U3483) );
  AOI211_X1 U13724 ( .C1(n14781), .C2(n11171), .A(n11170), .B(n11169), .ZN(
        n11175) );
  AOI22_X1 U13725 ( .A1(n14235), .A2(n11799), .B1(n14800), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n11172) );
  OAI21_X1 U13726 ( .B1(n11175), .B2(n14800), .A(n11172), .ZN(P1_U3535) );
  AOI22_X1 U13727 ( .A1(n11173), .A2(n11799), .B1(n14794), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n11174) );
  OAI21_X1 U13728 ( .B1(n11175), .B2(n14794), .A(n11174), .ZN(P1_U3480) );
  INV_X1 U13729 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11189) );
  OR2_X1 U13730 ( .A1(n11177), .A2(n11176), .ZN(n11178) );
  NAND2_X1 U13731 ( .A1(n11179), .A2(n11178), .ZN(n11254) );
  XNOR2_X1 U13732 ( .A(n11181), .B(n11180), .ZN(n11183) );
  AOI21_X1 U13733 ( .B1(n11183), .B2(n13540), .A(n11182), .ZN(n11257) );
  OAI21_X1 U13734 ( .B1(n11185), .B2(n11184), .A(n13528), .ZN(n11186) );
  NOR2_X1 U13735 ( .A1(n11186), .A2(n11270), .ZN(n11251) );
  AOI21_X1 U13736 ( .B1(n14918), .B2(n11250), .A(n11251), .ZN(n11187) );
  OAI211_X1 U13737 ( .C1(n11254), .C2(n14921), .A(n11257), .B(n11187), .ZN(
        n11190) );
  NAND2_X1 U13738 ( .A1(n11190), .A2(n14908), .ZN(n11188) );
  OAI21_X1 U13739 ( .B1(n14908), .B2(n11189), .A(n11188), .ZN(P2_U3457) );
  NAND2_X1 U13740 ( .A1(n11190), .A2(n14931), .ZN(n11191) );
  OAI21_X1 U13741 ( .B1(n14931), .B2(n10104), .A(n11191), .ZN(P2_U3508) );
  OAI211_X1 U13742 ( .C1(n6696), .C2(n11193), .A(n11192), .B(n14633), .ZN(
        n11200) );
  INV_X1 U13743 ( .A(n11266), .ZN(n11198) );
  NAND2_X1 U13744 ( .A1(n13227), .A2(n13518), .ZN(n11195) );
  NAND2_X1 U13745 ( .A1(n13225), .A2(n13516), .ZN(n11194) );
  NAND2_X1 U13746 ( .A1(n11195), .A2(n11194), .ZN(n11260) );
  INV_X1 U13747 ( .A(n11260), .ZN(n11196) );
  OAI22_X1 U13748 ( .A1(n13178), .A2(n11196), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7829), .ZN(n11197) );
  AOI21_X1 U13749 ( .B1(n11198), .B2(n9845), .A(n11197), .ZN(n11199) );
  OAI211_X1 U13750 ( .C1(n11269), .C2(n13183), .A(n11200), .B(n11199), .ZN(
        P2_U3189) );
  INV_X1 U13751 ( .A(n11201), .ZN(n11203) );
  OAI222_X1 U13752 ( .A1(P1_U3086), .A2(n14756), .B1(n14390), .B2(n11203), 
        .C1(n11202), .C2(n14384), .ZN(P1_U3337) );
  INV_X1 U13753 ( .A(n13283), .ZN(n13277) );
  OAI222_X1 U13754 ( .A1(n13736), .A2(n11204), .B1(n11298), .B2(n11203), .C1(
        n13277), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13755 ( .A(n11205), .ZN(n11207) );
  OR2_X1 U13756 ( .A1(n11782), .A2(n12345), .ZN(n11210) );
  NAND2_X1 U13757 ( .A1(n12362), .A2(n11783), .ZN(n11209) );
  NAND2_X1 U13758 ( .A1(n11210), .A2(n11209), .ZN(n11213) );
  OAI22_X1 U13759 ( .A1(n11782), .A2(n12305), .B1(n14774), .B2(n10522), .ZN(
        n11211) );
  XOR2_X1 U13760 ( .A(n12364), .B(n11211), .Z(n11228) );
  OAI22_X1 U13761 ( .A1(n11787), .A2(n6589), .B1(n11788), .B2(n10522), .ZN(
        n11215) );
  XNOR2_X1 U13762 ( .A(n11215), .B(n12364), .ZN(n11368) );
  OR2_X1 U13763 ( .A1(n11787), .A2(n12345), .ZN(n11217) );
  NAND2_X1 U13764 ( .A1(n11789), .A2(n12366), .ZN(n11216) );
  NAND2_X1 U13765 ( .A1(n11217), .A2(n11216), .ZN(n11369) );
  XNOR2_X1 U13766 ( .A(n11368), .B(n11369), .ZN(n11218) );
  XNOR2_X1 U13767 ( .A(n11370), .B(n11218), .ZN(n11225) );
  INV_X1 U13768 ( .A(n11219), .ZN(n11221) );
  OAI21_X1 U13769 ( .B1(n13887), .B2(n11221), .A(n11220), .ZN(n11223) );
  OAI22_X1 U13770 ( .A1(n11456), .A2(n13903), .B1(n13904), .B2(n11782), .ZN(
        n11222) );
  AOI211_X1 U13771 ( .C1(n11789), .C2(n13936), .A(n11223), .B(n11222), .ZN(
        n11224) );
  OAI21_X1 U13772 ( .B1(n11225), .B2(n13938), .A(n11224), .ZN(P1_U3227) );
  AOI211_X1 U13773 ( .C1(n11228), .C2(n11227), .A(n13938), .B(n11226), .ZN(
        n11235) );
  OAI22_X1 U13774 ( .A1(n13921), .A2(n14774), .B1(n13903), .B2(n11787), .ZN(
        n11234) );
  INV_X1 U13775 ( .A(n13887), .ZN(n13932) );
  NAND2_X1 U13776 ( .A1(n13932), .A2(n11229), .ZN(n11231) );
  OAI211_X1 U13777 ( .C1(n13904), .C2(n11232), .A(n11231), .B(n11230), .ZN(
        n11233) );
  OR3_X1 U13778 ( .A1(n11235), .A2(n11234), .A3(n11233), .ZN(P1_U3230) );
  NAND2_X1 U13779 ( .A1(n11241), .A2(n11236), .ZN(n11237) );
  XNOR2_X1 U13780 ( .A(n11240), .B(n12421), .ZN(n11463) );
  XNOR2_X1 U13781 ( .A(n11463), .B(n12610), .ZN(n11461) );
  XNOR2_X1 U13782 ( .A(n11462), .B(n11461), .ZN(n11239) );
  NAND2_X1 U13783 ( .A1(n11239), .A2(n14938), .ZN(n11245) );
  OAI22_X1 U13784 ( .A1(n11241), .A2(n12587), .B1(n14935), .B2(n11240), .ZN(
        n11242) );
  AOI211_X1 U13785 ( .C1(n14932), .C2(n12609), .A(n11243), .B(n11242), .ZN(
        n11244) );
  OAI211_X1 U13786 ( .C1(n11246), .C2(n12590), .A(n11245), .B(n11244), .ZN(
        P3_U3167) );
  OAI22_X1 U13787 ( .A1(n13557), .A2(n11248), .B1(n11247), .B2(n13573), .ZN(
        n11249) );
  AOI21_X1 U13788 ( .B1(n13577), .B2(n11250), .A(n11249), .ZN(n11253) );
  NAND2_X1 U13789 ( .A1(n11251), .A2(n13581), .ZN(n11252) );
  OAI211_X1 U13790 ( .C1(n11254), .C2(n13509), .A(n11253), .B(n11252), .ZN(
        n11255) );
  INV_X1 U13791 ( .A(n11255), .ZN(n11256) );
  OAI21_X1 U13792 ( .B1(n13552), .B2(n11257), .A(n11256), .ZN(P2_U3256) );
  XNOR2_X1 U13793 ( .A(n11259), .B(n11258), .ZN(n11261) );
  AOI21_X1 U13794 ( .B1(n11261), .B2(n13540), .A(n11260), .ZN(n11279) );
  OR2_X1 U13795 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  NAND2_X1 U13796 ( .A1(n11265), .A2(n11264), .ZN(n11280) );
  OAI22_X1 U13797 ( .A1(n13557), .A2(n11267), .B1(n11266), .B2(n13573), .ZN(
        n11268) );
  AOI21_X1 U13798 ( .B1(n11277), .B2(n13577), .A(n11268), .ZN(n11273) );
  OR2_X1 U13799 ( .A1(n11270), .A2(n11269), .ZN(n11271) );
  AND3_X1 U13800 ( .A1(n11349), .A2(n11271), .A3(n13528), .ZN(n11276) );
  NAND2_X1 U13801 ( .A1(n11276), .A2(n13581), .ZN(n11272) );
  OAI211_X1 U13802 ( .C1(n11280), .C2(n13509), .A(n11273), .B(n11272), .ZN(
        n11274) );
  INV_X1 U13803 ( .A(n11274), .ZN(n11275) );
  OAI21_X1 U13804 ( .B1(n13552), .B2(n11279), .A(n11275), .ZN(P2_U3255) );
  AOI21_X1 U13805 ( .B1(n14918), .B2(n11277), .A(n11276), .ZN(n11278) );
  OAI211_X1 U13806 ( .C1(n11280), .C2(n14921), .A(n11279), .B(n11278), .ZN(
        n11294) );
  NAND2_X1 U13807 ( .A1(n11294), .A2(n14908), .ZN(n11281) );
  OAI21_X1 U13808 ( .B1(n14908), .B2(n7827), .A(n11281), .ZN(P2_U3460) );
  NAND2_X1 U13809 ( .A1(n11282), .A2(n11283), .ZN(n15057) );
  XNOR2_X1 U13810 ( .A(n15057), .B(n15056), .ZN(n11288) );
  XNOR2_X1 U13811 ( .A(n11285), .B(n11284), .ZN(n15153) );
  INV_X1 U13812 ( .A(n15045), .ZN(n11684) );
  OAI22_X1 U13813 ( .A1(n11684), .A2(n15105), .B1(n11472), .B2(n15107), .ZN(
        n11286) );
  AOI21_X1 U13814 ( .B1(n15153), .B2(n15115), .A(n11286), .ZN(n11287) );
  OAI21_X1 U13815 ( .B1(n11288), .B2(n15110), .A(n11287), .ZN(n15151) );
  INV_X1 U13816 ( .A(n15151), .ZN(n11293) );
  NOR2_X1 U13817 ( .A1(n11471), .A2(n15098), .ZN(n15152) );
  INV_X1 U13818 ( .A(n11476), .ZN(n11289) );
  AOI22_X1 U13819 ( .A1(n15093), .A2(n15152), .B1(n15125), .B2(n11289), .ZN(
        n11290) );
  OAI21_X1 U13820 ( .B1(n9265), .B2(n15129), .A(n11290), .ZN(n11291) );
  AOI21_X1 U13821 ( .B1(n15153), .B2(n15126), .A(n11291), .ZN(n11292) );
  OAI21_X1 U13822 ( .B1(n11293), .B2(n15038), .A(n11292), .ZN(P3_U3226) );
  NAND2_X1 U13823 ( .A1(n11294), .A2(n14931), .ZN(n11295) );
  OAI21_X1 U13824 ( .B1(n14931), .B2(n10108), .A(n11295), .ZN(P2_U3509) );
  INV_X1 U13825 ( .A(n11296), .ZN(n11297) );
  OAI222_X1 U13826 ( .A1(n13992), .A2(P1_U3086), .B1(n14390), .B2(n11297), 
        .C1(n15248), .C2(n14384), .ZN(P1_U3336) );
  OAI222_X1 U13827 ( .A1(n13736), .A2(n11299), .B1(n11298), .B2(n11297), .C1(
        n13292), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U13828 ( .A(n11300), .ZN(n11321) );
  OAI222_X1 U13829 ( .A1(P1_U3086), .A2(n11925), .B1(n14390), .B2(n11321), 
        .C1(n11301), .C2(n14384), .ZN(P1_U3335) );
  OAI21_X1 U13830 ( .B1(n11303), .B2(n11946), .A(n11302), .ZN(n11423) );
  INV_X1 U13831 ( .A(n11423), .ZN(n11316) );
  INV_X1 U13832 ( .A(n11304), .ZN(n11305) );
  AOI21_X1 U13833 ( .B1(n11946), .B2(n11306), .A(n11305), .ZN(n11309) );
  AOI22_X1 U13834 ( .A1(n14174), .A2(n13952), .B1(n13950), .B2(n14172), .ZN(
        n11308) );
  NAND2_X1 U13835 ( .A1(n11423), .A2(n14076), .ZN(n11307) );
  OAI211_X1 U13836 ( .C1(n11309), .C2(n14110), .A(n11308), .B(n11307), .ZN(
        n11421) );
  NAND2_X1 U13837 ( .A1(n11421), .A2(n14529), .ZN(n11315) );
  INV_X1 U13838 ( .A(n11525), .ZN(n11310) );
  AOI211_X1 U13839 ( .C1(n11810), .C2(n11311), .A(n14252), .B(n11310), .ZN(
        n11422) );
  AOI22_X1 U13840 ( .A1(n14224), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11722), 
        .B2(n14222), .ZN(n11312) );
  OAI21_X1 U13841 ( .B1(n11725), .B2(n14525), .A(n11312), .ZN(n11313) );
  AOI21_X1 U13842 ( .B1(n11422), .B2(n14194), .A(n11313), .ZN(n11314) );
  OAI211_X1 U13843 ( .C1(n11316), .C2(n14517), .A(n11315), .B(n11314), .ZN(
        P1_U3284) );
  INV_X1 U13844 ( .A(n11317), .ZN(n11319) );
  OAI222_X1 U13845 ( .A1(n11320), .A2(P3_U3151), .B1(n13089), .B2(n11319), 
        .C1(n11318), .C2(n13092), .ZN(P3_U3271) );
  OAI222_X1 U13846 ( .A1(n13736), .A2(n11323), .B1(P2_U3088), .B2(n6771), .C1(
        n11298), .C2(n11321), .ZN(P2_U3307) );
  INV_X1 U13847 ( .A(n11629), .ZN(n11324) );
  OAI22_X1 U13848 ( .A1(n11632), .A2(n14525), .B1(n11324), .B2(n14526), .ZN(
        n11329) );
  OAI211_X1 U13849 ( .C1(n11760), .C2(n11326), .A(n11325), .B(n11627), .ZN(
        n11327) );
  MUX2_X1 U13850 ( .A(n11327), .B(P1_REG2_REG_8__SCAN_IN), .S(n14224), .Z(
        n11328) );
  AOI211_X1 U13851 ( .C1(n14233), .C2(n11330), .A(n11329), .B(n11328), .ZN(
        n11331) );
  INV_X1 U13852 ( .A(n11331), .ZN(P1_U3285) );
  INV_X1 U13853 ( .A(n11479), .ZN(n11340) );
  OAI21_X1 U13854 ( .B1(n11334), .B2(n11333), .A(n11429), .ZN(n11335) );
  NAND2_X1 U13855 ( .A1(n11335), .A2(n14633), .ZN(n11339) );
  INV_X1 U13856 ( .A(n11346), .ZN(n11337) );
  AOI22_X1 U13857 ( .A1(n13518), .A2(n13226), .B1(n13224), .B2(n13516), .ZN(
        n11342) );
  OAI22_X1 U13858 ( .A1(n13178), .A2(n11342), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15348), .ZN(n11336) );
  AOI21_X1 U13859 ( .B1(n11337), .B2(n9845), .A(n11336), .ZN(n11338) );
  OAI211_X1 U13860 ( .C1(n11340), .C2(n13183), .A(n11339), .B(n11338), .ZN(
        P2_U3208) );
  XOR2_X1 U13861 ( .A(n11341), .B(n11345), .Z(n11343) );
  OAI21_X1 U13862 ( .B1(n11343), .B2(n13562), .A(n11342), .ZN(n11477) );
  XOR2_X1 U13863 ( .A(n11345), .B(n11344), .Z(n11481) );
  OAI22_X1 U13864 ( .A1(n13557), .A2(n11347), .B1(n11346), .B2(n13573), .ZN(
        n11348) );
  AOI21_X1 U13865 ( .B1(n11479), .B2(n13577), .A(n11348), .ZN(n11352) );
  AOI21_X1 U13866 ( .B1(n11349), .B2(n11479), .A(n13564), .ZN(n11350) );
  AND2_X1 U13867 ( .A1(n11350), .A2(n11484), .ZN(n11478) );
  NAND2_X1 U13868 ( .A1(n11478), .A2(n13581), .ZN(n11351) );
  OAI211_X1 U13869 ( .C1(n11481), .C2(n13509), .A(n11352), .B(n11351), .ZN(
        n11353) );
  AOI21_X1 U13870 ( .B1(n13557), .B2(n11477), .A(n11353), .ZN(n11354) );
  INV_X1 U13871 ( .A(n11354), .ZN(P2_U3254) );
  NAND2_X1 U13872 ( .A1(n13270), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11355) );
  OAI21_X1 U13873 ( .B1(n13270), .B2(P2_REG2_REG_17__SCAN_IN), .A(n11355), 
        .ZN(n13263) );
  OAI21_X1 U13874 ( .B1(n13532), .B2(n11357), .A(n11356), .ZN(n13264) );
  XOR2_X1 U13875 ( .A(n13263), .B(n13264), .Z(n11367) );
  INV_X1 U13876 ( .A(n14857), .ZN(n14825) );
  AOI21_X1 U13877 ( .B1(n11359), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11358), 
        .ZN(n11361) );
  XNOR2_X1 U13878 ( .A(n13270), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11360) );
  NOR2_X1 U13879 ( .A1(n11361), .A2(n11360), .ZN(n13269) );
  AOI211_X1 U13880 ( .C1(n11361), .C2(n11360), .A(n14850), .B(n13269), .ZN(
        n11365) );
  NOR2_X1 U13881 ( .A1(n14862), .A2(n13267), .ZN(n11364) );
  NOR2_X1 U13882 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13141), .ZN(n11363) );
  AND2_X1 U13883 ( .A1(n14855), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n11362) );
  NOR4_X1 U13884 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11366) );
  OAI21_X1 U13885 ( .B1(n11367), .B2(n14825), .A(n11366), .ZN(P2_U3231) );
  NAND2_X1 U13886 ( .A1(n13954), .A2(n12366), .ZN(n11371) );
  OAI21_X1 U13887 ( .B1(n14779), .B2(n10522), .A(n11371), .ZN(n11372) );
  XNOR2_X1 U13888 ( .A(n11372), .B(n12343), .ZN(n11446) );
  OR2_X1 U13889 ( .A1(n14779), .A2(n12305), .ZN(n11374) );
  NAND2_X1 U13890 ( .A1(n10521), .A2(n13954), .ZN(n11373) );
  NAND2_X1 U13891 ( .A1(n11374), .A2(n11373), .ZN(n11443) );
  XNOR2_X1 U13892 ( .A(n11446), .B(n11443), .ZN(n11444) );
  XNOR2_X1 U13893 ( .A(n11445), .B(n11444), .ZN(n11381) );
  INV_X1 U13894 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11375) );
  OAI22_X1 U13895 ( .A1(n13887), .A2(n11376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11375), .ZN(n11379) );
  OAI22_X1 U13896 ( .A1(n11377), .A2(n13903), .B1(n13904), .B2(n11787), .ZN(
        n11378) );
  AOI211_X1 U13897 ( .C1(n11795), .C2(n13936), .A(n11379), .B(n11378), .ZN(
        n11380) );
  OAI21_X1 U13898 ( .B1(n11381), .B2(n13938), .A(n11380), .ZN(P1_U3239) );
  AOI21_X1 U13899 ( .B1(n9324), .B2(n11383), .A(n11538), .ZN(n11401) );
  INV_X1 U13900 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14426) );
  NOR2_X1 U13901 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11384), .ZN(n12554) );
  INV_X1 U13902 ( .A(n12554), .ZN(n11385) );
  OAI21_X1 U13903 ( .B1(n15008), .B2(n14426), .A(n11385), .ZN(n11394) );
  INV_X1 U13904 ( .A(n11386), .ZN(n11387) );
  NOR2_X1 U13905 ( .A1(n11388), .A2(n11387), .ZN(n11391) );
  MUX2_X1 U13906 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14941), .Z(n11546) );
  XNOR2_X1 U13907 ( .A(n11546), .B(n11389), .ZN(n11390) );
  NOR2_X1 U13908 ( .A1(n11391), .A2(n11390), .ZN(n11547) );
  AOI21_X1 U13909 ( .B1(n11391), .B2(n11390), .A(n11547), .ZN(n11392) );
  NOR2_X1 U13910 ( .A1(n11392), .A2(n15017), .ZN(n11393) );
  AOI211_X1 U13911 ( .C1(n14981), .C2(n11549), .A(n11394), .B(n11393), .ZN(
        n11400) );
  AOI21_X1 U13912 ( .B1(n9325), .B2(n11397), .A(n11544), .ZN(n11398) );
  OR2_X1 U13913 ( .A1(n11398), .A2(n15023), .ZN(n11399) );
  OAI211_X1 U13914 ( .C1(n11401), .C2(n15015), .A(n11400), .B(n11399), .ZN(
        P3_U3193) );
  INV_X1 U13915 ( .A(n11402), .ZN(n11403) );
  OAI222_X1 U13916 ( .A1(P3_U3151), .A2(n11404), .B1(n13092), .B2(n15435), 
        .C1(n13089), .C2(n11403), .ZN(P3_U3270) );
  INV_X1 U13917 ( .A(n11405), .ZN(n11409) );
  OAI222_X1 U13918 ( .A1(n13736), .A2(n11407), .B1(n11298), .B2(n11409), .C1(
        n11406), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13919 ( .A1(n8665), .A2(P1_U3086), .B1(n14390), .B2(n11409), .C1(
        n11408), .C2(n14384), .ZN(P1_U3334) );
  XNOR2_X1 U13920 ( .A(n11410), .B(n11413), .ZN(n11411) );
  AOI22_X1 U13921 ( .A1(n13518), .A2(n13224), .B1(n13222), .B2(n13516), .ZN(
        n11564) );
  OAI21_X1 U13922 ( .B1(n11411), .B2(n13562), .A(n11564), .ZN(n11569) );
  INV_X1 U13923 ( .A(n11569), .ZN(n11420) );
  XOR2_X1 U13924 ( .A(n11413), .B(n11412), .Z(n11571) );
  INV_X1 U13925 ( .A(n13565), .ZN(n11414) );
  AOI211_X1 U13926 ( .C1(n11575), .C2(n6957), .A(n9813), .B(n11414), .ZN(
        n11570) );
  NAND2_X1 U13927 ( .A1(n11570), .A2(n13581), .ZN(n11417) );
  INV_X1 U13928 ( .A(n11415), .ZN(n11566) );
  AOI22_X1 U13929 ( .A1(n13552), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11566), 
        .B2(n13544), .ZN(n11416) );
  OAI211_X1 U13930 ( .C1(n11572), .C2(n13486), .A(n11417), .B(n11416), .ZN(
        n11418) );
  AOI21_X1 U13931 ( .B1(n11571), .B2(n13579), .A(n11418), .ZN(n11419) );
  OAI21_X1 U13932 ( .B1(n13552), .B2(n11420), .A(n11419), .ZN(P2_U3252) );
  AOI211_X1 U13933 ( .C1(n14781), .C2(n11423), .A(n11422), .B(n11421), .ZN(
        n11428) );
  INV_X1 U13934 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11424) );
  OAI22_X1 U13935 ( .A1(n11725), .A2(n8752), .B1(n14796), .B2(n11424), .ZN(
        n11425) );
  INV_X1 U13936 ( .A(n11425), .ZN(n11426) );
  OAI21_X1 U13937 ( .B1(n11428), .B2(n14794), .A(n11426), .ZN(P1_U3486) );
  AOI22_X1 U13938 ( .A1(n11810), .A2(n14235), .B1(n14800), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n11427) );
  OAI21_X1 U13939 ( .B1(n11428), .B2(n14800), .A(n11427), .ZN(P1_U3537) );
  INV_X1 U13940 ( .A(n11429), .ZN(n11433) );
  INV_X1 U13941 ( .A(n11430), .ZN(n11432) );
  NOR3_X1 U13942 ( .A1(n11433), .A2(n11432), .A3(n11431), .ZN(n11436) );
  INV_X1 U13943 ( .A(n11434), .ZN(n11435) );
  OAI21_X1 U13944 ( .B1(n11436), .B2(n11435), .A(n14633), .ZN(n11442) );
  OAI22_X1 U13945 ( .A1(n11438), .A2(n13190), .B1(n11437), .B2(n13188), .ZN(
        n11490) );
  NOR2_X1 U13946 ( .A1(n14643), .A2(n13574), .ZN(n11439) );
  AOI211_X1 U13947 ( .C1(n14635), .C2(n11490), .A(n11440), .B(n11439), .ZN(
        n11441) );
  OAI211_X1 U13948 ( .C1(n6955), .C2(n13183), .A(n11442), .B(n11441), .ZN(
        P2_U3196) );
  INV_X1 U13949 ( .A(n11443), .ZN(n11447) );
  NAND2_X1 U13950 ( .A1(n11799), .A2(n12363), .ZN(n11450) );
  NAND2_X1 U13951 ( .A1(n13953), .A2(n12366), .ZN(n11449) );
  NAND2_X1 U13952 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  XNOR2_X1 U13953 ( .A(n11451), .B(n12364), .ZN(n11612) );
  AND2_X1 U13954 ( .A1(n10521), .A2(n13953), .ZN(n11452) );
  AOI21_X1 U13955 ( .B1(n11799), .B2(n12366), .A(n11452), .ZN(n11611) );
  XNOR2_X1 U13956 ( .A(n11612), .B(n11611), .ZN(n11614) );
  XNOR2_X1 U13957 ( .A(n11615), .B(n11614), .ZN(n11460) );
  INV_X1 U13958 ( .A(n11453), .ZN(n11455) );
  OAI21_X1 U13959 ( .B1(n13887), .B2(n11455), .A(n11454), .ZN(n11458) );
  OAI22_X1 U13960 ( .A1(n11719), .A2(n13903), .B1(n13904), .B2(n11456), .ZN(
        n11457) );
  AOI211_X1 U13961 ( .C1(n11799), .C2(n13936), .A(n11458), .B(n11457), .ZN(
        n11459) );
  OAI21_X1 U13962 ( .B1(n11460), .B2(n13938), .A(n11459), .ZN(P1_U3213) );
  INV_X1 U13963 ( .A(n12610), .ZN(n15086) );
  NAND2_X1 U13964 ( .A1(n15086), .A2(n11463), .ZN(n11464) );
  NAND2_X1 U13965 ( .A1(n11465), .A2(n11464), .ZN(n11509) );
  XNOR2_X1 U13966 ( .A(n15078), .B(n12462), .ZN(n11468) );
  XNOR2_X1 U13967 ( .A(n11468), .B(n12609), .ZN(n11510) );
  NAND2_X1 U13968 ( .A1(n11468), .A2(n12609), .ZN(n11469) );
  NAND2_X1 U13969 ( .A1(n11507), .A2(n11469), .ZN(n11470) );
  XNOR2_X1 U13970 ( .A(n15056), .B(n12421), .ZN(n11578) );
  NAND2_X1 U13971 ( .A1(n11470), .A2(n11578), .ZN(n11581) );
  OAI211_X1 U13972 ( .C1(n11470), .C2(n11578), .A(n11581), .B(n14938), .ZN(
        n11475) );
  AND2_X1 U13973 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n14977) );
  OAI22_X1 U13974 ( .A1(n11472), .A2(n12587), .B1(n14935), .B2(n11471), .ZN(
        n11473) );
  AOI211_X1 U13975 ( .C1(n14932), .C2(n15045), .A(n14977), .B(n11473), .ZN(
        n11474) );
  OAI211_X1 U13976 ( .C1(n11476), .C2(n12590), .A(n11475), .B(n11474), .ZN(
        P3_U3153) );
  AOI211_X1 U13977 ( .C1(n14918), .C2(n11479), .A(n11478), .B(n11477), .ZN(
        n11480) );
  OAI21_X1 U13978 ( .B1(n14921), .B2(n11481), .A(n11480), .ZN(n11498) );
  NAND2_X1 U13979 ( .A1(n11498), .A2(n14908), .ZN(n11482) );
  OAI21_X1 U13980 ( .B1(n14908), .B2(n7845), .A(n11482), .ZN(P2_U3463) );
  XNOR2_X1 U13981 ( .A(n11483), .B(n11489), .ZN(n13580) );
  NAND2_X1 U13982 ( .A1(n13578), .A2(n11484), .ZN(n11485) );
  NAND2_X1 U13983 ( .A1(n11485), .A2(n13528), .ZN(n11486) );
  NOR2_X1 U13984 ( .A1(n11487), .A2(n11486), .ZN(n13582) );
  XOR2_X1 U13985 ( .A(n11489), .B(n11488), .Z(n11492) );
  INV_X1 U13986 ( .A(n11490), .ZN(n11491) );
  OAI21_X1 U13987 ( .B1(n11492), .B2(n13562), .A(n11491), .ZN(n13572) );
  AOI211_X1 U13988 ( .C1(n14905), .C2(n13580), .A(n13582), .B(n13572), .ZN(
        n11497) );
  NAND2_X1 U13989 ( .A1(n14931), .A2(n14918), .ZN(n13629) );
  AOI22_X1 U13990 ( .A1(n13578), .A2(n13675), .B1(n14929), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11493) );
  OAI21_X1 U13991 ( .B1(n11497), .B2(n14929), .A(n11493), .ZN(P2_U3511) );
  INV_X1 U13992 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11494) );
  OAI22_X1 U13993 ( .A1(n6955), .A2(n13702), .B1(n14908), .B2(n11494), .ZN(
        n11495) );
  INV_X1 U13994 ( .A(n11495), .ZN(n11496) );
  OAI21_X1 U13995 ( .B1(n11497), .B2(n14924), .A(n11496), .ZN(P2_U3466) );
  NAND2_X1 U13996 ( .A1(n11498), .A2(n14931), .ZN(n11499) );
  OAI21_X1 U13997 ( .B1(n14931), .B2(n11500), .A(n11499), .ZN(P2_U3510) );
  INV_X1 U13998 ( .A(n11501), .ZN(n11503) );
  OAI222_X1 U13999 ( .A1(n11504), .A2(P3_U3151), .B1(n13089), .B2(n11503), 
        .C1(n11502), .C2(n13092), .ZN(P3_U3269) );
  INV_X1 U14000 ( .A(n12608), .ZN(n15072) );
  AOI22_X1 U14001 ( .A1(n12592), .A2(n11505), .B1(n12555), .B2(n12610), .ZN(
        n11506) );
  NAND2_X1 U14002 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14967) );
  OAI211_X1 U14003 ( .C1(n15072), .C2(n12575), .A(n11506), .B(n14967), .ZN(
        n11512) );
  INV_X1 U14004 ( .A(n11507), .ZN(n11508) );
  AOI211_X1 U14005 ( .C1(n11510), .C2(n11509), .A(n12594), .B(n11508), .ZN(
        n11511) );
  AOI211_X1 U14006 ( .C1(n15075), .C2(n12578), .A(n11512), .B(n11511), .ZN(
        n11513) );
  INV_X1 U14007 ( .A(n11513), .ZN(P3_U3179) );
  XNOR2_X1 U14008 ( .A(n13896), .B(n13949), .ZN(n11949) );
  XOR2_X1 U14009 ( .A(n11949), .B(n11514), .Z(n11604) );
  INV_X1 U14010 ( .A(n11604), .ZN(n11522) );
  XNOR2_X1 U14011 ( .A(n11515), .B(n11949), .ZN(n11516) );
  OAI222_X1 U14012 ( .A1(n14210), .A2(n12231), .B1(n11516), .B2(n14110), .C1(
        n14212), .C2(n12219), .ZN(n11602) );
  AOI211_X1 U14013 ( .C1(n13896), .C2(n11526), .A(n14252), .B(n14513), .ZN(
        n11603) );
  NAND2_X1 U14014 ( .A1(n11603), .A2(n14194), .ZN(n11519) );
  AOI22_X1 U14015 ( .A1(n14224), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11517), 
        .B2(n14222), .ZN(n11518) );
  OAI211_X1 U14016 ( .C1(n11607), .C2(n14525), .A(n11519), .B(n11518), .ZN(
        n11520) );
  AOI21_X1 U14017 ( .B1(n11602), .B2(n14529), .A(n11520), .ZN(n11521) );
  OAI21_X1 U14018 ( .B1(n14201), .B2(n11522), .A(n11521), .ZN(P1_U3282) );
  OAI21_X1 U14019 ( .B1(n11524), .B2(n11947), .A(n11523), .ZN(n14792) );
  AOI21_X1 U14020 ( .B1(n11525), .B2(n13768), .A(n14252), .ZN(n11527) );
  AOI22_X1 U14021 ( .A1(n11527), .A2(n11526), .B1(n14172), .B2(n13949), .ZN(
        n14787) );
  AOI22_X1 U14022 ( .A1(n14224), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n13777), 
        .B2(n14222), .ZN(n11529) );
  NAND2_X1 U14023 ( .A1(n13768), .A2(n14225), .ZN(n11528) );
  OAI211_X1 U14024 ( .C1(n14787), .C2(n14516), .A(n11529), .B(n11528), .ZN(
        n11535) );
  INV_X1 U14025 ( .A(n11530), .ZN(n11531) );
  AOI211_X1 U14026 ( .C1(n11947), .C2(n11532), .A(n14110), .B(n11531), .ZN(
        n14790) );
  INV_X1 U14027 ( .A(n14790), .ZN(n11533) );
  NAND2_X1 U14028 ( .A1(n13951), .A2(n14174), .ZN(n14786) );
  AOI21_X1 U14029 ( .B1(n11533), .B2(n14786), .A(n14224), .ZN(n11534) );
  AOI211_X1 U14030 ( .C1(n14233), .C2(n14792), .A(n11535), .B(n11534), .ZN(
        n11536) );
  INV_X1 U14031 ( .A(n11536), .ZN(P1_U3283) );
  NOR2_X1 U14032 ( .A1(n11549), .A2(n11537), .ZN(n11539) );
  NAND2_X1 U14033 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12619), .ZN(n11540) );
  OAI21_X1 U14034 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12619), .A(n11540), 
        .ZN(n11541) );
  AOI21_X1 U14035 ( .B1(n11542), .B2(n11541), .A(n12613), .ZN(n11558) );
  NAND2_X1 U14036 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12619), .ZN(n11545) );
  OAI21_X1 U14037 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12619), .A(n11545), 
        .ZN(n12617) );
  XNOR2_X1 U14038 ( .A(n12618), .B(n12617), .ZN(n11556) );
  INV_X1 U14039 ( .A(n11546), .ZN(n11548) );
  AOI21_X1 U14040 ( .B1(n11549), .B2(n11548), .A(n11547), .ZN(n11551) );
  MUX2_X1 U14041 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14941), .Z(n12622) );
  XNOR2_X1 U14042 ( .A(n12622), .B(n12625), .ZN(n11550) );
  NAND2_X1 U14043 ( .A1(n11551), .A2(n11550), .ZN(n12623) );
  OAI211_X1 U14044 ( .C1(n11551), .C2(n11550), .A(n12623), .B(n14999), .ZN(
        n11554) );
  INV_X1 U14045 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11552) );
  NOR2_X1 U14046 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11552), .ZN(n12487) );
  AOI21_X1 U14047 ( .B1(n14978), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12487), 
        .ZN(n11553) );
  OAI211_X1 U14048 ( .C1(n15007), .C2(n12619), .A(n11554), .B(n11553), .ZN(
        n11555) );
  AOI21_X1 U14049 ( .B1(n12732), .B2(n11556), .A(n11555), .ZN(n11557) );
  OAI21_X1 U14050 ( .B1(n11558), .B2(n15015), .A(n11557), .ZN(P3_U3194) );
  AOI21_X1 U14051 ( .B1(n11560), .B2(n11559), .A(n13202), .ZN(n11562) );
  NAND2_X1 U14052 ( .A1(n11562), .A2(n11561), .ZN(n11568) );
  OAI22_X1 U14053 ( .A1(n13178), .A2(n11564), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11563), .ZN(n11565) );
  AOI21_X1 U14054 ( .B1(n11566), .B2(n9845), .A(n11565), .ZN(n11567) );
  OAI211_X1 U14055 ( .C1(n11572), .C2(n13183), .A(n11568), .B(n11567), .ZN(
        P2_U3206) );
  AOI211_X1 U14056 ( .C1(n11571), .C2(n14905), .A(n11570), .B(n11569), .ZN(
        n11577) );
  OAI22_X1 U14057 ( .A1(n11572), .A2(n13702), .B1(n14908), .B2(n7881), .ZN(
        n11573) );
  INV_X1 U14058 ( .A(n11573), .ZN(n11574) );
  OAI21_X1 U14059 ( .B1(n11577), .B2(n14924), .A(n11574), .ZN(P2_U3469) );
  AOI22_X1 U14060 ( .A1(n11575), .A2(n13675), .B1(n14929), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11576) );
  OAI21_X1 U14061 ( .B1(n11577), .B2(n14929), .A(n11576), .ZN(P2_U3512) );
  INV_X1 U14062 ( .A(n11578), .ZN(n11579) );
  NAND2_X1 U14063 ( .A1(n11579), .A2(n12608), .ZN(n11580) );
  NAND2_X1 U14064 ( .A1(n11581), .A2(n11580), .ZN(n11583) );
  XNOR2_X1 U14065 ( .A(n15066), .B(n12462), .ZN(n11677) );
  XNOR2_X1 U14066 ( .A(n11677), .B(n15045), .ZN(n11582) );
  NAND2_X1 U14067 ( .A1(n11583), .A2(n11582), .ZN(n11680) );
  OAI211_X1 U14068 ( .C1(n11583), .C2(n11582), .A(n11680), .B(n14938), .ZN(
        n11587) );
  NAND2_X1 U14069 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15001) );
  INV_X1 U14070 ( .A(n15001), .ZN(n11585) );
  OAI22_X1 U14071 ( .A1(n15072), .A2(n12587), .B1(n14935), .B2(n12046), .ZN(
        n11584) );
  AOI211_X1 U14072 ( .C1(n14932), .C2(n12607), .A(n11585), .B(n11584), .ZN(
        n11586) );
  OAI211_X1 U14073 ( .C1(n12590), .C2(n15067), .A(n11587), .B(n11586), .ZN(
        P3_U3161) );
  INV_X1 U14074 ( .A(n11588), .ZN(n11590) );
  OAI222_X1 U14075 ( .A1(n13089), .A2(n11590), .B1(n13092), .B2(n11589), .C1(
        P3_U3151), .C2(n6550), .ZN(P3_U3268) );
  NAND2_X1 U14076 ( .A1(n11591), .A2(n15025), .ZN(n15064) );
  NAND2_X1 U14077 ( .A1(n15129), .A2(n15064), .ZN(n12869) );
  NAND2_X1 U14078 ( .A1(n14597), .A2(n12059), .ZN(n11592) );
  INV_X1 U14079 ( .A(n11593), .ZN(n12169) );
  XNOR2_X1 U14080 ( .A(n11592), .B(n12169), .ZN(n14612) );
  INV_X1 U14081 ( .A(n11594), .ZN(n11595) );
  OR2_X1 U14082 ( .A1(n11594), .A2(n11593), .ZN(n14587) );
  OAI211_X1 U14083 ( .C1(n11595), .C2(n12169), .A(n15039), .B(n14587), .ZN(
        n11597) );
  AOI22_X1 U14084 ( .A1(n15046), .A2(n12606), .B1(n12604), .B2(n15043), .ZN(
        n11596) );
  NAND2_X1 U14085 ( .A1(n11597), .A2(n11596), .ZN(n14614) );
  NAND2_X1 U14086 ( .A1(n14614), .A2(n15129), .ZN(n11601) );
  OAI22_X1 U14087 ( .A1(n15129), .A2(n11598), .B1(n12485), .B2(n15101), .ZN(
        n11599) );
  AOI21_X1 U14088 ( .B1(n12889), .B2(n12491), .A(n11599), .ZN(n11600) );
  OAI211_X1 U14089 ( .C1(n12869), .C2(n14612), .A(n11601), .B(n11600), .ZN(
        P3_U3221) );
  AOI211_X1 U14090 ( .C1(n11604), .C2(n14793), .A(n11603), .B(n11602), .ZN(
        n11610) );
  AOI22_X1 U14091 ( .A1(n13896), .A2(n14235), .B1(n14800), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11605) );
  OAI21_X1 U14092 ( .B1(n11610), .B2(n14800), .A(n11605), .ZN(P1_U3539) );
  INV_X1 U14093 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11606) );
  OAI22_X1 U14094 ( .A1(n11607), .A2(n8752), .B1(n14796), .B2(n11606), .ZN(
        n11608) );
  INV_X1 U14095 ( .A(n11608), .ZN(n11609) );
  OAI21_X1 U14096 ( .B1(n11610), .B2(n14794), .A(n11609), .ZN(P1_U3492) );
  INV_X1 U14097 ( .A(n11611), .ZN(n11613) );
  NAND2_X1 U14098 ( .A1(n11806), .A2(n12363), .ZN(n11617) );
  OR2_X1 U14099 ( .A1(n11719), .A2(n12305), .ZN(n11616) );
  NAND2_X1 U14100 ( .A1(n11617), .A2(n11616), .ZN(n11618) );
  XNOR2_X1 U14101 ( .A(n11618), .B(n12343), .ZN(n11621) );
  INV_X1 U14102 ( .A(n11621), .ZN(n11623) );
  NOR2_X1 U14103 ( .A1(n11719), .A2(n12345), .ZN(n11619) );
  AOI21_X1 U14104 ( .B1(n11806), .B2(n12366), .A(n11619), .ZN(n11620) );
  INV_X1 U14105 ( .A(n11620), .ZN(n11622) );
  AND2_X1 U14106 ( .A1(n11621), .A2(n11620), .ZN(n11711) );
  AOI21_X1 U14107 ( .B1(n11623), .B2(n11622), .A(n11711), .ZN(n11624) );
  OAI21_X1 U14108 ( .B1(n6694), .B2(n11624), .A(n11712), .ZN(n11625) );
  NAND2_X1 U14109 ( .A1(n11625), .A2(n13912), .ZN(n11631) );
  INV_X1 U14110 ( .A(n13795), .ZN(n13934) );
  OAI21_X1 U14111 ( .B1(n11627), .B2(n13934), .A(n11626), .ZN(n11628) );
  AOI21_X1 U14112 ( .B1(n11629), .B2(n13932), .A(n11628), .ZN(n11630) );
  OAI211_X1 U14113 ( .C1(n11632), .C2(n13921), .A(n11631), .B(n11630), .ZN(
        P1_U3221) );
  NAND2_X1 U14114 ( .A1(n11636), .A2(n11633), .ZN(n11634) );
  OAI211_X1 U14115 ( .C1(n11635), .C2(n14384), .A(n11634), .B(n11982), .ZN(
        P1_U3332) );
  NAND2_X1 U14116 ( .A1(n11636), .A2(n13727), .ZN(n11638) );
  OAI211_X1 U14117 ( .C1(n11639), .C2(n13736), .A(n11638), .B(n11637), .ZN(
        P2_U3304) );
  INV_X1 U14118 ( .A(n11640), .ZN(n11644) );
  INV_X1 U14119 ( .A(n11641), .ZN(n11642) );
  OAI222_X1 U14120 ( .A1(n13736), .A2(n15371), .B1(n11298), .B2(n11644), .C1(
        n11642), .C2(P2_U3088), .ZN(P2_U3303) );
  OAI222_X1 U14121 ( .A1(P1_U3086), .A2(n11645), .B1(n14390), .B2(n11644), 
        .C1(n11643), .C2(n14384), .ZN(P1_U3331) );
  XNOR2_X1 U14122 ( .A(n11646), .B(n7193), .ZN(n14648) );
  INV_X1 U14123 ( .A(n14648), .ZN(n11656) );
  OAI211_X1 U14124 ( .C1(n11648), .C2(n11951), .A(n11647), .B(n14522), .ZN(
        n11651) );
  OR2_X1 U14125 ( .A1(n13929), .A2(n14210), .ZN(n11650) );
  OR2_X1 U14126 ( .A1(n12231), .A2(n14212), .ZN(n11649) );
  AND2_X1 U14127 ( .A1(n11650), .A2(n11649), .ZN(n13866) );
  NAND2_X1 U14128 ( .A1(n11651), .A2(n13866), .ZN(n14646) );
  OAI211_X1 U14129 ( .C1(n14514), .C2(n14645), .A(n14512), .B(n11693), .ZN(
        n14644) );
  AOI22_X1 U14130 ( .A1(n14224), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n13864), 
        .B2(n14222), .ZN(n11653) );
  NAND2_X1 U14131 ( .A1(n13868), .A2(n14225), .ZN(n11652) );
  OAI211_X1 U14132 ( .C1(n14644), .C2(n14516), .A(n11653), .B(n11652), .ZN(
        n11654) );
  AOI21_X1 U14133 ( .B1(n14646), .B2(n14529), .A(n11654), .ZN(n11655) );
  OAI21_X1 U14134 ( .B1(n14201), .B2(n11656), .A(n11655), .ZN(P1_U3280) );
  OAI21_X1 U14135 ( .B1(n11658), .B2(n11657), .A(n13201), .ZN(n11659) );
  NAND2_X1 U14136 ( .A1(n11659), .A2(n14633), .ZN(n11663) );
  INV_X1 U14137 ( .A(n13555), .ZN(n11661) );
  AOI22_X1 U14138 ( .A1(n13519), .A2(n13516), .B1(n13223), .B2(n13518), .ZN(
        n13561) );
  OAI22_X1 U14139 ( .A1(n13178), .A2(n13561), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7900), .ZN(n11660) );
  AOI21_X1 U14140 ( .B1(n11661), .B2(n9845), .A(n11660), .ZN(n11662) );
  OAI211_X1 U14141 ( .C1(n7242), .C2(n13183), .A(n11663), .B(n11662), .ZN(
        P2_U3187) );
  XNOR2_X1 U14142 ( .A(n11664), .B(n6976), .ZN(n11665) );
  AOI222_X1 U14143 ( .A1(n15039), .A2(n11665), .B1(n12602), .B2(n15043), .C1(
        n12604), .C2(n15046), .ZN(n13005) );
  OAI22_X1 U14144 ( .A1(n15129), .A2(n11666), .B1(n12442), .B2(n15101), .ZN(
        n11667) );
  AOI21_X1 U14145 ( .B1(n13002), .B2(n12889), .A(n11667), .ZN(n11670) );
  XNOR2_X1 U14146 ( .A(n11668), .B(n12168), .ZN(n13003) );
  NAND2_X1 U14147 ( .A1(n13003), .A2(n15079), .ZN(n11669) );
  OAI211_X1 U14148 ( .C1(n13005), .C2(n15038), .A(n11670), .B(n11669), .ZN(
        P3_U3219) );
  INV_X1 U14149 ( .A(n11671), .ZN(n11675) );
  OAI222_X1 U14150 ( .A1(P1_U3086), .A2(n11673), .B1(n14390), .B2(n11675), 
        .C1(n11672), .C2(n14384), .ZN(P1_U3330) );
  OAI222_X1 U14151 ( .A1(n13736), .A2(n11676), .B1(n11298), .B2(n11675), .C1(
        n11674), .C2(P2_U3088), .ZN(P2_U3302) );
  XNOR2_X1 U14152 ( .A(n15052), .B(n12462), .ZN(n11700) );
  XNOR2_X1 U14153 ( .A(n11700), .B(n12607), .ZN(n11683) );
  INV_X1 U14154 ( .A(n11677), .ZN(n11678) );
  NAND2_X1 U14155 ( .A1(n11678), .A2(n15045), .ZN(n11679) );
  NAND2_X1 U14156 ( .A1(n11680), .A2(n11679), .ZN(n11682) );
  INV_X1 U14157 ( .A(n11703), .ZN(n11681) );
  AOI21_X1 U14158 ( .B1(n11683), .B2(n11682), .A(n11681), .ZN(n11689) );
  OAI22_X1 U14159 ( .A1(n11684), .A2(n12587), .B1(n14935), .B2(n15052), .ZN(
        n11685) );
  AOI211_X1 U14160 ( .C1(n14932), .C2(n15044), .A(n11686), .B(n11685), .ZN(
        n11688) );
  NAND2_X1 U14161 ( .A1(n12578), .A2(n15049), .ZN(n11687) );
  OAI211_X1 U14162 ( .C1(n11689), .C2(n12594), .A(n11688), .B(n11687), .ZN(
        P3_U3171) );
  XNOR2_X1 U14163 ( .A(n11690), .B(n7588), .ZN(n11691) );
  AOI222_X1 U14164 ( .A1(n13947), .A2(n14174), .B1(n13945), .B2(n14172), .C1(
        n14522), .C2(n11691), .ZN(n14335) );
  INV_X1 U14165 ( .A(n14220), .ZN(n11692) );
  AOI211_X1 U14166 ( .C1(n14329), .C2(n11693), .A(n14252), .B(n11692), .ZN(
        n14328) );
  INV_X1 U14167 ( .A(n14329), .ZN(n11695) );
  AOI22_X1 U14168 ( .A1(n14224), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n13749), 
        .B2(n14222), .ZN(n11694) );
  OAI21_X1 U14169 ( .B1(n11695), .B2(n14525), .A(n11694), .ZN(n11696) );
  AOI21_X1 U14170 ( .B1(n14328), .B2(n14194), .A(n11696), .ZN(n11699) );
  NAND2_X1 U14171 ( .A1(n11697), .A2(n11835), .ZN(n14331) );
  NAND3_X1 U14172 ( .A1(n14332), .A2(n14331), .A3(n14233), .ZN(n11698) );
  OAI211_X1 U14173 ( .C1(n14335), .C2(n14224), .A(n11699), .B(n11698), .ZN(
        P1_U3279) );
  INV_X1 U14174 ( .A(n12607), .ZN(n15063) );
  INV_X1 U14175 ( .A(n11700), .ZN(n11701) );
  NAND2_X1 U14176 ( .A1(n15063), .A2(n11701), .ZN(n11702) );
  XNOR2_X1 U14177 ( .A(n15033), .B(n12421), .ZN(n12387) );
  XNOR2_X1 U14178 ( .A(n12387), .B(n15044), .ZN(n11704) );
  OAI211_X1 U14179 ( .C1(n11705), .C2(n11704), .A(n12390), .B(n14938), .ZN(
        n11709) );
  OAI22_X1 U14180 ( .A1(n15063), .A2(n12587), .B1(n14935), .B2(n15033), .ZN(
        n11706) );
  AOI211_X1 U14181 ( .C1(n14932), .C2(n12606), .A(n11707), .B(n11706), .ZN(
        n11708) );
  OAI211_X1 U14182 ( .C1(n15034), .C2(n12590), .A(n11709), .B(n11708), .ZN(
        P3_U3157) );
  OAI22_X1 U14183 ( .A1(n11725), .A2(n10522), .B1(n13774), .B2(n12305), .ZN(
        n11710) );
  XOR2_X1 U14184 ( .A(n12364), .B(n11710), .Z(n11716) );
  NAND2_X1 U14185 ( .A1(n11810), .A2(n12366), .ZN(n11714) );
  OR2_X1 U14186 ( .A1(n13774), .A2(n12345), .ZN(n11713) );
  NAND2_X1 U14187 ( .A1(n11714), .A2(n11713), .ZN(n12216) );
  NAND2_X1 U14188 ( .A1(n11715), .A2(n11716), .ZN(n12222) );
  OAI21_X1 U14189 ( .B1(n11716), .B2(n11715), .A(n12222), .ZN(n11717) );
  NAND2_X1 U14190 ( .A1(n11717), .A2(n13912), .ZN(n11724) );
  INV_X1 U14191 ( .A(n11718), .ZN(n11721) );
  OAI22_X1 U14192 ( .A1(n12219), .A2(n13903), .B1(n13904), .B2(n11719), .ZN(
        n11720) );
  AOI211_X1 U14193 ( .C1(n11722), .C2(n13932), .A(n11721), .B(n11720), .ZN(
        n11723) );
  OAI211_X1 U14194 ( .C1(n11725), .C2(n13921), .A(n11724), .B(n11723), .ZN(
        P1_U3231) );
  INV_X1 U14195 ( .A(n13728), .ZN(n11727) );
  INV_X1 U14196 ( .A(n11728), .ZN(n11729) );
  OAI222_X1 U14197 ( .A1(n13092), .A2(n11730), .B1(n13089), .B2(n11729), .C1(
        n9623), .C2(P3_U3151), .ZN(P3_U3267) );
  INV_X1 U14198 ( .A(n11731), .ZN(n11733) );
  OAI222_X1 U14199 ( .A1(n13736), .A2(n11734), .B1(n11298), .B2(n11733), .C1(
        n11732), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14200 ( .A1(n14857), .A2(n11737), .ZN(n11735) );
  OAI211_X1 U14201 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14850), .A(n11735), .B(
        n14862), .ZN(n11739) );
  OAI22_X1 U14202 ( .A1(n14825), .A2(n11737), .B1(n11736), .B2(n14850), .ZN(
        n11738) );
  MUX2_X1 U14203 ( .A(n11739), .B(n11738), .S(n7656), .Z(n11743) );
  INV_X1 U14204 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n11741) );
  OAI22_X1 U14205 ( .A1(n14848), .A2(n11741), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11740), .ZN(n11742) );
  OR2_X1 U14206 ( .A1(n11743), .A2(n11742), .ZN(P2_U3214) );
  AOI21_X1 U14207 ( .B1(n13581), .B2(n11744), .A(n13577), .ZN(n11753) );
  INV_X1 U14208 ( .A(n11745), .ZN(n11750) );
  INV_X1 U14209 ( .A(n13395), .ZN(n11749) );
  AOI22_X1 U14210 ( .A1(n13557), .A2(n11746), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13544), .ZN(n11747) );
  OAI21_X1 U14211 ( .B1(n11737), .B2(n13557), .A(n11747), .ZN(n11748) );
  AOI21_X1 U14212 ( .B1(n11750), .B2(n11749), .A(n11748), .ZN(n11751) );
  OAI21_X1 U14213 ( .B1(n11753), .B2(n11752), .A(n11751), .ZN(P2_U3265) );
  INV_X1 U14214 ( .A(n13074), .ZN(n11754) );
  AOI22_X1 U14215 ( .A1(n11754), .A2(n11756), .B1(n15169), .B2(
        P3_REG0_REG_0__SCAN_IN), .ZN(n11755) );
  OAI21_X1 U14216 ( .B1(n11758), .B2(n15169), .A(n11755), .ZN(P3_U3390) );
  AOI22_X1 U14217 ( .A1(n12938), .A2(n11756), .B1(n15179), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n11757) );
  OAI21_X1 U14218 ( .B1(n11758), .B2(n15179), .A(n11757), .ZN(P3_U3459) );
  INV_X1 U14219 ( .A(n11759), .ZN(n11938) );
  XNOR2_X1 U14220 ( .A(n11760), .B(n11924), .ZN(n11908) );
  XNOR2_X1 U14221 ( .A(n11761), .B(n11921), .ZN(n11762) );
  OAI211_X1 U14222 ( .C1(n11935), .C2(n10282), .A(n11938), .B(n11762), .ZN(
        n11768) );
  NAND2_X1 U14223 ( .A1(n11768), .A2(n11767), .ZN(n11769) );
  NAND2_X1 U14224 ( .A1(n11769), .A2(n8335), .ZN(n11775) );
  NAND2_X1 U14225 ( .A1(n11921), .A2(n11770), .ZN(n11773) );
  NAND2_X1 U14226 ( .A1(n11911), .A2(n11771), .ZN(n11772) );
  NAND2_X1 U14227 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  NAND2_X1 U14228 ( .A1(n11775), .A2(n7608), .ZN(n11781) );
  MUX2_X1 U14229 ( .A(n11777), .B(n11776), .S(n11911), .Z(n11780) );
  OAI21_X1 U14230 ( .B1(n14774), .B2(n11782), .A(n11778), .ZN(n11779) );
  NAND3_X1 U14231 ( .A1(n11781), .A2(n11780), .A3(n11779), .ZN(n11786) );
  AOI21_X1 U14232 ( .B1(n11782), .B2(n11911), .A(n14774), .ZN(n11785) );
  AOI21_X1 U14233 ( .B1(n13956), .B2(n11921), .A(n11783), .ZN(n11784) );
  MUX2_X1 U14234 ( .A(n11788), .B(n11787), .S(n11911), .Z(n11791) );
  MUX2_X1 U14235 ( .A(n13955), .B(n11789), .S(n11911), .Z(n11790) );
  OAI21_X1 U14236 ( .B1(n11792), .B2(n11791), .A(n11790), .ZN(n11794) );
  NAND2_X1 U14237 ( .A1(n11792), .A2(n11791), .ZN(n11793) );
  MUX2_X1 U14238 ( .A(n13954), .B(n11795), .S(n11911), .Z(n11797) );
  MUX2_X1 U14239 ( .A(n13954), .B(n11795), .S(n11921), .Z(n11796) );
  INV_X1 U14240 ( .A(n11797), .ZN(n11798) );
  MUX2_X1 U14241 ( .A(n13953), .B(n11799), .S(n11921), .Z(n11802) );
  NAND2_X1 U14242 ( .A1(n11803), .A2(n11802), .ZN(n11801) );
  MUX2_X1 U14243 ( .A(n13953), .B(n11799), .S(n11911), .Z(n11800) );
  NAND2_X1 U14244 ( .A1(n11801), .A2(n11800), .ZN(n11805) );
  NAND2_X1 U14245 ( .A1(n11805), .A2(n11804), .ZN(n11809) );
  MUX2_X1 U14246 ( .A(n13952), .B(n11806), .S(n11911), .Z(n11808) );
  MUX2_X1 U14247 ( .A(n11806), .B(n13952), .S(n11911), .Z(n11807) );
  MUX2_X1 U14248 ( .A(n13951), .B(n11810), .S(n11921), .Z(n11814) );
  NAND2_X1 U14249 ( .A1(n11813), .A2(n11814), .ZN(n11812) );
  MUX2_X1 U14250 ( .A(n13951), .B(n11810), .S(n11911), .Z(n11811) );
  NAND2_X1 U14251 ( .A1(n11812), .A2(n11811), .ZN(n11818) );
  INV_X1 U14252 ( .A(n11814), .ZN(n11815) );
  NAND2_X1 U14253 ( .A1(n11816), .A2(n11815), .ZN(n11817) );
  MUX2_X1 U14254 ( .A(n13950), .B(n13768), .S(n11911), .Z(n11820) );
  MUX2_X1 U14255 ( .A(n13950), .B(n13768), .S(n11921), .Z(n11819) );
  INV_X1 U14256 ( .A(n11820), .ZN(n11821) );
  MUX2_X1 U14257 ( .A(n13949), .B(n13896), .S(n11921), .Z(n11824) );
  NAND2_X1 U14258 ( .A1(n11825), .A2(n11824), .ZN(n11823) );
  MUX2_X1 U14259 ( .A(n13949), .B(n13896), .S(n11911), .Z(n11822) );
  NAND2_X1 U14260 ( .A1(n11823), .A2(n11822), .ZN(n11827) );
  MUX2_X1 U14261 ( .A(n13948), .B(n12233), .S(n11911), .Z(n11829) );
  MUX2_X1 U14262 ( .A(n13948), .B(n12233), .S(n11921), .Z(n11828) );
  INV_X1 U14263 ( .A(n11829), .ZN(n11830) );
  MUX2_X1 U14264 ( .A(n13947), .B(n13868), .S(n11921), .Z(n11833) );
  MUX2_X1 U14265 ( .A(n13947), .B(n13868), .S(n11911), .Z(n11831) );
  INV_X1 U14266 ( .A(n11831), .ZN(n11832) );
  NAND2_X1 U14267 ( .A1(n11834), .A2(n11833), .ZN(n11836) );
  NAND2_X1 U14268 ( .A1(n11844), .A2(n6601), .ZN(n11840) );
  NAND2_X1 U14269 ( .A1(n11843), .A2(n11838), .ZN(n11839) );
  MUX2_X1 U14270 ( .A(n11840), .B(n11839), .S(n11911), .Z(n11841) );
  INV_X1 U14271 ( .A(n11841), .ZN(n11842) );
  MUX2_X1 U14272 ( .A(n11844), .B(n11843), .S(n11921), .Z(n11845) );
  MUX2_X1 U14273 ( .A(n13928), .B(n14365), .S(n11921), .Z(n11855) );
  NAND2_X1 U14274 ( .A1(n14310), .A2(n14211), .ZN(n11848) );
  NOR2_X1 U14275 ( .A1(n13928), .A2(n11911), .ZN(n11846) );
  AOI21_X1 U14276 ( .B1(n14206), .B2(n11911), .A(n11846), .ZN(n11847) );
  NAND3_X1 U14277 ( .A1(n11849), .A2(n11848), .A3(n11847), .ZN(n11856) );
  OAI21_X1 U14278 ( .B1(n11850), .B2(n11855), .A(n11856), .ZN(n11851) );
  NOR2_X1 U14279 ( .A1(n14211), .A2(n11921), .ZN(n11853) );
  OAI21_X1 U14280 ( .B1(n11911), .B2(n14175), .A(n14310), .ZN(n11852) );
  OAI21_X1 U14281 ( .B1(n11853), .B2(n14310), .A(n11852), .ZN(n11854) );
  OAI21_X1 U14282 ( .B1(n11856), .B2(n11855), .A(n11854), .ZN(n11857) );
  INV_X1 U14283 ( .A(n11857), .ZN(n11858) );
  NAND2_X1 U14284 ( .A1(n11859), .A2(n11858), .ZN(n11862) );
  XNOR2_X1 U14285 ( .A(n14163), .B(n11911), .ZN(n11861) );
  XNOR2_X1 U14286 ( .A(n14304), .B(n11921), .ZN(n11860) );
  NAND2_X1 U14287 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  OR2_X1 U14288 ( .A1(n14298), .A2(n13902), .ZN(n11866) );
  MUX2_X1 U14289 ( .A(n11866), .B(n11865), .S(n11911), .Z(n11867) );
  MUX2_X1 U14290 ( .A(n13785), .B(n8663), .S(n11921), .Z(n11869) );
  MUX2_X1 U14291 ( .A(n14164), .B(n14292), .S(n11911), .Z(n11868) );
  MUX2_X1 U14292 ( .A(n14140), .B(n14288), .S(n11911), .Z(n11871) );
  MUX2_X1 U14293 ( .A(n14140), .B(n14288), .S(n11921), .Z(n11870) );
  INV_X1 U14294 ( .A(n11871), .ZN(n11872) );
  INV_X1 U14295 ( .A(n13882), .ZN(n14284) );
  MUX2_X1 U14296 ( .A(n14092), .B(n14284), .S(n11921), .Z(n11875) );
  MUX2_X1 U14297 ( .A(n13763), .B(n13882), .S(n11911), .Z(n11873) );
  AOI21_X1 U14298 ( .B1(n11876), .B2(n11875), .A(n11873), .ZN(n11874) );
  NOR2_X1 U14299 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  MUX2_X1 U14300 ( .A(n14072), .B(n14276), .S(n11911), .Z(n11878) );
  MUX2_X1 U14301 ( .A(n14072), .B(n14276), .S(n11921), .Z(n11879) );
  MUX2_X1 U14302 ( .A(n14093), .B(n14266), .S(n11921), .Z(n11882) );
  MUX2_X1 U14303 ( .A(n14093), .B(n14266), .S(n11911), .Z(n11880) );
  NAND2_X1 U14304 ( .A1(n11881), .A2(n11880), .ZN(n11884) );
  MUX2_X1 U14305 ( .A(n14071), .B(n14259), .S(n11911), .Z(n11887) );
  MUX2_X1 U14306 ( .A(n14071), .B(n14259), .S(n11921), .Z(n11885) );
  INV_X1 U14307 ( .A(n11887), .ZN(n11888) );
  MUX2_X1 U14308 ( .A(n14053), .B(n12347), .S(n11921), .Z(n11890) );
  MUX2_X1 U14309 ( .A(n14053), .B(n12347), .S(n11911), .Z(n11889) );
  INV_X1 U14310 ( .A(n11890), .ZN(n11891) );
  MUX2_X1 U14311 ( .A(n13943), .B(n14248), .S(n11911), .Z(n11895) );
  MUX2_X1 U14312 ( .A(n13943), .B(n14248), .S(n11921), .Z(n11892) );
  NAND2_X1 U14313 ( .A1(n11893), .A2(n11892), .ZN(n11899) );
  INV_X1 U14314 ( .A(n11894), .ZN(n11897) );
  INV_X1 U14315 ( .A(n11895), .ZN(n11896) );
  NAND2_X1 U14316 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NAND2_X1 U14317 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  MUX2_X1 U14318 ( .A(n13942), .B(n14243), .S(n11921), .Z(n11901) );
  MUX2_X1 U14319 ( .A(n13942), .B(n14243), .S(n11911), .Z(n11902) );
  NAND2_X1 U14320 ( .A1(n8668), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U14321 ( .A1(n8669), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U14322 ( .A1(n11903), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11904) );
  OAI21_X1 U14323 ( .B1(n13999), .B2(n11925), .A(n13940), .ZN(n11907) );
  INV_X1 U14324 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14378) );
  MUX2_X1 U14325 ( .A(n11907), .B(n14344), .S(n11911), .Z(n11915) );
  INV_X1 U14326 ( .A(n13940), .ZN(n11910) );
  NOR2_X1 U14327 ( .A1(n11920), .A2(n11921), .ZN(n11922) );
  AOI21_X1 U14328 ( .B1(n11908), .B2(n8665), .A(n11922), .ZN(n11909) );
  OAI22_X1 U14329 ( .A1(n14344), .A2(n11911), .B1(n11910), .B2(n11909), .ZN(
        n11916) );
  INV_X1 U14330 ( .A(n12371), .ZN(n13941) );
  MUX2_X1 U14331 ( .A(n11912), .B(n13941), .S(n11911), .Z(n11913) );
  INV_X1 U14332 ( .A(n11915), .ZN(n11918) );
  INV_X1 U14333 ( .A(n11916), .ZN(n11917) );
  INV_X1 U14334 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12000) );
  NOR2_X1 U14335 ( .A1(n8356), .A2(n12000), .ZN(n11919) );
  MUX2_X1 U14336 ( .A(n11921), .B(n11920), .S(n14340), .Z(n11923) );
  AND2_X1 U14337 ( .A1(n11925), .A2(n11924), .ZN(n11927) );
  OAI21_X1 U14338 ( .B1(n11928), .B2(n11927), .A(n11926), .ZN(n11970) );
  NAND2_X1 U14339 ( .A1(n8665), .A2(n11929), .ZN(n11973) );
  NAND2_X1 U14340 ( .A1(n11970), .A2(n11973), .ZN(n11966) );
  NOR3_X1 U14341 ( .A1(n11932), .A2(n11969), .A3(n11966), .ZN(n11977) );
  XNOR2_X1 U14342 ( .A(n14340), .B(n13999), .ZN(n11968) );
  INV_X1 U14343 ( .A(n11968), .ZN(n11931) );
  INV_X1 U14344 ( .A(n11970), .ZN(n11930) );
  INV_X1 U14345 ( .A(n14344), .ZN(n11933) );
  XOR2_X1 U14346 ( .A(n13940), .B(n11933), .Z(n11964) );
  INV_X1 U14347 ( .A(n14129), .ZN(n14120) );
  NOR2_X1 U14348 ( .A1(n11935), .A2(n11934), .ZN(n11939) );
  NAND4_X1 U14349 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11941) );
  NOR2_X1 U14350 ( .A1(n11941), .A2(n11940), .ZN(n11943) );
  NAND4_X1 U14351 ( .A1(n8411), .A2(n11944), .A3(n11943), .A4(n11942), .ZN(
        n11945) );
  OR3_X1 U14352 ( .A1(n11947), .A2(n11946), .A3(n11945), .ZN(n11948) );
  NOR2_X1 U14353 ( .A1(n14519), .A2(n11948), .ZN(n11950) );
  NAND3_X1 U14354 ( .A1(n11951), .A2(n11950), .A3(n11949), .ZN(n11952) );
  NOR3_X1 U14355 ( .A1(n11953), .A2(n7588), .A3(n11952), .ZN(n11954) );
  NAND4_X1 U14356 ( .A1(n14182), .A2(n14189), .A3(n11954), .A4(n7183), .ZN(
        n11955) );
  NOR4_X1 U14357 ( .A1(n14120), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11958) );
  NAND4_X1 U14358 ( .A1(n8593), .A2(n8571), .A3(n11958), .A4(n14100), .ZN(
        n11959) );
  NOR3_X1 U14359 ( .A1(n14041), .A2(n11960), .A3(n11959), .ZN(n11961) );
  NAND4_X1 U14360 ( .A1(n11962), .A2(n11961), .A3(n14010), .A4(n14034), .ZN(
        n11963) );
  XNOR2_X1 U14361 ( .A(n11965), .B(n11760), .ZN(n11974) );
  INV_X1 U14362 ( .A(n11966), .ZN(n11967) );
  NAND2_X1 U14363 ( .A1(n11968), .A2(n11967), .ZN(n11971) );
  MUX2_X1 U14364 ( .A(n11971), .B(n11970), .S(n11969), .Z(n11972) );
  OAI21_X1 U14365 ( .B1(n11974), .B2(n11973), .A(n11972), .ZN(n11975) );
  NAND4_X1 U14366 ( .A1(n11979), .A2(n14174), .A3(n7145), .A4(n11978), .ZN(
        n11980) );
  OAI211_X1 U14367 ( .C1(n14393), .C2(n11982), .A(n11980), .B(P1_B_REG_SCAN_IN), .ZN(n11981) );
  OAI21_X1 U14368 ( .B1(n11983), .B2(n11982), .A(n11981), .ZN(P1_U3242) );
  INV_X1 U14369 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n15261) );
  INV_X1 U14370 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n15432) );
  OR2_X1 U14371 ( .A1(n11984), .A2(n15432), .ZN(n11987) );
  INV_X1 U14372 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n11985) );
  OR2_X1 U14373 ( .A1(n9369), .A2(n11985), .ZN(n11986) );
  OAI211_X1 U14374 ( .C1(n6558), .C2(n15261), .A(n11987), .B(n11986), .ZN(
        n11988) );
  INV_X1 U14375 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U14376 ( .A1(n11990), .A2(n11989), .ZN(n12596) );
  INV_X1 U14377 ( .A(n12596), .ZN(n12743) );
  INV_X1 U14378 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14379 ( .A1(n11993), .A2(n11992), .ZN(n11995) );
  NAND2_X1 U14380 ( .A1(n14381), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U14381 ( .A1(n11995), .A2(n11994), .ZN(n12003) );
  NAND2_X1 U14382 ( .A1(n14378), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U14383 ( .A1(n12214), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U14384 ( .A1(n11998), .A2(n11996), .ZN(n12002) );
  INV_X1 U14385 ( .A(n12002), .ZN(n11997) );
  NAND2_X1 U14386 ( .A1(n12003), .A2(n11997), .ZN(n11999) );
  XNOR2_X1 U14387 ( .A(n12000), .B(P1_DATAO_REG_31__SCAN_IN), .ZN(n12001) );
  INV_X1 U14388 ( .A(SI_31_), .ZN(n13080) );
  XNOR2_X1 U14389 ( .A(n12003), .B(n12002), .ZN(n12377) );
  NAND2_X1 U14390 ( .A1(n12377), .A2(n12004), .ZN(n12007) );
  INV_X1 U14391 ( .A(SI_30_), .ZN(n12378) );
  OR2_X1 U14392 ( .A1(n12005), .A2(n12378), .ZN(n12006) );
  INV_X1 U14393 ( .A(n13026), .ZN(n12149) );
  OAI22_X1 U14394 ( .A1(n13023), .A2(n12596), .B1(n12148), .B2(n12149), .ZN(
        n12179) );
  NAND2_X1 U14395 ( .A1(n12179), .A2(n12147), .ZN(n12156) );
  OAI21_X1 U14396 ( .B1(n15086), .B2(n12008), .A(n12036), .ZN(n12035) );
  AOI21_X1 U14397 ( .B1(n12039), .B2(n12009), .A(n12143), .ZN(n12040) );
  INV_X1 U14398 ( .A(n12018), .ZN(n12010) );
  AOI211_X1 U14399 ( .C1(n12014), .C2(n12011), .A(n12133), .B(n12010), .ZN(
        n12016) );
  INV_X1 U14400 ( .A(n12011), .ZN(n12013) );
  NOR3_X1 U14401 ( .A1(n13015), .A2(n12013), .A3(n12012), .ZN(n12015) );
  OAI22_X1 U14402 ( .A1(n12016), .A2(n12015), .B1(n12014), .B2(n13014), .ZN(
        n12020) );
  MUX2_X1 U14403 ( .A(n12018), .B(n12017), .S(n12143), .Z(n12019) );
  AND3_X1 U14404 ( .A1(n12020), .A2(n15109), .A3(n12019), .ZN(n12029) );
  NAND2_X1 U14405 ( .A1(n12026), .A2(n12021), .ZN(n12024) );
  NAND2_X1 U14406 ( .A1(n12025), .A2(n12022), .ZN(n12023) );
  MUX2_X1 U14407 ( .A(n12024), .B(n12023), .S(n12133), .Z(n12028) );
  MUX2_X1 U14408 ( .A(n12026), .B(n12025), .S(n12143), .Z(n12027) );
  OAI211_X1 U14409 ( .C1(n12029), .C2(n12028), .A(n15082), .B(n12027), .ZN(
        n12033) );
  MUX2_X1 U14410 ( .A(n12031), .B(n12030), .S(n12133), .Z(n12032) );
  AND3_X1 U14411 ( .A1(n12033), .A2(n12165), .A3(n12032), .ZN(n12034) );
  INV_X1 U14412 ( .A(n12036), .ZN(n12037) );
  AOI21_X1 U14413 ( .B1(n12037), .B2(n12133), .A(n15056), .ZN(n12038) );
  OAI21_X1 U14414 ( .B1(n12040), .B2(n12039), .A(n12038), .ZN(n12044) );
  MUX2_X1 U14415 ( .A(n12042), .B(n12041), .S(n12143), .Z(n12043) );
  OAI211_X1 U14416 ( .C1(n12045), .C2(n12044), .A(n15061), .B(n12043), .ZN(
        n12050) );
  INV_X1 U14417 ( .A(n15041), .ZN(n15050) );
  NAND2_X1 U14418 ( .A1(n15045), .A2(n12046), .ZN(n12047) );
  MUX2_X1 U14419 ( .A(n12048), .B(n12047), .S(n12133), .Z(n12049) );
  NAND3_X1 U14420 ( .A1(n12050), .A2(n15050), .A3(n12049), .ZN(n12054) );
  MUX2_X1 U14421 ( .A(n12052), .B(n12051), .S(n12143), .Z(n12053) );
  NAND3_X1 U14422 ( .A1(n12054), .A2(n12159), .A3(n12053), .ZN(n12058) );
  MUX2_X1 U14423 ( .A(n12056), .B(n12055), .S(n12133), .Z(n12057) );
  NAND2_X1 U14424 ( .A1(n12064), .A2(n12059), .ZN(n12062) );
  NAND2_X1 U14425 ( .A1(n12063), .A2(n12060), .ZN(n12061) );
  MUX2_X1 U14426 ( .A(n12062), .B(n12061), .S(n12133), .Z(n12066) );
  MUX2_X1 U14427 ( .A(n12064), .B(n12063), .S(n12143), .Z(n12065) );
  OAI21_X1 U14428 ( .B1(n12067), .B2(n12066), .A(n12065), .ZN(n12068) );
  NAND2_X1 U14429 ( .A1(n12070), .A2(n12075), .ZN(n14588) );
  INV_X1 U14430 ( .A(n14588), .ZN(n14584) );
  NAND2_X1 U14431 ( .A1(n12068), .A2(n14584), .ZN(n12069) );
  OAI211_X1 U14432 ( .C1(n12070), .C2(n12143), .A(n12069), .B(n6976), .ZN(
        n12079) );
  MUX2_X1 U14433 ( .A(n12071), .B(n12926), .S(n12143), .Z(n12072) );
  NAND2_X1 U14434 ( .A1(n12928), .A2(n12072), .ZN(n12076) );
  INV_X1 U14435 ( .A(n12076), .ZN(n12078) );
  OAI211_X1 U14436 ( .C1(n12076), .C2(n12075), .A(n12074), .B(n12073), .ZN(
        n12077) );
  AOI22_X1 U14437 ( .A1(n12079), .A2(n12078), .B1(n12143), .B2(n12077), .ZN(
        n12084) );
  INV_X1 U14438 ( .A(n12081), .ZN(n12083) );
  AND2_X1 U14439 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  OAI22_X1 U14440 ( .A1(n12084), .A2(n12083), .B1(n12082), .B2(n12143), .ZN(
        n12086) );
  INV_X1 U14441 ( .A(n12405), .ZN(n13071) );
  NAND3_X1 U14442 ( .A1(n13071), .A2(n12133), .A3(n12601), .ZN(n12085) );
  OAI211_X1 U14443 ( .C1(n6571), .C2(n12087), .A(n12095), .B(n12088), .ZN(
        n12093) );
  INV_X1 U14444 ( .A(n12088), .ZN(n12091) );
  OAI211_X1 U14445 ( .C1(n12091), .C2(n12090), .A(n12094), .B(n12089), .ZN(
        n12092) );
  MUX2_X1 U14446 ( .A(n12093), .B(n12092), .S(n12133), .Z(n12097) );
  MUX2_X1 U14447 ( .A(n12095), .B(n12094), .S(n12143), .Z(n12096) );
  OAI211_X1 U14448 ( .C1(n12098), .C2(n12097), .A(n12855), .B(n12096), .ZN(
        n12102) );
  NAND2_X1 U14449 ( .A1(n12866), .A2(n12872), .ZN(n12099) );
  MUX2_X1 U14450 ( .A(n12100), .B(n12099), .S(n12143), .Z(n12101) );
  NAND2_X1 U14451 ( .A1(n12102), .A2(n12101), .ZN(n12111) );
  INV_X1 U14452 ( .A(n12846), .ZN(n12110) );
  INV_X1 U14453 ( .A(n12105), .ZN(n12107) );
  MUX2_X1 U14454 ( .A(n12107), .B(n12106), .S(n12133), .Z(n12109) );
  INV_X1 U14455 ( .A(n12114), .ZN(n12108) );
  INV_X1 U14456 ( .A(n12835), .ZN(n12830) );
  AOI211_X1 U14457 ( .C1(n12111), .C2(n12110), .A(n12109), .B(n12830), .ZN(
        n12116) );
  INV_X1 U14458 ( .A(n12112), .ZN(n12113) );
  MUX2_X1 U14459 ( .A(n12114), .B(n12113), .S(n12143), .Z(n12115) );
  NAND3_X1 U14460 ( .A1(n12824), .A2(n12833), .A3(n12133), .ZN(n12117) );
  AOI21_X1 U14461 ( .B1(n12118), .B2(n12117), .A(n12807), .ZN(n12124) );
  AOI21_X1 U14462 ( .B1(n12120), .B2(n12119), .A(n12133), .ZN(n12122) );
  MUX2_X1 U14463 ( .A(n12133), .B(n12122), .S(n12121), .Z(n12123) );
  NOR3_X1 U14464 ( .A1(n12131), .A2(n12126), .A3(n12778), .ZN(n12128) );
  NOR2_X1 U14465 ( .A1(n12128), .A2(n12127), .ZN(n12135) );
  INV_X1 U14466 ( .A(n12129), .ZN(n12130) );
  NOR3_X1 U14467 ( .A1(n12131), .A2(n12130), .A3(n12778), .ZN(n12132) );
  NOR2_X1 U14468 ( .A1(n12132), .A2(n7497), .ZN(n12134) );
  MUX2_X1 U14469 ( .A(n12135), .B(n12134), .S(n12133), .Z(n12137) );
  INV_X1 U14470 ( .A(n12763), .ZN(n12136) );
  INV_X1 U14471 ( .A(n12142), .ZN(n12140) );
  NAND3_X1 U14472 ( .A1(n12140), .A2(n12139), .A3(n12138), .ZN(n12145) );
  INV_X1 U14473 ( .A(n12754), .ZN(n12175) );
  OAI21_X1 U14474 ( .B1(n12142), .B2(n12141), .A(n12175), .ZN(n12144) );
  INV_X1 U14475 ( .A(n12750), .ZN(n12466) );
  OAI21_X1 U14476 ( .B1(n12385), .B2(n12466), .A(n12146), .ZN(n12154) );
  INV_X1 U14477 ( .A(n12154), .ZN(n12153) );
  OR2_X1 U14478 ( .A1(n12147), .A2(n12743), .ZN(n12151) );
  NAND2_X1 U14479 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  NAND2_X1 U14480 ( .A1(n12151), .A2(n12150), .ZN(n12178) );
  AND2_X1 U14481 ( .A1(n12385), .A2(n12466), .ZN(n12152) );
  OAI22_X1 U14482 ( .A1(n12155), .A2(n12154), .B1(n13026), .B2(n12596), .ZN(
        n12158) );
  NAND3_X1 U14483 ( .A1(n15109), .A2(n15082), .A3(n12159), .ZN(n12160) );
  NOR4_X1 U14484 ( .A1(n12161), .A2(n9591), .A3(n12160), .A4(n13015), .ZN(
        n12166) );
  INV_X1 U14485 ( .A(n12162), .ZN(n12163) );
  NOR4_X1 U14486 ( .A1(n12163), .A2(n15056), .A3(n15041), .A4(n14937), .ZN(
        n12164) );
  NAND4_X1 U14487 ( .A1(n12166), .A2(n12165), .A3(n9339), .A4(n12164), .ZN(
        n12167) );
  NOR4_X1 U14488 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n14588), .ZN(
        n12170) );
  NAND4_X1 U14489 ( .A1(n12901), .A2(n12928), .A3(n12915), .A4(n12170), .ZN(
        n12171) );
  NOR4_X1 U14490 ( .A1(n12846), .A2(n9612), .A3(n6571), .A4(n12171), .ZN(
        n12172) );
  NAND4_X1 U14491 ( .A1(n12172), .A2(n12835), .A3(n12855), .A4(n12822), .ZN(
        n12173) );
  NOR4_X1 U14492 ( .A1(n12778), .A2(n12807), .A3(n12789), .A4(n12173), .ZN(
        n12174) );
  NAND4_X1 U14493 ( .A1(n12176), .A2(n12763), .A3(n12175), .A4(n12174), .ZN(
        n12177) );
  XNOR2_X1 U14494 ( .A(n12181), .B(n12180), .ZN(n12182) );
  NAND3_X1 U14495 ( .A1(n12188), .A2(n12187), .A3(n6550), .ZN(n12189) );
  OAI211_X1 U14496 ( .C1(n12190), .C2(n12192), .A(n12189), .B(P3_B_REG_SCAN_IN), .ZN(n12191) );
  OAI21_X1 U14497 ( .B1(n12193), .B2(n12192), .A(n12191), .ZN(P3_U3296) );
  INV_X1 U14498 ( .A(n12194), .ZN(n14382) );
  OAI222_X1 U14499 ( .A1(n11298), .A2(n14382), .B1(P2_U3088), .B2(n7627), .C1(
        n15334), .C2(n13736), .ZN(P2_U3298) );
  INV_X1 U14500 ( .A(n12196), .ZN(n12197) );
  OAI22_X1 U14501 ( .A1(n12199), .A2(n12198), .B1(n12197), .B2(n14526), .ZN(
        n12201) );
  NOR2_X1 U14502 ( .A1(n8747), .A2(n14525), .ZN(n12200) );
  AOI211_X1 U14503 ( .C1(n14224), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12201), 
        .B(n12200), .ZN(n12202) );
  OAI21_X1 U14504 ( .B1(n12203), .B2(n14516), .A(n12202), .ZN(n12204) );
  AOI21_X1 U14505 ( .B1(n12205), .B2(n14233), .A(n12204), .ZN(n12206) );
  OAI21_X1 U14506 ( .B1(n12195), .B2(n14224), .A(n12206), .ZN(P1_U3356) );
  NAND2_X1 U14507 ( .A1(n12207), .A2(n13912), .ZN(n12211) );
  AOI22_X1 U14508 ( .A1(n13936), .A2(n12209), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n12208), .ZN(n12210) );
  OAI211_X1 U14509 ( .C1(n12212), .C2(n13903), .A(n12211), .B(n12210), .ZN(
        P1_U3232) );
  INV_X1 U14510 ( .A(n12213), .ZN(n14379) );
  OAI222_X1 U14511 ( .A1(n11298), .A2(n14379), .B1(P2_U3088), .B2(n12215), 
        .C1(n12214), .C2(n13736), .ZN(P2_U3297) );
  INV_X1 U14512 ( .A(n12216), .ZN(n12217) );
  NAND2_X1 U14513 ( .A1(n12218), .A2(n12217), .ZN(n13771) );
  NOR2_X1 U14514 ( .A1(n12219), .A2(n12345), .ZN(n12220) );
  AOI21_X1 U14515 ( .B1(n13768), .B2(n12366), .A(n12220), .ZN(n12227) );
  AOI22_X1 U14516 ( .A1(n13768), .A2(n12363), .B1(n12362), .B2(n13950), .ZN(
        n12221) );
  XNOR2_X1 U14517 ( .A(n12221), .B(n12364), .ZN(n12228) );
  XOR2_X1 U14518 ( .A(n12227), .B(n12228), .Z(n13770) );
  NAND2_X1 U14519 ( .A1(n12222), .A2(n7603), .ZN(n13769) );
  NAND2_X1 U14520 ( .A1(n13896), .A2(n12363), .ZN(n12224) );
  OR2_X1 U14521 ( .A1(n13804), .A2(n12305), .ZN(n12223) );
  NAND2_X1 U14522 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  XNOR2_X1 U14523 ( .A(n12225), .B(n12343), .ZN(n12235) );
  NOR2_X1 U14524 ( .A1(n13804), .A2(n12345), .ZN(n12226) );
  AOI21_X1 U14525 ( .B1(n13896), .B2(n12366), .A(n12226), .ZN(n12234) );
  XNOR2_X1 U14526 ( .A(n12235), .B(n12234), .ZN(n13889) );
  NOR2_X1 U14527 ( .A1(n12228), .A2(n12227), .ZN(n13890) );
  NOR2_X1 U14528 ( .A1(n13889), .A2(n13890), .ZN(n12229) );
  NAND2_X1 U14529 ( .A1(n13769), .A2(n12229), .ZN(n13892) );
  OAI22_X1 U14530 ( .A1(n14538), .A2(n10522), .B1(n12231), .B2(n12305), .ZN(
        n12230) );
  XNOR2_X1 U14531 ( .A(n12230), .B(n12364), .ZN(n12236) );
  NOR2_X1 U14532 ( .A1(n12231), .A2(n12345), .ZN(n12232) );
  AOI21_X1 U14533 ( .B1(n12233), .B2(n12366), .A(n12232), .ZN(n12237) );
  XNOR2_X1 U14534 ( .A(n12236), .B(n12237), .ZN(n13802) );
  NAND2_X1 U14535 ( .A1(n12235), .A2(n12234), .ZN(n13800) );
  INV_X1 U14536 ( .A(n12236), .ZN(n12238) );
  OR2_X1 U14537 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  OAI22_X1 U14538 ( .A1(n14645), .A2(n10522), .B1(n13751), .B2(n12305), .ZN(
        n12240) );
  XNOR2_X1 U14539 ( .A(n12240), .B(n12364), .ZN(n12244) );
  AND2_X1 U14540 ( .A1(n10521), .A2(n13947), .ZN(n12241) );
  AOI21_X1 U14541 ( .B1(n13868), .B2(n12366), .A(n12241), .ZN(n12242) );
  XNOR2_X1 U14542 ( .A(n12244), .B(n12242), .ZN(n13862) );
  INV_X1 U14543 ( .A(n12242), .ZN(n12243) );
  NAND2_X1 U14544 ( .A1(n12244), .A2(n12243), .ZN(n12245) );
  NAND2_X1 U14545 ( .A1(n14329), .A2(n12363), .ZN(n12247) );
  OR2_X1 U14546 ( .A1(n13929), .A2(n12305), .ZN(n12246) );
  NAND2_X1 U14547 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  XNOR2_X1 U14548 ( .A(n12248), .B(n12343), .ZN(n12251) );
  NOR2_X1 U14549 ( .A1(n13929), .A2(n12345), .ZN(n12249) );
  AOI21_X1 U14550 ( .B1(n14329), .B2(n12366), .A(n12249), .ZN(n12250) );
  NAND2_X1 U14551 ( .A1(n12251), .A2(n12250), .ZN(n13922) );
  OAI21_X1 U14552 ( .B1(n12251), .B2(n12250), .A(n13922), .ZN(n13748) );
  INV_X1 U14553 ( .A(n13748), .ZN(n12252) );
  NAND2_X1 U14554 ( .A1(n14320), .A2(n12363), .ZN(n12254) );
  OR2_X1 U14555 ( .A1(n14213), .A2(n12305), .ZN(n12253) );
  NAND2_X1 U14556 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  XNOR2_X1 U14557 ( .A(n12255), .B(n12343), .ZN(n13925) );
  NOR2_X1 U14558 ( .A1(n14213), .A2(n12345), .ZN(n12256) );
  AOI21_X1 U14559 ( .B1(n14320), .B2(n12366), .A(n12256), .ZN(n13924) );
  INV_X1 U14560 ( .A(n13922), .ZN(n12257) );
  AOI21_X1 U14561 ( .B1(n13925), .B2(n13924), .A(n12257), .ZN(n12259) );
  NOR2_X1 U14562 ( .A1(n13925), .A2(n13924), .ZN(n12258) );
  NAND2_X1 U14563 ( .A1(n14206), .A2(n12363), .ZN(n12261) );
  OR2_X1 U14564 ( .A1(n13928), .A2(n12305), .ZN(n12260) );
  NAND2_X1 U14565 ( .A1(n12261), .A2(n12260), .ZN(n12262) );
  XNOR2_X1 U14566 ( .A(n12262), .B(n12343), .ZN(n12265) );
  INV_X1 U14567 ( .A(n12265), .ZN(n12267) );
  NOR2_X1 U14568 ( .A1(n13928), .A2(n12345), .ZN(n12263) );
  AOI21_X1 U14569 ( .B1(n14206), .B2(n12366), .A(n12263), .ZN(n12264) );
  INV_X1 U14570 ( .A(n12264), .ZN(n12266) );
  AOI21_X1 U14571 ( .B1(n12267), .B2(n12266), .A(n13833), .ZN(n13824) );
  NAND2_X1 U14572 ( .A1(n14310), .A2(n12363), .ZN(n12269) );
  OR2_X1 U14573 ( .A1(n14211), .A2(n12305), .ZN(n12268) );
  NAND2_X1 U14574 ( .A1(n12269), .A2(n12268), .ZN(n12270) );
  XNOR2_X1 U14575 ( .A(n12270), .B(n12343), .ZN(n12273) );
  NOR2_X1 U14576 ( .A1(n14211), .A2(n12345), .ZN(n12271) );
  AOI21_X1 U14577 ( .B1(n14310), .B2(n12366), .A(n12271), .ZN(n12272) );
  NAND2_X1 U14578 ( .A1(n12273), .A2(n12272), .ZN(n12276) );
  OR2_X1 U14579 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  AND2_X1 U14580 ( .A1(n12276), .A2(n12274), .ZN(n13832) );
  NAND2_X1 U14581 ( .A1(n13835), .A2(n12276), .ZN(n13899) );
  NAND2_X1 U14582 ( .A1(n14304), .A2(n12363), .ZN(n12278) );
  NAND2_X1 U14583 ( .A1(n14163), .A2(n12366), .ZN(n12277) );
  NAND2_X1 U14584 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  XNOR2_X1 U14585 ( .A(n12279), .B(n12364), .ZN(n12286) );
  AOI22_X1 U14586 ( .A1(n14304), .A2(n12366), .B1(n10521), .B2(n14163), .ZN(
        n12284) );
  XNOR2_X1 U14587 ( .A(n12286), .B(n12284), .ZN(n13900) );
  NAND2_X1 U14588 ( .A1(n14298), .A2(n12363), .ZN(n12281) );
  OR2_X1 U14589 ( .A1(n13902), .A2(n12305), .ZN(n12280) );
  NAND2_X1 U14590 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  XNOR2_X1 U14591 ( .A(n12282), .B(n12343), .ZN(n12289) );
  NOR2_X1 U14592 ( .A1(n13902), .A2(n12345), .ZN(n12283) );
  AOI21_X1 U14593 ( .B1(n14298), .B2(n12366), .A(n12283), .ZN(n12288) );
  XNOR2_X1 U14594 ( .A(n12289), .B(n12288), .ZN(n13780) );
  INV_X1 U14595 ( .A(n12284), .ZN(n12285) );
  NOR2_X1 U14596 ( .A1(n12286), .A2(n12285), .ZN(n13781) );
  NOR2_X1 U14597 ( .A1(n13780), .A2(n13781), .ZN(n12287) );
  OR2_X1 U14598 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  NAND2_X1 U14599 ( .A1(n14292), .A2(n12363), .ZN(n12292) );
  NAND2_X1 U14600 ( .A1(n14164), .A2(n12362), .ZN(n12291) );
  NAND2_X1 U14601 ( .A1(n12292), .A2(n12291), .ZN(n12293) );
  XNOR2_X1 U14602 ( .A(n12293), .B(n12364), .ZN(n12296) );
  AOI22_X1 U14603 ( .A1(n14292), .A2(n12366), .B1(n10521), .B2(n14164), .ZN(
        n12294) );
  XNOR2_X1 U14604 ( .A(n12296), .B(n12294), .ZN(n13855) );
  INV_X1 U14605 ( .A(n12294), .ZN(n12295) );
  NAND2_X1 U14606 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  NAND2_X1 U14607 ( .A1(n14288), .A2(n12363), .ZN(n12299) );
  NAND2_X1 U14608 ( .A1(n14140), .A2(n12366), .ZN(n12298) );
  NAND2_X1 U14609 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  XNOR2_X1 U14610 ( .A(n12300), .B(n12343), .ZN(n12303) );
  AND2_X1 U14611 ( .A1(n14140), .A2(n10521), .ZN(n12301) );
  AOI21_X1 U14612 ( .B1(n14288), .B2(n12366), .A(n12301), .ZN(n12302) );
  NAND2_X1 U14613 ( .A1(n12303), .A2(n12302), .ZN(n13871) );
  OAI21_X1 U14614 ( .B1(n12303), .B2(n12302), .A(n13871), .ZN(n13791) );
  INV_X1 U14615 ( .A(n13791), .ZN(n12304) );
  NAND2_X1 U14616 ( .A1(n13790), .A2(n13871), .ZN(n12314) );
  OAI22_X1 U14617 ( .A1(n13882), .A2(n10522), .B1(n13763), .B2(n12305), .ZN(
        n12306) );
  XNOR2_X1 U14618 ( .A(n12306), .B(n12343), .ZN(n12309) );
  OR2_X1 U14619 ( .A1(n13882), .A2(n12305), .ZN(n12308) );
  NAND2_X1 U14620 ( .A1(n14092), .A2(n10521), .ZN(n12307) );
  AND2_X1 U14621 ( .A1(n12308), .A2(n12307), .ZN(n12310) );
  NAND2_X1 U14622 ( .A1(n12309), .A2(n12310), .ZN(n13756) );
  INV_X1 U14623 ( .A(n12309), .ZN(n12312) );
  INV_X1 U14624 ( .A(n12310), .ZN(n12311) );
  NAND2_X1 U14625 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  NAND2_X1 U14626 ( .A1(n14276), .A2(n12363), .ZN(n12316) );
  NAND2_X1 U14627 ( .A1(n14072), .A2(n12362), .ZN(n12315) );
  NAND2_X1 U14628 ( .A1(n12316), .A2(n12315), .ZN(n12317) );
  XNOR2_X1 U14629 ( .A(n12317), .B(n12343), .ZN(n12319) );
  AND2_X1 U14630 ( .A1(n14072), .A2(n10521), .ZN(n12318) );
  AOI21_X1 U14631 ( .B1(n14276), .B2(n12366), .A(n12318), .ZN(n12320) );
  NAND2_X1 U14632 ( .A1(n12319), .A2(n12320), .ZN(n13843) );
  INV_X1 U14633 ( .A(n12319), .ZN(n12322) );
  INV_X1 U14634 ( .A(n12320), .ZN(n12321) );
  NAND2_X1 U14635 ( .A1(n12322), .A2(n12321), .ZN(n12323) );
  NAND2_X1 U14636 ( .A1(n14266), .A2(n12363), .ZN(n12326) );
  OR2_X1 U14637 ( .A1(n13817), .A2(n12305), .ZN(n12325) );
  NAND2_X1 U14638 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  XNOR2_X1 U14639 ( .A(n12327), .B(n12343), .ZN(n12330) );
  NOR2_X1 U14640 ( .A1(n13817), .A2(n12345), .ZN(n12328) );
  AOI21_X1 U14641 ( .B1(n14266), .B2(n12366), .A(n12328), .ZN(n12329) );
  NAND2_X1 U14642 ( .A1(n12330), .A2(n12329), .ZN(n13812) );
  OR2_X1 U14643 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  NAND2_X1 U14644 ( .A1(n14259), .A2(n12363), .ZN(n12333) );
  OR2_X1 U14645 ( .A1(n13914), .A2(n12305), .ZN(n12332) );
  NAND2_X1 U14646 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  XNOR2_X1 U14647 ( .A(n12334), .B(n12343), .ZN(n12337) );
  NOR2_X1 U14648 ( .A1(n13914), .A2(n12345), .ZN(n12335) );
  AOI21_X1 U14649 ( .B1(n14259), .B2(n12362), .A(n12335), .ZN(n12336) );
  NAND2_X1 U14650 ( .A1(n12337), .A2(n12336), .ZN(n12340) );
  OR2_X1 U14651 ( .A1(n12337), .A2(n12336), .ZN(n12338) );
  NAND2_X1 U14652 ( .A1(n12339), .A2(n13813), .ZN(n13814) );
  NAND2_X1 U14653 ( .A1(n12347), .A2(n12363), .ZN(n12342) );
  OR2_X1 U14654 ( .A1(n13818), .A2(n12305), .ZN(n12341) );
  NAND2_X1 U14655 ( .A1(n12342), .A2(n12341), .ZN(n12344) );
  XNOR2_X1 U14656 ( .A(n12344), .B(n12343), .ZN(n12349) );
  INV_X1 U14657 ( .A(n12349), .ZN(n12351) );
  NOR2_X1 U14658 ( .A1(n13818), .A2(n12345), .ZN(n12346) );
  AOI21_X1 U14659 ( .B1(n12347), .B2(n12362), .A(n12346), .ZN(n12348) );
  INV_X1 U14660 ( .A(n12348), .ZN(n12350) );
  AND2_X1 U14661 ( .A1(n12349), .A2(n12348), .ZN(n12352) );
  AOI21_X1 U14662 ( .B1(n12351), .B2(n12350), .A(n12352), .ZN(n13911) );
  INV_X1 U14663 ( .A(n12352), .ZN(n12353) );
  NAND2_X1 U14664 ( .A1(n14248), .A2(n12363), .ZN(n12355) );
  NAND2_X1 U14665 ( .A1(n13943), .A2(n12366), .ZN(n12354) );
  NAND2_X1 U14666 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  XNOR2_X1 U14667 ( .A(n12356), .B(n12364), .ZN(n12360) );
  NAND2_X1 U14668 ( .A1(n14248), .A2(n12362), .ZN(n12358) );
  NAND2_X1 U14669 ( .A1(n10521), .A2(n13943), .ZN(n12357) );
  NAND2_X1 U14670 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  NOR2_X1 U14671 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  AOI21_X1 U14672 ( .B1(n12360), .B2(n12359), .A(n12361), .ZN(n13740) );
  AOI22_X1 U14673 ( .A1(n14243), .A2(n12363), .B1(n12362), .B2(n13942), .ZN(
        n12365) );
  XNOR2_X1 U14674 ( .A(n12365), .B(n12364), .ZN(n12368) );
  AOI22_X1 U14675 ( .A1(n6879), .A2(n12366), .B1(n10521), .B2(n13942), .ZN(
        n12367) );
  XNOR2_X1 U14676 ( .A(n12368), .B(n12367), .ZN(n12369) );
  INV_X1 U14677 ( .A(n12370), .ZN(n14014) );
  OAI22_X1 U14678 ( .A1(n12372), .A2(n14212), .B1(n12371), .B2(n14210), .ZN(
        n14008) );
  AOI22_X1 U14679 ( .A1(n14008), .A2(n13795), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12373) );
  OAI21_X1 U14680 ( .B1(n14014), .B2(n13887), .A(n12373), .ZN(n12374) );
  AOI21_X1 U14681 ( .B1(n14243), .B2(n13936), .A(n12374), .ZN(n12375) );
  OAI21_X1 U14682 ( .B1(n12376), .B2(n13938), .A(n12375), .ZN(P1_U3220) );
  INV_X1 U14683 ( .A(n12377), .ZN(n12379) );
  OAI222_X1 U14684 ( .A1(P3_U3151), .A2(n12380), .B1(n13089), .B2(n12379), 
        .C1(n12378), .C2(n13092), .ZN(P3_U3265) );
  OR2_X1 U14685 ( .A1(n12381), .A2(n15101), .ZN(n12744) );
  OAI21_X1 U14686 ( .B1(n15129), .B2(n12382), .A(n12744), .ZN(n12384) );
  XNOR2_X1 U14687 ( .A(n13032), .B(n12462), .ZN(n12458) );
  XNOR2_X1 U14688 ( .A(n12458), .B(n12752), .ZN(n12460) );
  INV_X1 U14689 ( .A(n12387), .ZN(n12388) );
  NAND2_X1 U14690 ( .A1(n12388), .A2(n15044), .ZN(n12389) );
  XNOR2_X1 U14691 ( .A(n14610), .B(n12421), .ZN(n12482) );
  INV_X1 U14692 ( .A(n12605), .ZN(n14602) );
  XNOR2_X1 U14693 ( .A(n12391), .B(n12421), .ZN(n12480) );
  INV_X1 U14694 ( .A(n12480), .ZN(n12392) );
  INV_X1 U14695 ( .A(n12606), .ZN(n15029) );
  OAI22_X1 U14696 ( .A1(n12482), .A2(n14602), .B1(n12392), .B2(n15029), .ZN(
        n12396) );
  OAI21_X1 U14697 ( .B1(n12480), .B2(n12606), .A(n12605), .ZN(n12394) );
  NOR2_X1 U14698 ( .A1(n12605), .A2(n12606), .ZN(n12393) );
  AOI22_X1 U14699 ( .A1(n12394), .A2(n12482), .B1(n12393), .B2(n12392), .ZN(
        n12395) );
  XNOR2_X1 U14700 ( .A(n14592), .B(n12462), .ZN(n12536) );
  AND2_X1 U14701 ( .A1(n12536), .A2(n12439), .ZN(n12397) );
  INV_X1 U14702 ( .A(n12536), .ZN(n12398) );
  NAND2_X1 U14703 ( .A1(n12398), .A2(n12604), .ZN(n12399) );
  XNOR2_X1 U14704 ( .A(n13002), .B(n12462), .ZN(n12400) );
  XNOR2_X1 U14705 ( .A(n12400), .B(n12603), .ZN(n12437) );
  INV_X1 U14706 ( .A(n12400), .ZN(n12401) );
  NAND2_X1 U14707 ( .A1(n12401), .A2(n12603), .ZN(n12402) );
  XNOR2_X1 U14708 ( .A(n12930), .B(n12462), .ZN(n12403) );
  XNOR2_X1 U14709 ( .A(n12403), .B(n12912), .ZN(n12586) );
  NAND2_X1 U14710 ( .A1(n12403), .A2(n12912), .ZN(n12404) );
  XNOR2_X1 U14711 ( .A(n12405), .B(n12462), .ZN(n12406) );
  XNOR2_X1 U14712 ( .A(n12406), .B(n12601), .ZN(n12503) );
  NAND2_X1 U14713 ( .A1(n12504), .A2(n12503), .ZN(n12502) );
  INV_X1 U14714 ( .A(n12406), .ZN(n12407) );
  NAND2_X1 U14715 ( .A1(n12407), .A2(n12601), .ZN(n12408) );
  XNOR2_X1 U14716 ( .A(n12903), .B(n12462), .ZN(n12409) );
  XNOR2_X1 U14717 ( .A(n12409), .B(n12883), .ZN(n12509) );
  NAND2_X1 U14718 ( .A1(n12510), .A2(n12509), .ZN(n12412) );
  INV_X1 U14719 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14720 ( .A1(n12410), .A2(n12883), .ZN(n12411) );
  XNOR2_X1 U14721 ( .A(n12986), .B(n12462), .ZN(n12413) );
  NAND2_X1 U14722 ( .A1(n12413), .A2(n12900), .ZN(n12563) );
  INV_X1 U14723 ( .A(n12413), .ZN(n12414) );
  NAND2_X1 U14724 ( .A1(n12414), .A2(n12600), .ZN(n12564) );
  XNOR2_X1 U14725 ( .A(n13062), .B(n12462), .ZN(n12415) );
  XNOR2_X1 U14726 ( .A(n12415), .B(n12531), .ZN(n12452) );
  XNOR2_X1 U14727 ( .A(n12866), .B(n12462), .ZN(n12416) );
  XNOR2_X1 U14728 ( .A(n12416), .B(n12599), .ZN(n12528) );
  INV_X1 U14729 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U14730 ( .A1(n12417), .A2(n12599), .ZN(n12418) );
  NAND2_X1 U14731 ( .A1(n12527), .A2(n12418), .ZN(n12473) );
  XNOR2_X1 U14732 ( .A(n12848), .B(n12462), .ZN(n12419) );
  XNOR2_X1 U14733 ( .A(n12419), .B(n12834), .ZN(n12474) );
  NAND2_X1 U14734 ( .A1(n12419), .A2(n12834), .ZN(n12420) );
  XNOR2_X1 U14735 ( .A(n12837), .B(n12421), .ZN(n12422) );
  XNOR2_X2 U14736 ( .A(n12424), .B(n12422), .ZN(n12547) );
  INV_X1 U14737 ( .A(n12422), .ZN(n12423) );
  XNOR2_X1 U14738 ( .A(n12810), .B(n12462), .ZN(n12519) );
  XNOR2_X1 U14739 ( .A(n12824), .B(n12462), .ZN(n12426) );
  OAI22_X1 U14740 ( .A1(n12519), .A2(n12821), .B1(n12833), .B2(n12426), .ZN(
        n12428) );
  INV_X1 U14741 ( .A(n12426), .ZN(n12516) );
  OAI21_X1 U14742 ( .B1(n12516), .B2(n12803), .A(n12791), .ZN(n12427) );
  XNOR2_X1 U14743 ( .A(n13039), .B(n12462), .ZN(n12429) );
  XNOR2_X1 U14744 ( .A(n12429), .B(n12806), .ZN(n12495) );
  INV_X1 U14745 ( .A(n12429), .ZN(n12430) );
  XNOR2_X1 U14746 ( .A(n12579), .B(n12462), .ZN(n12431) );
  XNOR2_X1 U14747 ( .A(n12431), .B(n12765), .ZN(n12573) );
  XOR2_X1 U14748 ( .A(n12460), .B(n12461), .Z(n12436) );
  AOI22_X1 U14749 ( .A1(n12792), .A2(n12555), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12432) );
  OAI21_X1 U14750 ( .B1(n12766), .B2(n12575), .A(n12432), .ZN(n12434) );
  NOR2_X1 U14751 ( .A1(n13032), .A2(n14935), .ZN(n12433) );
  AOI211_X1 U14752 ( .C1(n12770), .C2(n12578), .A(n12434), .B(n12433), .ZN(
        n12435) );
  OAI21_X1 U14753 ( .B1(n12436), .B2(n12594), .A(n12435), .ZN(P3_U3154) );
  XNOR2_X1 U14754 ( .A(n12438), .B(n12437), .ZN(n12445) );
  NOR2_X1 U14755 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15366), .ZN(n12631) );
  NOR2_X1 U14756 ( .A1(n12439), .A2(n12587), .ZN(n12440) );
  AOI211_X1 U14757 ( .C1(n14932), .C2(n12602), .A(n12631), .B(n12440), .ZN(
        n12441) );
  OAI21_X1 U14758 ( .B1(n12442), .B2(n12590), .A(n12441), .ZN(n12443) );
  AOI21_X1 U14759 ( .B1(n12592), .B2(n13002), .A(n12443), .ZN(n12444) );
  OAI21_X1 U14760 ( .B1(n12445), .B2(n12594), .A(n12444), .ZN(P3_U3155) );
  XNOR2_X1 U14761 ( .A(n12518), .B(n12833), .ZN(n12450) );
  AOI22_X1 U14762 ( .A1(n12791), .A2(n14932), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12447) );
  NAND2_X1 U14763 ( .A1(n12578), .A2(n12825), .ZN(n12446) );
  OAI211_X1 U14764 ( .C1(n12845), .C2(n12587), .A(n12447), .B(n12446), .ZN(
        n12448) );
  AOI21_X1 U14765 ( .B1(n12824), .B2(n12592), .A(n12448), .ZN(n12449) );
  OAI21_X1 U14766 ( .B1(n12450), .B2(n12594), .A(n12449), .ZN(P3_U3156) );
  OAI211_X1 U14767 ( .C1(n12453), .C2(n12452), .A(n12451), .B(n14938), .ZN(
        n12457) );
  NAND2_X1 U14768 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12728)
         );
  OAI21_X1 U14769 ( .B1(n12872), .B2(n12575), .A(n12728), .ZN(n12455) );
  NOR2_X1 U14770 ( .A1(n12590), .A2(n12877), .ZN(n12454) );
  AOI211_X1 U14771 ( .C1(n12555), .C2(n12600), .A(n12455), .B(n12454), .ZN(
        n12456) );
  OAI211_X1 U14772 ( .C1(n14935), .C2(n13062), .A(n12457), .B(n12456), .ZN(
        P3_U3159) );
  INV_X1 U14773 ( .A(n12458), .ZN(n12459) );
  XOR2_X1 U14774 ( .A(n12462), .B(n12754), .Z(n12463) );
  XNOR2_X1 U14775 ( .A(n12464), .B(n12463), .ZN(n12470) );
  AOI22_X1 U14776 ( .A1(n12777), .A2(n12555), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12465) );
  OAI21_X1 U14777 ( .B1(n12466), .B2(n12575), .A(n12465), .ZN(n12468) );
  NOR2_X1 U14778 ( .A1(n13029), .A2(n14935), .ZN(n12467) );
  AOI211_X1 U14779 ( .C1(n12755), .C2(n12578), .A(n12468), .B(n12467), .ZN(
        n12469) );
  OAI21_X1 U14780 ( .B1(n12470), .B2(n12594), .A(n12469), .ZN(P3_U3160) );
  INV_X1 U14781 ( .A(n12471), .ZN(n12472) );
  AOI21_X1 U14782 ( .B1(n12474), .B2(n12473), .A(n12472), .ZN(n12479) );
  NOR2_X1 U14783 ( .A1(n12845), .A2(n12575), .ZN(n12476) );
  OAI22_X1 U14784 ( .A1(n12872), .A2(n12587), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15291), .ZN(n12475) );
  AOI211_X1 U14785 ( .C1(n12849), .C2(n12578), .A(n12476), .B(n12475), .ZN(
        n12478) );
  NAND2_X1 U14786 ( .A1(n12848), .A2(n12592), .ZN(n12477) );
  OAI211_X1 U14787 ( .C1(n12479), .C2(n12594), .A(n12478), .B(n12477), .ZN(
        P3_U3163) );
  XNOR2_X1 U14788 ( .A(n12481), .B(n12480), .ZN(n12559) );
  NOR2_X1 U14789 ( .A1(n12559), .A2(n15029), .ZN(n12558) );
  AOI21_X1 U14790 ( .B1(n12481), .B2(n12480), .A(n12558), .ZN(n12484) );
  XNOR2_X1 U14791 ( .A(n12482), .B(n14602), .ZN(n12483) );
  XNOR2_X1 U14792 ( .A(n12484), .B(n12483), .ZN(n12493) );
  INV_X1 U14793 ( .A(n12485), .ZN(n12486) );
  NAND2_X1 U14794 ( .A1(n12578), .A2(n12486), .ZN(n12489) );
  AOI21_X1 U14795 ( .B1(n12604), .B2(n14932), .A(n12487), .ZN(n12488) );
  OAI211_X1 U14796 ( .C1(n15029), .C2(n12587), .A(n12489), .B(n12488), .ZN(
        n12490) );
  AOI21_X1 U14797 ( .B1(n12592), .B2(n12491), .A(n12490), .ZN(n12492) );
  OAI21_X1 U14798 ( .B1(n12493), .B2(n12594), .A(n12492), .ZN(P3_U3164) );
  XOR2_X1 U14799 ( .A(n12495), .B(n12494), .Z(n12501) );
  AOI22_X1 U14800 ( .A1(n12791), .A2(n12555), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12497) );
  NAND2_X1 U14801 ( .A1(n12578), .A2(n12797), .ZN(n12496) );
  OAI211_X1 U14802 ( .C1(n12765), .C2(n12575), .A(n12497), .B(n12496), .ZN(
        n12498) );
  AOI21_X1 U14803 ( .B1(n12499), .B2(n12592), .A(n12498), .ZN(n12500) );
  OAI21_X1 U14804 ( .B1(n12501), .B2(n12594), .A(n12500), .ZN(P3_U3165) );
  OAI211_X1 U14805 ( .C1(n12504), .C2(n12503), .A(n12502), .B(n14938), .ZN(
        n12508) );
  NAND2_X1 U14806 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12654)
         );
  OAI21_X1 U14807 ( .B1(n12913), .B2(n12575), .A(n12654), .ZN(n12506) );
  NOR2_X1 U14808 ( .A1(n12590), .A2(n12917), .ZN(n12505) );
  AOI211_X1 U14809 ( .C1(n12555), .C2(n12602), .A(n12506), .B(n12505), .ZN(
        n12507) );
  OAI211_X1 U14810 ( .C1(n13071), .C2(n14935), .A(n12508), .B(n12507), .ZN(
        P3_U3166) );
  XNOR2_X1 U14811 ( .A(n12510), .B(n12509), .ZN(n12515) );
  NAND2_X1 U14812 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12677)
         );
  OAI21_X1 U14813 ( .B1(n12900), .B2(n12575), .A(n12677), .ZN(n12511) );
  AOI21_X1 U14814 ( .B1(n12555), .B2(n12601), .A(n12511), .ZN(n12512) );
  OAI21_X1 U14815 ( .B1(n12904), .B2(n12590), .A(n12512), .ZN(n12513) );
  AOI21_X1 U14816 ( .B1(n12903), .B2(n12592), .A(n12513), .ZN(n12514) );
  OAI21_X1 U14817 ( .B1(n12515), .B2(n12594), .A(n12514), .ZN(P3_U3168) );
  OAI22_X1 U14818 ( .A1(n12518), .A2(n12803), .B1(n12517), .B2(n12516), .ZN(
        n12521) );
  XNOR2_X1 U14819 ( .A(n12519), .B(n12821), .ZN(n12520) );
  XNOR2_X1 U14820 ( .A(n12521), .B(n12520), .ZN(n12526) );
  AOI22_X1 U14821 ( .A1(n12803), .A2(n12555), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12523) );
  NAND2_X1 U14822 ( .A1(n12578), .A2(n12811), .ZN(n12522) );
  OAI211_X1 U14823 ( .C1(n12806), .C2(n12575), .A(n12523), .B(n12522), .ZN(
        n12524) );
  AOI21_X1 U14824 ( .B1(n12810), .B2(n12592), .A(n12524), .ZN(n12525) );
  OAI21_X1 U14825 ( .B1(n12526), .B2(n12594), .A(n12525), .ZN(P3_U3169) );
  INV_X1 U14826 ( .A(n12866), .ZN(n13058) );
  OAI211_X1 U14827 ( .C1(n12529), .C2(n12528), .A(n12527), .B(n14938), .ZN(
        n12535) );
  AOI22_X1 U14828 ( .A1(n12860), .A2(n14932), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12530) );
  OAI21_X1 U14829 ( .B1(n12531), .B2(n12587), .A(n12530), .ZN(n12532) );
  AOI21_X1 U14830 ( .B1(n12533), .B2(n12578), .A(n12532), .ZN(n12534) );
  OAI211_X1 U14831 ( .C1(n13058), .C2(n14935), .A(n12535), .B(n12534), .ZN(
        P3_U3173) );
  XNOR2_X1 U14832 ( .A(n12536), .B(n12604), .ZN(n12537) );
  XNOR2_X1 U14833 ( .A(n12538), .B(n12537), .ZN(n12545) );
  AND2_X1 U14834 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15021) );
  AOI21_X1 U14835 ( .B1(n12603), .B2(n14932), .A(n15021), .ZN(n12543) );
  NAND2_X1 U14836 ( .A1(n14592), .A2(n12592), .ZN(n12542) );
  INV_X1 U14837 ( .A(n12539), .ZN(n14594) );
  NAND2_X1 U14838 ( .A1(n12578), .A2(n14594), .ZN(n12541) );
  NAND2_X1 U14839 ( .A1(n12605), .A2(n12555), .ZN(n12540) );
  NAND4_X1 U14840 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12544) );
  AOI21_X1 U14841 ( .B1(n12545), .B2(n14938), .A(n12544), .ZN(n12546) );
  INV_X1 U14842 ( .A(n12546), .ZN(P3_U3174) );
  XNOR2_X1 U14843 ( .A(n12547), .B(n12818), .ZN(n12552) );
  AOI22_X1 U14844 ( .A1(n12860), .A2(n12555), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12549) );
  NAND2_X1 U14845 ( .A1(n12578), .A2(n12838), .ZN(n12548) );
  OAI211_X1 U14846 ( .C1(n12833), .C2(n12575), .A(n12549), .B(n12548), .ZN(
        n12550) );
  AOI21_X1 U14847 ( .B1(n12837), .B2(n12592), .A(n12550), .ZN(n12551) );
  OAI21_X1 U14848 ( .B1(n12552), .B2(n12594), .A(n12551), .ZN(P3_U3175) );
  INV_X1 U14849 ( .A(n12553), .ZN(n14604) );
  AOI21_X1 U14850 ( .B1(n12605), .B2(n14932), .A(n12554), .ZN(n12557) );
  NAND2_X1 U14851 ( .A1(n15044), .A2(n12555), .ZN(n12556) );
  OAI211_X1 U14852 ( .C1(n14935), .C2(n14603), .A(n12557), .B(n12556), .ZN(
        n12561) );
  AOI211_X1 U14853 ( .C1(n15029), .C2(n12559), .A(n12594), .B(n12558), .ZN(
        n12560) );
  AOI211_X1 U14854 ( .C1(n14604), .C2(n12578), .A(n12561), .B(n12560), .ZN(
        n12562) );
  INV_X1 U14855 ( .A(n12562), .ZN(P3_U3176) );
  NAND2_X1 U14856 ( .A1(n12564), .A2(n12563), .ZN(n12566) );
  XOR2_X1 U14857 ( .A(n12566), .B(n6797), .Z(n12571) );
  NOR2_X1 U14858 ( .A1(n15273), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12700) );
  NOR2_X1 U14859 ( .A1(n12913), .A2(n12587), .ZN(n12567) );
  AOI211_X1 U14860 ( .C1(n14932), .C2(n12884), .A(n12700), .B(n12567), .ZN(
        n12568) );
  OAI21_X1 U14861 ( .B1(n12886), .B2(n12590), .A(n12568), .ZN(n12569) );
  AOI21_X1 U14862 ( .B1(n12986), .B2(n12592), .A(n12569), .ZN(n12570) );
  OAI21_X1 U14863 ( .B1(n12571), .B2(n12594), .A(n12570), .ZN(P3_U3178) );
  XOR2_X1 U14864 ( .A(n12573), .B(n12572), .Z(n12582) );
  OAI22_X1 U14865 ( .A1(n12806), .A2(n12587), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12574), .ZN(n12577) );
  NOR2_X1 U14866 ( .A1(n12752), .A2(n12575), .ZN(n12576) );
  AOI211_X1 U14867 ( .C1(n12783), .C2(n12578), .A(n12577), .B(n12576), .ZN(
        n12581) );
  NAND2_X1 U14868 ( .A1(n12579), .A2(n12592), .ZN(n12580) );
  INV_X1 U14869 ( .A(n12583), .ZN(n12584) );
  AOI21_X1 U14870 ( .B1(n12586), .B2(n12585), .A(n12584), .ZN(n12595) );
  INV_X1 U14871 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15413) );
  NOR2_X1 U14872 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15413), .ZN(n14578) );
  NOR2_X1 U14873 ( .A1(n14591), .A2(n12587), .ZN(n12588) );
  AOI211_X1 U14874 ( .C1(n14932), .C2(n12601), .A(n14578), .B(n12588), .ZN(
        n12589) );
  OAI21_X1 U14875 ( .B1(n12931), .B2(n12590), .A(n12589), .ZN(n12591) );
  AOI21_X1 U14876 ( .B1(n12592), .B2(n12930), .A(n12591), .ZN(n12593) );
  OAI21_X1 U14877 ( .B1(n12595), .B2(n12594), .A(n12593), .ZN(P3_U3181) );
  MUX2_X1 U14878 ( .A(n12596), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12598), .Z(
        P3_U3522) );
  MUX2_X1 U14879 ( .A(n12750), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12598), .Z(
        P3_U3520) );
  MUX2_X1 U14880 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12597), .S(n12612), .Z(
        P3_U3519) );
  MUX2_X1 U14881 ( .A(n12792), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12598), .Z(
        P3_U3517) );
  INV_X1 U14882 ( .A(n12806), .ZN(n12776) );
  MUX2_X1 U14883 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12776), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14884 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12791), .S(n12612), .Z(
        P3_U3515) );
  MUX2_X1 U14885 ( .A(n12803), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12598), .Z(
        P3_U3514) );
  MUX2_X1 U14886 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12818), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14887 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12860), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14888 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12599), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12884), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12600), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14891 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12883), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12601), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14893 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12602), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12603), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14895 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12604), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12605), .S(n12612), .Z(
        P3_U3503) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12606), .S(n12612), .Z(
        P3_U3502) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n15044), .S(n12612), .Z(
        P3_U3501) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12607), .S(n12612), .Z(
        P3_U3500) );
  MUX2_X1 U14900 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15045), .S(n12612), .Z(
        P3_U3499) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12608), .S(n12612), .Z(
        P3_U3498) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12609), .S(n12612), .Z(
        P3_U3497) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12610), .S(n12612), .Z(
        P3_U3496) );
  MUX2_X1 U14904 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12611), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14905 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n9585), .S(n12612), .Z(
        P3_U3494) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13008), .S(n12612), .Z(
        P3_U3493) );
  MUX2_X1 U14907 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15104), .S(n12612), .Z(
        P3_U3492) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13009), .S(n12612), .Z(
        P3_U3491) );
  NOR2_X1 U14909 ( .A1(n12620), .A2(n12614), .ZN(n12615) );
  NAND2_X1 U14910 ( .A1(n12634), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12645) );
  OAI21_X1 U14911 ( .B1(n12634), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12645), 
        .ZN(n12627) );
  AOI21_X1 U14912 ( .B1(n12616), .B2(n12627), .A(n12639), .ZN(n12638) );
  NAND2_X1 U14913 ( .A1(n12634), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12656) );
  OAI21_X1 U14914 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12634), .A(n12656), 
        .ZN(n12657) );
  XNOR2_X1 U14915 ( .A(n12658), .B(n12657), .ZN(n12636) );
  INV_X1 U14916 ( .A(n12622), .ZN(n12624) );
  OAI21_X1 U14917 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n15011) );
  MUX2_X1 U14918 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14941), .Z(n12626) );
  XNOR2_X1 U14919 ( .A(n12626), .B(n15006), .ZN(n15012) );
  NOR2_X1 U14920 ( .A1(n15011), .A2(n15012), .ZN(n15010) );
  NOR2_X1 U14921 ( .A1(n12626), .A2(n15006), .ZN(n12629) );
  MUX2_X1 U14922 ( .A(n12657), .B(n12627), .S(n6550), .Z(n12628) );
  OAI21_X1 U14923 ( .B1(n15010), .B2(n12629), .A(n12628), .ZN(n12630) );
  NAND3_X1 U14924 ( .A1(n12630), .A2(n14999), .A3(n12647), .ZN(n12633) );
  AOI21_X1 U14925 ( .B1(n14978), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12631), 
        .ZN(n12632) );
  OAI211_X1 U14926 ( .C1(n15007), .C2(n12634), .A(n12633), .B(n12632), .ZN(
        n12635) );
  AOI21_X1 U14927 ( .B1(n12732), .B2(n12636), .A(n12635), .ZN(n12637) );
  OAI21_X1 U14928 ( .B1(n12638), .B2(n15015), .A(n12637), .ZN(P3_U3196) );
  AND2_X1 U14929 ( .A1(n14566), .A2(n12640), .ZN(n12641) );
  NAND2_X1 U14930 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12674), .ZN(n12642) );
  OAI21_X1 U14931 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n12674), .A(n12642), 
        .ZN(n12643) );
  AOI21_X1 U14932 ( .B1(n12644), .B2(n12643), .A(n12671), .ZN(n12670) );
  MUX2_X1 U14933 ( .A(n12656), .B(n12645), .S(n6550), .Z(n12646) );
  NAND2_X1 U14934 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  INV_X1 U14935 ( .A(n12648), .ZN(n12649) );
  XNOR2_X1 U14936 ( .A(n12648), .B(n14566), .ZN(n14569) );
  MUX2_X1 U14937 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n14941), .Z(n14570) );
  NOR2_X1 U14938 ( .A1(n14569), .A2(n14570), .ZN(n14568) );
  AOI21_X1 U14939 ( .B1(n12649), .B2(n12660), .A(n14568), .ZN(n12681) );
  MUX2_X1 U14940 ( .A(n12918), .B(n12996), .S(n6550), .Z(n12650) );
  NOR2_X1 U14941 ( .A1(n12650), .A2(n12653), .ZN(n12680) );
  INV_X1 U14942 ( .A(n12680), .ZN(n12651) );
  NAND2_X1 U14943 ( .A1(n12650), .A2(n12653), .ZN(n12679) );
  NAND2_X1 U14944 ( .A1(n12651), .A2(n12679), .ZN(n12652) );
  XNOR2_X1 U14945 ( .A(n12681), .B(n12652), .ZN(n12668) );
  INV_X1 U14946 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U14947 ( .A1(n14981), .A2(n12653), .ZN(n12655) );
  OAI211_X1 U14948 ( .C1(n15245), .C2(n15008), .A(n12655), .B(n12654), .ZN(
        n12667) );
  INV_X1 U14949 ( .A(n12656), .ZN(n12659) );
  XNOR2_X1 U14950 ( .A(n12661), .B(n12660), .ZN(n14564) );
  NAND2_X1 U14951 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12674), .ZN(n12662) );
  OAI21_X1 U14952 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12674), .A(n12662), 
        .ZN(n12663) );
  AOI21_X1 U14953 ( .B1(n12664), .B2(n12663), .A(n12673), .ZN(n12665) );
  NOR2_X1 U14954 ( .A1(n12665), .A2(n15023), .ZN(n12666) );
  AOI211_X1 U14955 ( .C1(n14999), .C2(n12668), .A(n12667), .B(n12666), .ZN(
        n12669) );
  OAI21_X1 U14956 ( .B1(n12670), .B2(n15015), .A(n12669), .ZN(P3_U3198) );
  XNOR2_X1 U14957 ( .A(n12706), .B(n12705), .ZN(n12672) );
  AOI21_X1 U14958 ( .B1(n12992), .B2(n12672), .A(n12704), .ZN(n12687) );
  XNOR2_X1 U14959 ( .A(n12692), .B(n12705), .ZN(n12675) );
  NAND2_X1 U14960 ( .A1(n14978), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12676) );
  OAI211_X1 U14961 ( .C1(n15023), .C2(n12678), .A(n12677), .B(n12676), .ZN(
        n12685) );
  MUX2_X1 U14962 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6550), .Z(n12689) );
  XOR2_X1 U14963 ( .A(n12705), .B(n12689), .Z(n12683) );
  OAI21_X1 U14964 ( .B1(n12681), .B2(n12680), .A(n12679), .ZN(n12682) );
  NOR2_X1 U14965 ( .A1(n12682), .A2(n12683), .ZN(n12688) );
  AOI211_X1 U14966 ( .C1(n12683), .C2(n12682), .A(n15017), .B(n12688), .ZN(
        n12684) );
  AOI211_X1 U14967 ( .C1(n14981), .C2(n12705), .A(n12685), .B(n12684), .ZN(
        n12686) );
  OAI21_X1 U14968 ( .B1(n12687), .B2(n15015), .A(n12686), .ZN(P3_U3199) );
  MUX2_X1 U14969 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6550), .Z(n12691) );
  AOI21_X1 U14970 ( .B1(n12689), .B2(n12695), .A(n12688), .ZN(n12717) );
  XNOR2_X1 U14971 ( .A(n12717), .B(n12716), .ZN(n12690) );
  NOR2_X1 U14972 ( .A1(n12690), .A2(n12691), .ZN(n12715) );
  AOI21_X1 U14973 ( .B1(n12691), .B2(n12690), .A(n12715), .ZN(n12714) );
  INV_X1 U14974 ( .A(n12692), .ZN(n12694) );
  OR2_X1 U14975 ( .A1(n12716), .A2(n12887), .ZN(n12721) );
  NAND2_X1 U14976 ( .A1(n12716), .A2(n12887), .ZN(n12696) );
  NAND2_X1 U14977 ( .A1(n12721), .A2(n12696), .ZN(n12697) );
  NOR2_X1 U14978 ( .A1(n12698), .A2(n12697), .ZN(n12723) );
  NOR2_X1 U14979 ( .A1(n12723), .A2(n12699), .ZN(n12702) );
  AOI21_X1 U14980 ( .B1(n14978), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12700), 
        .ZN(n12701) );
  OAI21_X1 U14981 ( .B1(n15023), .B2(n12702), .A(n12701), .ZN(n12703) );
  OR2_X1 U14982 ( .A1(n12706), .A2(n12705), .ZN(n12710) );
  INV_X1 U14983 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12707) );
  OR2_X1 U14984 ( .A1(n12716), .A2(n12707), .ZN(n12733) );
  NAND2_X1 U14985 ( .A1(n12716), .A2(n12707), .ZN(n12708) );
  NAND2_X1 U14986 ( .A1(n12733), .A2(n12708), .ZN(n12709) );
  AND3_X1 U14987 ( .A1(n7119), .A2(n12710), .A3(n12709), .ZN(n12711) );
  OAI21_X1 U14988 ( .B1(n12734), .B2(n12711), .A(n12737), .ZN(n12712) );
  OAI211_X1 U14989 ( .C1(n12714), .C2(n15017), .A(n12713), .B(n12712), .ZN(
        P3_U3200) );
  AOI21_X1 U14990 ( .B1(n12717), .B2(n12716), .A(n12715), .ZN(n12720) );
  XNOR2_X1 U14991 ( .A(n6555), .B(n12878), .ZN(n12724) );
  XNOR2_X1 U14992 ( .A(n6555), .B(n12984), .ZN(n12735) );
  MUX2_X1 U14993 ( .A(n12724), .B(n12735), .S(n14941), .Z(n12719) );
  XNOR2_X1 U14994 ( .A(n12720), .B(n12719), .ZN(n12741) );
  INV_X1 U14995 ( .A(n12721), .ZN(n12722) );
  NOR2_X1 U14996 ( .A1(n12723), .A2(n12722), .ZN(n12726) );
  INV_X1 U14997 ( .A(n12724), .ZN(n12725) );
  NOR2_X1 U14998 ( .A1(n15007), .A2(n6555), .ZN(n12731) );
  OAI21_X1 U14999 ( .B1(n15008), .B2(n12729), .A(n12728), .ZN(n12730) );
  INV_X1 U15000 ( .A(n12735), .ZN(n12736) );
  NAND2_X1 U15001 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  OAI211_X1 U15002 ( .C1(n12741), .C2(n15017), .A(n12740), .B(n12739), .ZN(
        P3_U3201) );
  NOR2_X1 U15003 ( .A1(n12743), .A2(n12742), .ZN(n13021) );
  INV_X1 U15004 ( .A(n13021), .ZN(n12939) );
  OAI21_X1 U15005 ( .B1(n12939), .B2(n15038), .A(n12744), .ZN(n12746) );
  AOI21_X1 U15006 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15038), .A(n12746), 
        .ZN(n12745) );
  OAI21_X1 U15007 ( .B1(n13023), .B2(n12934), .A(n12745), .ZN(P3_U3202) );
  AOI21_X1 U15008 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15038), .A(n12746), 
        .ZN(n12747) );
  OAI21_X1 U15009 ( .B1(n13026), .B2(n12934), .A(n12747), .ZN(P3_U3203) );
  OAI211_X1 U15010 ( .C1(n12749), .C2(n12754), .A(n12748), .B(n15039), .ZN(
        n12751) );
  INV_X1 U15011 ( .A(n12943), .ZN(n12759) );
  AOI22_X1 U15012 ( .A1(n12755), .A2(n15125), .B1(n15038), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12756) );
  OAI21_X1 U15013 ( .B1(n13029), .B2(n12934), .A(n12756), .ZN(n12757) );
  AOI21_X1 U15014 ( .B1(n12944), .B2(n15079), .A(n12757), .ZN(n12758) );
  OAI21_X1 U15015 ( .B1(n12759), .B2(n15038), .A(n12758), .ZN(P3_U3205) );
  AOI21_X1 U15016 ( .B1(n12763), .B2(n12761), .A(n12760), .ZN(n12769) );
  OAI22_X1 U15017 ( .A1(n12766), .A2(n15105), .B1(n12765), .B2(n15107), .ZN(
        n12767) );
  AOI21_X1 U15018 ( .B1(n12948), .B2(n15115), .A(n12767), .ZN(n12768) );
  INV_X1 U15019 ( .A(n12947), .ZN(n12774) );
  AOI22_X1 U15020 ( .A1(n12770), .A2(n15125), .B1(n15038), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12771) );
  OAI21_X1 U15021 ( .B1(n13032), .B2(n12934), .A(n12771), .ZN(n12772) );
  AOI21_X1 U15022 ( .B1(n12948), .B2(n15126), .A(n12772), .ZN(n12773) );
  OAI21_X1 U15023 ( .B1(n12774), .B2(n15038), .A(n12773), .ZN(P3_U3206) );
  XNOR2_X1 U15024 ( .A(n12775), .B(n12778), .ZN(n12782) );
  AOI22_X1 U15025 ( .A1(n12777), .A2(n15043), .B1(n12776), .B2(n15046), .ZN(
        n12781) );
  XNOR2_X1 U15026 ( .A(n12779), .B(n12778), .ZN(n12952) );
  NAND2_X1 U15027 ( .A1(n12952), .A2(n15115), .ZN(n12780) );
  INV_X1 U15028 ( .A(n12951), .ZN(n12787) );
  AOI22_X1 U15029 ( .A1(n12783), .A2(n15125), .B1(n15038), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12784) );
  OAI21_X1 U15030 ( .B1(n13036), .B2(n12934), .A(n12784), .ZN(n12785) );
  AOI21_X1 U15031 ( .B1(n12952), .B2(n15126), .A(n12785), .ZN(n12786) );
  OAI21_X1 U15032 ( .B1(n12787), .B2(n15038), .A(n12786), .ZN(P3_U3207) );
  OAI211_X1 U15033 ( .C1(n12790), .C2(n12789), .A(n12788), .B(n15039), .ZN(
        n12794) );
  AOI22_X1 U15034 ( .A1(n12792), .A2(n15043), .B1(n12791), .B2(n15046), .ZN(
        n12793) );
  AND2_X1 U15035 ( .A1(n12794), .A2(n12793), .ZN(n12957) );
  XNOR2_X1 U15036 ( .A(n12796), .B(n12795), .ZN(n12955) );
  AOI22_X1 U15037 ( .A1(n12797), .A2(n15125), .B1(n15038), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12798) );
  OAI21_X1 U15038 ( .B1(n13039), .B2(n12934), .A(n12798), .ZN(n12799) );
  AOI21_X1 U15039 ( .B1(n12955), .B2(n15079), .A(n12799), .ZN(n12800) );
  OAI21_X1 U15040 ( .B1(n12957), .B2(n15038), .A(n12800), .ZN(P3_U3208) );
  OAI211_X1 U15041 ( .C1(n12807), .C2(n12802), .A(n12801), .B(n15039), .ZN(
        n12805) );
  NAND2_X1 U15042 ( .A1(n12803), .A2(n15046), .ZN(n12804) );
  OAI211_X1 U15043 ( .C1(n12806), .C2(n15105), .A(n12805), .B(n12804), .ZN(
        n12960) );
  INV_X1 U15044 ( .A(n12960), .ZN(n12815) );
  OAI21_X1 U15045 ( .B1(n12809), .B2(n9529), .A(n12808), .ZN(n12961) );
  INV_X1 U15046 ( .A(n12810), .ZN(n13042) );
  AOI22_X1 U15047 ( .A1(n15038), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12811), 
        .B2(n15125), .ZN(n12812) );
  OAI21_X1 U15048 ( .B1(n13042), .B2(n12934), .A(n12812), .ZN(n12813) );
  AOI21_X1 U15049 ( .B1(n12961), .B2(n15079), .A(n12813), .ZN(n12814) );
  OAI21_X1 U15050 ( .B1(n12815), .B2(n15038), .A(n12814), .ZN(P3_U3209) );
  OAI211_X1 U15051 ( .C1(n9618), .C2(n12817), .A(n12816), .B(n15039), .ZN(
        n12820) );
  NAND2_X1 U15052 ( .A1(n12818), .A2(n15046), .ZN(n12819) );
  OAI211_X1 U15053 ( .C1(n12821), .C2(n15105), .A(n12820), .B(n12819), .ZN(
        n12964) );
  INV_X1 U15054 ( .A(n12964), .ZN(n12829) );
  XOR2_X1 U15055 ( .A(n12823), .B(n12822), .Z(n12965) );
  INV_X1 U15056 ( .A(n12824), .ZN(n13046) );
  AOI22_X1 U15057 ( .A1(n15038), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15125), 
        .B2(n12825), .ZN(n12826) );
  OAI21_X1 U15058 ( .B1(n13046), .B2(n12934), .A(n12826), .ZN(n12827) );
  AOI21_X1 U15059 ( .B1(n12965), .B2(n15079), .A(n12827), .ZN(n12828) );
  OAI21_X1 U15060 ( .B1(n12829), .B2(n15038), .A(n12828), .ZN(P3_U3210) );
  XNOR2_X1 U15061 ( .A(n12831), .B(n12830), .ZN(n12832) );
  OAI222_X1 U15062 ( .A1(n15107), .A2(n12834), .B1(n15105), .B2(n12833), .C1(
        n12832), .C2(n15110), .ZN(n12968) );
  INV_X1 U15063 ( .A(n12968), .ZN(n12842) );
  XNOR2_X1 U15064 ( .A(n12836), .B(n12835), .ZN(n12969) );
  INV_X1 U15065 ( .A(n12837), .ZN(n13050) );
  AOI22_X1 U15066 ( .A1(n15038), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15125), 
        .B2(n12838), .ZN(n12839) );
  OAI21_X1 U15067 ( .B1(n13050), .B2(n12934), .A(n12839), .ZN(n12840) );
  AOI21_X1 U15068 ( .B1(n12969), .B2(n15079), .A(n12840), .ZN(n12841) );
  OAI21_X1 U15069 ( .B1(n12842), .B2(n15038), .A(n12841), .ZN(P3_U3211) );
  XNOR2_X1 U15070 ( .A(n12843), .B(n12846), .ZN(n12844) );
  OAI222_X1 U15071 ( .A1(n15105), .A2(n12845), .B1(n15107), .B2(n12872), .C1(
        n15110), .C2(n12844), .ZN(n12972) );
  INV_X1 U15072 ( .A(n12972), .ZN(n12853) );
  XNOR2_X1 U15073 ( .A(n12847), .B(n12846), .ZN(n12973) );
  INV_X1 U15074 ( .A(n12848), .ZN(n13054) );
  AOI22_X1 U15075 ( .A1(n15038), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15125), 
        .B2(n12849), .ZN(n12850) );
  OAI21_X1 U15076 ( .B1(n13054), .B2(n12934), .A(n12850), .ZN(n12851) );
  AOI21_X1 U15077 ( .B1(n12973), .B2(n15079), .A(n12851), .ZN(n12852) );
  OAI21_X1 U15078 ( .B1(n12853), .B2(n15038), .A(n12852), .ZN(P3_U3212) );
  OAI21_X1 U15079 ( .B1(n12856), .B2(n12855), .A(n12854), .ZN(n12976) );
  OAI211_X1 U15080 ( .C1(n12859), .C2(n12858), .A(n12857), .B(n15039), .ZN(
        n12862) );
  AOI22_X1 U15081 ( .A1(n15046), .A2(n12884), .B1(n12860), .B2(n15043), .ZN(
        n12861) );
  NAND2_X1 U15082 ( .A1(n12862), .A2(n12861), .ZN(n12977) );
  NAND2_X1 U15083 ( .A1(n12977), .A2(n15129), .ZN(n12868) );
  OAI22_X1 U15084 ( .A1(n15129), .A2(n12864), .B1(n12863), .B2(n15101), .ZN(
        n12865) );
  AOI21_X1 U15085 ( .B1(n12866), .B2(n12889), .A(n12865), .ZN(n12867) );
  OAI211_X1 U15086 ( .C1(n12976), .C2(n12869), .A(n12868), .B(n12867), .ZN(
        P3_U3213) );
  AOI21_X1 U15087 ( .B1(n12870), .B2(n12871), .A(n15110), .ZN(n12875) );
  OAI22_X1 U15088 ( .A1(n12900), .A2(n15107), .B1(n12872), .B2(n15105), .ZN(
        n12873) );
  AOI21_X1 U15089 ( .B1(n12875), .B2(n12874), .A(n12873), .ZN(n12983) );
  XNOR2_X1 U15090 ( .A(n12876), .B(n9612), .ZN(n12981) );
  NOR2_X1 U15091 ( .A1(n13062), .A2(n12934), .ZN(n12880) );
  OAI22_X1 U15092 ( .A1(n15129), .A2(n12878), .B1(n12877), .B2(n15101), .ZN(
        n12879) );
  AOI211_X1 U15093 ( .C1(n12981), .C2(n15079), .A(n12880), .B(n12879), .ZN(
        n12881) );
  OAI21_X1 U15094 ( .B1(n12983), .B2(n15038), .A(n12881), .ZN(P3_U3214) );
  OAI21_X1 U15095 ( .B1(n7597), .B2(n6571), .A(n12882), .ZN(n12885) );
  AOI222_X1 U15096 ( .A1(n15039), .A2(n12885), .B1(n12884), .B2(n15043), .C1(
        n12883), .C2(n15046), .ZN(n12989) );
  OAI22_X1 U15097 ( .A1(n15129), .A2(n12887), .B1(n12886), .B2(n15101), .ZN(
        n12888) );
  AOI21_X1 U15098 ( .B1(n12986), .B2(n12889), .A(n12888), .ZN(n12894) );
  INV_X1 U15099 ( .A(n12890), .ZN(n12891) );
  AOI21_X1 U15100 ( .B1(n6571), .B2(n12892), .A(n12891), .ZN(n12987) );
  NAND2_X1 U15101 ( .A1(n12987), .A2(n15079), .ZN(n12893) );
  OAI211_X1 U15102 ( .C1(n12989), .C2(n15038), .A(n12894), .B(n12893), .ZN(
        P3_U3215) );
  OAI211_X1 U15103 ( .C1(n12897), .C2(n12896), .A(n12895), .B(n15039), .ZN(
        n12899) );
  OR2_X1 U15104 ( .A1(n12925), .A2(n15107), .ZN(n12898) );
  OAI211_X1 U15105 ( .C1(n12900), .C2(n15105), .A(n12899), .B(n12898), .ZN(
        n12990) );
  INV_X1 U15106 ( .A(n12990), .ZN(n12909) );
  XNOR2_X1 U15107 ( .A(n12902), .B(n12901), .ZN(n12991) );
  INV_X1 U15108 ( .A(n12903), .ZN(n13067) );
  NOR2_X1 U15109 ( .A1(n13067), .A2(n12934), .ZN(n12907) );
  OAI22_X1 U15110 ( .A1(n15129), .A2(n12905), .B1(n12904), .B2(n15101), .ZN(
        n12906) );
  AOI211_X1 U15111 ( .C1(n12991), .C2(n15079), .A(n12907), .B(n12906), .ZN(
        n12908) );
  OAI21_X1 U15112 ( .B1(n12909), .B2(n15038), .A(n12908), .ZN(P3_U3216) );
  XNOR2_X1 U15113 ( .A(n12910), .B(n12915), .ZN(n12911) );
  OAI222_X1 U15114 ( .A1(n15105), .A2(n12913), .B1(n15107), .B2(n12912), .C1(
        n15110), .C2(n12911), .ZN(n12994) );
  INV_X1 U15115 ( .A(n12994), .ZN(n12922) );
  OAI21_X1 U15116 ( .B1(n12916), .B2(n12915), .A(n12914), .ZN(n12995) );
  NOR2_X1 U15117 ( .A1(n13071), .A2(n12934), .ZN(n12920) );
  OAI22_X1 U15118 ( .A1(n15129), .A2(n12918), .B1(n12917), .B2(n15101), .ZN(
        n12919) );
  AOI211_X1 U15119 ( .C1(n12995), .C2(n15079), .A(n12920), .B(n12919), .ZN(
        n12921) );
  OAI21_X1 U15120 ( .B1(n12922), .B2(n15038), .A(n12921), .ZN(P3_U3217) );
  XOR2_X1 U15121 ( .A(n12928), .B(n12923), .Z(n12924) );
  OAI222_X1 U15122 ( .A1(n15105), .A2(n12925), .B1(n15107), .B2(n14591), .C1(
        n12924), .C2(n15110), .ZN(n12998) );
  INV_X1 U15123 ( .A(n12998), .ZN(n12937) );
  NAND2_X1 U15124 ( .A1(n12927), .A2(n12926), .ZN(n12929) );
  XNOR2_X1 U15125 ( .A(n12929), .B(n12928), .ZN(n12999) );
  INV_X1 U15126 ( .A(n12930), .ZN(n13075) );
  INV_X1 U15127 ( .A(n12931), .ZN(n12932) );
  AOI22_X1 U15128 ( .A1(n15038), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15125), 
        .B2(n12932), .ZN(n12933) );
  OAI21_X1 U15129 ( .B1(n13075), .B2(n12934), .A(n12933), .ZN(n12935) );
  AOI21_X1 U15130 ( .B1(n12999), .B2(n15079), .A(n12935), .ZN(n12936) );
  OAI21_X1 U15131 ( .B1(n12937), .B2(n15038), .A(n12936), .ZN(P3_U3218) );
  NOR2_X1 U15132 ( .A1(n12939), .A2(n15179), .ZN(n12941) );
  AOI21_X1 U15133 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15179), .A(n12941), 
        .ZN(n12940) );
  OAI21_X1 U15134 ( .B1(n13023), .B2(n13001), .A(n12940), .ZN(P3_U3490) );
  AOI21_X1 U15135 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15179), .A(n12941), 
        .ZN(n12942) );
  OAI21_X1 U15136 ( .B1(n13026), .B2(n13001), .A(n12942), .ZN(P3_U3489) );
  INV_X1 U15137 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12949) );
  MUX2_X1 U15138 ( .A(n12949), .B(n13030), .S(n15181), .Z(n12950) );
  MUX2_X1 U15139 ( .A(n12953), .B(n13033), .S(n15181), .Z(n12954) );
  OAI21_X1 U15140 ( .B1(n13036), .B2(n13001), .A(n12954), .ZN(P3_U3485) );
  INV_X1 U15141 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12958) );
  NAND2_X1 U15142 ( .A1(n12955), .A2(n15162), .ZN(n12956) );
  AND2_X1 U15143 ( .A1(n12957), .A2(n12956), .ZN(n13037) );
  MUX2_X1 U15144 ( .A(n12958), .B(n13037), .S(n15181), .Z(n12959) );
  OAI21_X1 U15145 ( .B1(n13039), .B2(n13001), .A(n12959), .ZN(P3_U3484) );
  INV_X1 U15146 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12962) );
  AOI21_X1 U15147 ( .B1(n15162), .B2(n12961), .A(n12960), .ZN(n13040) );
  MUX2_X1 U15148 ( .A(n12962), .B(n13040), .S(n15181), .Z(n12963) );
  OAI21_X1 U15149 ( .B1(n13042), .B2(n13001), .A(n12963), .ZN(P3_U3483) );
  INV_X1 U15150 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12966) );
  AOI21_X1 U15151 ( .B1(n12965), .B2(n15162), .A(n12964), .ZN(n13043) );
  MUX2_X1 U15152 ( .A(n12966), .B(n13043), .S(n15181), .Z(n12967) );
  OAI21_X1 U15153 ( .B1(n13046), .B2(n13001), .A(n12967), .ZN(P3_U3482) );
  INV_X1 U15154 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12970) );
  AOI21_X1 U15155 ( .B1(n12969), .B2(n15162), .A(n12968), .ZN(n13047) );
  MUX2_X1 U15156 ( .A(n12970), .B(n13047), .S(n15181), .Z(n12971) );
  OAI21_X1 U15157 ( .B1(n13050), .B2(n13001), .A(n12971), .ZN(P3_U3481) );
  AOI21_X1 U15158 ( .B1(n12973), .B2(n15162), .A(n12972), .ZN(n13051) );
  MUX2_X1 U15159 ( .A(n12974), .B(n13051), .S(n15181), .Z(n12975) );
  OAI21_X1 U15160 ( .B1(n13054), .B2(n13001), .A(n12975), .ZN(P3_U3480) );
  INV_X1 U15161 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12979) );
  INV_X1 U15162 ( .A(n12976), .ZN(n12978) );
  AOI21_X1 U15163 ( .B1(n12978), .B2(n15162), .A(n12977), .ZN(n13055) );
  MUX2_X1 U15164 ( .A(n12979), .B(n13055), .S(n15181), .Z(n12980) );
  OAI21_X1 U15165 ( .B1(n13058), .B2(n13001), .A(n12980), .ZN(P3_U3479) );
  NAND2_X1 U15166 ( .A1(n12981), .A2(n15162), .ZN(n12982) );
  AND2_X1 U15167 ( .A1(n12983), .A2(n12982), .ZN(n13059) );
  MUX2_X1 U15168 ( .A(n12984), .B(n13059), .S(n15181), .Z(n12985) );
  OAI21_X1 U15169 ( .B1(n13001), .B2(n13062), .A(n12985), .ZN(P3_U3478) );
  AOI22_X1 U15170 ( .A1(n12987), .A2(n15162), .B1(n15065), .B2(n12986), .ZN(
        n12988) );
  NAND2_X1 U15171 ( .A1(n12989), .A2(n12988), .ZN(n13063) );
  MUX2_X1 U15172 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13063), .S(n15181), .Z(
        P3_U3477) );
  AOI21_X1 U15173 ( .B1(n12991), .B2(n15162), .A(n12990), .ZN(n13064) );
  MUX2_X1 U15174 ( .A(n12992), .B(n13064), .S(n15181), .Z(n12993) );
  OAI21_X1 U15175 ( .B1(n13067), .B2(n13001), .A(n12993), .ZN(P3_U3476) );
  AOI21_X1 U15176 ( .B1(n15162), .B2(n12995), .A(n12994), .ZN(n13068) );
  MUX2_X1 U15177 ( .A(n12996), .B(n13068), .S(n15181), .Z(n12997) );
  OAI21_X1 U15178 ( .B1(n13071), .B2(n13001), .A(n12997), .ZN(P3_U3475) );
  AOI21_X1 U15179 ( .B1(n12999), .B2(n15162), .A(n12998), .ZN(n13072) );
  MUX2_X1 U15180 ( .A(n14573), .B(n13072), .S(n15181), .Z(n13000) );
  OAI21_X1 U15181 ( .B1(n13075), .B2(n13001), .A(n13000), .ZN(P3_U3474) );
  AOI22_X1 U15182 ( .A1(n13003), .A2(n15162), .B1(n15065), .B2(n13002), .ZN(
        n13004) );
  NAND2_X1 U15183 ( .A1(n13005), .A2(n13004), .ZN(n13076) );
  MUX2_X1 U15184 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13076), .S(n15181), .Z(
        P3_U3473) );
  OAI21_X1 U15185 ( .B1(n13007), .B2(n13015), .A(n13006), .ZN(n13013) );
  NAND2_X1 U15186 ( .A1(n13008), .A2(n15043), .ZN(n13011) );
  NAND2_X1 U15187 ( .A1(n13009), .A2(n15046), .ZN(n13010) );
  NAND2_X1 U15188 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  AOI21_X1 U15189 ( .B1(n13013), .B2(n15039), .A(n13012), .ZN(n13017) );
  XNOR2_X1 U15190 ( .A(n13014), .B(n13015), .ZN(n15127) );
  NAND2_X1 U15191 ( .A1(n15127), .A2(n15115), .ZN(n13016) );
  AND2_X1 U15192 ( .A1(n13017), .A2(n13016), .ZN(n15121) );
  NOR2_X1 U15193 ( .A1(n13018), .A2(n15098), .ZN(n15124) );
  AOI21_X1 U15194 ( .B1(n15127), .B2(n15168), .A(n15124), .ZN(n13019) );
  AND2_X1 U15195 ( .A1(n15121), .A2(n13019), .ZN(n15131) );
  INV_X1 U15196 ( .A(n15131), .ZN(n13020) );
  MUX2_X1 U15197 ( .A(n13020), .B(P3_REG1_REG_1__SCAN_IN), .S(n15179), .Z(
        P3_U3460) );
  NAND2_X1 U15198 ( .A1(n13021), .A2(n15170), .ZN(n13025) );
  NAND2_X1 U15199 ( .A1(n15169), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13022) );
  OAI211_X1 U15200 ( .C1(n13023), .C2(n13074), .A(n13025), .B(n13022), .ZN(
        P3_U3458) );
  NAND2_X1 U15201 ( .A1(n15169), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13024) );
  OAI211_X1 U15202 ( .C1(n13026), .C2(n13074), .A(n13025), .B(n13024), .ZN(
        P3_U3457) );
  INV_X1 U15203 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13028) );
  MUX2_X1 U15204 ( .A(n15289), .B(n13030), .S(n15170), .Z(n13031) );
  INV_X1 U15205 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13034) );
  MUX2_X1 U15206 ( .A(n13034), .B(n13033), .S(n15170), .Z(n13035) );
  OAI21_X1 U15207 ( .B1(n13036), .B2(n13074), .A(n13035), .ZN(P3_U3453) );
  INV_X1 U15208 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n15233) );
  MUX2_X1 U15209 ( .A(n13037), .B(n15233), .S(n15169), .Z(n13038) );
  OAI21_X1 U15210 ( .B1(n13039), .B2(n13074), .A(n13038), .ZN(P3_U3452) );
  INV_X1 U15211 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n15306) );
  MUX2_X1 U15212 ( .A(n15306), .B(n13040), .S(n15170), .Z(n13041) );
  OAI21_X1 U15213 ( .B1(n13042), .B2(n13074), .A(n13041), .ZN(P3_U3451) );
  INV_X1 U15214 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13044) );
  MUX2_X1 U15215 ( .A(n13044), .B(n13043), .S(n15170), .Z(n13045) );
  OAI21_X1 U15216 ( .B1(n13046), .B2(n13074), .A(n13045), .ZN(P3_U3450) );
  MUX2_X1 U15217 ( .A(n13048), .B(n13047), .S(n15170), .Z(n13049) );
  OAI21_X1 U15218 ( .B1(n13050), .B2(n13074), .A(n13049), .ZN(P3_U3449) );
  MUX2_X1 U15219 ( .A(n13052), .B(n13051), .S(n15170), .Z(n13053) );
  OAI21_X1 U15220 ( .B1(n13054), .B2(n13074), .A(n13053), .ZN(P3_U3448) );
  MUX2_X1 U15221 ( .A(n13056), .B(n13055), .S(n15170), .Z(n13057) );
  OAI21_X1 U15222 ( .B1(n13058), .B2(n13074), .A(n13057), .ZN(P3_U3447) );
  INV_X1 U15223 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13060) );
  MUX2_X1 U15224 ( .A(n13060), .B(n13059), .S(n15170), .Z(n13061) );
  OAI21_X1 U15225 ( .B1(n13074), .B2(n13062), .A(n13061), .ZN(P3_U3446) );
  MUX2_X1 U15226 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13063), .S(n15170), .Z(
        P3_U3444) );
  INV_X1 U15227 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13065) );
  MUX2_X1 U15228 ( .A(n13065), .B(n13064), .S(n15170), .Z(n13066) );
  OAI21_X1 U15229 ( .B1(n13067), .B2(n13074), .A(n13066), .ZN(P3_U3441) );
  INV_X1 U15230 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13069) );
  MUX2_X1 U15231 ( .A(n13069), .B(n13068), .S(n15170), .Z(n13070) );
  OAI21_X1 U15232 ( .B1(n13071), .B2(n13074), .A(n13070), .ZN(P3_U3438) );
  MUX2_X1 U15233 ( .A(n15434), .B(n13072), .S(n15170), .Z(n13073) );
  OAI21_X1 U15234 ( .B1(n13075), .B2(n13074), .A(n13073), .ZN(P3_U3435) );
  MUX2_X1 U15235 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13076), .S(n15170), .Z(
        P3_U3432) );
  MUX2_X1 U15236 ( .A(n13077), .B(P3_D_REG_1__SCAN_IN), .S(n13078), .Z(
        P3_U3377) );
  MUX2_X1 U15237 ( .A(n13079), .B(P3_D_REG_0__SCAN_IN), .S(n13078), .Z(
        P3_U3376) );
  NAND3_X1 U15238 ( .A1(n9165), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13081) );
  OAI22_X1 U15239 ( .A1(n13082), .A2(n13081), .B1(n13080), .B2(n13092), .ZN(
        n13083) );
  AOI21_X1 U15240 ( .B1(n13085), .B2(n13084), .A(n13083), .ZN(n13086) );
  INV_X1 U15241 ( .A(n13086), .ZN(P3_U3264) );
  INV_X1 U15242 ( .A(n13087), .ZN(n13088) );
  OAI222_X1 U15243 ( .A1(n13092), .A2(n13091), .B1(P3_U3151), .B2(n13090), 
        .C1(n13089), .C2(n13088), .ZN(P3_U3266) );
  MUX2_X1 U15244 ( .A(n13093), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15245 ( .A(n13094), .B(n13095), .ZN(n13102) );
  OR2_X1 U15246 ( .A1(n13096), .A2(n13188), .ZN(n13098) );
  NAND2_X1 U15247 ( .A1(n13212), .A2(n13518), .ZN(n13097) );
  NAND2_X1 U15248 ( .A1(n13098), .A2(n13097), .ZN(n13337) );
  AOI22_X1 U15249 ( .A1(n14635), .A2(n13337), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13099) );
  OAI21_X1 U15250 ( .B1(n13344), .B2(n14643), .A(n13099), .ZN(n13100) );
  AOI21_X1 U15251 ( .B1(n13347), .B2(n14638), .A(n13100), .ZN(n13101) );
  OAI21_X1 U15252 ( .B1(n13102), .B2(n13202), .A(n13101), .ZN(P2_U3186) );
  XNOR2_X1 U15253 ( .A(n13104), .B(n13103), .ZN(n13110) );
  NAND2_X1 U15254 ( .A1(n13216), .A2(n13518), .ZN(n13106) );
  NAND2_X1 U15255 ( .A1(n13214), .A2(n13516), .ZN(n13105) );
  NAND2_X1 U15256 ( .A1(n13106), .A2(n13105), .ZN(n13403) );
  AOI22_X1 U15257 ( .A1(n13403), .A2(n14635), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13107) );
  OAI21_X1 U15258 ( .B1(n13409), .B2(n14643), .A(n13107), .ZN(n13108) );
  AOI21_X1 U15259 ( .B1(n13408), .B2(n14638), .A(n13108), .ZN(n13109) );
  OAI21_X1 U15260 ( .B1(n13110), .B2(n13202), .A(n13109), .ZN(P2_U3188) );
  INV_X1 U15261 ( .A(n13647), .ZN(n13476) );
  OAI21_X1 U15262 ( .B1(n13113), .B2(n13112), .A(n13111), .ZN(n13114) );
  NAND2_X1 U15263 ( .A1(n13114), .A2(n14633), .ZN(n13118) );
  INV_X1 U15264 ( .A(n13115), .ZN(n13474) );
  AOI22_X1 U15265 ( .A1(n13218), .A2(n13516), .B1(n13518), .B2(n13220), .ZN(
        n13470) );
  NAND2_X1 U15266 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13295)
         );
  OAI21_X1 U15267 ( .B1(n13470), .B2(n13178), .A(n13295), .ZN(n13116) );
  AOI21_X1 U15268 ( .B1(n13474), .B2(n9845), .A(n13116), .ZN(n13117) );
  OAI211_X1 U15269 ( .C1(n13476), .C2(n13183), .A(n13118), .B(n13117), .ZN(
        P2_U3191) );
  XNOR2_X1 U15270 ( .A(n13120), .B(n13119), .ZN(n13126) );
  OAI22_X1 U15271 ( .A1(n13122), .A2(n13188), .B1(n13121), .B2(n13190), .ZN(
        n13448) );
  AOI22_X1 U15272 ( .A1(n13448), .A2(n14635), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13123) );
  OAI21_X1 U15273 ( .B1(n13439), .B2(n14643), .A(n13123), .ZN(n13124) );
  AOI21_X1 U15274 ( .B1(n13636), .B2(n14638), .A(n13124), .ZN(n13125) );
  OAI21_X1 U15275 ( .B1(n13126), .B2(n13202), .A(n13125), .ZN(P2_U3195) );
  XNOR2_X1 U15276 ( .A(n13128), .B(n13127), .ZN(n13134) );
  NAND2_X1 U15277 ( .A1(n13214), .A2(n13518), .ZN(n13130) );
  NAND2_X1 U15278 ( .A1(n13212), .A2(n13516), .ZN(n13129) );
  NAND2_X1 U15279 ( .A1(n13130), .A2(n13129), .ZN(n13370) );
  AOI22_X1 U15280 ( .A1(n14635), .A2(n13370), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13131) );
  OAI21_X1 U15281 ( .B1(n13375), .B2(n14643), .A(n13131), .ZN(n13132) );
  AOI21_X1 U15282 ( .B1(n13696), .B2(n14638), .A(n13132), .ZN(n13133) );
  OAI21_X1 U15283 ( .B1(n13134), .B2(n13202), .A(n13133), .ZN(P2_U3197) );
  OAI21_X1 U15284 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(n13138) );
  NAND2_X1 U15285 ( .A1(n13138), .A2(n14633), .ZN(n13146) );
  INV_X1 U15286 ( .A(n13501), .ZN(n13144) );
  OAI22_X1 U15287 ( .A1(n13140), .A2(n13188), .B1(n13139), .B2(n13190), .ZN(
        n13496) );
  INV_X1 U15288 ( .A(n13496), .ZN(n13142) );
  OAI22_X1 U15289 ( .A1(n13178), .A2(n13142), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13141), .ZN(n13143) );
  AOI21_X1 U15290 ( .B1(n13144), .B2(n9845), .A(n13143), .ZN(n13145) );
  OAI211_X1 U15291 ( .C1(n13504), .C2(n13183), .A(n13146), .B(n13145), .ZN(
        P2_U3200) );
  XNOR2_X1 U15292 ( .A(n13148), .B(n13147), .ZN(n13153) );
  OAI22_X1 U15293 ( .A1(n13149), .A2(n13190), .B1(n13191), .B2(n13188), .ZN(
        n13388) );
  AOI22_X1 U15294 ( .A1(n13388), .A2(n14635), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13150) );
  OAI21_X1 U15295 ( .B1(n13391), .B2(n14643), .A(n13150), .ZN(n13151) );
  AOI21_X1 U15296 ( .B1(n13620), .B2(n14638), .A(n13151), .ZN(n13152) );
  OAI21_X1 U15297 ( .B1(n13153), .B2(n13202), .A(n13152), .ZN(P2_U3201) );
  INV_X1 U15298 ( .A(n13154), .ZN(n13156) );
  NAND2_X1 U15299 ( .A1(n13156), .A2(n13155), .ZN(n13157) );
  XNOR2_X1 U15300 ( .A(n13158), .B(n13157), .ZN(n13163) );
  AOI22_X1 U15301 ( .A1(n13217), .A2(n13516), .B1(n13518), .B2(n13219), .ZN(
        n13456) );
  OAI22_X1 U15302 ( .A1(n13456), .A2(n13178), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13159), .ZN(n13160) );
  AOI21_X1 U15303 ( .B1(n13461), .B2(n9845), .A(n13160), .ZN(n13162) );
  NAND2_X1 U15304 ( .A1(n13642), .A2(n14638), .ZN(n13161) );
  OAI211_X1 U15305 ( .C1(n13163), .C2(n13202), .A(n13162), .B(n13161), .ZN(
        P2_U3205) );
  XNOR2_X1 U15306 ( .A(n13165), .B(n13164), .ZN(n13171) );
  NOR2_X1 U15307 ( .A1(n14643), .A2(n13429), .ZN(n13169) );
  AND2_X1 U15308 ( .A1(n13217), .A2(n13518), .ZN(n13166) );
  AOI21_X1 U15309 ( .B1(n13215), .B2(n13516), .A(n13166), .ZN(n13420) );
  OAI22_X1 U15310 ( .A1(n13420), .A2(n13178), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13167), .ZN(n13168) );
  AOI211_X1 U15311 ( .C1(n13705), .C2(n14638), .A(n13169), .B(n13168), .ZN(
        n13170) );
  OAI21_X1 U15312 ( .B1(n13171), .B2(n13202), .A(n13170), .ZN(P2_U3207) );
  INV_X1 U15313 ( .A(n13651), .ZN(n13487) );
  AOI21_X1 U15314 ( .B1(n13173), .B2(n13172), .A(n13202), .ZN(n13175) );
  NAND2_X1 U15315 ( .A1(n13175), .A2(n13174), .ZN(n13182) );
  OAI22_X1 U15316 ( .A1(n13177), .A2(n13188), .B1(n13176), .B2(n13190), .ZN(
        n13481) );
  INV_X1 U15317 ( .A(n13481), .ZN(n13179) );
  OAI22_X1 U15318 ( .A1(n13179), .A2(n13178), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15292), .ZN(n13180) );
  AOI21_X1 U15319 ( .B1(n13484), .B2(n9845), .A(n13180), .ZN(n13181) );
  OAI211_X1 U15320 ( .C1(n13487), .C2(n13183), .A(n13182), .B(n13181), .ZN(
        P2_U3210) );
  INV_X1 U15321 ( .A(n13184), .ZN(n13185) );
  AOI21_X1 U15322 ( .B1(n13187), .B2(n13186), .A(n13185), .ZN(n13195) );
  OAI22_X1 U15323 ( .A1(n13191), .A2(n13190), .B1(n13189), .B2(n13188), .ZN(
        n13358) );
  AOI22_X1 U15324 ( .A1(n14635), .A2(n13358), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13192) );
  OAI21_X1 U15325 ( .B1(n13353), .B2(n14643), .A(n13192), .ZN(n13193) );
  AOI21_X1 U15326 ( .B1(n13361), .B2(n14638), .A(n13193), .ZN(n13194) );
  OAI21_X1 U15327 ( .B1(n13195), .B2(n13202), .A(n13194), .ZN(P2_U3212) );
  NAND2_X1 U15328 ( .A1(n13221), .A2(n13516), .ZN(n13197) );
  NAND2_X1 U15329 ( .A1(n13222), .A2(n13518), .ZN(n13196) );
  NAND2_X1 U15330 ( .A1(n13197), .A2(n13196), .ZN(n13665) );
  NAND2_X1 U15331 ( .A1(n14635), .A2(n13665), .ZN(n13198) );
  NAND2_X1 U15332 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14849)
         );
  OAI211_X1 U15333 ( .C1(n14643), .C2(n13538), .A(n13198), .B(n14849), .ZN(
        n13206) );
  INV_X1 U15334 ( .A(n13199), .ZN(n13200) );
  NAND2_X1 U15335 ( .A1(n13201), .A2(n13200), .ZN(n14625) );
  XNOR2_X1 U15336 ( .A(n14625), .B(n14626), .ZN(n13204) );
  NOR2_X1 U15337 ( .A1(n13204), .A2(n13203), .ZN(n14627) );
  AOI211_X1 U15338 ( .C1(n13204), .C2(n13203), .A(n13202), .B(n14627), .ZN(
        n13205) );
  AOI211_X1 U15339 ( .C1(n13715), .C2(n14638), .A(n13206), .B(n13205), .ZN(
        n13207) );
  INV_X1 U15340 ( .A(n13207), .ZN(P2_U3213) );
  MUX2_X1 U15341 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13302), .S(n6554), .Z(
        P2_U3562) );
  MUX2_X1 U15342 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13208), .S(n6554), .Z(
        P2_U3561) );
  MUX2_X1 U15343 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13209), .S(n6554), .Z(
        P2_U3560) );
  MUX2_X1 U15344 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13210), .S(n6554), .Z(
        P2_U3559) );
  MUX2_X1 U15345 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13211), .S(n6554), .Z(
        P2_U3558) );
  MUX2_X1 U15346 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13212), .S(n6554), .Z(
        P2_U3557) );
  MUX2_X1 U15347 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13213), .S(n6554), .Z(
        P2_U3556) );
  MUX2_X1 U15348 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13214), .S(n6554), .Z(
        P2_U3555) );
  MUX2_X1 U15349 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13215), .S(n6554), .Z(
        P2_U3554) );
  MUX2_X1 U15350 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13216), .S(n6554), .Z(
        P2_U3553) );
  MUX2_X1 U15351 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13217), .S(n6554), .Z(
        P2_U3552) );
  MUX2_X1 U15352 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13218), .S(n6554), .Z(
        P2_U3551) );
  MUX2_X1 U15353 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13219), .S(n6554), .Z(
        P2_U3550) );
  MUX2_X1 U15354 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13220), .S(n6554), .Z(
        P2_U3549) );
  MUX2_X1 U15355 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13517), .S(n6554), .Z(
        P2_U3548) );
  MUX2_X1 U15356 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13221), .S(n6554), .Z(
        P2_U3547) );
  MUX2_X1 U15357 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13519), .S(n6554), .Z(
        P2_U3546) );
  MUX2_X1 U15358 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13222), .S(n6554), .Z(
        P2_U3545) );
  MUX2_X1 U15359 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13223), .S(n6554), .Z(
        P2_U3544) );
  MUX2_X1 U15360 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13224), .S(n6554), .Z(
        P2_U3543) );
  MUX2_X1 U15361 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13225), .S(n6554), .Z(
        P2_U3542) );
  MUX2_X1 U15362 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13226), .S(n6554), .Z(
        P2_U3541) );
  MUX2_X1 U15363 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13227), .S(n6554), .Z(
        P2_U3540) );
  MUX2_X1 U15364 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13228), .S(n6554), .Z(
        P2_U3539) );
  MUX2_X1 U15365 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13229), .S(n6554), .Z(
        P2_U3538) );
  MUX2_X1 U15366 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13230), .S(n6554), .Z(
        P2_U3537) );
  MUX2_X1 U15367 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13231), .S(n6554), .Z(
        P2_U3536) );
  MUX2_X1 U15368 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13232), .S(n6554), .Z(
        P2_U3535) );
  MUX2_X1 U15369 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13233), .S(n6554), .Z(
        P2_U3534) );
  MUX2_X1 U15370 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13234), .S(n6554), .Z(
        P2_U3533) );
  MUX2_X1 U15371 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8764), .S(n6554), .Z(
        P2_U3532) );
  MUX2_X1 U15372 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n7655), .S(n6554), .Z(
        P2_U3531) );
  INV_X1 U15373 ( .A(n13235), .ZN(n13236) );
  AOI21_X1 U15374 ( .B1(n14855), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n13236), .ZN(
        n13248) );
  OAI211_X1 U15375 ( .C1(n13239), .C2(n13238), .A(n14833), .B(n13237), .ZN(
        n13247) );
  NAND2_X1 U15376 ( .A1(n14838), .A2(n13240), .ZN(n13246) );
  MUX2_X1 U15377 ( .A(n11136), .B(P2_REG2_REG_7__SCAN_IN), .S(n13240), .Z(
        n13241) );
  NAND3_X1 U15378 ( .A1(n13243), .A2(n13242), .A3(n13241), .ZN(n13244) );
  NAND3_X1 U15379 ( .A1(n14857), .A2(n13255), .A3(n13244), .ZN(n13245) );
  NAND4_X1 U15380 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        P2_U3221) );
  AND2_X1 U15381 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13249) );
  AOI21_X1 U15382 ( .B1(n14855), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n13249), .ZN(
        n13262) );
  OAI211_X1 U15383 ( .C1(n13252), .C2(n13251), .A(n14833), .B(n13250), .ZN(
        n13261) );
  MUX2_X1 U15384 ( .A(n11105), .B(P2_REG2_REG_8__SCAN_IN), .S(n13258), .Z(
        n13253) );
  NAND3_X1 U15385 ( .A1(n13255), .A2(n13254), .A3(n13253), .ZN(n13256) );
  NAND3_X1 U15386 ( .A1(n14857), .A2(n13257), .A3(n13256), .ZN(n13260) );
  NAND2_X1 U15387 ( .A1(n14838), .A2(n13258), .ZN(n13259) );
  NAND4_X1 U15388 ( .A1(n13262), .A2(n13261), .A3(n13260), .A4(n13259), .ZN(
        P2_U3222) );
  INV_X1 U15389 ( .A(n13263), .ZN(n13265) );
  NAND2_X1 U15390 ( .A1(n13265), .A2(n13264), .ZN(n13266) );
  OAI21_X1 U15391 ( .B1(n13502), .B2(n13267), .A(n13266), .ZN(n13282) );
  XNOR2_X1 U15392 ( .A(n13283), .B(n13282), .ZN(n13268) );
  NOR2_X1 U15393 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13268), .ZN(n13284) );
  AOI21_X1 U15394 ( .B1(n13268), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13284), 
        .ZN(n13276) );
  NOR2_X1 U15395 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15292), .ZN(n13273) );
  AOI21_X1 U15396 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n13270), .A(n13269), 
        .ZN(n13278) );
  XNOR2_X1 U15397 ( .A(n13277), .B(n13278), .ZN(n13271) );
  NOR2_X1 U15398 ( .A1(n15350), .A2(n13271), .ZN(n13280) );
  AOI211_X1 U15399 ( .C1(n13271), .C2(n15350), .A(n13280), .B(n14850), .ZN(
        n13272) );
  AOI211_X1 U15400 ( .C1(n14838), .C2(n13283), .A(n13273), .B(n13272), .ZN(
        n13275) );
  NAND2_X1 U15401 ( .A1(n14855), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13274) );
  OAI211_X1 U15402 ( .C1(n13276), .C2(n14825), .A(n13275), .B(n13274), .ZN(
        P2_U3232) );
  NOR2_X1 U15403 ( .A1(n13278), .A2(n13277), .ZN(n13279) );
  NOR2_X1 U15404 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  XOR2_X1 U15405 ( .A(n13281), .B(n15450), .Z(n13291) );
  NOR2_X1 U15406 ( .A1(n13283), .A2(n13282), .ZN(n13285) );
  NOR2_X1 U15407 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  XNOR2_X1 U15408 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13286), .ZN(n13289) );
  NAND2_X1 U15409 ( .A1(n13289), .A2(n14857), .ZN(n13287) );
  OAI211_X1 U15410 ( .C1(n13291), .C2(n14850), .A(n14862), .B(n13287), .ZN(
        n13288) );
  INV_X1 U15411 ( .A(n13288), .ZN(n13294) );
  INV_X1 U15412 ( .A(n13289), .ZN(n13290) );
  AOI22_X1 U15413 ( .A1(n13291), .A2(n14833), .B1(n14857), .B2(n13290), .ZN(
        n13293) );
  MUX2_X1 U15414 ( .A(n13294), .B(n13293), .S(n13292), .Z(n13296) );
  OAI211_X1 U15415 ( .C1(n13297), .C2(n14848), .A(n13296), .B(n13295), .ZN(
        P2_U3233) );
  INV_X1 U15416 ( .A(n13298), .ZN(n13307) );
  NAND2_X1 U15417 ( .A1(n13307), .A2(n13684), .ZN(n13306) );
  XNOR2_X1 U15418 ( .A(n13299), .B(n13306), .ZN(n13300) );
  NOR2_X2 U15419 ( .A1(n13300), .A2(n9813), .ZN(n13588) );
  NAND2_X1 U15420 ( .A1(n13588), .A2(n13581), .ZN(n13305) );
  INV_X1 U15421 ( .A(n13301), .ZN(n13303) );
  AND2_X1 U15422 ( .A1(n13303), .A2(n13302), .ZN(n13587) );
  INV_X1 U15423 ( .A(n13587), .ZN(n13591) );
  NOR2_X1 U15424 ( .A1(n13552), .A2(n13591), .ZN(n13309) );
  AOI21_X1 U15425 ( .B1(n13552), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13309), 
        .ZN(n13304) );
  OAI211_X1 U15426 ( .C1(n13680), .C2(n13486), .A(n13305), .B(n13304), .ZN(
        P2_U3234) );
  OAI211_X1 U15427 ( .C1(n13307), .C2(n13684), .A(n13528), .B(n13306), .ZN(
        n13592) );
  NOR2_X1 U15428 ( .A1(n13557), .A2(n13308), .ZN(n13310) );
  AOI211_X1 U15429 ( .C1(n13311), .C2(n13577), .A(n13310), .B(n13309), .ZN(
        n13312) );
  OAI21_X1 U15430 ( .B1(n13592), .B2(n13549), .A(n13312), .ZN(P2_U3235) );
  OAI22_X1 U15431 ( .A1(n13557), .A2(n13314), .B1(n13573), .B2(n13313), .ZN(
        n13315) );
  AOI21_X1 U15432 ( .B1(n13316), .B2(n13577), .A(n13315), .ZN(n13317) );
  OAI21_X1 U15433 ( .B1(n13318), .B2(n13549), .A(n13317), .ZN(n13319) );
  AOI21_X1 U15434 ( .B1(n13320), .B2(n13579), .A(n13319), .ZN(n13321) );
  OAI21_X1 U15435 ( .B1(n13322), .B2(n13552), .A(n13321), .ZN(P2_U3236) );
  AOI21_X1 U15436 ( .B1(n13323), .B2(n13330), .A(n13562), .ZN(n13326) );
  AOI21_X1 U15437 ( .B1(n13326), .B2(n13325), .A(n13324), .ZN(n13600) );
  AOI211_X1 U15438 ( .C1(n13598), .C2(n6954), .A(n9813), .B(n13327), .ZN(
        n13597) );
  AOI22_X1 U15439 ( .A1(n13552), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n9846), 
        .B2(n13544), .ZN(n13329) );
  OAI21_X1 U15440 ( .B1(n7422), .B2(n13486), .A(n13329), .ZN(n13333) );
  XNOR2_X1 U15441 ( .A(n13331), .B(n13330), .ZN(n13601) );
  NOR2_X1 U15442 ( .A1(n13601), .A2(n13509), .ZN(n13332) );
  AOI211_X1 U15443 ( .C1(n13581), .C2(n13597), .A(n13333), .B(n13332), .ZN(
        n13334) );
  OAI21_X1 U15444 ( .B1(n13600), .B2(n13552), .A(n13334), .ZN(P2_U3237) );
  INV_X1 U15445 ( .A(n13337), .ZN(n13338) );
  OAI21_X1 U15446 ( .B1(n13339), .B2(n13562), .A(n13338), .ZN(n13603) );
  INV_X1 U15447 ( .A(n13603), .ZN(n13351) );
  XOR2_X1 U15448 ( .A(n13341), .B(n13340), .Z(n13605) );
  OAI21_X1 U15449 ( .B1(n13689), .B2(n13364), .A(n13528), .ZN(n13342) );
  OR2_X1 U15450 ( .A1(n13343), .A2(n13342), .ZN(n13602) );
  OAI22_X1 U15451 ( .A1(n13557), .A2(n13345), .B1(n13344), .B2(n13573), .ZN(
        n13346) );
  AOI21_X1 U15452 ( .B1(n13347), .B2(n13577), .A(n13346), .ZN(n13348) );
  OAI21_X1 U15453 ( .B1(n13602), .B2(n13549), .A(n13348), .ZN(n13349) );
  AOI21_X1 U15454 ( .B1(n13605), .B2(n13579), .A(n13349), .ZN(n13350) );
  OAI21_X1 U15455 ( .B1(n13351), .B2(n13552), .A(n13350), .ZN(P2_U3238) );
  XNOR2_X1 U15456 ( .A(n13352), .B(n13356), .ZN(n13610) );
  NAND2_X1 U15457 ( .A1(n13610), .A2(n13579), .ZN(n13368) );
  OAI22_X1 U15458 ( .A1(n13557), .A2(n13354), .B1(n13353), .B2(n13573), .ZN(
        n13355) );
  AOI21_X1 U15459 ( .B1(n13361), .B2(n13577), .A(n13355), .ZN(n13367) );
  XNOR2_X1 U15460 ( .A(n13357), .B(n13356), .ZN(n13360) );
  INV_X1 U15461 ( .A(n13358), .ZN(n13359) );
  OAI21_X1 U15462 ( .B1(n13360), .B2(n13562), .A(n13359), .ZN(n13608) );
  NAND2_X1 U15463 ( .A1(n13608), .A2(n13557), .ZN(n13366) );
  NAND2_X1 U15464 ( .A1(n6614), .A2(n13361), .ZN(n13362) );
  NAND2_X1 U15465 ( .A1(n13362), .A2(n13528), .ZN(n13363) );
  NOR2_X1 U15466 ( .A1(n13364), .A2(n13363), .ZN(n13609) );
  NAND2_X1 U15467 ( .A1(n13609), .A2(n13581), .ZN(n13365) );
  NAND4_X1 U15468 ( .A1(n13368), .A2(n13367), .A3(n13366), .A4(n13365), .ZN(
        P2_U3239) );
  XNOR2_X1 U15469 ( .A(n13369), .B(n13372), .ZN(n13371) );
  AOI21_X1 U15470 ( .B1(n13371), .B2(n13540), .A(n13370), .ZN(n13615) );
  XNOR2_X1 U15471 ( .A(n13373), .B(n13372), .ZN(n13613) );
  AOI21_X1 U15472 ( .B1(n13390), .B2(n13696), .A(n9813), .ZN(n13374) );
  NAND2_X1 U15473 ( .A1(n13374), .A2(n6614), .ZN(n13614) );
  OAI22_X1 U15474 ( .A1(n13557), .A2(n13376), .B1(n13375), .B2(n13573), .ZN(
        n13377) );
  AOI21_X1 U15475 ( .B1(n13696), .B2(n13577), .A(n13377), .ZN(n13378) );
  OAI21_X1 U15476 ( .B1(n13614), .B2(n13549), .A(n13378), .ZN(n13379) );
  AOI21_X1 U15477 ( .B1(n13613), .B2(n13579), .A(n13379), .ZN(n13380) );
  OAI21_X1 U15478 ( .B1(n13552), .B2(n13615), .A(n13380), .ZN(P2_U3240) );
  OAI21_X1 U15479 ( .B1(n13383), .B2(n13382), .A(n13381), .ZN(n13389) );
  NOR2_X1 U15480 ( .A1(n13623), .A2(n6794), .ZN(n13387) );
  AOI211_X1 U15481 ( .C1(n13620), .C2(n13406), .A(n9813), .B(n6952), .ZN(
        n13619) );
  INV_X1 U15482 ( .A(n13620), .ZN(n13394) );
  INV_X1 U15483 ( .A(n13391), .ZN(n13392) );
  AOI22_X1 U15484 ( .A1(n13552), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n13392), 
        .B2(n13544), .ZN(n13393) );
  OAI21_X1 U15485 ( .B1(n13394), .B2(n13486), .A(n13393), .ZN(n13397) );
  NOR2_X1 U15486 ( .A1(n13623), .A2(n13395), .ZN(n13396) );
  AOI211_X1 U15487 ( .C1(n13619), .C2(n13581), .A(n13397), .B(n13396), .ZN(
        n13398) );
  OAI21_X1 U15488 ( .B1(n13622), .B2(n13552), .A(n13398), .ZN(P2_U3241) );
  XNOR2_X1 U15489 ( .A(n13399), .B(n13401), .ZN(n13626) );
  INV_X1 U15490 ( .A(n13626), .ZN(n13415) );
  OAI211_X1 U15491 ( .C1(n13402), .C2(n13401), .A(n13400), .B(n13540), .ZN(
        n13405) );
  INV_X1 U15492 ( .A(n13403), .ZN(n13404) );
  NAND2_X1 U15493 ( .A1(n13405), .A2(n13404), .ZN(n13625) );
  INV_X1 U15494 ( .A(n13406), .ZN(n13407) );
  AOI211_X1 U15495 ( .C1(n13408), .C2(n13426), .A(n9813), .B(n13407), .ZN(
        n13624) );
  NAND2_X1 U15496 ( .A1(n13624), .A2(n13581), .ZN(n13412) );
  INV_X1 U15497 ( .A(n13409), .ZN(n13410) );
  AOI22_X1 U15498 ( .A1(n13410), .A2(n13544), .B1(n13552), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13411) );
  OAI211_X1 U15499 ( .C1(n6939), .C2(n13486), .A(n13412), .B(n13411), .ZN(
        n13413) );
  AOI21_X1 U15500 ( .B1(n13557), .B2(n13625), .A(n13413), .ZN(n13414) );
  OAI21_X1 U15501 ( .B1(n13415), .B2(n13509), .A(n13414), .ZN(P2_U3242) );
  NAND2_X1 U15502 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  NAND3_X1 U15503 ( .A1(n13419), .A2(n13540), .A3(n13418), .ZN(n13421) );
  AND2_X1 U15504 ( .A1(n13421), .A2(n13420), .ZN(n13631) );
  NAND2_X1 U15505 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  NAND2_X1 U15506 ( .A1(n13425), .A2(n13424), .ZN(n13632) );
  INV_X1 U15507 ( .A(n13632), .ZN(n13433) );
  AOI21_X1 U15508 ( .B1(n13705), .B2(n13436), .A(n9813), .ZN(n13427) );
  NAND2_X1 U15509 ( .A1(n13427), .A2(n13426), .ZN(n13630) );
  INV_X1 U15510 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13428) );
  OAI22_X1 U15511 ( .A1(n13429), .A2(n13573), .B1(n13557), .B2(n13428), .ZN(
        n13430) );
  AOI21_X1 U15512 ( .B1(n13705), .B2(n13577), .A(n13430), .ZN(n13431) );
  OAI21_X1 U15513 ( .B1(n13630), .B2(n13549), .A(n13431), .ZN(n13432) );
  AOI21_X1 U15514 ( .B1(n13433), .B2(n13579), .A(n13432), .ZN(n13434) );
  OAI21_X1 U15515 ( .B1(n13552), .B2(n13631), .A(n13434), .ZN(P2_U3243) );
  XOR2_X1 U15516 ( .A(n13447), .B(n13435), .Z(n13639) );
  INV_X1 U15517 ( .A(n13460), .ZN(n13438) );
  INV_X1 U15518 ( .A(n13436), .ZN(n13437) );
  AOI211_X1 U15519 ( .C1(n13636), .C2(n13438), .A(n9813), .B(n13437), .ZN(
        n13635) );
  INV_X1 U15520 ( .A(n13439), .ZN(n13440) );
  AOI22_X1 U15521 ( .A1(n13552), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13440), 
        .B2(n13544), .ZN(n13441) );
  OAI21_X1 U15522 ( .B1(n13442), .B2(n13486), .A(n13441), .ZN(n13451) );
  OAI21_X1 U15523 ( .B1(n13455), .B2(n13454), .A(n13445), .ZN(n13446) );
  XOR2_X1 U15524 ( .A(n13447), .B(n13446), .Z(n13449) );
  AOI21_X1 U15525 ( .B1(n13449), .B2(n13540), .A(n13448), .ZN(n13638) );
  NOR2_X1 U15526 ( .A1(n13638), .A2(n13552), .ZN(n13450) );
  AOI211_X1 U15527 ( .C1(n13635), .C2(n13581), .A(n13451), .B(n13450), .ZN(
        n13452) );
  OAI21_X1 U15528 ( .B1(n13509), .B2(n13639), .A(n13452), .ZN(P2_U3244) );
  XNOR2_X1 U15529 ( .A(n13453), .B(n13454), .ZN(n13644) );
  XOR2_X1 U15530 ( .A(n13455), .B(n13454), .Z(n13457) );
  OAI21_X1 U15531 ( .B1(n13457), .B2(n13562), .A(n13456), .ZN(n13640) );
  INV_X1 U15532 ( .A(n13642), .ZN(n13464) );
  NAND2_X1 U15533 ( .A1(n13472), .A2(n13642), .ZN(n13458) );
  NAND2_X1 U15534 ( .A1(n13458), .A2(n13528), .ZN(n13459) );
  NOR2_X1 U15535 ( .A1(n13460), .A2(n13459), .ZN(n13641) );
  NAND2_X1 U15536 ( .A1(n13641), .A2(n13581), .ZN(n13463) );
  AOI22_X1 U15537 ( .A1(n13552), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13461), 
        .B2(n13544), .ZN(n13462) );
  OAI211_X1 U15538 ( .C1(n13464), .C2(n13486), .A(n13463), .B(n13462), .ZN(
        n13465) );
  AOI21_X1 U15539 ( .B1(n13640), .B2(n13557), .A(n13465), .ZN(n13466) );
  OAI21_X1 U15540 ( .B1(n13644), .B2(n13509), .A(n13466), .ZN(P2_U3245) );
  XNOR2_X1 U15541 ( .A(n13467), .B(n13468), .ZN(n13649) );
  XOR2_X1 U15542 ( .A(n13469), .B(n13468), .Z(n13471) );
  OAI21_X1 U15543 ( .B1(n13471), .B2(n13562), .A(n13470), .ZN(n13645) );
  NAND2_X1 U15544 ( .A1(n13645), .A2(n13557), .ZN(n13479) );
  INV_X1 U15545 ( .A(n13472), .ZN(n13473) );
  AOI211_X1 U15546 ( .C1(n13647), .C2(n13483), .A(n9813), .B(n13473), .ZN(
        n13646) );
  AOI22_X1 U15547 ( .A1(n13552), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13474), 
        .B2(n13544), .ZN(n13475) );
  OAI21_X1 U15548 ( .B1(n13476), .B2(n13486), .A(n13475), .ZN(n13477) );
  AOI21_X1 U15549 ( .B1(n13646), .B2(n13581), .A(n13477), .ZN(n13478) );
  OAI211_X1 U15550 ( .C1(n13509), .C2(n13649), .A(n13479), .B(n13478), .ZN(
        P2_U3246) );
  XNOR2_X1 U15551 ( .A(n13480), .B(n13491), .ZN(n13482) );
  AOI21_X1 U15552 ( .B1(n13482), .B2(n13540), .A(n13481), .ZN(n13653) );
  AOI211_X1 U15553 ( .C1(n13651), .C2(n13506), .A(n9813), .B(n6935), .ZN(
        n13650) );
  AOI22_X1 U15554 ( .A1(n13552), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13484), 
        .B2(n13544), .ZN(n13485) );
  OAI21_X1 U15555 ( .B1(n13487), .B2(n13486), .A(n13485), .ZN(n13493) );
  INV_X1 U15556 ( .A(n13488), .ZN(n13489) );
  AOI21_X1 U15557 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(n13654) );
  NOR2_X1 U15558 ( .A1(n13654), .A2(n13509), .ZN(n13492) );
  AOI211_X1 U15559 ( .C1(n13650), .C2(n13581), .A(n13493), .B(n13492), .ZN(
        n13494) );
  OAI21_X1 U15560 ( .B1(n13552), .B2(n13653), .A(n13494), .ZN(P2_U3247) );
  XNOR2_X1 U15561 ( .A(n13495), .B(n13499), .ZN(n13497) );
  AOI21_X1 U15562 ( .B1(n13497), .B2(n13540), .A(n13496), .ZN(n13658) );
  OAI21_X1 U15563 ( .B1(n13500), .B2(n13499), .A(n13498), .ZN(n13659) );
  OAI22_X1 U15564 ( .A1(n13557), .A2(n13502), .B1(n13501), .B2(n13573), .ZN(
        n13503) );
  AOI21_X1 U15565 ( .B1(n13656), .B2(n13577), .A(n13503), .ZN(n13508) );
  OR2_X1 U15566 ( .A1(n13504), .A2(n13531), .ZN(n13505) );
  AND3_X1 U15567 ( .A1(n13506), .A2(n13505), .A3(n13528), .ZN(n13655) );
  NAND2_X1 U15568 ( .A1(n13655), .A2(n13581), .ZN(n13507) );
  OAI211_X1 U15569 ( .C1(n13659), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        n13510) );
  INV_X1 U15570 ( .A(n13510), .ZN(n13511) );
  OAI21_X1 U15571 ( .B1(n13552), .B2(n13658), .A(n13511), .ZN(P2_U3248) );
  NAND2_X1 U15572 ( .A1(n13513), .A2(n13512), .ZN(n13514) );
  NAND3_X1 U15573 ( .A1(n13515), .A2(n13540), .A3(n13514), .ZN(n13523) );
  NAND2_X1 U15574 ( .A1(n13517), .A2(n13516), .ZN(n13521) );
  NAND2_X1 U15575 ( .A1(n13519), .A2(n13518), .ZN(n13520) );
  NAND2_X1 U15576 ( .A1(n13521), .A2(n13520), .ZN(n14636) );
  INV_X1 U15577 ( .A(n14636), .ZN(n13522) );
  AND2_X1 U15578 ( .A1(n13523), .A2(n13522), .ZN(n13661) );
  NAND2_X1 U15579 ( .A1(n13525), .A2(n13524), .ZN(n13526) );
  NAND2_X1 U15580 ( .A1(n13527), .A2(n13526), .ZN(n13662) );
  INV_X1 U15581 ( .A(n13662), .ZN(n13536) );
  NAND2_X1 U15582 ( .A1(n14637), .A2(n6594), .ZN(n13529) );
  NAND2_X1 U15583 ( .A1(n13529), .A2(n13528), .ZN(n13530) );
  OR2_X1 U15584 ( .A1(n13531), .A2(n13530), .ZN(n13660) );
  OAI22_X1 U15585 ( .A1(n13557), .A2(n13532), .B1(n14642), .B2(n13573), .ZN(
        n13533) );
  AOI21_X1 U15586 ( .B1(n14637), .B2(n13577), .A(n13533), .ZN(n13534) );
  OAI21_X1 U15587 ( .B1(n13660), .B2(n13549), .A(n13534), .ZN(n13535) );
  AOI21_X1 U15588 ( .B1(n13536), .B2(n13579), .A(n13535), .ZN(n13537) );
  OAI21_X1 U15589 ( .B1(n13552), .B2(n13661), .A(n13537), .ZN(P2_U3249) );
  INV_X1 U15590 ( .A(n13538), .ZN(n13543) );
  XNOR2_X1 U15591 ( .A(n13539), .B(n13545), .ZN(n13541) );
  NAND2_X1 U15592 ( .A1(n13541), .A2(n13540), .ZN(n13668) );
  INV_X1 U15593 ( .A(n13668), .ZN(n13542) );
  AOI211_X1 U15594 ( .C1(n13544), .C2(n13543), .A(n13665), .B(n13542), .ZN(
        n13553) );
  XNOR2_X1 U15595 ( .A(n13546), .B(n13545), .ZN(n13670) );
  AOI21_X1 U15596 ( .B1(n13715), .B2(n13566), .A(n9813), .ZN(n13547) );
  NAND2_X1 U15597 ( .A1(n13547), .A2(n6594), .ZN(n13666) );
  AOI22_X1 U15598 ( .A1(n13715), .A2(n13577), .B1(n13552), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n13548) );
  OAI21_X1 U15599 ( .B1(n13666), .B2(n13549), .A(n13548), .ZN(n13550) );
  AOI21_X1 U15600 ( .B1(n13670), .B2(n13579), .A(n13550), .ZN(n13551) );
  OAI21_X1 U15601 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(P2_U3250) );
  XOR2_X1 U15602 ( .A(n13559), .B(n13554), .Z(n13674) );
  NAND2_X1 U15603 ( .A1(n13674), .A2(n13579), .ZN(n13571) );
  OAI22_X1 U15604 ( .A1(n13557), .A2(n13556), .B1(n13555), .B2(n13573), .ZN(
        n13558) );
  AOI21_X1 U15605 ( .B1(n13718), .B2(n13577), .A(n13558), .ZN(n13570) );
  XNOR2_X1 U15606 ( .A(n13560), .B(n13559), .ZN(n13563) );
  OAI21_X1 U15607 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13672) );
  NAND2_X1 U15608 ( .A1(n13672), .A2(n13557), .ZN(n13569) );
  AOI21_X1 U15609 ( .B1(n13718), .B2(n13565), .A(n13564), .ZN(n13567) );
  AND2_X1 U15610 ( .A1(n13567), .A2(n13566), .ZN(n13673) );
  NAND2_X1 U15611 ( .A1(n13673), .A2(n13581), .ZN(n13568) );
  NAND4_X1 U15612 ( .A1(n13571), .A2(n13570), .A3(n13569), .A4(n13568), .ZN(
        P2_U3251) );
  NAND2_X1 U15613 ( .A1(n13572), .A2(n13557), .ZN(n13586) );
  OAI22_X1 U15614 ( .A1(n13557), .A2(n13575), .B1(n13574), .B2(n13573), .ZN(
        n13576) );
  AOI21_X1 U15615 ( .B1(n13578), .B2(n13577), .A(n13576), .ZN(n13585) );
  NAND2_X1 U15616 ( .A1(n13580), .A2(n13579), .ZN(n13584) );
  NAND2_X1 U15617 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  NAND4_X1 U15618 ( .A1(n13586), .A2(n13585), .A3(n13584), .A4(n13583), .ZN(
        P2_U3253) );
  NOR2_X1 U15619 ( .A1(n13588), .A2(n13587), .ZN(n13677) );
  MUX2_X1 U15620 ( .A(n13589), .B(n13677), .S(n14931), .Z(n13590) );
  OAI21_X1 U15621 ( .B1(n13680), .B2(n13629), .A(n13590), .ZN(P2_U3530) );
  AND2_X1 U15622 ( .A1(n13592), .A2(n13591), .ZN(n13681) );
  MUX2_X1 U15623 ( .A(n13593), .B(n13681), .S(n14931), .Z(n13594) );
  OAI21_X1 U15624 ( .B1(n13684), .B2(n13629), .A(n13594), .ZN(P2_U3529) );
  AOI21_X1 U15625 ( .B1(n14918), .B2(n13598), .A(n13597), .ZN(n13599) );
  OAI211_X1 U15626 ( .C1(n13601), .C2(n14921), .A(n13600), .B(n13599), .ZN(
        n13685) );
  MUX2_X1 U15627 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13685), .S(n14931), .Z(
        P2_U3527) );
  INV_X1 U15628 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13606) );
  INV_X1 U15629 ( .A(n13602), .ZN(n13604) );
  MUX2_X1 U15630 ( .A(n13606), .B(n13686), .S(n14931), .Z(n13607) );
  OAI21_X1 U15631 ( .B1(n13689), .B2(n13629), .A(n13607), .ZN(P2_U3526) );
  AOI211_X1 U15632 ( .C1(n13610), .C2(n14905), .A(n13609), .B(n13608), .ZN(
        n13690) );
  MUX2_X1 U15633 ( .A(n13611), .B(n13690), .S(n14931), .Z(n13612) );
  OAI21_X1 U15634 ( .B1(n13693), .B2(n13629), .A(n13612), .ZN(P2_U3525) );
  NAND2_X1 U15635 ( .A1(n13613), .A2(n14905), .ZN(n13616) );
  NAND3_X1 U15636 ( .A1(n13616), .A2(n13615), .A3(n13614), .ZN(n13694) );
  MUX2_X1 U15637 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13694), .S(n14931), .Z(
        n13617) );
  AOI21_X1 U15638 ( .B1(n13675), .B2(n13696), .A(n13617), .ZN(n13618) );
  INV_X1 U15639 ( .A(n13618), .ZN(P2_U3524) );
  AOI21_X1 U15640 ( .B1(n14918), .B2(n13620), .A(n13619), .ZN(n13621) );
  OAI211_X1 U15641 ( .C1(n13623), .C2(n8756), .A(n13622), .B(n13621), .ZN(
        n13698) );
  MUX2_X1 U15642 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13698), .S(n14931), .Z(
        P2_U3523) );
  AOI211_X1 U15643 ( .C1(n14905), .C2(n13626), .A(n13625), .B(n13624), .ZN(
        n13699) );
  MUX2_X1 U15644 ( .A(n13627), .B(n13699), .S(n14931), .Z(n13628) );
  OAI21_X1 U15645 ( .B1(n6939), .B2(n13629), .A(n13628), .ZN(P2_U3522) );
  OAI211_X1 U15646 ( .C1(n13632), .C2(n14921), .A(n13631), .B(n13630), .ZN(
        n13703) );
  MUX2_X1 U15647 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13703), .S(n14931), .Z(
        n13633) );
  AOI21_X1 U15648 ( .B1(n13675), .B2(n13705), .A(n13633), .ZN(n13634) );
  INV_X1 U15649 ( .A(n13634), .ZN(P2_U3521) );
  AOI21_X1 U15650 ( .B1(n14918), .B2(n13636), .A(n13635), .ZN(n13637) );
  OAI211_X1 U15651 ( .C1(n13639), .C2(n14921), .A(n13638), .B(n13637), .ZN(
        n13707) );
  MUX2_X1 U15652 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13707), .S(n14931), .Z(
        P2_U3520) );
  AOI211_X1 U15653 ( .C1(n14918), .C2(n13642), .A(n13641), .B(n13640), .ZN(
        n13643) );
  OAI21_X1 U15654 ( .B1(n14921), .B2(n13644), .A(n13643), .ZN(n13708) );
  MUX2_X1 U15655 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13708), .S(n14931), .Z(
        P2_U3519) );
  AOI211_X1 U15656 ( .C1(n14918), .C2(n13647), .A(n13646), .B(n13645), .ZN(
        n13648) );
  OAI21_X1 U15657 ( .B1(n14921), .B2(n13649), .A(n13648), .ZN(n13709) );
  MUX2_X1 U15658 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13709), .S(n14931), .Z(
        P2_U3518) );
  AOI21_X1 U15659 ( .B1(n14918), .B2(n13651), .A(n13650), .ZN(n13652) );
  OAI211_X1 U15660 ( .C1(n13654), .C2(n14921), .A(n13653), .B(n13652), .ZN(
        n13710) );
  MUX2_X1 U15661 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13710), .S(n14931), .Z(
        P2_U3517) );
  AOI21_X1 U15662 ( .B1(n14918), .B2(n13656), .A(n13655), .ZN(n13657) );
  OAI211_X1 U15663 ( .C1(n13659), .C2(n14921), .A(n13658), .B(n13657), .ZN(
        n13711) );
  MUX2_X1 U15664 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13711), .S(n14931), .Z(
        P2_U3516) );
  OAI211_X1 U15665 ( .C1(n13662), .C2(n14921), .A(n13661), .B(n13660), .ZN(
        n13712) );
  MUX2_X1 U15666 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13712), .S(n14931), .Z(
        n13663) );
  AOI21_X1 U15667 ( .B1(n13675), .B2(n14637), .A(n13663), .ZN(n13664) );
  INV_X1 U15668 ( .A(n13664), .ZN(P2_U3515) );
  INV_X1 U15669 ( .A(n13665), .ZN(n13667) );
  NAND3_X1 U15670 ( .A1(n13668), .A2(n13667), .A3(n13666), .ZN(n13669) );
  AOI21_X1 U15671 ( .B1(n13670), .B2(n14905), .A(n13669), .ZN(n13717) );
  AOI22_X1 U15672 ( .A1(n13715), .A2(n13675), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n14929), .ZN(n13671) );
  OAI21_X1 U15673 ( .B1(n13717), .B2(n14929), .A(n13671), .ZN(P2_U3514) );
  AOI211_X1 U15674 ( .C1(n13674), .C2(n14905), .A(n13673), .B(n13672), .ZN(
        n13720) );
  AOI22_X1 U15675 ( .A1(n13718), .A2(n13675), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n14929), .ZN(n13676) );
  OAI21_X1 U15676 ( .B1(n13720), .B2(n14929), .A(n13676), .ZN(P2_U3513) );
  MUX2_X1 U15677 ( .A(n13678), .B(n13677), .S(n14908), .Z(n13679) );
  OAI21_X1 U15678 ( .B1(n13680), .B2(n13702), .A(n13679), .ZN(P2_U3498) );
  MUX2_X1 U15679 ( .A(n13682), .B(n13681), .S(n14908), .Z(n13683) );
  OAI21_X1 U15680 ( .B1(n13684), .B2(n13702), .A(n13683), .ZN(P2_U3497) );
  MUX2_X1 U15681 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13685), .S(n14908), .Z(
        P2_U3495) );
  MUX2_X1 U15682 ( .A(n13687), .B(n13686), .S(n14908), .Z(n13688) );
  OAI21_X1 U15683 ( .B1(n13689), .B2(n13702), .A(n13688), .ZN(P2_U3494) );
  INV_X1 U15684 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13691) );
  MUX2_X1 U15685 ( .A(n13691), .B(n13690), .S(n14908), .Z(n13692) );
  OAI21_X1 U15686 ( .B1(n13693), .B2(n13702), .A(n13692), .ZN(P2_U3493) );
  MUX2_X1 U15687 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13694), .S(n14908), .Z(
        n13695) );
  AOI21_X1 U15688 ( .B1(n8282), .B2(n13696), .A(n13695), .ZN(n13697) );
  INV_X1 U15689 ( .A(n13697), .ZN(P2_U3492) );
  MUX2_X1 U15690 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13698), .S(n14908), .Z(
        P2_U3491) );
  INV_X1 U15691 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13700) );
  MUX2_X1 U15692 ( .A(n13700), .B(n13699), .S(n14908), .Z(n13701) );
  OAI21_X1 U15693 ( .B1(n6939), .B2(n13702), .A(n13701), .ZN(P2_U3490) );
  MUX2_X1 U15694 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13703), .S(n14908), .Z(
        n13704) );
  AOI21_X1 U15695 ( .B1(n8282), .B2(n13705), .A(n13704), .ZN(n13706) );
  INV_X1 U15696 ( .A(n13706), .ZN(P2_U3489) );
  MUX2_X1 U15697 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13707), .S(n14908), .Z(
        P2_U3488) );
  MUX2_X1 U15698 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13708), .S(n14908), .Z(
        P2_U3487) );
  MUX2_X1 U15699 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13709), .S(n14908), .Z(
        P2_U3486) );
  MUX2_X1 U15700 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13710), .S(n14908), .Z(
        P2_U3484) );
  MUX2_X1 U15701 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13711), .S(n14908), .Z(
        P2_U3481) );
  MUX2_X1 U15702 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13712), .S(n14908), .Z(
        n13713) );
  AOI21_X1 U15703 ( .B1(n8282), .B2(n14637), .A(n13713), .ZN(n13714) );
  INV_X1 U15704 ( .A(n13714), .ZN(P2_U3478) );
  AOI22_X1 U15705 ( .A1(n13715), .A2(n8282), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n14924), .ZN(n13716) );
  OAI21_X1 U15706 ( .B1(n13717), .B2(n14924), .A(n13716), .ZN(P2_U3475) );
  AOI22_X1 U15707 ( .A1(n13718), .A2(n8282), .B1(P2_REG0_REG_14__SCAN_IN), 
        .B2(n14924), .ZN(n13719) );
  OAI21_X1 U15708 ( .B1(n13720), .B2(n14924), .A(n13719), .ZN(P2_U3472) );
  INV_X1 U15709 ( .A(n13721), .ZN(n14377) );
  NAND3_X1 U15710 ( .A1(n13723), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13724) );
  INV_X1 U15711 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n15386) );
  OAI22_X1 U15712 ( .A1(n13722), .A2(n13724), .B1(n15386), .B2(n13736), .ZN(
        n13725) );
  INV_X1 U15713 ( .A(n13725), .ZN(n13726) );
  OAI21_X1 U15714 ( .B1(n14377), .B2(n11298), .A(n13726), .ZN(P2_U3296) );
  NAND2_X1 U15715 ( .A1(n13728), .A2(n13727), .ZN(n13730) );
  OAI211_X1 U15716 ( .C1(n13736), .C2(n13731), .A(n13730), .B(n13729), .ZN(
        P2_U3299) );
  INV_X1 U15717 ( .A(n13732), .ZN(n14386) );
  OAI222_X1 U15718 ( .A1(n13736), .A2(n13734), .B1(n11298), .B2(n14386), .C1(
        n13733), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15719 ( .A(n13735), .ZN(n14389) );
  OAI222_X1 U15720 ( .A1(n13737), .A2(P2_U3088), .B1(n11298), .B2(n14389), 
        .C1(n15264), .C2(n13736), .ZN(P2_U3301) );
  INV_X1 U15721 ( .A(n13738), .ZN(n13739) );
  MUX2_X1 U15722 ( .A(n13739), .B(n6810), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  OAI22_X1 U15723 ( .A1(n13818), .A2(n14212), .B1(n13741), .B2(n14210), .ZN(
        n14025) );
  AOI22_X1 U15724 ( .A1(n14025), .A2(n13795), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13744) );
  NAND2_X1 U15725 ( .A1(n14248), .A2(n13936), .ZN(n13743) );
  NAND2_X1 U15726 ( .A1(n13932), .A2(n14028), .ZN(n13742) );
  NAND4_X1 U15727 ( .A1(n13745), .A2(n13744), .A3(n13743), .A4(n13742), .ZN(
        P1_U3214) );
  INV_X1 U15728 ( .A(n13923), .ZN(n13746) );
  AOI21_X1 U15729 ( .B1(n13748), .B2(n13747), .A(n13746), .ZN(n13755) );
  INV_X1 U15730 ( .A(n13749), .ZN(n13750) );
  NAND2_X1 U15731 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14697)
         );
  OAI21_X1 U15732 ( .B1(n13887), .B2(n13750), .A(n14697), .ZN(n13753) );
  OAI22_X1 U15733 ( .A1(n13751), .A2(n13904), .B1(n13903), .B2(n14213), .ZN(
        n13752) );
  AOI211_X1 U15734 ( .C1(n14329), .C2(n13936), .A(n13753), .B(n13752), .ZN(
        n13754) );
  OAI21_X1 U15735 ( .B1(n13755), .B2(n13938), .A(n13754), .ZN(P1_U3215) );
  INV_X1 U15736 ( .A(n13756), .ZN(n13757) );
  NOR2_X1 U15737 ( .A1(n13758), .A2(n13757), .ZN(n13762) );
  INV_X1 U15738 ( .A(n13760), .ZN(n13761) );
  AOI21_X1 U15739 ( .B1(n13762), .B2(n13759), .A(n13761), .ZN(n13767) );
  OAI22_X1 U15740 ( .A1(n13887), .A2(n14096), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15336), .ZN(n13765) );
  OAI22_X1 U15741 ( .A1(n13763), .A2(n13904), .B1(n13903), .B2(n13817), .ZN(
        n13764) );
  AOI211_X1 U15742 ( .C1(n14276), .C2(n13936), .A(n13765), .B(n13764), .ZN(
        n13766) );
  OAI21_X1 U15743 ( .B1(n13767), .B2(n13938), .A(n13766), .ZN(P1_U3216) );
  INV_X1 U15744 ( .A(n13768), .ZN(n14789) );
  INV_X1 U15745 ( .A(n13769), .ZN(n13891) );
  AOI21_X1 U15746 ( .B1(n12222), .B2(n13771), .A(n13770), .ZN(n13772) );
  INV_X1 U15747 ( .A(n13773), .ZN(n13776) );
  OAI22_X1 U15748 ( .A1(n13804), .A2(n13903), .B1(n13904), .B2(n13774), .ZN(
        n13775) );
  AOI211_X1 U15749 ( .C1(n13932), .C2(n13777), .A(n13776), .B(n13775), .ZN(
        n13778) );
  OAI211_X1 U15750 ( .C1(n14789), .C2(n13921), .A(n13779), .B(n13778), .ZN(
        P1_U3217) );
  INV_X1 U15751 ( .A(n14298), .ZN(n14159) );
  INV_X1 U15752 ( .A(n13898), .ZN(n13782) );
  OAI21_X1 U15753 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n13784) );
  NAND3_X1 U15754 ( .A1(n13784), .A2(n13912), .A3(n13783), .ZN(n13789) );
  AND2_X1 U15755 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13993) );
  OAI22_X1 U15756 ( .A1(n13786), .A2(n13904), .B1(n13903), .B2(n13785), .ZN(
        n13787) );
  AOI211_X1 U15757 ( .C1(n13932), .C2(n14157), .A(n13993), .B(n13787), .ZN(
        n13788) );
  OAI211_X1 U15758 ( .C1(n14159), .C2(n13921), .A(n13789), .B(n13788), .ZN(
        P1_U3219) );
  INV_X1 U15759 ( .A(n13790), .ZN(n13874) );
  AOI21_X1 U15760 ( .B1(n13792), .B2(n13791), .A(n13874), .ZN(n13799) );
  NAND2_X1 U15761 ( .A1(n14092), .A2(n14172), .ZN(n13794) );
  NAND2_X1 U15762 ( .A1(n14164), .A2(n14174), .ZN(n13793) );
  NAND2_X1 U15763 ( .A1(n13794), .A2(n13793), .ZN(n14121) );
  AOI22_X1 U15764 ( .A1(n14121), .A2(n13795), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13796) );
  OAI21_X1 U15765 ( .B1(n14124), .B2(n13887), .A(n13796), .ZN(n13797) );
  AOI21_X1 U15766 ( .B1(n14288), .B2(n13936), .A(n13797), .ZN(n13798) );
  OAI21_X1 U15767 ( .B1(n13799), .B2(n13938), .A(n13798), .ZN(P1_U3223) );
  AND2_X1 U15768 ( .A1(n13892), .A2(n13800), .ZN(n13803) );
  OAI211_X1 U15769 ( .C1(n13803), .C2(n13802), .A(n13912), .B(n13801), .ZN(
        n13811) );
  OR2_X1 U15770 ( .A1(n13804), .A2(n14212), .ZN(n13806) );
  NAND2_X1 U15771 ( .A1(n13947), .A2(n14172), .ZN(n13805) );
  AND2_X1 U15772 ( .A1(n13806), .A2(n13805), .ZN(n14536) );
  OAI21_X1 U15773 ( .B1(n13934), .B2(n14536), .A(n13807), .ZN(n13808) );
  AOI21_X1 U15774 ( .B1(n13809), .B2(n13932), .A(n13808), .ZN(n13810) );
  OAI211_X1 U15775 ( .C1(n14538), .C2(n13921), .A(n13811), .B(n13810), .ZN(
        P1_U3224) );
  NOR2_X1 U15776 ( .A1(n13813), .A2(n7360), .ZN(n13816) );
  INV_X1 U15777 ( .A(n13814), .ZN(n13815) );
  AOI21_X1 U15778 ( .B1(n13816), .B2(n13845), .A(n13815), .ZN(n13822) );
  INV_X1 U15779 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15263) );
  OAI22_X1 U15780 ( .A1(n13887), .A2(n14060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15263), .ZN(n13820) );
  OAI22_X1 U15781 ( .A1(n13818), .A2(n13903), .B1(n13904), .B2(n13817), .ZN(
        n13819) );
  AOI211_X1 U15782 ( .C1(n14259), .C2(n13936), .A(n13820), .B(n13819), .ZN(
        n13821) );
  OAI21_X1 U15783 ( .B1(n13822), .B2(n13938), .A(n13821), .ZN(P1_U3225) );
  OAI21_X1 U15784 ( .B1(n13824), .B2(n13823), .A(n13831), .ZN(n13825) );
  NAND2_X1 U15785 ( .A1(n13825), .A2(n13912), .ZN(n13830) );
  NAND2_X1 U15786 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14727)
         );
  INV_X1 U15787 ( .A(n14727), .ZN(n13827) );
  OAI22_X1 U15788 ( .A1(n14211), .A2(n13903), .B1(n13904), .B2(n14213), .ZN(
        n13826) );
  AOI211_X1 U15789 ( .C1(n13932), .C2(n13828), .A(n13827), .B(n13826), .ZN(
        n13829) );
  OAI211_X1 U15790 ( .C1(n14365), .C2(n13921), .A(n13830), .B(n13829), .ZN(
        P1_U3226) );
  INV_X1 U15791 ( .A(n14310), .ZN(n14198) );
  INV_X1 U15792 ( .A(n13831), .ZN(n13834) );
  NOR3_X1 U15793 ( .A1(n13834), .A2(n13833), .A3(n13832), .ZN(n13837) );
  INV_X1 U15794 ( .A(n13835), .ZN(n13836) );
  OAI21_X1 U15795 ( .B1(n13837), .B2(n13836), .A(n13912), .ZN(n13842) );
  OR2_X1 U15796 ( .A1(n13928), .A2(n14212), .ZN(n13839) );
  NAND2_X1 U15797 ( .A1(n14163), .A2(n14172), .ZN(n13838) );
  AND2_X1 U15798 ( .A1(n13839), .A2(n13838), .ZN(n14190) );
  NAND2_X1 U15799 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14742)
         );
  OAI21_X1 U15800 ( .B1(n13934), .B2(n14190), .A(n14742), .ZN(n13840) );
  AOI21_X1 U15801 ( .B1(n14195), .B2(n13932), .A(n13840), .ZN(n13841) );
  OAI211_X1 U15802 ( .C1(n14198), .C2(n13921), .A(n13842), .B(n13841), .ZN(
        P1_U3228) );
  NOR2_X1 U15803 ( .A1(n13844), .A2(n7363), .ZN(n13847) );
  INV_X1 U15804 ( .A(n13845), .ZN(n13846) );
  AOI21_X1 U15805 ( .B1(n13847), .B2(n13760), .A(n13846), .ZN(n13854) );
  INV_X1 U15806 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13848) );
  OAI22_X1 U15807 ( .A1(n13887), .A2(n13849), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13848), .ZN(n13852) );
  OAI22_X1 U15808 ( .A1(n13850), .A2(n13904), .B1(n13903), .B2(n13914), .ZN(
        n13851) );
  AOI211_X1 U15809 ( .C1(n14266), .C2(n13936), .A(n13852), .B(n13851), .ZN(
        n13853) );
  OAI21_X1 U15810 ( .B1(n13854), .B2(n13938), .A(n13853), .ZN(P1_U3229) );
  XNOR2_X1 U15811 ( .A(n13856), .B(n13855), .ZN(n13861) );
  OAI22_X1 U15812 ( .A1(n13887), .A2(n14143), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15252), .ZN(n13859) );
  OAI22_X1 U15813 ( .A1(n13857), .A2(n13903), .B1(n13904), .B2(n13902), .ZN(
        n13858) );
  AOI211_X1 U15814 ( .C1(n14292), .C2(n13936), .A(n13859), .B(n13858), .ZN(
        n13860) );
  OAI21_X1 U15815 ( .B1(n13861), .B2(n13938), .A(n13860), .ZN(P1_U3233) );
  XNOR2_X1 U15816 ( .A(n13863), .B(n13862), .ZN(n13870) );
  NAND2_X1 U15817 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14682)
         );
  NAND2_X1 U15818 ( .A1(n13932), .A2(n13864), .ZN(n13865) );
  OAI211_X1 U15819 ( .C1(n13934), .C2(n13866), .A(n14682), .B(n13865), .ZN(
        n13867) );
  AOI21_X1 U15820 ( .B1(n13868), .B2(n13936), .A(n13867), .ZN(n13869) );
  OAI21_X1 U15821 ( .B1(n13870), .B2(n13938), .A(n13869), .ZN(P1_U3234) );
  INV_X1 U15822 ( .A(n13871), .ZN(n13873) );
  NOR3_X1 U15823 ( .A1(n13874), .A2(n13873), .A3(n13872), .ZN(n13876) );
  INV_X1 U15824 ( .A(n13759), .ZN(n13875) );
  OAI21_X1 U15825 ( .B1(n13876), .B2(n13875), .A(n13912), .ZN(n13881) );
  INV_X1 U15826 ( .A(n14114), .ZN(n13879) );
  AOI22_X1 U15827 ( .A1(n14072), .A2(n14172), .B1(n14140), .B2(n14174), .ZN(
        n14109) );
  INV_X1 U15828 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13877) );
  OAI22_X1 U15829 ( .A1(n14109), .A2(n13934), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13877), .ZN(n13878) );
  AOI21_X1 U15830 ( .B1(n13879), .B2(n13932), .A(n13878), .ZN(n13880) );
  OAI211_X1 U15831 ( .C1(n13921), .C2(n13882), .A(n13881), .B(n13880), .ZN(
        P1_U3235) );
  AOI22_X1 U15832 ( .A1(n13884), .A2(n13948), .B1(n13883), .B2(n13950), .ZN(
        n13886) );
  OAI211_X1 U15833 ( .C1(n13888), .C2(n13887), .A(n13886), .B(n13885), .ZN(
        n13895) );
  OAI21_X1 U15834 ( .B1(n13891), .B2(n13890), .A(n13889), .ZN(n13893) );
  AOI21_X1 U15835 ( .B1(n13893), .B2(n13892), .A(n13938), .ZN(n13894) );
  AOI211_X1 U15836 ( .C1(n13896), .C2(n13936), .A(n13895), .B(n13894), .ZN(
        n13897) );
  INV_X1 U15837 ( .A(n13897), .ZN(P1_U3236) );
  INV_X1 U15838 ( .A(n14304), .ZN(n14180) );
  OAI21_X1 U15839 ( .B1(n13900), .B2(n13899), .A(n13898), .ZN(n13901) );
  NAND2_X1 U15840 ( .A1(n13901), .A2(n13912), .ZN(n13908) );
  NAND2_X1 U15841 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14759)
         );
  INV_X1 U15842 ( .A(n14759), .ZN(n13906) );
  OAI22_X1 U15843 ( .A1(n14211), .A2(n13904), .B1(n13903), .B2(n13902), .ZN(
        n13905) );
  AOI211_X1 U15844 ( .C1(n13932), .C2(n14178), .A(n13906), .B(n13905), .ZN(
        n13907) );
  OAI211_X1 U15845 ( .C1(n14180), .C2(n13921), .A(n13908), .B(n13907), .ZN(
        P1_U3238) );
  OAI21_X1 U15846 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n13913) );
  NAND2_X1 U15847 ( .A1(n13913), .A2(n13912), .ZN(n13920) );
  OR2_X1 U15848 ( .A1(n13914), .A2(n14212), .ZN(n13916) );
  NAND2_X1 U15849 ( .A1(n13943), .A2(n14172), .ZN(n13915) );
  AND2_X1 U15850 ( .A1(n13916), .A2(n13915), .ZN(n14043) );
  OAI22_X1 U15851 ( .A1(n13934), .A2(n14043), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13917), .ZN(n13918) );
  AOI21_X1 U15852 ( .B1(n14046), .B2(n13932), .A(n13918), .ZN(n13919) );
  OAI211_X1 U15853 ( .C1(n14350), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        P1_U3240) );
  NAND2_X1 U15854 ( .A1(n13923), .A2(n13922), .ZN(n13927) );
  XNOR2_X1 U15855 ( .A(n13925), .B(n13924), .ZN(n13926) );
  XNOR2_X1 U15856 ( .A(n13927), .B(n13926), .ZN(n13939) );
  OR2_X1 U15857 ( .A1(n13928), .A2(n14210), .ZN(n13931) );
  OR2_X1 U15858 ( .A1(n13929), .A2(n14212), .ZN(n13930) );
  AND2_X1 U15859 ( .A1(n13931), .A2(n13930), .ZN(n14322) );
  NAND2_X1 U15860 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14712)
         );
  NAND2_X1 U15861 ( .A1(n13932), .A2(n14223), .ZN(n13933) );
  OAI211_X1 U15862 ( .C1(n13934), .C2(n14322), .A(n14712), .B(n13933), .ZN(
        n13935) );
  AOI21_X1 U15863 ( .B1(n14320), .B2(n13936), .A(n13935), .ZN(n13937) );
  OAI21_X1 U15864 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(P1_U3241) );
  MUX2_X1 U15865 ( .A(n13999), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13959), .Z(
        P1_U3591) );
  MUX2_X1 U15866 ( .A(n13940), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13959), .Z(
        P1_U3590) );
  MUX2_X1 U15867 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13941), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15868 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13942), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15869 ( .A(n13943), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13959), .Z(
        P1_U3587) );
  MUX2_X1 U15870 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14053), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15871 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14071), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15872 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14093), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15873 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14072), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15874 ( .A(n14092), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13959), .Z(
        P1_U3582) );
  MUX2_X1 U15875 ( .A(n14140), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13959), .Z(
        P1_U3581) );
  MUX2_X1 U15876 ( .A(n14164), .B(P1_DATAO_REG_20__SCAN_IN), .S(n13959), .Z(
        P1_U3580) );
  MUX2_X1 U15877 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14173), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15878 ( .A(n14163), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13959), .Z(
        P1_U3578) );
  MUX2_X1 U15879 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14175), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15880 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13944), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15881 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13945), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15882 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13946), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15883 ( .A(n13947), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13959), .Z(
        P1_U3573) );
  MUX2_X1 U15884 ( .A(n13948), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13959), .Z(
        P1_U3572) );
  MUX2_X1 U15885 ( .A(n13949), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13959), .Z(
        P1_U3571) );
  MUX2_X1 U15886 ( .A(n13950), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13959), .Z(
        P1_U3570) );
  MUX2_X1 U15887 ( .A(n13951), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13959), .Z(
        P1_U3569) );
  MUX2_X1 U15888 ( .A(n13952), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13959), .Z(
        P1_U3568) );
  MUX2_X1 U15889 ( .A(n13953), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13959), .Z(
        P1_U3567) );
  MUX2_X1 U15890 ( .A(n13954), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13959), .Z(
        P1_U3566) );
  MUX2_X1 U15891 ( .A(n13955), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13959), .Z(
        P1_U3565) );
  MUX2_X1 U15892 ( .A(n13956), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13959), .Z(
        P1_U3564) );
  MUX2_X1 U15893 ( .A(n13957), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13959), .Z(
        P1_U3563) );
  MUX2_X1 U15894 ( .A(n13958), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13959), .Z(
        P1_U3562) );
  MUX2_X1 U15895 ( .A(n13960), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13959), .Z(
        P1_U3561) );
  MUX2_X1 U15896 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13961), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U15897 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13963) );
  NOR2_X1 U15898 ( .A1(n14725), .A2(n13963), .ZN(n13962) );
  AOI21_X1 U15899 ( .B1(n14725), .B2(n13963), .A(n13962), .ZN(n14721) );
  NAND2_X1 U15900 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n14681), .ZN(n13964) );
  OAI21_X1 U15901 ( .B1(n14681), .B2(P1_REG2_REG_13__SCAN_IN), .A(n13964), 
        .ZN(n14677) );
  NOR2_X1 U15902 ( .A1(n14677), .A2(n14678), .ZN(n14676) );
  INV_X1 U15903 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13966) );
  MUX2_X1 U15904 ( .A(n13966), .B(P1_REG2_REG_14__SCAN_IN), .S(n13980), .Z(
        n14687) );
  NAND2_X1 U15905 ( .A1(n13967), .A2(n14710), .ZN(n13969) );
  XNOR2_X1 U15906 ( .A(n14710), .B(n13968), .ZN(n14702) );
  INV_X1 U15907 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14701) );
  NAND2_X1 U15908 ( .A1(n14702), .A2(n14701), .ZN(n14700) );
  NAND2_X1 U15909 ( .A1(n13969), .A2(n14700), .ZN(n14722) );
  INV_X1 U15910 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13970) );
  OR2_X1 U15911 ( .A1(n13984), .A2(n13970), .ZN(n13972) );
  NAND2_X1 U15912 ( .A1(n13984), .A2(n13970), .ZN(n13971) );
  AND2_X1 U15913 ( .A1(n13972), .A2(n13971), .ZN(n14732) );
  NOR2_X1 U15914 ( .A1(n13973), .A2(n14756), .ZN(n13974) );
  INV_X1 U15915 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14746) );
  XNOR2_X1 U15916 ( .A(n14756), .B(n13973), .ZN(n14747) );
  NOR2_X1 U15917 ( .A1(n14746), .A2(n14747), .ZN(n14745) );
  NOR2_X1 U15918 ( .A1(n13974), .A2(n14745), .ZN(n13975) );
  XNOR2_X1 U15919 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13975), .ZN(n13991) );
  INV_X1 U15920 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15249) );
  XNOR2_X1 U15921 ( .A(n14725), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n14717) );
  INV_X1 U15922 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13976) );
  XNOR2_X1 U15923 ( .A(n13980), .B(n13976), .ZN(n14691) );
  OAI21_X1 U15924 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n13978), .A(n13977), 
        .ZN(n14675) );
  INV_X1 U15925 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13979) );
  MUX2_X1 U15926 ( .A(n13979), .B(P1_REG1_REG_13__SCAN_IN), .S(n14681), .Z(
        n14674) );
  NOR2_X1 U15927 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  NAND2_X1 U15928 ( .A1(n14691), .A2(n14690), .ZN(n14689) );
  OAI21_X1 U15929 ( .B1(n13980), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14689), 
        .ZN(n13981) );
  NAND2_X1 U15930 ( .A1(n14710), .A2(n13981), .ZN(n13983) );
  INV_X1 U15931 ( .A(n13981), .ZN(n13982) );
  INV_X1 U15932 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14705) );
  NAND2_X1 U15933 ( .A1(n14706), .A2(n14705), .ZN(n14704) );
  NAND2_X1 U15934 ( .A1(n13983), .A2(n14704), .ZN(n14718) );
  XNOR2_X1 U15935 ( .A(n13984), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U15936 ( .A1(n13985), .A2(n14756), .ZN(n13986) );
  NOR2_X1 U15937 ( .A1(n14750), .A2(n13986), .ZN(n13988) );
  INV_X1 U15938 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13987) );
  INV_X1 U15939 ( .A(n13993), .ZN(n13994) );
  XNOR2_X1 U15940 ( .A(n14340), .B(n14002), .ZN(n13997) );
  NAND2_X1 U15941 ( .A1(n13997), .A2(n14512), .ZN(n14236) );
  NAND2_X1 U15942 ( .A1(n13999), .A2(n13998), .ZN(n14238) );
  NOR2_X1 U15943 ( .A1(n14224), .A2(n14238), .ZN(n14005) );
  NOR2_X1 U15944 ( .A1(n14340), .A2(n14525), .ZN(n14000) );
  AOI211_X1 U15945 ( .C1(n14224), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14005), 
        .B(n14000), .ZN(n14001) );
  OAI21_X1 U15946 ( .B1(n14236), .B2(n14516), .A(n14001), .ZN(P1_U3263) );
  OAI211_X1 U15947 ( .C1(n14344), .C2(n14003), .A(n14002), .B(n14512), .ZN(
        n14239) );
  NOR2_X1 U15948 ( .A1(n14344), .A2(n14525), .ZN(n14004) );
  AOI211_X1 U15949 ( .C1(n14224), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14005), 
        .B(n14004), .ZN(n14006) );
  OAI21_X1 U15950 ( .B1(n14516), .B2(n14239), .A(n14006), .ZN(P1_U3264) );
  XNOR2_X1 U15951 ( .A(n14007), .B(n14010), .ZN(n14009) );
  AOI21_X1 U15952 ( .B1(n14009), .B2(n14522), .A(n14008), .ZN(n14245) );
  NAND2_X1 U15953 ( .A1(n14011), .A2(n14010), .ZN(n14012) );
  NAND2_X1 U15954 ( .A1(n14013), .A2(n14012), .ZN(n14246) );
  INV_X1 U15955 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14015) );
  OAI22_X1 U15956 ( .A1(n14529), .A2(n14015), .B1(n14014), .B2(n14526), .ZN(
        n14016) );
  AOI21_X1 U15957 ( .B1(n14243), .B2(n14225), .A(n14016), .ZN(n14021) );
  AOI21_X1 U15958 ( .B1(n6879), .B2(n14027), .A(n14252), .ZN(n14019) );
  AND2_X1 U15959 ( .A1(n14019), .A2(n14018), .ZN(n14242) );
  NAND2_X1 U15960 ( .A1(n14242), .A2(n14194), .ZN(n14020) );
  OAI211_X1 U15961 ( .C1(n14246), .C2(n14201), .A(n14021), .B(n14020), .ZN(
        n14022) );
  INV_X1 U15962 ( .A(n14022), .ZN(n14023) );
  OAI21_X1 U15963 ( .B1(n14245), .B2(n14224), .A(n14023), .ZN(P1_U3265) );
  XNOR2_X1 U15964 ( .A(n14024), .B(n14034), .ZN(n14026) );
  AOI21_X1 U15965 ( .B1(n14026), .B2(n14522), .A(n14025), .ZN(n14250) );
  AOI211_X1 U15966 ( .C1(n14248), .C2(n14045), .A(n14252), .B(n14017), .ZN(
        n14247) );
  INV_X1 U15967 ( .A(n14248), .ZN(n14030) );
  AOI22_X1 U15968 ( .A1(n14224), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14028), 
        .B2(n14222), .ZN(n14029) );
  OAI21_X1 U15969 ( .B1(n14030), .B2(n14525), .A(n14029), .ZN(n14035) );
  INV_X1 U15970 ( .A(n14031), .ZN(n14032) );
  OAI21_X1 U15971 ( .B1(n14224), .B2(n14250), .A(n14036), .ZN(P1_U3266) );
  NAND2_X1 U15972 ( .A1(n14261), .A2(n14037), .ZN(n14038) );
  NAND2_X1 U15973 ( .A1(n14038), .A2(n14041), .ZN(n14040) );
  OR2_X1 U15974 ( .A1(n14038), .A2(n14041), .ZN(n14039) );
  NAND2_X1 U15975 ( .A1(n14040), .A2(n14039), .ZN(n14254) );
  XNOR2_X1 U15976 ( .A(n14042), .B(n14041), .ZN(n14044) );
  OAI21_X1 U15977 ( .B1(n14044), .B2(n14110), .A(n14043), .ZN(n14256) );
  NAND2_X1 U15978 ( .A1(n14256), .A2(n14529), .ZN(n14051) );
  OAI21_X1 U15979 ( .B1(n14056), .B2(n14350), .A(n14045), .ZN(n14253) );
  INV_X1 U15980 ( .A(n14253), .ZN(n14049) );
  AOI22_X1 U15981 ( .A1(n14224), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14046), 
        .B2(n14222), .ZN(n14047) );
  OAI21_X1 U15982 ( .B1(n14350), .B2(n14525), .A(n14047), .ZN(n14048) );
  AOI21_X1 U15983 ( .B1(n14049), .B2(n14168), .A(n14048), .ZN(n14050) );
  OAI211_X1 U15984 ( .C1(n14201), .C2(n14254), .A(n14051), .B(n14050), .ZN(
        P1_U3267) );
  OAI21_X1 U15985 ( .B1(n7601), .B2(n14058), .A(n14052), .ZN(n14054) );
  AOI222_X1 U15986 ( .A1(n14522), .A2(n14054), .B1(n14053), .B2(n14172), .C1(
        n14093), .C2(n14174), .ZN(n14265) );
  NAND2_X1 U15987 ( .A1(n14081), .A2(n14259), .ZN(n14055) );
  NAND2_X1 U15988 ( .A1(n14055), .A2(n14512), .ZN(n14057) );
  OR2_X1 U15989 ( .A1(n14057), .A2(n14056), .ZN(n14262) );
  NAND2_X1 U15990 ( .A1(n14059), .A2(n14058), .ZN(n14260) );
  NAND3_X1 U15991 ( .A1(n14261), .A2(n14260), .A3(n14233), .ZN(n14064) );
  INV_X1 U15992 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14061) );
  OAI22_X1 U15993 ( .A1(n14529), .A2(n14061), .B1(n14060), .B2(n14526), .ZN(
        n14062) );
  AOI21_X1 U15994 ( .B1(n14259), .B2(n14225), .A(n14062), .ZN(n14063) );
  OAI211_X1 U15995 ( .C1(n14262), .C2(n14516), .A(n14064), .B(n14063), .ZN(
        n14065) );
  INV_X1 U15996 ( .A(n14065), .ZN(n14066) );
  OAI21_X1 U15997 ( .B1(n14265), .B2(n14224), .A(n14066), .ZN(P1_U3268) );
  NAND2_X1 U15998 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  NAND3_X1 U15999 ( .A1(n14070), .A2(n14522), .A3(n14069), .ZN(n14079) );
  AOI22_X1 U16000 ( .A1(n14072), .A2(n14174), .B1(n14172), .B2(n14071), .ZN(
        n14078) );
  NAND2_X1 U16001 ( .A1(n14073), .A2(n8593), .ZN(n14074) );
  NAND2_X1 U16002 ( .A1(n14075), .A2(n14074), .ZN(n14267) );
  NAND2_X1 U16003 ( .A1(n14267), .A2(n14076), .ZN(n14077) );
  NAND3_X1 U16004 ( .A1(n14079), .A2(n14078), .A3(n14077), .ZN(n14272) );
  INV_X1 U16005 ( .A(n14272), .ZN(n14089) );
  AOI21_X1 U16006 ( .B1(n14095), .B2(n14266), .A(n14252), .ZN(n14082) );
  NAND2_X1 U16007 ( .A1(n14082), .A2(n14081), .ZN(n14268) );
  AOI22_X1 U16008 ( .A1(n14224), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14083), 
        .B2(n14222), .ZN(n14085) );
  NAND2_X1 U16009 ( .A1(n14266), .A2(n14225), .ZN(n14084) );
  OAI211_X1 U16010 ( .C1(n14268), .C2(n14516), .A(n14085), .B(n14084), .ZN(
        n14086) );
  AOI21_X1 U16011 ( .B1(n14267), .B2(n14087), .A(n14086), .ZN(n14088) );
  OAI21_X1 U16012 ( .B1(n14089), .B2(n14224), .A(n14088), .ZN(P1_U3269) );
  OAI21_X1 U16013 ( .B1(n14091), .B2(n14100), .A(n14090), .ZN(n14094) );
  AOI222_X1 U16014 ( .A1(n14522), .A2(n14094), .B1(n14093), .B2(n14172), .C1(
        n14092), .C2(n14174), .ZN(n14281) );
  AOI211_X1 U16015 ( .C1(n14276), .C2(n14112), .A(n14252), .B(n14080), .ZN(
        n14275) );
  NOR2_X1 U16016 ( .A1(n6864), .A2(n14525), .ZN(n14099) );
  OAI22_X1 U16017 ( .A1(n14529), .A2(n14097), .B1(n14096), .B2(n14526), .ZN(
        n14098) );
  AOI211_X1 U16018 ( .C1(n14275), .C2(n14194), .A(n14099), .B(n14098), .ZN(
        n14103) );
  NAND2_X1 U16019 ( .A1(n14101), .A2(n14100), .ZN(n14277) );
  NAND3_X1 U16020 ( .A1(n14278), .A2(n14277), .A3(n14233), .ZN(n14102) );
  OAI211_X1 U16021 ( .C1(n14281), .C2(n14224), .A(n14103), .B(n14102), .ZN(
        P1_U3270) );
  XNOR2_X1 U16022 ( .A(n14104), .B(n8571), .ZN(n14286) );
  INV_X1 U16023 ( .A(n14105), .ZN(n14106) );
  AOI21_X1 U16024 ( .B1(n14108), .B2(n14107), .A(n14106), .ZN(n14111) );
  OAI21_X1 U16025 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14282) );
  INV_X1 U16026 ( .A(n14112), .ZN(n14113) );
  AOI211_X1 U16027 ( .C1(n14284), .C2(n6868), .A(n14252), .B(n14113), .ZN(
        n14283) );
  INV_X1 U16028 ( .A(n14283), .ZN(n14115) );
  OAI22_X1 U16029 ( .A1(n14115), .A2(n11760), .B1(n14526), .B2(n14114), .ZN(
        n14116) );
  OAI21_X1 U16030 ( .B1(n14282), .B2(n14116), .A(n14529), .ZN(n14118) );
  AOI22_X1 U16031 ( .A1(n14284), .A2(n14225), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14224), .ZN(n14117) );
  OAI211_X1 U16032 ( .C1(n14201), .C2(n14286), .A(n14118), .B(n14117), .ZN(
        P1_U3271) );
  XNOR2_X1 U16033 ( .A(n14119), .B(n14120), .ZN(n14122) );
  AOI21_X1 U16034 ( .B1(n14122), .B2(n14522), .A(n14121), .ZN(n14290) );
  AOI211_X1 U16035 ( .C1(n14288), .C2(n14146), .A(n14252), .B(n14123), .ZN(
        n14287) );
  INV_X1 U16036 ( .A(n14288), .ZN(n14127) );
  INV_X1 U16037 ( .A(n14124), .ZN(n14125) );
  AOI22_X1 U16038 ( .A1(n14224), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14125), 
        .B2(n14222), .ZN(n14126) );
  OAI21_X1 U16039 ( .B1(n14127), .B2(n14525), .A(n14126), .ZN(n14131) );
  AOI21_X1 U16040 ( .B1(n14129), .B2(n14128), .A(n6580), .ZN(n14291) );
  NOR2_X1 U16041 ( .A1(n14291), .A2(n14201), .ZN(n14130) );
  AOI211_X1 U16042 ( .C1(n14287), .C2(n14194), .A(n14131), .B(n14130), .ZN(
        n14132) );
  OAI21_X1 U16043 ( .B1(n14224), .B2(n14290), .A(n14132), .ZN(P1_U3272) );
  NAND2_X1 U16044 ( .A1(n14134), .A2(n14133), .ZN(n14135) );
  NAND2_X1 U16045 ( .A1(n14135), .A2(n7159), .ZN(n14136) );
  NAND2_X1 U16046 ( .A1(n14137), .A2(n14136), .ZN(n14295) );
  XNOR2_X1 U16047 ( .A(n14138), .B(n7159), .ZN(n14139) );
  NAND2_X1 U16048 ( .A1(n14139), .A2(n14522), .ZN(n14142) );
  AOI22_X1 U16049 ( .A1(n14140), .A2(n14172), .B1(n14174), .B2(n14173), .ZN(
        n14141) );
  NAND2_X1 U16050 ( .A1(n14142), .A2(n14141), .ZN(n14297) );
  NAND2_X1 U16051 ( .A1(n14297), .A2(n14529), .ZN(n14151) );
  INV_X1 U16052 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14144) );
  OAI22_X1 U16053 ( .A1(n14529), .A2(n14144), .B1(n14143), .B2(n14526), .ZN(
        n14149) );
  INV_X1 U16054 ( .A(n14145), .ZN(n14156) );
  AOI21_X1 U16055 ( .B1(n14156), .B2(n14292), .A(n14252), .ZN(n14147) );
  NAND2_X1 U16056 ( .A1(n14147), .A2(n14146), .ZN(n14294) );
  NOR2_X1 U16057 ( .A1(n14294), .A2(n14516), .ZN(n14148) );
  AOI211_X1 U16058 ( .C1(n14225), .C2(n14292), .A(n14149), .B(n14148), .ZN(
        n14150) );
  OAI211_X1 U16059 ( .C1(n14201), .C2(n14295), .A(n14151), .B(n14150), .ZN(
        P1_U3273) );
  OR2_X1 U16060 ( .A1(n14181), .A2(n14152), .ZN(n14154) );
  NAND2_X1 U16061 ( .A1(n14154), .A2(n14153), .ZN(n14155) );
  XNOR2_X1 U16062 ( .A(n14155), .B(n14161), .ZN(n14302) );
  AOI21_X1 U16063 ( .B1(n14298), .B2(n14176), .A(n14145), .ZN(n14299) );
  AOI22_X1 U16064 ( .A1(n14224), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14157), 
        .B2(n14222), .ZN(n14158) );
  OAI21_X1 U16065 ( .B1(n14159), .B2(n14525), .A(n14158), .ZN(n14167) );
  OAI21_X1 U16066 ( .B1(n14162), .B2(n14161), .A(n14160), .ZN(n14165) );
  AOI222_X1 U16067 ( .A1(n14522), .A2(n14165), .B1(n14164), .B2(n14172), .C1(
        n14163), .C2(n14174), .ZN(n14301) );
  NOR2_X1 U16068 ( .A1(n14301), .A2(n14224), .ZN(n14166) );
  AOI211_X1 U16069 ( .C1(n14299), .C2(n14168), .A(n14167), .B(n14166), .ZN(
        n14169) );
  OAI21_X1 U16070 ( .B1(n14201), .B2(n14302), .A(n14169), .ZN(P1_U3274) );
  XOR2_X1 U16071 ( .A(n14170), .B(n14182), .Z(n14171) );
  AOI222_X1 U16072 ( .A1(n14175), .A2(n14174), .B1(n14173), .B2(n14172), .C1(
        n14522), .C2(n14171), .ZN(n14306) );
  INV_X1 U16073 ( .A(n14176), .ZN(n14177) );
  AOI211_X1 U16074 ( .C1(n14304), .C2(n14192), .A(n14252), .B(n14177), .ZN(
        n14303) );
  AOI22_X1 U16075 ( .A1(n14224), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14178), 
        .B2(n14222), .ZN(n14179) );
  OAI21_X1 U16076 ( .B1(n14180), .B2(n14525), .A(n14179), .ZN(n14184) );
  XOR2_X1 U16077 ( .A(n14182), .B(n14181), .Z(n14307) );
  NOR2_X1 U16078 ( .A1(n14307), .A2(n14201), .ZN(n14183) );
  AOI211_X1 U16079 ( .C1(n14303), .C2(n14194), .A(n14184), .B(n14183), .ZN(
        n14185) );
  OAI21_X1 U16080 ( .B1(n14306), .B2(n14224), .A(n14185), .ZN(P1_U3275) );
  XNOR2_X1 U16081 ( .A(n14186), .B(n14189), .ZN(n14312) );
  OAI211_X1 U16082 ( .C1(n14189), .C2(n14188), .A(n14187), .B(n14522), .ZN(
        n14191) );
  NAND2_X1 U16083 ( .A1(n14191), .A2(n14190), .ZN(n14308) );
  AOI21_X1 U16084 ( .B1(n14310), .B2(n14203), .A(n14252), .ZN(n14193) );
  AND2_X1 U16085 ( .A1(n14193), .A2(n14192), .ZN(n14309) );
  NAND2_X1 U16086 ( .A1(n14309), .A2(n14194), .ZN(n14197) );
  AOI22_X1 U16087 ( .A1(n14224), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14195), 
        .B2(n14222), .ZN(n14196) );
  OAI211_X1 U16088 ( .C1(n14198), .C2(n14525), .A(n14197), .B(n14196), .ZN(
        n14199) );
  AOI21_X1 U16089 ( .B1(n14308), .B2(n14529), .A(n14199), .ZN(n14200) );
  OAI21_X1 U16090 ( .B1(n14201), .B2(n14312), .A(n14200), .ZN(P1_U3276) );
  XNOR2_X1 U16091 ( .A(n14202), .B(n14208), .ZN(n14314) );
  OAI211_X1 U16092 ( .C1(n14365), .C2(n6693), .A(n14512), .B(n14203), .ZN(
        n14315) );
  OAI22_X1 U16093 ( .A1(n14529), .A2(n13963), .B1(n14204), .B2(n14526), .ZN(
        n14205) );
  AOI21_X1 U16094 ( .B1(n14206), .B2(n14225), .A(n14205), .ZN(n14207) );
  OAI21_X1 U16095 ( .B1(n14315), .B2(n14516), .A(n14207), .ZN(n14217) );
  XNOR2_X1 U16096 ( .A(n14209), .B(n14208), .ZN(n14215) );
  OAI22_X1 U16097 ( .A1(n14213), .A2(n14212), .B1(n14211), .B2(n14210), .ZN(
        n14214) );
  AOI21_X1 U16098 ( .B1(n14215), .B2(n14522), .A(n14214), .ZN(n14317) );
  NOR2_X1 U16099 ( .A1(n14317), .A2(n14224), .ZN(n14216) );
  AOI211_X1 U16100 ( .C1(n14314), .C2(n14233), .A(n14217), .B(n14216), .ZN(
        n14218) );
  INV_X1 U16101 ( .A(n14218), .ZN(P1_U3277) );
  XNOR2_X1 U16102 ( .A(n14219), .B(n14228), .ZN(n14325) );
  XOR2_X1 U16103 ( .A(n14220), .B(n14320), .Z(n14221) );
  NAND2_X1 U16104 ( .A1(n14221), .A2(n14512), .ZN(n14321) );
  AOI22_X1 U16105 ( .A1(n14224), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14223), 
        .B2(n14222), .ZN(n14227) );
  NAND2_X1 U16106 ( .A1(n14320), .A2(n14225), .ZN(n14226) );
  OAI211_X1 U16107 ( .C1(n14321), .C2(n14516), .A(n14227), .B(n14226), .ZN(
        n14232) );
  XNOR2_X1 U16108 ( .A(n14229), .B(n14228), .ZN(n14230) );
  NAND2_X1 U16109 ( .A1(n14230), .A2(n14522), .ZN(n14323) );
  AOI21_X1 U16110 ( .B1(n14323), .B2(n14322), .A(n14224), .ZN(n14231) );
  AOI211_X1 U16111 ( .C1(n14325), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14234) );
  INV_X1 U16112 ( .A(n14234), .ZN(P1_U3278) );
  INV_X1 U16113 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15320) );
  MUX2_X1 U16114 ( .A(n15320), .B(n14337), .S(n14803), .Z(n14237) );
  OAI21_X1 U16115 ( .B1(n14340), .B2(n14327), .A(n14237), .ZN(P1_U3559) );
  AND2_X1 U16116 ( .A1(n14239), .A2(n14238), .ZN(n14342) );
  MUX2_X1 U16117 ( .A(n14342), .B(n14240), .S(n14800), .Z(n14241) );
  OAI21_X1 U16118 ( .B1(n14344), .B2(n14327), .A(n14241), .ZN(P1_U3558) );
  AOI21_X1 U16119 ( .B1(n14330), .B2(n14243), .A(n14242), .ZN(n14244) );
  OAI211_X1 U16120 ( .C1(n14313), .C2(n14246), .A(n14245), .B(n14244), .ZN(
        n14345) );
  MUX2_X1 U16121 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14345), .S(n14803), .Z(
        P1_U3556) );
  AOI21_X1 U16122 ( .B1(n14330), .B2(n14248), .A(n14247), .ZN(n14249) );
  OAI211_X1 U16123 ( .C1(n14251), .C2(n14313), .A(n14250), .B(n14249), .ZN(
        n14346) );
  MUX2_X1 U16124 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14346), .S(n14803), .Z(
        P1_U3555) );
  INV_X1 U16125 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14257) );
  OAI22_X1 U16126 ( .A1(n14254), .A2(n14313), .B1(n14253), .B2(n14252), .ZN(
        n14255) );
  NOR2_X1 U16127 ( .A1(n14256), .A2(n14255), .ZN(n14347) );
  MUX2_X1 U16128 ( .A(n14257), .B(n14347), .S(n14803), .Z(n14258) );
  OAI21_X1 U16129 ( .B1(n14350), .B2(n14327), .A(n14258), .ZN(P1_U3554) );
  NAND2_X1 U16130 ( .A1(n14259), .A2(n14330), .ZN(n14264) );
  NAND3_X1 U16131 ( .A1(n14261), .A2(n14793), .A3(n14260), .ZN(n14263) );
  NAND4_X1 U16132 ( .A1(n14265), .A2(n14264), .A3(n14263), .A4(n14262), .ZN(
        n14351) );
  MUX2_X1 U16133 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14351), .S(n14803), .Z(
        P1_U3553) );
  INV_X1 U16134 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14273) );
  INV_X1 U16135 ( .A(n14266), .ZN(n14270) );
  NAND2_X1 U16136 ( .A1(n14267), .A2(n14781), .ZN(n14269) );
  OAI211_X1 U16137 ( .C1(n14270), .C2(n14788), .A(n14269), .B(n14268), .ZN(
        n14271) );
  NOR2_X1 U16138 ( .A1(n14272), .A2(n14271), .ZN(n14352) );
  MUX2_X1 U16139 ( .A(n14273), .B(n14352), .S(n14803), .Z(n14274) );
  INV_X1 U16140 ( .A(n14274), .ZN(P1_U3552) );
  AOI21_X1 U16141 ( .B1(n14330), .B2(n14276), .A(n14275), .ZN(n14280) );
  NAND3_X1 U16142 ( .A1(n14278), .A2(n14277), .A3(n14793), .ZN(n14279) );
  NAND3_X1 U16143 ( .A1(n14281), .A2(n14280), .A3(n14279), .ZN(n14355) );
  MUX2_X1 U16144 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14355), .S(n14803), .Z(
        P1_U3551) );
  AOI211_X1 U16145 ( .C1(n14330), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n14285) );
  OAI21_X1 U16146 ( .B1(n14313), .B2(n14286), .A(n14285), .ZN(n14356) );
  MUX2_X1 U16147 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14356), .S(n14803), .Z(
        P1_U3550) );
  AOI21_X1 U16148 ( .B1(n14330), .B2(n14288), .A(n14287), .ZN(n14289) );
  OAI211_X1 U16149 ( .C1(n14313), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        n14357) );
  MUX2_X1 U16150 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14357), .S(n14803), .Z(
        P1_U3549) );
  NAND2_X1 U16151 ( .A1(n14292), .A2(n14330), .ZN(n14293) );
  OAI211_X1 U16152 ( .C1(n14295), .C2(n14313), .A(n14294), .B(n14293), .ZN(
        n14296) );
  MUX2_X1 U16153 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14358), .S(n14803), .Z(
        P1_U3548) );
  AOI22_X1 U16154 ( .A1(n14299), .A2(n14512), .B1(n14330), .B2(n14298), .ZN(
        n14300) );
  OAI211_X1 U16155 ( .C1(n14313), .C2(n14302), .A(n14301), .B(n14300), .ZN(
        n14359) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14359), .S(n14803), .Z(
        P1_U3547) );
  AOI21_X1 U16157 ( .B1(n14330), .B2(n14304), .A(n14303), .ZN(n14305) );
  OAI211_X1 U16158 ( .C1(n14313), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        n14360) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14360), .S(n14803), .Z(
        P1_U3546) );
  AOI211_X1 U16160 ( .C1(n14330), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        n14311) );
  OAI21_X1 U16161 ( .B1(n14313), .B2(n14312), .A(n14311), .ZN(n14361) );
  MUX2_X1 U16162 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14361), .S(n14803), .Z(
        P1_U3545) );
  INV_X1 U16163 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14318) );
  NAND2_X1 U16164 ( .A1(n14314), .A2(n14793), .ZN(n14316) );
  AND3_X1 U16165 ( .A1(n14317), .A2(n14316), .A3(n14315), .ZN(n14362) );
  MUX2_X1 U16166 ( .A(n14318), .B(n14362), .S(n14803), .Z(n14319) );
  OAI21_X1 U16167 ( .B1(n14365), .B2(n14327), .A(n14319), .ZN(P1_U3544) );
  INV_X1 U16168 ( .A(n14320), .ZN(n14369) );
  NAND3_X1 U16169 ( .A1(n14323), .A2(n14322), .A3(n14321), .ZN(n14324) );
  AOI21_X1 U16170 ( .B1(n14325), .B2(n14793), .A(n14324), .ZN(n14366) );
  MUX2_X1 U16171 ( .A(n14705), .B(n14366), .S(n14803), .Z(n14326) );
  OAI21_X1 U16172 ( .B1(n14369), .B2(n14327), .A(n14326), .ZN(P1_U3543) );
  AOI21_X1 U16173 ( .B1(n14330), .B2(n14329), .A(n14328), .ZN(n14334) );
  NAND3_X1 U16174 ( .A1(n14332), .A2(n14331), .A3(n14793), .ZN(n14333) );
  NAND3_X1 U16175 ( .A1(n14335), .A2(n14334), .A3(n14333), .ZN(n14370) );
  MUX2_X1 U16176 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14370), .S(n14803), .Z(
        P1_U3542) );
  MUX2_X1 U16177 ( .A(n14336), .B(P1_REG1_REG_0__SCAN_IN), .S(n14800), .Z(
        P1_U3528) );
  INV_X1 U16178 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14338) );
  MUX2_X1 U16179 ( .A(n14338), .B(n14337), .S(n14796), .Z(n14339) );
  OAI21_X1 U16180 ( .B1(n14340), .B2(n8752), .A(n14339), .ZN(P1_U3527) );
  INV_X1 U16181 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14341) );
  MUX2_X1 U16182 ( .A(n14342), .B(n14341), .S(n14794), .Z(n14343) );
  OAI21_X1 U16183 ( .B1(n14344), .B2(n8752), .A(n14343), .ZN(P1_U3526) );
  MUX2_X1 U16184 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14345), .S(n14796), .Z(
        P1_U3524) );
  MUX2_X1 U16185 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14346), .S(n14796), .Z(
        P1_U3523) );
  INV_X1 U16186 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14348) );
  MUX2_X1 U16187 ( .A(n14348), .B(n14347), .S(n14796), .Z(n14349) );
  OAI21_X1 U16188 ( .B1(n14350), .B2(n8752), .A(n14349), .ZN(P1_U3522) );
  MUX2_X1 U16189 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14351), .S(n14796), .Z(
        P1_U3521) );
  INV_X1 U16190 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14353) );
  MUX2_X1 U16191 ( .A(n14353), .B(n14352), .S(n14796), .Z(n14354) );
  INV_X1 U16192 ( .A(n14354), .ZN(P1_U3520) );
  MUX2_X1 U16193 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14355), .S(n14796), .Z(
        P1_U3519) );
  MUX2_X1 U16194 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14356), .S(n14796), .Z(
        P1_U3518) );
  MUX2_X1 U16195 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14357), .S(n14796), .Z(
        P1_U3517) );
  MUX2_X1 U16196 ( .A(n14358), .B(P1_REG0_REG_20__SCAN_IN), .S(n14794), .Z(
        P1_U3516) );
  MUX2_X1 U16197 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14359), .S(n14796), .Z(
        P1_U3515) );
  MUX2_X1 U16198 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14360), .S(n14796), .Z(
        P1_U3513) );
  MUX2_X1 U16199 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14361), .S(n14796), .Z(
        P1_U3510) );
  INV_X1 U16200 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14363) );
  MUX2_X1 U16201 ( .A(n14363), .B(n14362), .S(n14796), .Z(n14364) );
  OAI21_X1 U16202 ( .B1(n14365), .B2(n8752), .A(n14364), .ZN(P1_U3507) );
  INV_X1 U16203 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14367) );
  MUX2_X1 U16204 ( .A(n14367), .B(n14366), .S(n14796), .Z(n14368) );
  OAI21_X1 U16205 ( .B1(n14369), .B2(n8752), .A(n14368), .ZN(P1_U3504) );
  MUX2_X1 U16206 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n14370), .S(n14796), .Z(
        P1_U3501) );
  NOR4_X1 U16207 ( .A1(n14373), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14371), .ZN(n14374) );
  AOI21_X1 U16208 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14375), .A(n14374), 
        .ZN(n14376) );
  OAI21_X1 U16209 ( .B1(n14377), .B2(n14390), .A(n14376), .ZN(P1_U3324) );
  OAI222_X1 U16210 ( .A1(P1_U3086), .A2(n14380), .B1(n14390), .B2(n14379), 
        .C1(n14378), .C2(n14384), .ZN(P1_U3325) );
  OAI222_X1 U16211 ( .A1(P1_U3086), .A2(n14383), .B1(n14390), .B2(n14382), 
        .C1(n14381), .C2(n14384), .ZN(P1_U3326) );
  OAI222_X1 U16212 ( .A1(P1_U3086), .A2(n6705), .B1(n14390), .B2(n14386), .C1(
        n14385), .C2(n14384), .ZN(P1_U3328) );
  OAI222_X1 U16213 ( .A1(n14391), .A2(P1_U3086), .B1(n14390), .B2(n14389), 
        .C1(n14388), .C2(n14384), .ZN(P1_U3329) );
  MUX2_X1 U16214 ( .A(n14393), .B(n14392), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16215 ( .A(n14394), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16216 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14684) );
  INV_X1 U16217 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14472) );
  INV_X1 U16218 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14411) );
  XNOR2_X1 U16219 ( .A(n14411), .B(n14395), .ZN(n14463) );
  NAND2_X1 U16220 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n15377), .ZN(n14396) );
  XOR2_X1 U16221 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14434) );
  NOR2_X1 U16222 ( .A1(n14402), .A2(n14401), .ZN(n14404) );
  NOR2_X1 U16223 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n15395), .ZN(n14405) );
  INV_X1 U16224 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14969) );
  NOR2_X1 U16225 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14406), .ZN(n14408) );
  XNOR2_X1 U16226 ( .A(n14406), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14456) );
  XNOR2_X1 U16227 ( .A(n15003), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14429) );
  NAND2_X1 U16228 ( .A1(n14463), .A2(n14462), .ZN(n14410) );
  NOR2_X1 U16229 ( .A1(n14412), .A2(n14466), .ZN(n14414) );
  INV_X1 U16230 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U16231 ( .A1(n14412), .A2(n14466), .ZN(n14413) );
  NAND2_X1 U16232 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14426), .ZN(n14415) );
  AND2_X1 U16233 ( .A1(n14472), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n14417) );
  INV_X1 U16234 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U16235 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15009), .ZN(n14418) );
  INV_X1 U16236 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U16237 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n14699), .ZN(n14419) );
  INV_X1 U16238 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U16239 ( .A1(n14480), .A2(n14419), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14479), .ZN(n14484) );
  INV_X1 U16240 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U16241 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14567), .ZN(n14483) );
  NOR2_X1 U16242 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14567), .ZN(n14420) );
  AOI21_X1 U16243 ( .B1(n14484), .B2(n14483), .A(n14420), .ZN(n14491) );
  INV_X1 U16244 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14729) );
  NAND2_X1 U16245 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14729), .ZN(n14421) );
  AOI22_X1 U16246 ( .A1(n14491), .A2(n14421), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n15245), .ZN(n14422) );
  INV_X1 U16247 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14744) );
  NAND2_X1 U16248 ( .A1(n14422), .A2(n14744), .ZN(n14424) );
  XOR2_X1 U16249 ( .A(n14744), .B(n14422), .Z(n14493) );
  NAND2_X1 U16250 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14493), .ZN(n14423) );
  NAND2_X1 U16251 ( .A1(n14424), .A2(n14423), .ZN(n14554) );
  INV_X1 U16252 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14557) );
  NOR2_X1 U16253 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14557), .ZN(n14425) );
  AOI21_X1 U16254 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14557), .A(n14425), 
        .ZN(n14555) );
  XNOR2_X1 U16255 ( .A(n14554), .B(n14555), .ZN(n14550) );
  INV_X1 U16256 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14494) );
  INV_X1 U16257 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14492) );
  INV_X1 U16258 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14847) );
  INV_X1 U16259 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14471) );
  XNOR2_X1 U16260 ( .A(n14426), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n14427) );
  XOR2_X1 U16261 ( .A(n14428), .B(n14427), .Z(n14653) );
  INV_X1 U16262 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14465) );
  XOR2_X1 U16263 ( .A(n14430), .B(n14429), .Z(n14461) );
  NAND2_X1 U16264 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14432), .ZN(n14444) );
  XNOR2_X1 U16265 ( .A(n14434), .B(n14433), .ZN(n14440) );
  XNOR2_X1 U16266 ( .A(n14435), .B(n14436), .ZN(n14437) );
  NAND2_X1 U16267 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14437), .ZN(n14438) );
  AOI21_X1 U16268 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14952), .A(n14436), .ZN(
        n15474) );
  NOR2_X1 U16269 ( .A1(n15474), .A2(n11741), .ZN(n15482) );
  NOR2_X1 U16270 ( .A1(n14440), .A2(n14439), .ZN(n14498) );
  XOR2_X1 U16271 ( .A(n14442), .B(n14441), .Z(n15478) );
  NAND2_X1 U16272 ( .A1(n15479), .A2(n15478), .ZN(n14443) );
  NOR2_X1 U16273 ( .A1(n15479), .A2(n15478), .ZN(n15477) );
  NOR2_X1 U16274 ( .A1(n14448), .A2(n14447), .ZN(n14450) );
  NOR2_X1 U16275 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15473), .ZN(n14449) );
  NAND2_X1 U16276 ( .A1(n14451), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14454) );
  XNOR2_X1 U16277 ( .A(n15395), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n14452) );
  XNOR2_X1 U16278 ( .A(n14453), .B(n14452), .ZN(n14500) );
  NAND2_X1 U16279 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14455), .ZN(n14459) );
  INV_X1 U16280 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15301) );
  XOR2_X1 U16281 ( .A(n14457), .B(n14456), .Z(n15475) );
  NAND2_X1 U16282 ( .A1(n15476), .A2(n15475), .ZN(n14458) );
  XNOR2_X1 U16283 ( .A(n14463), .B(n14462), .ZN(n14504) );
  NAND2_X1 U16284 ( .A1(n14505), .A2(n14504), .ZN(n14464) );
  XNOR2_X1 U16285 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14466), .ZN(n14467) );
  XOR2_X1 U16286 ( .A(n14468), .B(n14467), .Z(n14509) );
  INV_X1 U16287 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U16288 ( .A1(n14508), .A2(n14509), .ZN(n14507) );
  XOR2_X1 U16289 ( .A(n14472), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14474) );
  XOR2_X1 U16290 ( .A(n14474), .B(n14473), .Z(n14657) );
  XNOR2_X1 U16291 ( .A(n15009), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14475) );
  XOR2_X1 U16292 ( .A(n14476), .B(n14475), .Z(n14477) );
  NOR2_X1 U16293 ( .A1(n14478), .A2(n14477), .ZN(n14660) );
  XOR2_X1 U16294 ( .A(n14479), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14481) );
  XOR2_X1 U16295 ( .A(n14481), .B(n14480), .Z(n14664) );
  NAND2_X1 U16296 ( .A1(n14663), .A2(n14664), .ZN(n14482) );
  OAI21_X1 U16297 ( .B1(n14567), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n14483), 
        .ZN(n14485) );
  XOR2_X1 U16298 ( .A(n14485), .B(n14484), .Z(n14487) );
  NOR2_X1 U16299 ( .A1(n14486), .A2(n14487), .ZN(n14667) );
  NAND2_X1 U16300 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15245), .ZN(n14489) );
  OAI21_X1 U16301 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n15245), .A(n14489), 
        .ZN(n14490) );
  XNOR2_X1 U16302 ( .A(n14491), .B(n14490), .ZN(n14671) );
  XNOR2_X1 U16303 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14493), .ZN(n14546) );
  XNOR2_X1 U16304 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14549), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16305 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14495) );
  OAI21_X1 U16306 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14495), 
        .ZN(U28) );
  AOI21_X1 U16307 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14496) );
  OAI21_X1 U16308 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14496), 
        .ZN(U29) );
  NOR2_X1 U16309 ( .A1(n14498), .A2(n14497), .ZN(n14499) );
  XOR2_X1 U16310 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n14499), .Z(SUB_1596_U61) );
  XOR2_X1 U16311 ( .A(n14501), .B(n14500), .Z(SUB_1596_U57) );
  XNOR2_X1 U16312 ( .A(n14502), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U16313 ( .B1(n14505), .B2(n14504), .A(n14503), .ZN(n14506) );
  XOR2_X1 U16314 ( .A(n14506), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI21_X1 U16315 ( .B1(n14509), .B2(n14508), .A(n14507), .ZN(n14510) );
  XOR2_X1 U16316 ( .A(n14510), .B(n14832), .Z(SUB_1596_U70) );
  INV_X1 U16317 ( .A(n14519), .ZN(n14511) );
  XNOR2_X1 U16318 ( .A(n6689), .B(n14511), .ZN(n14535) );
  OAI21_X1 U16319 ( .B1(n14513), .B2(n14538), .A(n14512), .ZN(n14515) );
  OR2_X1 U16320 ( .A1(n14515), .A2(n14514), .ZN(n14537) );
  OAI22_X1 U16321 ( .A1(n14535), .A2(n14517), .B1(n14516), .B2(n14537), .ZN(
        n14518) );
  INV_X1 U16322 ( .A(n14518), .ZN(n14534) );
  NAND2_X1 U16323 ( .A1(n14520), .A2(n14519), .ZN(n14521) );
  NAND3_X1 U16324 ( .A1(n14523), .A2(n14522), .A3(n14521), .ZN(n14539) );
  OAI211_X1 U16325 ( .C1(n14535), .C2(n14524), .A(n14536), .B(n14539), .ZN(
        n14532) );
  NOR2_X1 U16326 ( .A1(n14538), .A2(n14525), .ZN(n14531) );
  INV_X1 U16327 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n14528) );
  OAI22_X1 U16328 ( .A1(n14529), .A2(n14528), .B1(n14527), .B2(n14526), .ZN(
        n14530) );
  AOI211_X1 U16329 ( .C1(n14532), .C2(n14529), .A(n14531), .B(n14530), .ZN(
        n14533) );
  NAND2_X1 U16330 ( .A1(n14534), .A2(n14533), .ZN(P1_U3281) );
  INV_X1 U16331 ( .A(n14535), .ZN(n14542) );
  OAI211_X1 U16332 ( .C1(n14538), .C2(n14788), .A(n14537), .B(n14536), .ZN(
        n14541) );
  INV_X1 U16333 ( .A(n14539), .ZN(n14540) );
  AOI211_X1 U16334 ( .C1(n14793), .C2(n14542), .A(n14541), .B(n14540), .ZN(
        n14544) );
  INV_X1 U16335 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14543) );
  AOI22_X1 U16336 ( .A1(n14796), .A2(n14544), .B1(n14543), .B2(n14794), .ZN(
        P1_U3495) );
  AOI22_X1 U16337 ( .A1(n14803), .A2(n14544), .B1(n10950), .B2(n14800), .ZN(
        P1_U3540) );
  AOI21_X1 U16338 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14548) );
  XOR2_X1 U16339 ( .A(n14548), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16340 ( .A1(n14551), .A2(n14550), .ZN(n14552) );
  NAND2_X1 U16341 ( .A1(n14555), .A2(n14554), .ZN(n14556) );
  OAI21_X1 U16342 ( .B1(n14557), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14556), 
        .ZN(n14560) );
  XNOR2_X1 U16343 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14558) );
  XNOR2_X1 U16344 ( .A(n14558), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14559) );
  XNOR2_X1 U16345 ( .A(n14560), .B(n14559), .ZN(n14561) );
  XNOR2_X1 U16346 ( .A(n14562), .B(n14561), .ZN(SUB_1596_U4) );
  AOI21_X1 U16347 ( .B1(n14565), .B2(n14564), .A(n14563), .ZN(n14580) );
  OAI22_X1 U16348 ( .A1(n14567), .A2(n15008), .B1(n15007), .B2(n14566), .ZN(
        n14577) );
  AOI21_X1 U16349 ( .B1(n14570), .B2(n14569), .A(n14568), .ZN(n14575) );
  AOI21_X1 U16350 ( .B1(n14573), .B2(n14572), .A(n14571), .ZN(n14574) );
  OAI22_X1 U16351 ( .A1(n14575), .A2(n15017), .B1(n14574), .B2(n15015), .ZN(
        n14576) );
  NOR3_X1 U16352 ( .A1(n14578), .A2(n14577), .A3(n14576), .ZN(n14579) );
  OAI21_X1 U16353 ( .B1(n14580), .B2(n15023), .A(n14579), .ZN(P3_U3197) );
  NAND2_X1 U16354 ( .A1(n14597), .A2(n14581), .ZN(n14583) );
  AND2_X1 U16355 ( .A1(n14583), .A2(n14582), .ZN(n14585) );
  XNOR2_X1 U16356 ( .A(n14585), .B(n14584), .ZN(n14609) );
  NAND2_X1 U16357 ( .A1(n14587), .A2(n14586), .ZN(n14589) );
  XNOR2_X1 U16358 ( .A(n14589), .B(n14588), .ZN(n14590) );
  OAI222_X1 U16359 ( .A1(n15105), .A2(n14591), .B1(n15107), .B2(n14602), .C1(
        n14590), .C2(n15110), .ZN(n14607) );
  AOI21_X1 U16360 ( .B1(n14609), .B2(n15064), .A(n14607), .ZN(n14596) );
  INV_X1 U16361 ( .A(n14592), .ZN(n14593) );
  NOR2_X1 U16362 ( .A1(n14593), .A2(n15098), .ZN(n14608) );
  AOI22_X1 U16363 ( .A1(n14608), .A2(n15093), .B1(n15125), .B2(n14594), .ZN(
        n14595) );
  OAI221_X1 U16364 ( .B1(n15038), .B2(n14596), .C1(n15129), .C2(n9368), .A(
        n14595), .ZN(P3_U3220) );
  OAI21_X1 U16365 ( .B1(n7602), .B2(n9339), .A(n14597), .ZN(n14618) );
  INV_X1 U16366 ( .A(n15044), .ZN(n14601) );
  XNOR2_X1 U16367 ( .A(n6746), .B(n14598), .ZN(n14600) );
  OAI222_X1 U16368 ( .A1(n15105), .A2(n14602), .B1(n15107), .B2(n14601), .C1(
        n14600), .C2(n15110), .ZN(n14616) );
  AOI21_X1 U16369 ( .B1(n15064), .B2(n14618), .A(n14616), .ZN(n14606) );
  NOR2_X1 U16370 ( .A1(n14603), .A2(n15098), .ZN(n14617) );
  AOI22_X1 U16371 ( .A1(n14617), .A2(n15093), .B1(n14604), .B2(n15125), .ZN(
        n14605) );
  OAI221_X1 U16372 ( .B1(n15038), .B2(n14606), .C1(n15129), .C2(n9325), .A(
        n14605), .ZN(P3_U3222) );
  AOI211_X1 U16373 ( .C1(n14609), .C2(n15162), .A(n14608), .B(n14607), .ZN(
        n14620) );
  AOI22_X1 U16374 ( .A1(n15181), .A2(n14620), .B1(n9365), .B2(n15179), .ZN(
        P3_U3472) );
  OAI22_X1 U16375 ( .A1(n14612), .A2(n14611), .B1(n14610), .B2(n15098), .ZN(
        n14613) );
  NOR2_X1 U16376 ( .A1(n14614), .A2(n14613), .ZN(n14622) );
  AOI22_X1 U16377 ( .A1(n15181), .A2(n14622), .B1(n14615), .B2(n15179), .ZN(
        P3_U3471) );
  AOI211_X1 U16378 ( .C1(n15162), .C2(n14618), .A(n14617), .B(n14616), .ZN(
        n14624) );
  AOI22_X1 U16379 ( .A1(n15181), .A2(n14624), .B1(n9324), .B2(n15179), .ZN(
        P3_U3470) );
  INV_X1 U16380 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14619) );
  AOI22_X1 U16381 ( .A1(n15170), .A2(n14620), .B1(n14619), .B2(n15169), .ZN(
        P3_U3429) );
  INV_X1 U16382 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U16383 ( .A1(n15170), .A2(n14622), .B1(n14621), .B2(n15169), .ZN(
        P3_U3426) );
  INV_X1 U16384 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U16385 ( .A1(n15170), .A2(n14624), .B1(n14623), .B2(n15169), .ZN(
        P3_U3423) );
  INV_X1 U16386 ( .A(n14625), .ZN(n14629) );
  INV_X1 U16387 ( .A(n14626), .ZN(n14628) );
  AOI21_X1 U16388 ( .B1(n14629), .B2(n14628), .A(n14627), .ZN(n14632) );
  OAI21_X1 U16389 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14634) );
  AOI222_X1 U16390 ( .A1(n14638), .A2(n14637), .B1(n14636), .B2(n14635), .C1(
        n14634), .C2(n14633), .ZN(n14641) );
  INV_X1 U16391 ( .A(n14639), .ZN(n14640) );
  OAI211_X1 U16392 ( .C1(n14643), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        P2_U3198) );
  OAI21_X1 U16393 ( .B1(n14645), .B2(n14788), .A(n14644), .ZN(n14647) );
  AOI211_X1 U16394 ( .C1(n14648), .C2(n14793), .A(n14647), .B(n14646), .ZN(
        n14650) );
  AOI22_X1 U16395 ( .A1(n14803), .A2(n14650), .B1(n13979), .B2(n14800), .ZN(
        P1_U3541) );
  INV_X1 U16396 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U16397 ( .A1(n14796), .A2(n14650), .B1(n14649), .B2(n14794), .ZN(
        P1_U3498) );
  AOI21_X1 U16398 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14654) );
  XOR2_X1 U16399 ( .A(n14654), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16400 ( .B1(n14657), .B2(n14656), .A(n14655), .ZN(n14658) );
  XOR2_X1 U16401 ( .A(n14658), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  NOR2_X1 U16402 ( .A1(n14660), .A2(n14659), .ZN(n14661) );
  XOR2_X1 U16403 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14661), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16404 ( .B1(n14664), .B2(n14663), .A(n14662), .ZN(n14665) );
  XOR2_X1 U16405 ( .A(n14665), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  INV_X1 U16406 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15453) );
  NOR2_X1 U16407 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  XNOR2_X1 U16408 ( .A(n15453), .B(n14668), .ZN(SUB_1596_U65) );
  AOI21_X1 U16409 ( .B1(n14671), .B2(n14670), .A(n14669), .ZN(n14672) );
  XOR2_X1 U16410 ( .A(n14672), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI211_X1 U16411 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14715), .ZN(
        n14680) );
  AOI211_X1 U16412 ( .C1(n14678), .C2(n14677), .A(n14676), .B(n14719), .ZN(
        n14679) );
  AOI211_X1 U16413 ( .C1(n14726), .C2(n14681), .A(n14680), .B(n14679), .ZN(
        n14683) );
  OAI211_X1 U16414 ( .C1(n14684), .C2(n14761), .A(n14683), .B(n14682), .ZN(
        P1_U3256) );
  AOI21_X1 U16415 ( .B1(n14687), .B2(n14686), .A(n14685), .ZN(n14688) );
  NAND2_X1 U16416 ( .A1(n14749), .A2(n14688), .ZN(n14694) );
  OAI21_X1 U16417 ( .B1(n14691), .B2(n14690), .A(n14689), .ZN(n14692) );
  NAND2_X1 U16418 ( .A1(n14753), .A2(n14692), .ZN(n14693) );
  OAI211_X1 U16419 ( .C1(n14757), .C2(n14695), .A(n14694), .B(n14693), .ZN(
        n14696) );
  INV_X1 U16420 ( .A(n14696), .ZN(n14698) );
  OAI211_X1 U16421 ( .C1(n14699), .C2(n14761), .A(n14698), .B(n14697), .ZN(
        P1_U3257) );
  INV_X1 U16422 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14714) );
  OAI21_X1 U16423 ( .B1(n14702), .B2(n14701), .A(n14700), .ZN(n14703) );
  NAND2_X1 U16424 ( .A1(n14749), .A2(n14703), .ZN(n14709) );
  OAI21_X1 U16425 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14707) );
  NAND2_X1 U16426 ( .A1(n14753), .A2(n14707), .ZN(n14708) );
  OAI211_X1 U16427 ( .C1(n14757), .C2(n14710), .A(n14709), .B(n14708), .ZN(
        n14711) );
  INV_X1 U16428 ( .A(n14711), .ZN(n14713) );
  OAI211_X1 U16429 ( .C1(n14714), .C2(n14761), .A(n14713), .B(n14712), .ZN(
        P1_U3258) );
  AOI211_X1 U16430 ( .C1(n14718), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        n14724) );
  AOI211_X1 U16431 ( .C1(n14722), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        n14723) );
  AOI211_X1 U16432 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14728) );
  OAI211_X1 U16433 ( .C1(n14729), .C2(n14761), .A(n14728), .B(n14727), .ZN(
        P1_U3259) );
  AOI21_X1 U16434 ( .B1(n14732), .B2(n14731), .A(n14730), .ZN(n14733) );
  NAND2_X1 U16435 ( .A1(n14749), .A2(n14733), .ZN(n14739) );
  AOI21_X1 U16436 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n14737) );
  NAND2_X1 U16437 ( .A1(n14753), .A2(n14737), .ZN(n14738) );
  OAI211_X1 U16438 ( .C1(n14757), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14741) );
  INV_X1 U16439 ( .A(n14741), .ZN(n14743) );
  OAI211_X1 U16440 ( .C1(n14744), .C2(n14761), .A(n14743), .B(n14742), .ZN(
        P1_U3260) );
  INV_X1 U16441 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14762) );
  AOI21_X1 U16442 ( .B1(n14747), .B2(n14746), .A(n14745), .ZN(n14748) );
  NAND2_X1 U16443 ( .A1(n14749), .A2(n14748), .ZN(n14755) );
  AOI21_X1 U16444 ( .B1(n14751), .B2(n15249), .A(n14750), .ZN(n14752) );
  NAND2_X1 U16445 ( .A1(n14753), .A2(n14752), .ZN(n14754) );
  OAI211_X1 U16446 ( .C1(n14757), .C2(n14756), .A(n14755), .B(n14754), .ZN(
        n14758) );
  INV_X1 U16447 ( .A(n14758), .ZN(n14760) );
  OAI211_X1 U16448 ( .C1(n14762), .C2(n14761), .A(n14760), .B(n14759), .ZN(
        P1_U3261) );
  INV_X1 U16449 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15444) );
  NOR2_X1 U16450 ( .A1(n14763), .A2(n15444), .ZN(P1_U3294) );
  AND2_X1 U16451 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14764), .ZN(P1_U3295) );
  AND2_X1 U16452 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14764), .ZN(P1_U3296) );
  AND2_X1 U16453 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14764), .ZN(P1_U3297) );
  AND2_X1 U16454 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14764), .ZN(P1_U3298) );
  AND2_X1 U16455 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14764), .ZN(P1_U3299) );
  AND2_X1 U16456 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14764), .ZN(P1_U3300) );
  INV_X1 U16457 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15318) );
  NOR2_X1 U16458 ( .A1(n14763), .A2(n15318), .ZN(P1_U3301) );
  AND2_X1 U16459 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14764), .ZN(P1_U3302) );
  AND2_X1 U16460 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14764), .ZN(P1_U3303) );
  AND2_X1 U16461 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14764), .ZN(P1_U3304) );
  AND2_X1 U16462 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14764), .ZN(P1_U3305) );
  AND2_X1 U16463 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14764), .ZN(P1_U3306) );
  INV_X1 U16464 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15372) );
  NOR2_X1 U16465 ( .A1(n14763), .A2(n15372), .ZN(P1_U3307) );
  AND2_X1 U16466 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14764), .ZN(P1_U3308) );
  INV_X1 U16467 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15310) );
  NOR2_X1 U16468 ( .A1(n14763), .A2(n15310), .ZN(P1_U3309) );
  AND2_X1 U16469 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14764), .ZN(P1_U3310) );
  INV_X1 U16470 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15410) );
  NOR2_X1 U16471 ( .A1(n14763), .A2(n15410), .ZN(P1_U3311) );
  INV_X1 U16472 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15275) );
  NOR2_X1 U16473 ( .A1(n14763), .A2(n15275), .ZN(P1_U3312) );
  INV_X1 U16474 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15356) );
  NOR2_X1 U16475 ( .A1(n14763), .A2(n15356), .ZN(P1_U3313) );
  AND2_X1 U16476 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14764), .ZN(P1_U3314) );
  AND2_X1 U16477 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14764), .ZN(P1_U3315) );
  AND2_X1 U16478 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14764), .ZN(P1_U3316) );
  AND2_X1 U16479 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14764), .ZN(P1_U3317) );
  AND2_X1 U16480 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14764), .ZN(P1_U3318) );
  AND2_X1 U16481 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14764), .ZN(P1_U3319) );
  AND2_X1 U16482 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14764), .ZN(P1_U3320) );
  AND2_X1 U16483 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14764), .ZN(P1_U3321) );
  AND2_X1 U16484 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14764), .ZN(P1_U3322) );
  AND2_X1 U16485 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14764), .ZN(P1_U3323) );
  OAI21_X1 U16486 ( .B1(n14766), .B2(n14788), .A(n14765), .ZN(n14767) );
  AOI21_X1 U16487 ( .B1(n14768), .B2(n14781), .A(n14767), .ZN(n14769) );
  AND2_X1 U16488 ( .A1(n14770), .A2(n14769), .ZN(n14797) );
  INV_X1 U16489 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14771) );
  AOI22_X1 U16490 ( .A1(n14796), .A2(n14797), .B1(n14771), .B2(n14794), .ZN(
        P1_U3465) );
  OAI211_X1 U16491 ( .C1(n14774), .C2(n14788), .A(n14773), .B(n14772), .ZN(
        n14775) );
  AOI21_X1 U16492 ( .B1(n14793), .B2(n14776), .A(n14775), .ZN(n14798) );
  INV_X1 U16493 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U16494 ( .A1(n14796), .A2(n14798), .B1(n14777), .B2(n14794), .ZN(
        P1_U3471) );
  OAI21_X1 U16495 ( .B1(n14779), .B2(n14788), .A(n14778), .ZN(n14780) );
  AOI21_X1 U16496 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n14783) );
  AND2_X1 U16497 ( .A1(n14784), .A2(n14783), .ZN(n14799) );
  INV_X1 U16498 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14785) );
  AOI22_X1 U16499 ( .A1(n14796), .A2(n14799), .B1(n14785), .B2(n14794), .ZN(
        P1_U3477) );
  OAI211_X1 U16500 ( .C1(n14789), .C2(n14788), .A(n14787), .B(n14786), .ZN(
        n14791) );
  AOI211_X1 U16501 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14802) );
  INV_X1 U16502 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14795) );
  AOI22_X1 U16503 ( .A1(n14796), .A2(n14802), .B1(n14795), .B2(n14794), .ZN(
        P1_U3489) );
  AOI22_X1 U16504 ( .A1(n14803), .A2(n14797), .B1(n10190), .B2(n14800), .ZN(
        P1_U3530) );
  AOI22_X1 U16505 ( .A1(n14803), .A2(n14798), .B1(n10192), .B2(n14800), .ZN(
        P1_U3532) );
  AOI22_X1 U16506 ( .A1(n14803), .A2(n14799), .B1(n10193), .B2(n14800), .ZN(
        P1_U3534) );
  INV_X1 U16507 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16508 ( .A1(n14803), .A2(n14802), .B1(n14801), .B2(n14800), .ZN(
        P1_U3538) );
  NOR2_X1 U16509 ( .A1(n14855), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16510 ( .A1(n14855), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14812) );
  OAI211_X1 U16511 ( .C1(n14806), .C2(n14805), .A(n14833), .B(n14804), .ZN(
        n14811) );
  NAND2_X1 U16512 ( .A1(n14838), .A2(n14807), .ZN(n14810) );
  NAND2_X1 U16513 ( .A1(P2_U3088), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n14809) );
  AND4_X1 U16514 ( .A1(n14812), .A2(n14811), .A3(n14810), .A4(n14809), .ZN(
        n14817) );
  OAI211_X1 U16515 ( .C1(n14815), .C2(n14814), .A(n14857), .B(n14813), .ZN(
        n14816) );
  NAND2_X1 U16516 ( .A1(n14817), .A2(n14816), .ZN(P2_U3216) );
  NOR2_X1 U16517 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7829), .ZN(n14823) );
  INV_X1 U16518 ( .A(n14818), .ZN(n14819) );
  AOI211_X1 U16519 ( .C1(n14821), .C2(n14820), .A(n14850), .B(n14819), .ZN(
        n14822) );
  AOI211_X1 U16520 ( .C1(n14838), .C2(n14824), .A(n14823), .B(n14822), .ZN(
        n14831) );
  AOI21_X1 U16521 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14829) );
  NAND2_X1 U16522 ( .A1(n14829), .A2(n14828), .ZN(n14830) );
  OAI211_X1 U16523 ( .C1(n14848), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        P2_U3224) );
  OAI21_X1 U16524 ( .B1(n14835), .B2(n14834), .A(n14833), .ZN(n14841) );
  NOR2_X1 U16525 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7900), .ZN(n14836) );
  AOI21_X1 U16526 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14839) );
  OAI21_X1 U16527 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n14842) );
  INV_X1 U16528 ( .A(n14842), .ZN(n14846) );
  OAI211_X1 U16529 ( .C1(n14844), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14857), 
        .B(n14843), .ZN(n14845) );
  OAI211_X1 U16530 ( .C1(n14848), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        P2_U3228) );
  INV_X1 U16531 ( .A(n14849), .ZN(n14854) );
  AOI211_X1 U16532 ( .C1(n14852), .C2(n15235), .A(n14851), .B(n14850), .ZN(
        n14853) );
  AOI211_X1 U16533 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14855), .A(n14854), 
        .B(n14853), .ZN(n14860) );
  OAI211_X1 U16534 ( .C1(n14858), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14857), 
        .B(n14856), .ZN(n14859) );
  OAI211_X1 U16535 ( .C1(n14862), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        P2_U3229) );
  INV_X1 U16536 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15431) );
  NOR2_X1 U16537 ( .A1(n14888), .A2(n15431), .ZN(P2_U3266) );
  INV_X1 U16538 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16539 ( .A1(n14888), .A2(n15347), .ZN(P2_U3267) );
  INV_X1 U16540 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n14864) );
  NOR2_X1 U16541 ( .A1(n14888), .A2(n14864), .ZN(P2_U3268) );
  INV_X1 U16542 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n14865) );
  NOR2_X1 U16543 ( .A1(n14884), .A2(n14865), .ZN(P2_U3269) );
  INV_X1 U16544 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n14866) );
  NOR2_X1 U16545 ( .A1(n14884), .A2(n14866), .ZN(P2_U3270) );
  INV_X1 U16546 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n14867) );
  NOR2_X1 U16547 ( .A1(n14884), .A2(n14867), .ZN(P2_U3271) );
  INV_X1 U16548 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n14868) );
  NOR2_X1 U16549 ( .A1(n14884), .A2(n14868), .ZN(P2_U3272) );
  INV_X1 U16550 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n14869) );
  NOR2_X1 U16551 ( .A1(n14884), .A2(n14869), .ZN(P2_U3273) );
  INV_X1 U16552 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n14870) );
  NOR2_X1 U16553 ( .A1(n14884), .A2(n14870), .ZN(P2_U3274) );
  INV_X1 U16554 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n14871) );
  NOR2_X1 U16555 ( .A1(n14884), .A2(n14871), .ZN(P2_U3275) );
  INV_X1 U16556 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n14872) );
  NOR2_X1 U16557 ( .A1(n14884), .A2(n14872), .ZN(P2_U3276) );
  INV_X1 U16558 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n14873) );
  NOR2_X1 U16559 ( .A1(n14884), .A2(n14873), .ZN(P2_U3277) );
  INV_X1 U16560 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U16561 ( .A1(n14888), .A2(n15362), .ZN(P2_U3278) );
  INV_X1 U16562 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n14874) );
  NOR2_X1 U16563 ( .A1(n14888), .A2(n14874), .ZN(P2_U3279) );
  INV_X1 U16564 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14875) );
  NOR2_X1 U16565 ( .A1(n14888), .A2(n14875), .ZN(P2_U3280) );
  INV_X1 U16566 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15385) );
  NOR2_X1 U16567 ( .A1(n14888), .A2(n15385), .ZN(P2_U3281) );
  INV_X1 U16568 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U16569 ( .A1(n14888), .A2(n15329), .ZN(P2_U3282) );
  INV_X1 U16570 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n14876) );
  NOR2_X1 U16571 ( .A1(n14888), .A2(n14876), .ZN(P2_U3283) );
  INV_X1 U16572 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n14877) );
  NOR2_X1 U16573 ( .A1(n14888), .A2(n14877), .ZN(P2_U3284) );
  INV_X1 U16574 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U16575 ( .A1(n14888), .A2(n14878), .ZN(P2_U3285) );
  INV_X1 U16576 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14879) );
  NOR2_X1 U16577 ( .A1(n14888), .A2(n14879), .ZN(P2_U3286) );
  INV_X1 U16578 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U16579 ( .A1(n14888), .A2(n15357), .ZN(P2_U3287) );
  INV_X1 U16580 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n14880) );
  NOR2_X1 U16581 ( .A1(n14888), .A2(n14880), .ZN(P2_U3288) );
  INV_X1 U16582 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15279) );
  NOR2_X1 U16583 ( .A1(n14888), .A2(n15279), .ZN(P2_U3289) );
  INV_X1 U16584 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n14881) );
  NOR2_X1 U16585 ( .A1(n14884), .A2(n14881), .ZN(P2_U3290) );
  INV_X1 U16586 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n14882) );
  NOR2_X1 U16587 ( .A1(n14888), .A2(n14882), .ZN(P2_U3291) );
  INV_X1 U16588 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n14883) );
  NOR2_X1 U16589 ( .A1(n14884), .A2(n14883), .ZN(P2_U3292) );
  INV_X1 U16590 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n14885) );
  NOR2_X1 U16591 ( .A1(n14888), .A2(n14885), .ZN(P2_U3293) );
  INV_X1 U16592 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14886) );
  NOR2_X1 U16593 ( .A1(n14888), .A2(n14886), .ZN(P2_U3294) );
  INV_X1 U16594 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14887) );
  NOR2_X1 U16595 ( .A1(n14888), .A2(n14887), .ZN(P2_U3295) );
  AOI22_X1 U16596 ( .A1(n14891), .A2(n14890), .B1(n14889), .B2(n14893), .ZN(
        P2_U3416) );
  AOI21_X1 U16597 ( .B1(n14893), .B2(n15401), .A(n14892), .ZN(P2_U3417) );
  INV_X1 U16598 ( .A(n14894), .ZN(n14895) );
  OAI21_X1 U16599 ( .B1(n6561), .B2(n14902), .A(n14895), .ZN(n14898) );
  INV_X1 U16600 ( .A(n14896), .ZN(n14897) );
  AOI211_X1 U16601 ( .C1(n14899), .C2(n14905), .A(n14898), .B(n14897), .ZN(
        n14926) );
  INV_X1 U16602 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U16603 ( .A1(n14908), .A2(n14926), .B1(n14900), .B2(n14924), .ZN(
        P2_U3433) );
  OAI21_X1 U16604 ( .B1(n6938), .B2(n14902), .A(n14901), .ZN(n14904) );
  AOI211_X1 U16605 ( .C1(n14906), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14927) );
  INV_X1 U16606 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16607 ( .A1(n14908), .A2(n14927), .B1(n14907), .B2(n14924), .ZN(
        P2_U3445) );
  AOI21_X1 U16608 ( .B1(n14918), .B2(n14910), .A(n14909), .ZN(n14911) );
  OAI211_X1 U16609 ( .C1(n8756), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        n14914) );
  INV_X1 U16610 ( .A(n14914), .ZN(n14928) );
  INV_X1 U16611 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U16612 ( .A1(n14908), .A2(n14928), .B1(n14915), .B2(n14924), .ZN(
        P2_U3448) );
  AOI21_X1 U16613 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14919) );
  OAI211_X1 U16614 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14923) );
  INV_X1 U16615 ( .A(n14923), .ZN(n14930) );
  INV_X1 U16616 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16617 ( .A1(n14908), .A2(n14930), .B1(n14925), .B2(n14924), .ZN(
        P2_U3451) );
  AOI22_X1 U16618 ( .A1(n14931), .A2(n14926), .B1(n7631), .B2(n14929), .ZN(
        P2_U3500) );
  AOI22_X1 U16619 ( .A1(n14931), .A2(n14927), .B1(n9948), .B2(n14929), .ZN(
        P2_U3504) );
  AOI22_X1 U16620 ( .A1(n14931), .A2(n14928), .B1(n7749), .B2(n14929), .ZN(
        P2_U3505) );
  AOI22_X1 U16621 ( .A1(n14931), .A2(n14930), .B1(n7770), .B2(n14929), .ZN(
        P2_U3506) );
  NOR2_X1 U16622 ( .A1(P3_U3897), .A2(n14978), .ZN(P3_U3150) );
  NAND2_X1 U16623 ( .A1(n15104), .A2(n14932), .ZN(n14933) );
  OAI21_X1 U16624 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n14936) );
  AOI21_X1 U16625 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14939) );
  OAI21_X1 U16626 ( .B1(n14940), .B2(n14947), .A(n14939), .ZN(P3_U3172) );
  NAND3_X1 U16627 ( .A1(n15023), .A2(n15015), .A3(n15017), .ZN(n14946) );
  MUX2_X1 U16628 ( .A(n14942), .B(n10366), .S(n6550), .Z(n14944) );
  OAI21_X1 U16629 ( .B1(P3_IR_REG_0__SCAN_IN), .B2(n14944), .A(n14943), .ZN(
        n14945) );
  NAND2_X1 U16630 ( .A1(n14946), .A2(n14945), .ZN(n14951) );
  OAI22_X1 U16631 ( .A1(n15007), .A2(n14948), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14947), .ZN(n14949) );
  INV_X1 U16632 ( .A(n14949), .ZN(n14950) );
  OAI211_X1 U16633 ( .C1(n14952), .C2(n15008), .A(n14951), .B(n14950), .ZN(
        P3_U3182) );
  XNOR2_X1 U16634 ( .A(n14954), .B(n14953), .ZN(n14966) );
  AOI21_X1 U16635 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14958) );
  NOR2_X1 U16636 ( .A1(n14958), .A2(n15023), .ZN(n14965) );
  AOI21_X1 U16637 ( .B1(n14961), .B2(n14960), .A(n14959), .ZN(n14963) );
  OAI22_X1 U16638 ( .A1(n15015), .A2(n14963), .B1(n15007), .B2(n14962), .ZN(
        n14964) );
  AOI211_X1 U16639 ( .C1(n14966), .C2(n14999), .A(n14965), .B(n14964), .ZN(
        n14968) );
  OAI211_X1 U16640 ( .C1(n14969), .C2(n15008), .A(n14968), .B(n14967), .ZN(
        P3_U3188) );
  AOI21_X1 U16641 ( .B1(n9261), .B2(n14971), .A(n14970), .ZN(n14975) );
  AOI21_X1 U16642 ( .B1(n9265), .B2(n14973), .A(n14972), .ZN(n14974) );
  OAI22_X1 U16643 ( .A1(n14975), .A2(n15015), .B1(n14974), .B2(n15023), .ZN(
        n14976) );
  AOI211_X1 U16644 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14978), .A(n14977), .B(
        n14976), .ZN(n14985) );
  XNOR2_X1 U16645 ( .A(n14980), .B(n14979), .ZN(n14983) );
  AOI22_X1 U16646 ( .A1(n14983), .A2(n14999), .B1(n14982), .B2(n14981), .ZN(
        n14984) );
  NAND2_X1 U16647 ( .A1(n14985), .A2(n14984), .ZN(P3_U3189) );
  XNOR2_X1 U16648 ( .A(n14987), .B(n14986), .ZN(n15000) );
  NAND2_X1 U16649 ( .A1(n14989), .A2(n14988), .ZN(n14990) );
  AOI21_X1 U16650 ( .B1(n14991), .B2(n14990), .A(n15015), .ZN(n14998) );
  INV_X1 U16651 ( .A(n14992), .ZN(n14993) );
  AOI21_X1 U16652 ( .B1(n6695), .B2(n14994), .A(n14993), .ZN(n14996) );
  OAI22_X1 U16653 ( .A1(n14996), .A2(n15023), .B1(n14995), .B2(n15007), .ZN(
        n14997) );
  AOI211_X1 U16654 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15002) );
  OAI211_X1 U16655 ( .C1(n15003), .C2(n15008), .A(n15002), .B(n15001), .ZN(
        P3_U3190) );
  AOI21_X1 U16656 ( .B1(n9368), .B2(n15005), .A(n15004), .ZN(n15024) );
  OAI22_X1 U16657 ( .A1(n15009), .A2(n15008), .B1(n15007), .B2(n15006), .ZN(
        n15020) );
  AOI21_X1 U16658 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(n15018) );
  AOI21_X1 U16659 ( .B1(n9365), .B2(n15014), .A(n15013), .ZN(n15016) );
  OAI22_X1 U16660 ( .A1(n15018), .A2(n15017), .B1(n15016), .B2(n15015), .ZN(
        n15019) );
  NOR3_X1 U16661 ( .A1(n15021), .A2(n15020), .A3(n15019), .ZN(n15022) );
  OAI21_X1 U16662 ( .B1(n15024), .B2(n15023), .A(n15022), .ZN(P3_U3195) );
  INV_X1 U16663 ( .A(n15025), .ZN(n15118) );
  XNOR2_X1 U16664 ( .A(n15026), .B(n15027), .ZN(n15167) );
  XNOR2_X1 U16665 ( .A(n15028), .B(n15027), .ZN(n15032) );
  OAI22_X1 U16666 ( .A1(n15063), .A2(n15107), .B1(n15029), .B2(n15105), .ZN(
        n15030) );
  AOI21_X1 U16667 ( .B1(n15167), .B2(n15115), .A(n15030), .ZN(n15031) );
  OAI21_X1 U16668 ( .B1(n15032), .B2(n15110), .A(n15031), .ZN(n15165) );
  AOI21_X1 U16669 ( .B1(n15118), .B2(n15167), .A(n15165), .ZN(n15037) );
  NOR2_X1 U16670 ( .A1(n15033), .A2(n15098), .ZN(n15166) );
  INV_X1 U16671 ( .A(n15034), .ZN(n15035) );
  AOI22_X1 U16672 ( .A1(n15093), .A2(n15166), .B1(n15125), .B2(n15035), .ZN(
        n15036) );
  OAI221_X1 U16673 ( .B1(n15038), .B2(n15037), .C1(n15129), .C2(n10859), .A(
        n15036), .ZN(P3_U3223) );
  OAI211_X1 U16674 ( .C1(n15042), .C2(n15041), .A(n15040), .B(n15039), .ZN(
        n15048) );
  AOI22_X1 U16675 ( .A1(n15046), .A2(n15045), .B1(n15044), .B2(n15043), .ZN(
        n15047) );
  AND2_X1 U16676 ( .A1(n15048), .A2(n15047), .ZN(n15159) );
  AOI22_X1 U16677 ( .A1(n15038), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n15125), 
        .B2(n15049), .ZN(n15054) );
  XNOR2_X1 U16678 ( .A(n15051), .B(n15050), .ZN(n15163) );
  NOR2_X1 U16679 ( .A1(n15052), .A2(n15098), .ZN(n15161) );
  AOI22_X1 U16680 ( .A1(n15163), .A2(n15079), .B1(n15093), .B2(n15161), .ZN(
        n15053) );
  OAI211_X1 U16681 ( .C1(n15038), .C2(n15159), .A(n15054), .B(n15053), .ZN(
        P3_U3224) );
  XNOR2_X1 U16682 ( .A(n15055), .B(n15061), .ZN(n15157) );
  NAND2_X1 U16683 ( .A1(n15057), .A2(n15056), .ZN(n15059) );
  NAND2_X1 U16684 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  AOI21_X1 U16685 ( .B1(n15061), .B2(n15060), .A(n6686), .ZN(n15062) );
  OAI222_X1 U16686 ( .A1(n15105), .A2(n15063), .B1(n15107), .B2(n15072), .C1(
        n15110), .C2(n15062), .ZN(n15155) );
  AOI21_X1 U16687 ( .B1(n15064), .B2(n15157), .A(n15155), .ZN(n15070) );
  AND2_X1 U16688 ( .A1(n15066), .A2(n15065), .ZN(n15156) );
  INV_X1 U16689 ( .A(n15067), .ZN(n15068) );
  AOI22_X1 U16690 ( .A1(n15093), .A2(n15156), .B1(n15068), .B2(n15125), .ZN(
        n15069) );
  OAI221_X1 U16691 ( .B1(n15038), .B2(n15070), .C1(n15129), .C2(n10817), .A(
        n15069), .ZN(P3_U3225) );
  AOI21_X1 U16692 ( .B1(n15071), .B2(n15076), .A(n15110), .ZN(n15074) );
  OAI22_X1 U16693 ( .A1(n15086), .A2(n15107), .B1(n15072), .B2(n15105), .ZN(
        n15073) );
  AOI21_X1 U16694 ( .B1(n15074), .B2(n11282), .A(n15073), .ZN(n15147) );
  AOI22_X1 U16695 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n15038), .B1(n15125), 
        .B2(n15075), .ZN(n15081) );
  XNOR2_X1 U16696 ( .A(n15076), .B(n6783), .ZN(n15150) );
  NOR2_X1 U16697 ( .A1(n15078), .A2(n15098), .ZN(n15149) );
  AOI22_X1 U16698 ( .A1(n15150), .A2(n15079), .B1(n15093), .B2(n15149), .ZN(
        n15080) );
  OAI211_X1 U16699 ( .C1(n15038), .C2(n15147), .A(n15081), .B(n15080), .ZN(
        P3_U3227) );
  XNOR2_X1 U16700 ( .A(n15082), .B(n15083), .ZN(n15141) );
  XNOR2_X1 U16701 ( .A(n15085), .B(n15084), .ZN(n15089) );
  OAI22_X1 U16702 ( .A1(n15106), .A2(n15107), .B1(n15086), .B2(n15105), .ZN(
        n15087) );
  AOI21_X1 U16703 ( .B1(n15141), .B2(n15115), .A(n15087), .ZN(n15088) );
  OAI21_X1 U16704 ( .B1(n15110), .B2(n15089), .A(n15088), .ZN(n15139) );
  AOI21_X1 U16705 ( .B1(n15118), .B2(n15141), .A(n15139), .ZN(n15095) );
  NOR2_X1 U16706 ( .A1(n15090), .A2(n15098), .ZN(n15140) );
  INV_X1 U16707 ( .A(n15091), .ZN(n15092) );
  AOI22_X1 U16708 ( .A1(n15093), .A2(n15140), .B1(n15125), .B2(n15092), .ZN(
        n15094) );
  OAI221_X1 U16709 ( .B1(n15038), .B2(n15095), .C1(n15129), .C2(n10361), .A(
        n15094), .ZN(P3_U3229) );
  OAI21_X1 U16710 ( .B1(n15097), .B2(n15109), .A(n15096), .ZN(n15134) );
  NOR2_X1 U16711 ( .A1(n15099), .A2(n15098), .ZN(n15133) );
  INV_X1 U16712 ( .A(n15133), .ZN(n15103) );
  OAI22_X1 U16713 ( .A1(n15103), .A2(n15102), .B1(n15101), .B2(n15100), .ZN(
        n15117) );
  OAI22_X1 U16714 ( .A1(n6796), .A2(n15107), .B1(n15106), .B2(n15105), .ZN(
        n15114) );
  NAND3_X1 U16715 ( .A1(n13006), .A2(n15109), .A3(n15108), .ZN(n15111) );
  AOI21_X1 U16716 ( .B1(n15112), .B2(n15111), .A(n15110), .ZN(n15113) );
  AOI211_X1 U16717 ( .C1(n15115), .C2(n15134), .A(n15114), .B(n15113), .ZN(
        n15116) );
  INV_X1 U16718 ( .A(n15116), .ZN(n15132) );
  AOI211_X1 U16719 ( .C1(n15118), .C2(n15134), .A(n15117), .B(n15132), .ZN(
        n15119) );
  AOI22_X1 U16720 ( .A1(n15038), .A2(n15120), .B1(n15119), .B2(n15129), .ZN(
        P3_U3231) );
  INV_X1 U16721 ( .A(n15121), .ZN(n15122) );
  AOI21_X1 U16722 ( .B1(n15124), .B2(n15123), .A(n15122), .ZN(n15130) );
  AOI22_X1 U16723 ( .A1(n15127), .A2(n15126), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15125), .ZN(n15128) );
  OAI221_X1 U16724 ( .B1(n15038), .B2(n15130), .C1(n15129), .C2(n10330), .A(
        n15128), .ZN(P3_U3232) );
  AOI22_X1 U16725 ( .A1(n15170), .A2(n15131), .B1(n9176), .B2(n15169), .ZN(
        P3_U3393) );
  AOI211_X1 U16726 ( .C1(n15168), .C2(n15134), .A(n15133), .B(n15132), .ZN(
        n15171) );
  AOI22_X1 U16727 ( .A1(n15170), .A2(n15171), .B1(n9194), .B2(n15169), .ZN(
        P3_U3396) );
  AOI211_X1 U16728 ( .C1(n15137), .C2(n15168), .A(n15136), .B(n15135), .ZN(
        n15172) );
  INV_X1 U16729 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15138) );
  AOI22_X1 U16730 ( .A1(n15170), .A2(n15172), .B1(n15138), .B2(n15169), .ZN(
        P3_U3399) );
  AOI211_X1 U16731 ( .C1(n15141), .C2(n15168), .A(n15140), .B(n15139), .ZN(
        n15173) );
  INV_X1 U16732 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15142) );
  AOI22_X1 U16733 ( .A1(n15170), .A2(n15173), .B1(n15142), .B2(n15169), .ZN(
        P3_U3402) );
  AOI211_X1 U16734 ( .C1(n15145), .C2(n15168), .A(n15144), .B(n15143), .ZN(
        n15174) );
  INV_X1 U16735 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15146) );
  AOI22_X1 U16736 ( .A1(n15170), .A2(n15174), .B1(n15146), .B2(n15169), .ZN(
        P3_U3405) );
  INV_X1 U16737 ( .A(n15147), .ZN(n15148) );
  AOI211_X1 U16738 ( .C1(n15150), .C2(n15162), .A(n15149), .B(n15148), .ZN(
        n15175) );
  AOI22_X1 U16739 ( .A1(n15170), .A2(n15175), .B1(n9245), .B2(n15169), .ZN(
        P3_U3408) );
  AOI211_X1 U16740 ( .C1(n15153), .C2(n15168), .A(n15152), .B(n15151), .ZN(
        n15176) );
  INV_X1 U16741 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U16742 ( .A1(n15170), .A2(n15176), .B1(n15154), .B2(n15169), .ZN(
        P3_U3411) );
  AOI211_X1 U16743 ( .C1(n15162), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        n15177) );
  INV_X1 U16744 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15158) );
  AOI22_X1 U16745 ( .A1(n15170), .A2(n15177), .B1(n15158), .B2(n15169), .ZN(
        P3_U3414) );
  INV_X1 U16746 ( .A(n15159), .ZN(n15160) );
  AOI211_X1 U16747 ( .C1(n15163), .C2(n15162), .A(n15161), .B(n15160), .ZN(
        n15178) );
  INV_X1 U16748 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15164) );
  AOI22_X1 U16749 ( .A1(n15170), .A2(n15178), .B1(n15164), .B2(n15169), .ZN(
        P3_U3417) );
  AOI211_X1 U16750 ( .C1(n15168), .C2(n15167), .A(n15166), .B(n15165), .ZN(
        n15180) );
  INV_X1 U16751 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U16752 ( .A1(n15170), .A2(n15180), .B1(n15391), .B2(n15169), .ZN(
        P3_U3420) );
  AOI22_X1 U16753 ( .A1(n15181), .A2(n15171), .B1(n10368), .B2(n15179), .ZN(
        P3_U3461) );
  AOI22_X1 U16754 ( .A1(n15181), .A2(n15172), .B1(n10340), .B2(n15179), .ZN(
        P3_U3462) );
  AOI22_X1 U16755 ( .A1(n15181), .A2(n15173), .B1(n10372), .B2(n15179), .ZN(
        P3_U3463) );
  AOI22_X1 U16756 ( .A1(n15181), .A2(n15174), .B1(n9229), .B2(n15179), .ZN(
        P3_U3464) );
  AOI22_X1 U16757 ( .A1(n15181), .A2(n15175), .B1(n9244), .B2(n15179), .ZN(
        P3_U3465) );
  AOI22_X1 U16758 ( .A1(n15181), .A2(n15176), .B1(n9261), .B2(n15179), .ZN(
        P3_U3466) );
  AOI22_X1 U16759 ( .A1(n15181), .A2(n15177), .B1(n10795), .B2(n15179), .ZN(
        P3_U3467) );
  AOI22_X1 U16760 ( .A1(n15181), .A2(n15178), .B1(n15236), .B2(n15179), .ZN(
        P3_U3468) );
  AOI22_X1 U16761 ( .A1(n15181), .A2(n15180), .B1(n10858), .B2(n15179), .ZN(
        P3_U3469) );
  NOR4_X1 U16762 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .A3(P2_REG3_REG_10__SCAN_IN), .A4(P3_REG0_REG_31__SCAN_IN), .ZN(n15191) );
  NOR4_X1 U16763 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P2_D_REG_1__SCAN_IN), 
        .A3(P3_REG1_REG_31__SCAN_IN), .A4(P3_DATAO_REG_27__SCAN_IN), .ZN(
        n15190) );
  NAND4_X1 U16764 ( .A1(SI_13_), .A2(P2_REG3_REG_14__SCAN_IN), .A3(
        P2_REG2_REG_4__SCAN_IN), .A4(P2_REG0_REG_3__SCAN_IN), .ZN(n15188) );
  NAND4_X1 U16765 ( .A1(SI_10_), .A2(SI_0_), .A3(P2_D_REG_16__SCAN_IN), .A4(
        P2_REG0_REG_8__SCAN_IN), .ZN(n15187) );
  NOR4_X1 U16766 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_REG3_REG_6__SCAN_IN), 
        .A3(P3_REG1_REG_9__SCAN_IN), .A4(P3_REG0_REG_0__SCAN_IN), .ZN(n15185)
         );
  NOR4_X1 U16767 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P2_DATAO_REG_4__SCAN_IN), 
        .A3(P3_REG0_REG_10__SCAN_IN), .A4(P3_REG0_REG_25__SCAN_IN), .ZN(n15184) );
  NOR4_X1 U16768 ( .A1(SI_16_), .A2(SI_15_), .A3(P2_IR_REG_13__SCAN_IN), .A4(
        P2_REG2_REG_3__SCAN_IN), .ZN(n15183) );
  NOR4_X1 U16769 ( .A1(SI_3_), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_REG1_REG_19__SCAN_IN), .ZN(n15182) );
  NAND4_X1 U16770 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15186) );
  NOR3_X1 U16771 ( .A1(n15188), .A2(n15187), .A3(n15186), .ZN(n15189) );
  NAND3_X1 U16772 ( .A1(n15191), .A2(n15190), .A3(n15189), .ZN(n15230) );
  NOR4_X1 U16773 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(P1_DATAO_REG_24__SCAN_IN), .A3(P2_DATAO_REG_22__SCAN_IN), .A4(P1_DATAO_REG_29__SCAN_IN), .ZN(n15195) );
  NOR4_X1 U16774 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG2_REG_26__SCAN_IN), 
        .A3(P2_REG1_REG_18__SCAN_IN), .A4(P2_REG2_REG_14__SCAN_IN), .ZN(n15194) );
  NOR4_X1 U16775 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(SI_22_), .A3(
        P2_REG2_REG_13__SCAN_IN), .A4(P2_REG3_REG_1__SCAN_IN), .ZN(n15193) );
  NOR4_X1 U16776 ( .A1(P3_REG3_REG_26__SCAN_IN), .A2(P3_REG0_REG_24__SCAN_IN), 
        .A3(P3_REG0_REG_15__SCAN_IN), .A4(P1_DATAO_REG_31__SCAN_IN), .ZN(
        n15192) );
  NAND4_X1 U16777 ( .A1(n15195), .A2(n15194), .A3(n15193), .A4(n15192), .ZN(
        n15229) );
  NOR4_X1 U16778 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n15199) );
  NOR4_X1 U16779 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(P2_REG3_REG_2__SCAN_IN), 
        .A3(P1_REG3_REG_25__SCAN_IN), .A4(P1_REG3_REG_23__SCAN_IN), .ZN(n15198) );
  NOR4_X1 U16780 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(P1_REG3_REG_24__SCAN_IN), .A4(P1_REG2_REG_11__SCAN_IN), .ZN(n15197) );
  NOR4_X1 U16781 ( .A1(SI_14_), .A2(P1_REG3_REG_5__SCAN_IN), .A3(
        P1_REG1_REG_17__SCAN_IN), .A4(P1_REG2_REG_9__SCAN_IN), .ZN(n15196) );
  NAND4_X1 U16782 ( .A1(n15199), .A2(n15198), .A3(n15197), .A4(n15196), .ZN(
        n15228) );
  NAND4_X1 U16783 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n15203) );
  NAND4_X1 U16784 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), 
        .A3(P1_REG1_REG_28__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n15202) );
  NAND4_X1 U16785 ( .A1(SI_18_), .A2(P1_IR_REG_30__SCAN_IN), .A3(
        P1_REG3_REG_20__SCAN_IN), .A4(P2_ADDR_REG_15__SCAN_IN), .ZN(n15201) );
  NAND4_X1 U16786 ( .A1(SI_25_), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_REG1_REG_18__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n15200) );
  NOR4_X1 U16787 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        n15226) );
  NAND4_X1 U16788 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(P2_ADDR_REG_5__SCAN_IN), .A4(n15301), .ZN(n15204) );
  NOR2_X1 U16789 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n15204), .ZN(n15214) );
  INV_X1 U16790 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n15205) );
  NAND2_X1 U16791 ( .A1(n15206), .A2(n15205), .ZN(n15207) );
  NOR2_X1 U16792 ( .A1(n15208), .A2(n15207), .ZN(n15212) );
  NAND3_X1 U16793 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), 
        .A3(n10127), .ZN(n15209) );
  NOR2_X1 U16794 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  AND4_X1 U16795 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        n15225) );
  NAND4_X1 U16796 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P2_DATAO_REG_9__SCAN_IN), 
        .A3(P2_DATAO_REG_7__SCAN_IN), .A4(P3_REG0_REG_6__SCAN_IN), .ZN(n15218)
         );
  NAND4_X1 U16797 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P2_IR_REG_16__SCAN_IN), .A4(P2_D_REG_0__SCAN_IN), .ZN(n15217) );
  NAND4_X1 U16798 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_REG1_REG_26__SCAN_IN), .ZN(n15216) );
  NAND4_X1 U16799 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(
        P2_DATAO_REG_10__SCAN_IN), .A3(P3_REG2_REG_9__SCAN_IN), .A4(
        P3_REG1_REG_5__SCAN_IN), .ZN(n15215) );
  NOR4_X1 U16800 ( .A1(n15218), .A2(n15217), .A3(n15216), .A4(n15215), .ZN(
        n15224) );
  NAND4_X1 U16801 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .A3(
        P2_DATAO_REG_19__SCAN_IN), .A4(SI_28_), .ZN(n15222) );
  NAND4_X1 U16802 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_REG0_REG_18__SCAN_IN), 
        .A3(P2_REG2_REG_15__SCAN_IN), .A4(P1_REG3_REG_17__SCAN_IN), .ZN(n15221) );
  NAND4_X1 U16803 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(SI_17_), .A3(
        P2_REG3_REG_18__SCAN_IN), .A4(P1_REG3_REG_18__SCAN_IN), .ZN(n15220) );
  NAND4_X1 U16804 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(SI_20_), .A3(
        P1_IR_REG_15__SCAN_IN), .A4(P3_ADDR_REG_16__SCAN_IN), .ZN(n15219) );
  NOR4_X1 U16805 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15223) );
  NAND4_X1 U16806 ( .A1(n15226), .A2(n15225), .A3(n15224), .A4(n15223), .ZN(
        n15227) );
  NOR4_X1 U16807 ( .A1(n15230), .A2(n15229), .A3(n15228), .A4(n15227), .ZN(
        n15470) );
  AOI22_X1 U16808 ( .A1(n15233), .A2(keyinput7), .B1(n15232), .B2(keyinput87), 
        .ZN(n15231) );
  OAI221_X1 U16809 ( .B1(n15233), .B2(keyinput7), .C1(n15232), .C2(keyinput87), 
        .A(n15231), .ZN(n15243) );
  AOI22_X1 U16810 ( .A1(n15236), .A2(keyinput123), .B1(keyinput39), .B2(n15235), .ZN(n15234) );
  OAI221_X1 U16811 ( .B1(n15236), .B2(keyinput123), .C1(n15235), .C2(
        keyinput39), .A(n15234), .ZN(n15242) );
  XNOR2_X1 U16812 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput73), .ZN(n15240)
         );
  XNOR2_X1 U16813 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput76), .ZN(n15239)
         );
  XNOR2_X1 U16814 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput34), .ZN(n15238) );
  XNOR2_X1 U16815 ( .A(SI_22_), .B(keyinput25), .ZN(n15237) );
  NAND4_X1 U16816 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15241) );
  NOR3_X1 U16817 ( .A1(n15243), .A2(n15242), .A3(n15241), .ZN(n15287) );
  AOI22_X1 U16818 ( .A1(n15246), .A2(keyinput66), .B1(keyinput31), .B2(n15245), 
        .ZN(n15244) );
  OAI221_X1 U16819 ( .B1(n15246), .B2(keyinput66), .C1(n15245), .C2(keyinput31), .A(n15244), .ZN(n15258) );
  AOI22_X1 U16820 ( .A1(n15249), .A2(keyinput59), .B1(n15248), .B2(keyinput62), 
        .ZN(n15247) );
  OAI221_X1 U16821 ( .B1(n15249), .B2(keyinput59), .C1(n15248), .C2(keyinput62), .A(n15247), .ZN(n15257) );
  AOI22_X1 U16822 ( .A1(n15252), .A2(keyinput90), .B1(n15251), .B2(keyinput117), .ZN(n15250) );
  OAI221_X1 U16823 ( .B1(n15252), .B2(keyinput90), .C1(n15251), .C2(
        keyinput117), .A(n15250), .ZN(n15256) );
  XNOR2_X1 U16824 ( .A(P1_REG3_REG_17__SCAN_IN), .B(keyinput69), .ZN(n15254)
         );
  XNOR2_X1 U16825 ( .A(SI_3_), .B(keyinput38), .ZN(n15253) );
  NAND2_X1 U16826 ( .A1(n15254), .A2(n15253), .ZN(n15255) );
  NOR4_X1 U16827 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15286) );
  AOI22_X1 U16828 ( .A1(n15261), .A2(keyinput43), .B1(keyinput77), .B2(n15260), 
        .ZN(n15259) );
  OAI221_X1 U16829 ( .B1(n15261), .B2(keyinput43), .C1(n15260), .C2(keyinput77), .A(n15259), .ZN(n15271) );
  AOI22_X1 U16830 ( .A1(n15264), .A2(keyinput93), .B1(keyinput88), .B2(n15263), 
        .ZN(n15262) );
  OAI221_X1 U16831 ( .B1(n15264), .B2(keyinput93), .C1(n15263), .C2(keyinput88), .A(n15262), .ZN(n15270) );
  XNOR2_X1 U16832 ( .A(SI_0_), .B(keyinput44), .ZN(n15268) );
  XNOR2_X1 U16833 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput64), .ZN(n15267)
         );
  XNOR2_X1 U16834 ( .A(P3_REG2_REG_29__SCAN_IN), .B(keyinput11), .ZN(n15266)
         );
  XNOR2_X1 U16835 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput118), .ZN(n15265)
         );
  NAND4_X1 U16836 ( .A1(n15268), .A2(n15267), .A3(n15266), .A4(n15265), .ZN(
        n15269) );
  NOR3_X1 U16837 ( .A1(n15271), .A2(n15270), .A3(n15269), .ZN(n15285) );
  AOI22_X1 U16838 ( .A1(n15273), .A2(keyinput2), .B1(keyinput68), .B2(n10226), 
        .ZN(n15272) );
  OAI221_X1 U16839 ( .B1(n15273), .B2(keyinput2), .C1(n10226), .C2(keyinput68), 
        .A(n15272), .ZN(n15283) );
  AOI22_X1 U16840 ( .A1(n7900), .A2(keyinput110), .B1(keyinput55), .B2(n15275), 
        .ZN(n15274) );
  OAI221_X1 U16841 ( .B1(n7900), .B2(keyinput110), .C1(n15275), .C2(keyinput55), .A(n15274), .ZN(n15282) );
  XNOR2_X1 U16842 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput18), .ZN(n15278)
         );
  XNOR2_X1 U16843 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput13), .ZN(n15277) );
  XNOR2_X1 U16844 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput75), .ZN(n15276) );
  NAND3_X1 U16845 ( .A1(n15278), .A2(n15277), .A3(n15276), .ZN(n15281) );
  XNOR2_X1 U16846 ( .A(n15279), .B(keyinput52), .ZN(n15280) );
  NOR4_X1 U16847 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n15284) );
  NAND4_X1 U16848 ( .A1(n15287), .A2(n15286), .A3(n15285), .A4(n15284), .ZN(
        n15465) );
  AOI22_X1 U16849 ( .A1(n15289), .A2(keyinput37), .B1(keyinput121), .B2(n11066), .ZN(n15288) );
  OAI221_X1 U16850 ( .B1(n15289), .B2(keyinput37), .C1(n11066), .C2(
        keyinput121), .A(n15288), .ZN(n15299) );
  AOI22_X1 U16851 ( .A1(n15292), .A2(keyinput107), .B1(n15291), .B2(keyinput50), .ZN(n15290) );
  OAI221_X1 U16852 ( .B1(n15292), .B2(keyinput107), .C1(n15291), .C2(
        keyinput50), .A(n15290), .ZN(n15298) );
  XNOR2_X1 U16853 ( .A(SI_20_), .B(keyinput71), .ZN(n15296) );
  XNOR2_X1 U16854 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput97), .ZN(n15295) );
  XNOR2_X1 U16855 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput127), .ZN(n15294) );
  XNOR2_X1 U16856 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput89), .ZN(n15293)
         );
  NAND4_X1 U16857 ( .A1(n15296), .A2(n15295), .A3(n15294), .A4(n15293), .ZN(
        n15297) );
  NOR3_X1 U16858 ( .A1(n15299), .A2(n15298), .A3(n15297), .ZN(n15345) );
  AOI22_X1 U16859 ( .A1(n11083), .A2(keyinput101), .B1(keyinput126), .B2(
        n15301), .ZN(n15300) );
  OAI221_X1 U16860 ( .B1(n11083), .B2(keyinput101), .C1(n15301), .C2(
        keyinput126), .A(n15300), .ZN(n15314) );
  AOI22_X1 U16861 ( .A1(n15304), .A2(keyinput9), .B1(keyinput85), .B2(n15303), 
        .ZN(n15302) );
  OAI221_X1 U16862 ( .B1(n15304), .B2(keyinput9), .C1(n15303), .C2(keyinput85), 
        .A(n15302), .ZN(n15313) );
  AOI22_X1 U16863 ( .A1(n15307), .A2(keyinput29), .B1(n15306), .B2(keyinput99), 
        .ZN(n15305) );
  OAI221_X1 U16864 ( .B1(n15307), .B2(keyinput29), .C1(n15306), .C2(keyinput99), .A(n15305), .ZN(n15312) );
  AOI22_X1 U16865 ( .A1(n15310), .A2(keyinput14), .B1(n15309), .B2(keyinput78), 
        .ZN(n15308) );
  OAI221_X1 U16866 ( .B1(n15310), .B2(keyinput14), .C1(n15309), .C2(keyinput78), .A(n15308), .ZN(n15311) );
  NOR4_X1 U16867 ( .A1(n15314), .A2(n15313), .A3(n15312), .A4(n15311), .ZN(
        n15344) );
  INV_X1 U16868 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15316) );
  AOI22_X1 U16869 ( .A1(n15316), .A2(keyinput47), .B1(n9226), .B2(keyinput20), 
        .ZN(n15315) );
  OAI221_X1 U16870 ( .B1(n15316), .B2(keyinput47), .C1(n9226), .C2(keyinput20), 
        .A(n15315), .ZN(n15326) );
  AOI22_X1 U16871 ( .A1(n15318), .A2(keyinput108), .B1(keyinput96), .B2(n14097), .ZN(n15317) );
  OAI221_X1 U16872 ( .B1(n15318), .B2(keyinput108), .C1(n14097), .C2(
        keyinput96), .A(n15317), .ZN(n15325) );
  AOI22_X1 U16873 ( .A1(n15320), .A2(keyinput95), .B1(n7674), .B2(keyinput106), 
        .ZN(n15319) );
  OAI221_X1 U16874 ( .B1(n15320), .B2(keyinput95), .C1(n7674), .C2(keyinput106), .A(n15319), .ZN(n15324) );
  XOR2_X1 U16875 ( .A(n13848), .B(keyinput103), .Z(n15322) );
  XNOR2_X1 U16876 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput102), .ZN(n15321) );
  NAND2_X1 U16877 ( .A1(n15322), .A2(n15321), .ZN(n15323) );
  NOR4_X1 U16878 ( .A1(n15326), .A2(n15325), .A3(n15324), .A4(n15323), .ZN(
        n15343) );
  INV_X1 U16879 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U16880 ( .A1(n15329), .A2(keyinput53), .B1(keyinput104), .B2(n15328), .ZN(n15327) );
  OAI221_X1 U16881 ( .B1(n15329), .B2(keyinput53), .C1(n15328), .C2(
        keyinput104), .A(n15327), .ZN(n15341) );
  INV_X1 U16882 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U16883 ( .A1(n15332), .A2(keyinput63), .B1(n15331), .B2(keyinput41), 
        .ZN(n15330) );
  OAI221_X1 U16884 ( .B1(n15332), .B2(keyinput63), .C1(n15331), .C2(keyinput41), .A(n15330), .ZN(n15340) );
  AOI22_X1 U16885 ( .A1(n9183), .A2(keyinput10), .B1(n15334), .B2(keyinput83), 
        .ZN(n15333) );
  OAI221_X1 U16886 ( .B1(n9183), .B2(keyinput10), .C1(n15334), .C2(keyinput83), 
        .A(n15333), .ZN(n15339) );
  AOI22_X1 U16887 ( .A1(n15337), .A2(keyinput40), .B1(keyinput6), .B2(n15336), 
        .ZN(n15335) );
  OAI221_X1 U16888 ( .B1(n15337), .B2(keyinput40), .C1(n15336), .C2(keyinput6), 
        .A(n15335), .ZN(n15338) );
  NOR4_X1 U16889 ( .A1(n15341), .A2(n15340), .A3(n15339), .A4(n15338), .ZN(
        n15342) );
  NAND4_X1 U16890 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15464) );
  AOI22_X1 U16891 ( .A1(n15348), .A2(keyinput112), .B1(n15347), .B2(
        keyinput109), .ZN(n15346) );
  OAI221_X1 U16892 ( .B1(n15348), .B2(keyinput112), .C1(n15347), .C2(
        keyinput109), .A(n15346), .ZN(n15355) );
  AOI22_X1 U16893 ( .A1(n10761), .A2(keyinput120), .B1(n15350), .B2(keyinput98), .ZN(n15349) );
  OAI221_X1 U16894 ( .B1(n10761), .B2(keyinput120), .C1(n15350), .C2(
        keyinput98), .A(n15349), .ZN(n15354) );
  XNOR2_X1 U16895 ( .A(n15351), .B(keyinput105), .ZN(n15353) );
  XOR2_X1 U16896 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput86), .Z(n15352) );
  OR4_X1 U16897 ( .A1(n15355), .A2(n15354), .A3(n15353), .A4(n15352), .ZN(
        n15360) );
  XNOR2_X1 U16898 ( .A(n15356), .B(keyinput111), .ZN(n15359) );
  XNOR2_X1 U16899 ( .A(n15357), .B(keyinput60), .ZN(n15358) );
  NOR3_X1 U16900 ( .A1(n15360), .A2(n15359), .A3(n15358), .ZN(n15408) );
  AOI22_X1 U16901 ( .A1(n15363), .A2(keyinput115), .B1(n15362), .B2(keyinput42), .ZN(n15361) );
  OAI221_X1 U16902 ( .B1(n15363), .B2(keyinput115), .C1(n15362), .C2(
        keyinput42), .A(n15361), .ZN(n15369) );
  AOI22_X1 U16903 ( .A1(n15366), .A2(keyinput8), .B1(keyinput24), .B2(n15365), 
        .ZN(n15364) );
  OAI221_X1 U16904 ( .B1(n15366), .B2(keyinput8), .C1(n15365), .C2(keyinput24), 
        .A(n15364), .ZN(n15368) );
  XOR2_X1 U16905 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput45), .Z(n15367) );
  OR3_X1 U16906 ( .A1(n15369), .A2(n15368), .A3(n15367), .ZN(n15375) );
  AOI22_X1 U16907 ( .A1(n15371), .A2(keyinput80), .B1(keyinput36), .B2(n7829), 
        .ZN(n15370) );
  OAI221_X1 U16908 ( .B1(n15371), .B2(keyinput80), .C1(n7829), .C2(keyinput36), 
        .A(n15370), .ZN(n15374) );
  XNOR2_X1 U16909 ( .A(n15372), .B(keyinput91), .ZN(n15373) );
  NOR3_X1 U16910 ( .A1(n15375), .A2(n15374), .A3(n15373), .ZN(n15407) );
  AOI22_X1 U16911 ( .A1(n15377), .A2(keyinput22), .B1(n13354), .B2(keyinput1), 
        .ZN(n15376) );
  OAI221_X1 U16912 ( .B1(n15377), .B2(keyinput22), .C1(n13354), .C2(keyinput1), 
        .A(n15376), .ZN(n15381) );
  XOR2_X1 U16913 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput56), .Z(n15380) );
  XNOR2_X1 U16914 ( .A(n15378), .B(keyinput113), .ZN(n15379) );
  OR3_X1 U16915 ( .A1(n15381), .A2(n15380), .A3(n15379), .ZN(n15389) );
  AOI22_X1 U16916 ( .A1(n15383), .A2(keyinput12), .B1(n11730), .B2(keyinput100), .ZN(n15382) );
  OAI221_X1 U16917 ( .B1(n15383), .B2(keyinput12), .C1(n11730), .C2(
        keyinput100), .A(n15382), .ZN(n15388) );
  AOI22_X1 U16918 ( .A1(n15386), .A2(keyinput54), .B1(n15385), .B2(keyinput46), 
        .ZN(n15384) );
  OAI221_X1 U16919 ( .B1(n15386), .B2(keyinput54), .C1(n15385), .C2(keyinput46), .A(n15384), .ZN(n15387) );
  NOR3_X1 U16920 ( .A1(n15389), .A2(n15388), .A3(n15387), .ZN(n15406) );
  AOI22_X1 U16921 ( .A1(n15391), .A2(keyinput82), .B1(keyinput124), .B2(n7793), 
        .ZN(n15390) );
  OAI221_X1 U16922 ( .B1(n15391), .B2(keyinput82), .C1(n7793), .C2(keyinput124), .A(n15390), .ZN(n15404) );
  AOI22_X1 U16923 ( .A1(n15392), .A2(keyinput72), .B1(keyinput30), .B2(n15394), 
        .ZN(n15393) );
  OAI221_X1 U16924 ( .B1(n15392), .B2(keyinput72), .C1(n15394), .C2(keyinput30), .A(n15393), .ZN(n15399) );
  XNOR2_X1 U16925 ( .A(n15395), .B(keyinput79), .ZN(n15398) );
  XNOR2_X1 U16926 ( .A(n15396), .B(keyinput67), .ZN(n15397) );
  OR3_X1 U16927 ( .A1(n15399), .A2(n15398), .A3(n15397), .ZN(n15403) );
  AOI22_X1 U16928 ( .A1(n10127), .A2(keyinput119), .B1(n15401), .B2(keyinput70), .ZN(n15400) );
  OAI221_X1 U16929 ( .B1(n10127), .B2(keyinput119), .C1(n15401), .C2(
        keyinput70), .A(n15400), .ZN(n15402) );
  NOR3_X1 U16930 ( .A1(n15404), .A2(n15403), .A3(n15402), .ZN(n15405) );
  NAND4_X1 U16931 ( .A1(n15408), .A2(n15407), .A3(n15406), .A4(n15405), .ZN(
        n15463) );
  AOI22_X1 U16932 ( .A1(n15410), .A2(keyinput0), .B1(n13556), .B2(keyinput26), 
        .ZN(n15409) );
  OAI221_X1 U16933 ( .B1(n15410), .B2(keyinput0), .C1(n13556), .C2(keyinput26), 
        .A(n15409), .ZN(n15420) );
  INV_X1 U16934 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U16935 ( .A1(n15412), .A2(keyinput5), .B1(n8542), .B2(keyinput81), 
        .ZN(n15411) );
  OAI221_X1 U16936 ( .B1(n15412), .B2(keyinput5), .C1(n8542), .C2(keyinput81), 
        .A(n15411), .ZN(n15419) );
  XOR2_X1 U16937 ( .A(n15413), .B(keyinput49), .Z(n15417) );
  XOR2_X1 U16938 ( .A(n7278), .B(keyinput35), .Z(n15416) );
  XNOR2_X1 U16939 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput15), .ZN(n15415)
         );
  XNOR2_X1 U16940 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput28), .ZN(n15414) );
  NAND4_X1 U16941 ( .A1(n15417), .A2(n15416), .A3(n15415), .A4(n15414), .ZN(
        n15418) );
  NOR3_X1 U16942 ( .A1(n15420), .A2(n15419), .A3(n15418), .ZN(n15461) );
  AOI22_X1 U16943 ( .A1(n9245), .A2(keyinput58), .B1(keyinput116), .B2(n7947), 
        .ZN(n15421) );
  OAI221_X1 U16944 ( .B1(n9245), .B2(keyinput58), .C1(n7947), .C2(keyinput116), 
        .A(n15421), .ZN(n15429) );
  XOR2_X1 U16945 ( .A(P3_IR_REG_18__SCAN_IN), .B(keyinput4), .Z(n15428) );
  XNOR2_X1 U16946 ( .A(keyinput48), .B(n10235), .ZN(n15427) );
  XNOR2_X1 U16947 ( .A(SI_13_), .B(keyinput92), .ZN(n15425) );
  XNOR2_X1 U16948 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput94), .ZN(n15424)
         );
  XNOR2_X1 U16949 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput16), .ZN(n15423) );
  XNOR2_X1 U16950 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput23), .ZN(n15422)
         );
  NAND4_X1 U16951 ( .A1(n15425), .A2(n15424), .A3(n15423), .A4(n15422), .ZN(
        n15426) );
  NOR4_X1 U16952 ( .A1(n15429), .A2(n15428), .A3(n15427), .A4(n15426), .ZN(
        n15460) );
  AOI22_X1 U16953 ( .A1(n15432), .A2(keyinput27), .B1(n15431), .B2(keyinput51), 
        .ZN(n15430) );
  OAI221_X1 U16954 ( .B1(n15432), .B2(keyinput27), .C1(n15431), .C2(keyinput51), .A(n15430), .ZN(n15442) );
  AOI22_X1 U16955 ( .A1(n15435), .A2(keyinput122), .B1(n15434), .B2(keyinput61), .ZN(n15433) );
  OAI221_X1 U16956 ( .B1(n15435), .B2(keyinput122), .C1(n15434), .C2(
        keyinput61), .A(n15433), .ZN(n15441) );
  XOR2_X1 U16957 ( .A(n9979), .B(keyinput17), .Z(n15439) );
  XNOR2_X1 U16958 ( .A(keyinput33), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15438)
         );
  XNOR2_X1 U16959 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput57), .ZN(n15437) );
  XNOR2_X1 U16960 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput114), .ZN(n15436) );
  NAND4_X1 U16961 ( .A1(n15439), .A2(n15438), .A3(n15437), .A4(n15436), .ZN(
        n15440) );
  NOR3_X1 U16962 ( .A1(n15442), .A2(n15441), .A3(n15440), .ZN(n15459) );
  AOI22_X1 U16963 ( .A1(n15445), .A2(keyinput125), .B1(keyinput74), .B2(n15444), .ZN(n15443) );
  OAI221_X1 U16964 ( .B1(n15445), .B2(keyinput125), .C1(n15444), .C2(
        keyinput74), .A(n15443), .ZN(n15457) );
  INV_X1 U16965 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n15447) );
  AOI22_X1 U16966 ( .A1(n15448), .A2(keyinput65), .B1(n15447), .B2(keyinput84), 
        .ZN(n15446) );
  OAI221_X1 U16967 ( .B1(n15448), .B2(keyinput65), .C1(n15447), .C2(keyinput84), .A(n15446), .ZN(n15456) );
  AOI22_X1 U16968 ( .A1(n15450), .A2(keyinput3), .B1(n9229), .B2(keyinput19), 
        .ZN(n15449) );
  OAI221_X1 U16969 ( .B1(n15450), .B2(keyinput3), .C1(n9229), .C2(keyinput19), 
        .A(n15449), .ZN(n15455) );
  AOI22_X1 U16970 ( .A1(n15453), .A2(keyinput21), .B1(n15452), .B2(keyinput32), 
        .ZN(n15451) );
  OAI221_X1 U16971 ( .B1(n15453), .B2(keyinput21), .C1(n15452), .C2(keyinput32), .A(n15451), .ZN(n15454) );
  NOR4_X1 U16972 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15458) );
  NAND4_X1 U16973 ( .A1(n15461), .A2(n15460), .A3(n15459), .A4(n15458), .ZN(
        n15462) );
  NOR4_X1 U16974 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        n15468) );
  NAND2_X1 U16975 ( .A1(n15466), .A2(P3_D_REG_4__SCAN_IN), .ZN(n15467) );
  XOR2_X1 U16976 ( .A(n15468), .B(n15467), .Z(n15469) );
  XNOR2_X1 U16977 ( .A(n15470), .B(n15469), .ZN(P3_U3261) );
  XOR2_X1 U16978 ( .A(n15471), .B(n15472), .Z(SUB_1596_U59) );
  XOR2_X1 U16979 ( .A(n9979), .B(n15473), .Z(SUB_1596_U58) );
  AOI21_X1 U16980 ( .B1(n15474), .B2(n11741), .A(n15482), .ZN(SUB_1596_U53) );
  XOR2_X1 U16981 ( .A(n15476), .B(n15475), .Z(SUB_1596_U56) );
  AOI21_X1 U16982 ( .B1(n15479), .B2(n15478), .A(n15477), .ZN(n15480) );
  XOR2_X1 U16983 ( .A(n15480), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U16984 ( .A(n15481), .B(n15482), .Z(SUB_1596_U5) );
  NAND2_X1 U7633 ( .A1(n7275), .A2(n14454), .ZN(n14455) );
  NAND2_X1 U9630 ( .A1(n14458), .A2(n14459), .ZN(n14460) );
  XNOR2_X1 U10614 ( .A(n8961), .B(n8960), .ZN(n12194) );
  OAI21_X1 U9556 ( .B1(n7021), .B2(n7020), .A(n11914), .ZN(n7019) );
  NOR3_X1 U9322 ( .A1(n11968), .A2(n11964), .A3(n11963), .ZN(n11965) );
  CLKBUF_X2 U7301 ( .A(n8414), .Z(n8417) );
  CLKBUF_X1 U7309 ( .A(n11448), .Z(n12363) );
  CLKBUF_X1 U7344 ( .A(n6589), .Z(n12305) );
  CLKBUF_X1 U7365 ( .A(n9203), .Z(n6558) );
  CLKBUF_X1 U7368 ( .A(n9714), .Z(n13564) );
  CLKBUF_X1 U7378 ( .A(n12727), .Z(n6555) );
  CLKBUF_X1 U7390 ( .A(n10499), .Z(n6548) );
  XNOR2_X1 U7417 ( .A(n14460), .B(n14461), .ZN(n14502) );
  BUF_X4 U7425 ( .A(n9903), .Z(n6568) );
endmodule

