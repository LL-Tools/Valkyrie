

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040;

  BUF_X1 U2379 ( .A(n2978), .Z(n3148) );
  CLKBUF_X2 U2380 ( .A(n2516), .Z(n2555) );
  NAND2_X1 U2381 ( .A1(n2805), .A2(n2770), .ZN(n2819) );
  NAND4_X1 U2383 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n4154)
         );
  INV_X2 U2386 ( .A(n3146), .ZN(n3142) );
  NAND2_X1 U2387 ( .A1(n2879), .A2(n2878), .ZN(n2972) );
  OAI21_X1 U2388 ( .B1(n3457), .B2(n2207), .A(n2204), .ZN(n3521) );
  CLKBUF_X3 U2389 ( .A(n2472), .Z(n2143) );
  INV_X1 U2390 ( .A(IR_REG_3__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U2391 ( .A1(n2431), .A2(n2429), .ZN(n3883) );
  BUF_X1 U2392 ( .A(n2518), .Z(n2750) );
  NAND2_X1 U2393 ( .A1(n4170), .A2(n2902), .ZN(n4168) );
  INV_X1 U2394 ( .A(n4498), .ZN(n4459) );
  NOR2_X1 U2395 ( .A1(n4338), .A2(n4315), .ZN(n4316) );
  INV_X1 U2396 ( .A(n2827), .ZN(n2878) );
  INV_X2 U2397 ( .A(n4724), .ZN(n4726) );
  NOR2_X2 U2398 ( .A1(n4430), .A2(n3088), .ZN(n4409) );
  NOR2_X2 U2399 ( .A1(n2916), .A2(n4190), .ZN(n2918) );
  OAI21_X2 U2400 ( .B1(n4711), .B2(n2328), .A(n2327), .ZN(n4190) );
  OAI21_X2 U2401 ( .B1(n3941), .B2(n2410), .A(n2220), .ZN(n3906) );
  OAI21_X2 U2402 ( .B1(n3771), .B2(n2212), .A(n2209), .ZN(n3941) );
  XNOR2_X2 U2403 ( .A(n2891), .B(n4689), .ZN(n3350) );
  NAND2_X1 U2404 ( .A1(n2875), .A2(n2874), .ZN(n2368) );
  NAND2_X1 U2405 ( .A1(n2284), .A2(n2285), .ZN(n4440) );
  NAND2_X1 U2406 ( .A1(n2428), .A2(n2427), .ZN(n3457) );
  NAND2_X2 U2407 ( .A1(n2828), .A2(n4492), .ZN(n4724) );
  INV_X1 U2408 ( .A(n3437), .ZN(n3571) );
  INV_X2 U2409 ( .A(n2988), .ZN(n2998) );
  OR2_X1 U2410 ( .A1(n2978), .A2(n4611), .ZN(n3008) );
  AND2_X1 U2411 ( .A1(n2478), .A2(n2477), .ZN(n2178) );
  CLKBUF_X3 U2412 ( .A(n2541), .Z(n3837) );
  AND2_X1 U2413 ( .A1(n2298), .A2(n2299), .ZN(n2300) );
  BUF_X2 U2414 ( .A(n2544), .Z(n3833) );
  AND2_X1 U2415 ( .A1(n2476), .A2(n3271), .ZN(n2545) );
  AND2_X2 U2416 ( .A1(n2476), .A2(n2475), .ZN(n2544) );
  NAND2_X1 U2417 ( .A1(n2490), .A2(n2452), .ZN(n2513) );
  OAI21_X1 U2418 ( .B1(n2832), .B2(n2831), .A(n4724), .ZN(n2885) );
  OR2_X1 U2419 ( .A1(n3226), .A2(n4754), .ZN(n3223) );
  OR2_X1 U2420 ( .A1(n3226), .A2(n4749), .ZN(n3229) );
  NAND2_X1 U2421 ( .A1(n4440), .A2(n4103), .ZN(n4425) );
  OAI21_X1 U2422 ( .B1(n4362), .B2(n2868), .A(n2867), .ZN(n4349) );
  NAND2_X1 U2423 ( .A1(n2346), .A2(n2345), .ZN(n4362) );
  XNOR2_X1 U2424 ( .A(n2907), .B(n4683), .ZN(n4180) );
  CLKBUF_X1 U2425 ( .A(n4455), .Z(n2140) );
  AND2_X1 U2426 ( .A1(n4316), .A2(n2195), .ZN(n4241) );
  NAND2_X1 U2427 ( .A1(n2275), .A2(n2273), .ZN(n3668) );
  NAND2_X1 U2428 ( .A1(n3755), .A2(n2858), .ZN(n4463) );
  NAND2_X1 U2429 ( .A1(n2307), .A2(n2306), .ZN(n4170) );
  AOI21_X1 U2430 ( .B1(n2420), .B2(n2422), .A(n2170), .ZN(n2417) );
  OAI21_X1 U2431 ( .B1(n2424), .B2(n2422), .A(n3561), .ZN(n2421) );
  AND2_X1 U2432 ( .A1(n2205), .A2(n3017), .ZN(n2204) );
  AOI21_X1 U2433 ( .B1(n2277), .B2(n2280), .A(n2274), .ZN(n2273) );
  AND2_X1 U2434 ( .A1(n3009), .A2(n3003), .ZN(n2427) );
  AND2_X1 U2435 ( .A1(n2405), .A2(n2278), .ZN(n2277) );
  OAI21_X1 U2436 ( .B1(n2351), .B2(n2352), .A(n2171), .ZN(n2350) );
  NOR2_X1 U2437 ( .A1(n2283), .A2(n2282), .ZN(n2281) );
  NAND2_X2 U2438 ( .A1(n4751), .A2(n4611), .ZN(n4674) );
  AND2_X1 U2439 ( .A1(n4088), .A2(n2163), .ZN(n2352) );
  NAND2_X2 U2440 ( .A1(n2178), .A2(n2300), .ZN(n4153) );
  INV_X1 U2441 ( .A(n3043), .ZN(n3774) );
  INV_X1 U2442 ( .A(n3596), .ZN(n3599) );
  NAND4_X2 U2443 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), .ZN(n3596)
         );
  AND4_X1 U2444 ( .A1(n2562), .A2(n2561), .A3(n2560), .A4(n2559), .ZN(n3685)
         );
  OR2_X1 U2445 ( .A1(n2608), .A2(n2607), .ZN(n4597) );
  OR2_X1 U2446 ( .A1(n2331), .A2(n2333), .ZN(n3525) );
  OAI21_X2 U2447 ( .B1(n2555), .B2(n2540), .A(n2539), .ZN(n3592) );
  AND2_X4 U2448 ( .A1(n3233), .A2(n4729), .ZN(U4043) );
  AND4_X2 U2449 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n3573)
         );
  AND4_X1 U2450 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n3732)
         );
  NAND2_X1 U2451 ( .A1(n2555), .A2(n2538), .ZN(n2539) );
  AND2_X2 U2452 ( .A1(n2972), .A2(n3174), .ZN(n3146) );
  INV_X1 U2453 ( .A(n2972), .ZN(n2970) );
  INV_X1 U2454 ( .A(n3432), .ZN(n3364) );
  BUF_X4 U2455 ( .A(n2555), .Z(n3832) );
  INV_X1 U2456 ( .A(n3005), .ZN(n3553) );
  AND2_X2 U2457 ( .A1(n3367), .A2(n2879), .ZN(n4611) );
  NAND2_X1 U2458 ( .A1(n2208), .A2(n4679), .ZN(n2971) );
  AND2_X1 U2459 ( .A1(n2975), .A2(n2827), .ZN(n3367) );
  NAND2_X1 U2460 ( .A1(n3294), .A2(n2890), .ZN(n2891) );
  CLKBUF_X3 U2461 ( .A(n2545), .Z(n3834) );
  NOR2_X1 U2462 ( .A1(n2819), .A2(n2820), .ZN(n2208) );
  AND2_X1 U2463 ( .A1(n2759), .A2(n2655), .ZN(n4681) );
  NAND2_X1 U2464 ( .A1(n3295), .A2(REG1_REG_3__SCAN_IN), .ZN(n3294) );
  XNOR2_X1 U2465 ( .A(n2800), .B(IR_REG_25__SCAN_IN), .ZN(n4679) );
  MUX2_X1 U2466 ( .A(IR_REG_31__SCAN_IN), .B(n2763), .S(IR_REG_21__SCAN_IN), 
        .Z(n2766) );
  MUX2_X1 U2467 ( .A(IR_REG_31__SCAN_IN), .B(n2804), .S(IR_REG_26__SCAN_IN), 
        .Z(n2805) );
  XNOR2_X1 U2468 ( .A(n2767), .B(n2794), .ZN(n2975) );
  NAND2_X1 U2469 ( .A1(n2799), .A2(IR_REG_31__SCAN_IN), .ZN(n2800) );
  AND2_X1 U2470 ( .A1(n2799), .A2(n2793), .ZN(n2798) );
  OR2_X1 U2471 ( .A1(n2795), .A2(n2651), .ZN(n2767) );
  NAND2_X1 U2472 ( .A1(n2773), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  NAND2_X2 U2473 ( .A1(n2494), .A2(n2493), .ZN(n3329) );
  INV_X1 U2474 ( .A(n2513), .ZN(n2453) );
  AND3_X1 U2475 ( .A1(n2762), .A2(n2438), .A3(n2164), .ZN(n2471) );
  AND4_X1 U2476 ( .A1(n2459), .A2(n2458), .A3(n2457), .A4(n2456), .ZN(n2762)
         );
  NOR2_X1 U2477 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2460)
         );
  INV_X1 U2478 ( .A(IR_REG_23__SCAN_IN), .ZN(n2822) );
  INV_X1 U2479 ( .A(IR_REG_22__SCAN_IN), .ZN(n2794) );
  INV_X1 U2480 ( .A(IR_REG_27__SCAN_IN), .ZN(n2470) );
  INV_X1 U2481 ( .A(IR_REG_2__SCAN_IN), .ZN(n2452) );
  NOR2_X2 U2482 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2490)
         );
  NOR2_X2 U2483 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n4784)
         );
  INV_X1 U2484 ( .A(IR_REG_21__SCAN_IN), .ZN(n2764) );
  NOR2_X1 U2485 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2456)
         );
  NOR2_X1 U2486 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2457)
         );
  NOR2_X1 U2487 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2458)
         );
  NOR2_X1 U2488 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2459)
         );
  OR2_X1 U2489 ( .A1(n4623), .A2(n4674), .ZN(n2138) );
  NAND2_X1 U2490 ( .A1(n2138), .A2(n4622), .ZN(U3513) );
  AOI22_X1 U2491 ( .A1(n4313), .A2(n2870), .B1(n4315), .B2(n4293), .ZN(n2139)
         );
  INV_X1 U2492 ( .A(n2476), .ZN(n2141) );
  AOI22_X1 U2493 ( .A1(n4313), .A2(n2870), .B1(n4315), .B2(n4293), .ZN(n4286)
         );
  AOI21_X1 U2494 ( .B1(n4463), .B2(n2860), .A(n2859), .ZN(n4455) );
  XNOR2_X1 U2495 ( .A(n2334), .B(IR_REG_30__SCAN_IN), .ZN(n3278) );
  NOR2_X4 U2496 ( .A1(n2575), .A2(n2161), .ZN(n2472) );
  NAND2_X1 U2497 ( .A1(n3392), .A2(n2990), .ZN(n4000) );
  NOR2_X2 U2498 ( .A1(n3930), .A2(n3931), .ZN(n3929) );
  OAI22_X2 U2499 ( .A1(n3087), .A2(n2197), .B1(n2199), .B2(n2184), .ZN(n3930)
         );
  BUF_X4 U2500 ( .A(n3008), .Z(n2142) );
  OAI21_X1 U2501 ( .B1(n4256), .B2(n2390), .A(n2387), .ZN(n2758) );
  AOI21_X1 U2502 ( .B1(n4256), .B2(n4121), .A(n4052), .ZN(n4239) );
  OR2_X1 U2503 ( .A1(n4304), .A2(n4305), .ZN(n4326) );
  MUX2_X2 U2504 ( .A(n4621), .B(n4620), .S(n4751), .Z(n4622) );
  NAND2_X2 U2505 ( .A1(n2165), .A2(n2453), .ZN(n2575) );
  AND4_X2 U2506 ( .A1(n4784), .A2(n2451), .A3(n2450), .A4(n2511), .ZN(n2165)
         );
  MUX2_X2 U2507 ( .A(n4837), .B(n4624), .S(n4751), .Z(n4625) );
  MUX2_X2 U2508 ( .A(n4839), .B(n4624), .S(n4756), .Z(n4516) );
  XNOR2_X2 U2509 ( .A(n4237), .B(n4238), .ZN(n4512) );
  NAND2_X2 U2510 ( .A1(n2141), .A2(n2475), .ZN(n2541) );
  INV_X2 U2511 ( .A(n2518), .ZN(n2501) );
  OAI21_X2 U2512 ( .B1(n3658), .B2(n2853), .A(n2852), .ZN(n3669) );
  NAND2_X1 U2513 ( .A1(n3278), .A2(n3271), .ZN(n2518) );
  OR2_X1 U2514 ( .A1(n2415), .A2(n3872), .ZN(n2410) );
  AOI21_X1 U2515 ( .B1(n2414), .B2(n2413), .A(n2192), .ZN(n2412) );
  INV_X1 U2516 ( .A(IR_REG_17__SCAN_IN), .ZN(n2648) );
  INV_X1 U2517 ( .A(IR_REG_20__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U2518 ( .A1(n2759), .A2(IR_REG_31__SCAN_IN), .ZN(n2761) );
  OR2_X1 U2519 ( .A1(n2975), .A2(n4681), .ZN(n3174) );
  NAND2_X1 U2520 ( .A1(n2949), .A2(n2948), .ZN(n2950) );
  INV_X1 U2521 ( .A(n2391), .ZN(n2390) );
  AOI21_X1 U2522 ( .B1(n2391), .B2(n2389), .A(n2388), .ZN(n2387) );
  AND2_X1 U2523 ( .A1(n2392), .A2(n4051), .ZN(n2391) );
  INV_X1 U2524 ( .A(n2185), .ZN(n2396) );
  AND2_X1 U2525 ( .A1(n2710), .A2(n2254), .ZN(n2741) );
  NOR2_X1 U2526 ( .A1(n2255), .A2(n2258), .ZN(n2254) );
  OR2_X1 U2527 ( .A1(n2257), .A2(n2256), .ZN(n2255) );
  INV_X1 U2528 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2258) );
  INV_X1 U2529 ( .A(n2338), .ZN(n2337) );
  OAI21_X1 U2530 ( .B1(n4454), .B2(n2339), .A(n2862), .ZN(n2338) );
  NAND2_X1 U2531 ( .A1(n2281), .A2(n2279), .ZN(n2278) );
  AND2_X1 U2532 ( .A1(n4020), .A2(n4011), .ZN(n2405) );
  INV_X1 U2533 ( .A(n4012), .ZN(n2279) );
  INV_X1 U2534 ( .A(n2281), .ZN(n2280) );
  INV_X1 U2535 ( .A(IR_REG_15__SCAN_IN), .ZN(n2643) );
  INV_X1 U2536 ( .A(n2421), .ZN(n2420) );
  NAND2_X1 U2537 ( .A1(n3480), .A2(n3481), .ZN(n2428) );
  OR2_X1 U2538 ( .A1(n2201), .A2(n2184), .ZN(n2197) );
  INV_X1 U2539 ( .A(n2200), .ZN(n2199) );
  AOI21_X1 U2540 ( .B1(n2211), .B2(n2213), .A(n2210), .ZN(n2209) );
  INV_X1 U2541 ( .A(n2213), .ZN(n2212) );
  INV_X1 U2542 ( .A(n2217), .ZN(n2211) );
  OR2_X1 U2543 ( .A1(n2617), .A2(n3987), .ZN(n2627) );
  NOR2_X1 U2544 ( .A1(n3310), .A2(n2437), .ZN(n2894) );
  NOR2_X1 U2545 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2451)
         );
  NAND2_X1 U2546 ( .A1(n3535), .A2(n2900), .ZN(n2308) );
  OR2_X1 U2547 ( .A1(n3533), .A2(n2897), .ZN(n2900) );
  AOI21_X1 U2548 ( .B1(n2317), .B2(REG1_REG_12__SCAN_IN), .A(n4685), .ZN(n2314) );
  AND2_X1 U2549 ( .A1(n2363), .A2(n2362), .ZN(n2361) );
  NOR2_X1 U2550 ( .A1(n2180), .A2(n2366), .ZN(n2365) );
  INV_X1 U2551 ( .A(n2367), .ZN(n2366) );
  AND2_X1 U2552 ( .A1(n2734), .A2(n4255), .ZN(n4121) );
  AOI21_X1 U2553 ( .B1(n2286), .B2(n2400), .A(n4454), .ZN(n2285) );
  NAND2_X1 U2554 ( .A1(n3195), .A2(n2445), .ZN(n3196) );
  INV_X1 U2555 ( .A(n3868), .ZN(n4511) );
  NAND2_X1 U2556 ( .A1(n2769), .A2(n2768), .ZN(n4590) );
  AND2_X1 U2557 ( .A1(n3367), .A2(n4680), .ZN(n4540) );
  NOR2_X1 U2558 ( .A1(n2672), .A2(n2649), .ZN(n2650) );
  OR2_X1 U2559 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2649)
         );
  NOR2_X1 U2560 ( .A1(n2526), .A2(IR_REG_5__SCAN_IN), .ZN(n2537) );
  INV_X1 U2561 ( .A(n4681), .ZN(n4211) );
  XNOR2_X1 U2562 ( .A(n2928), .B(n3568), .ZN(n4164) );
  NAND2_X1 U2563 ( .A1(n3331), .A2(n3332), .ZN(n3330) );
  NOR3_X1 U2564 ( .A1(n4094), .A2(n4348), .A3(n4454), .ZN(n2270) );
  INV_X1 U2565 ( .A(n3080), .ZN(n3074) );
  OR2_X1 U2566 ( .A1(n4363), .A2(n2685), .ZN(n4109) );
  INV_X1 U2567 ( .A(n2348), .ZN(n2347) );
  OAI21_X1 U2568 ( .B1(n2863), .B2(n2349), .A(n2866), .ZN(n2348) );
  INV_X1 U2569 ( .A(n2865), .ZN(n2349) );
  INV_X1 U2570 ( .A(n4412), .ZN(n2863) );
  INV_X1 U2571 ( .A(n4003), .ZN(n2386) );
  AND2_X1 U2572 ( .A1(n2156), .A2(n4266), .ZN(n2409) );
  AND2_X1 U2573 ( .A1(n4399), .A2(n4376), .ZN(n2408) );
  INV_X1 U2574 ( .A(n4417), .ZN(n3088) );
  AND2_X1 U2575 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2464)
         );
  AND2_X1 U2576 ( .A1(n2762), .A2(n2438), .ZN(n2461) );
  AND2_X1 U2577 ( .A1(n2143), .A2(n2166), .ZN(n2795) );
  INV_X1 U2578 ( .A(n2642), .ZN(n2646) );
  NAND2_X1 U2579 ( .A1(n2455), .A2(n2454), .ZN(n2642) );
  INV_X1 U2580 ( .A(IR_REG_12__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U2581 ( .A1(n2426), .A2(n2425), .ZN(n2424) );
  INV_X1 U2582 ( .A(n3518), .ZN(n2426) );
  INV_X1 U2583 ( .A(n3519), .ZN(n2425) );
  NAND2_X1 U2584 ( .A1(n3518), .A2(n3519), .ZN(n2423) );
  NAND2_X1 U2585 ( .A1(n3942), .A2(n3057), .ZN(n2416) );
  NAND2_X1 U2586 ( .A1(n2434), .A2(n2433), .ZN(n3262) );
  NAND2_X1 U2587 ( .A1(n3702), .A2(n3042), .ZN(n3771) );
  INV_X1 U2588 ( .A(n3472), .ZN(n2207) );
  AND2_X1 U2589 ( .A1(n3853), .A2(n3126), .ZN(n3127) );
  NAND2_X1 U2590 ( .A1(n2579), .A2(n2149), .ZN(n2617) );
  INV_X1 U2591 ( .A(n4133), .ZN(n2271) );
  NAND2_X1 U2592 ( .A1(n2267), .A2(n2827), .ZN(n2266) );
  OAI211_X1 U2593 ( .C1(n2750), .C2(n3603), .A(n2546), .B(n2547), .ZN(n2331)
         );
  OR2_X1 U2594 ( .A1(n2541), .A2(n2479), .ZN(n2482) );
  NAND2_X1 U2595 ( .A1(n2791), .A2(n2452), .ZN(n2492) );
  NAND2_X1 U2596 ( .A1(n3334), .A2(n3335), .ZN(n3333) );
  AND2_X1 U2597 ( .A1(n3333), .A2(n2305), .ZN(n2889) );
  NAND2_X1 U2598 ( .A1(n4690), .A2(REG1_REG_2__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2599 ( .A1(n3330), .A2(n2931), .ZN(n2243) );
  NAND2_X1 U2600 ( .A1(n2228), .A2(n2226), .ZN(n2939) );
  INV_X1 U2601 ( .A(n2229), .ZN(n2228) );
  OAI21_X1 U2602 ( .B1(n2936), .B2(n2230), .A(n2938), .ZN(n2229) );
  NAND2_X1 U2603 ( .A1(n2311), .A2(n2896), .ZN(n2310) );
  OR2_X1 U2604 ( .A1(n3374), .A2(n4796), .ZN(n2896) );
  NAND2_X1 U2605 ( .A1(n3376), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U2606 ( .A1(n2240), .A2(n2238), .ZN(n2954) );
  INV_X1 U2607 ( .A(n2239), .ZN(n2238) );
  OAI21_X1 U2608 ( .B1(n2951), .B2(n2378), .A(n2953), .ZN(n2239) );
  XNOR2_X1 U2609 ( .A(n2954), .B(n3792), .ZN(n3790) );
  OAI21_X1 U2610 ( .B1(n3810), .B2(n2957), .A(n2958), .ZN(n2959) );
  AND2_X1 U2611 ( .A1(n2960), .A2(n2385), .ZN(n4693) );
  INV_X1 U2612 ( .A(n4694), .ZN(n2385) );
  OR2_X1 U2613 ( .A1(n2741), .A2(n2736), .ZN(n4245) );
  NAND2_X1 U2614 ( .A1(n2664), .A2(n2272), .ZN(n2700) );
  AND2_X1 U2615 ( .A1(n2157), .A2(n2194), .ZN(n2272) );
  NOR2_X1 U2616 ( .A1(n2700), .A2(n3885), .ZN(n2710) );
  AOI21_X1 U2617 ( .B1(n2153), .B2(n2342), .A(n2188), .ZN(n2341) );
  INV_X1 U2618 ( .A(n2179), .ZN(n2342) );
  NAND2_X1 U2619 ( .A1(n2664), .A2(n2157), .ZN(n2694) );
  NOR2_X1 U2620 ( .A1(n2627), .A2(n4855), .ZN(n2664) );
  AOI21_X1 U2621 ( .B1(n2337), .B2(n2339), .A(n2169), .ZN(n2335) );
  NAND2_X1 U2622 ( .A1(n2864), .A2(n2863), .ZN(n4406) );
  AOI21_X1 U2623 ( .B1(n2399), .B2(n3756), .A(n2287), .ZN(n2286) );
  INV_X1 U2624 ( .A(n4017), .ZN(n2287) );
  INV_X1 U2625 ( .A(n4462), .ZN(n2626) );
  NAND2_X1 U2626 ( .A1(n2354), .A2(n2144), .ZN(n2353) );
  NAND2_X1 U2627 ( .A1(n2353), .A2(n2352), .ZN(n4488) );
  AND2_X1 U2628 ( .A1(n2549), .A2(n4012), .ZN(n2282) );
  INV_X1 U2629 ( .A(n4013), .ZN(n2283) );
  NAND2_X1 U2630 ( .A1(n3590), .A2(n4012), .ZN(n2276) );
  AND3_X1 U2631 ( .A1(n3554), .A2(n2175), .A3(n3631), .ZN(n2403) );
  NAND2_X1 U2632 ( .A1(n3209), .A2(n2785), .ZN(n4217) );
  NAND2_X1 U2633 ( .A1(n4316), .A2(n2409), .ZN(n4265) );
  INV_X1 U2634 ( .A(n4744), .ZN(n4607) );
  INV_X1 U2635 ( .A(n4590), .ZN(n4485) );
  NAND2_X1 U2636 ( .A1(n3554), .A2(n3553), .ZN(n3552) );
  INV_X1 U2637 ( .A(n4544), .ZN(n4598) );
  AND3_X1 U2638 ( .A1(n3206), .A2(n3205), .A3(n3204), .ZN(n3214) );
  AND2_X1 U2639 ( .A1(n2625), .A2(n2632), .ZN(n2962) );
  OR2_X1 U2640 ( .A1(n2513), .A2(n2512), .ZN(n2526) );
  INV_X1 U2641 ( .A(IR_REG_5__SCAN_IN), .ZN(n2514) );
  INV_X1 U2642 ( .A(IR_REG_1__SCAN_IN), .ZN(n2236) );
  AOI21_X1 U2643 ( .B1(n3964), .B2(n3966), .A(n3965), .ZN(n3864) );
  AND2_X1 U2644 ( .A1(n2430), .A2(n3119), .ZN(n2429) );
  NAND2_X1 U2645 ( .A1(n3457), .A2(n3012), .ZN(n3473) );
  AND2_X1 U2646 ( .A1(n2707), .A2(n2706), .ZN(n4332) );
  NAND2_X1 U2647 ( .A1(n2224), .A2(n3262), .ZN(n2223) );
  NAND2_X1 U2648 ( .A1(n2432), .A2(n2225), .ZN(n2224) );
  INV_X1 U2649 ( .A(n3263), .ZN(n2225) );
  NAND2_X1 U2650 ( .A1(n2434), .A2(n2183), .ZN(n2432) );
  OR2_X1 U2651 ( .A1(n3183), .A2(n3179), .ZN(n3984) );
  AND2_X1 U2652 ( .A1(n3181), .A2(n4492), .ZN(n3986) );
  INV_X1 U2653 ( .A(n4576), .ZN(n4482) );
  OR2_X1 U2654 ( .A1(n3183), .A2(n3182), .ZN(n3988) );
  NAND2_X1 U2655 ( .A1(n2253), .A2(n2749), .ZN(n3868) );
  OR2_X1 U2656 ( .A1(n4226), .A2(n2750), .ZN(n2253) );
  NAND2_X1 U2657 ( .A1(n2733), .A2(n2732), .ZN(n4508) );
  OAI21_X1 U2658 ( .B1(n4421), .B2(n2750), .A(n2662), .ZN(n4561) );
  NAND4_X1 U2659 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4149)
         );
  INV_X1 U2660 ( .A(n3685), .ZN(n3691) );
  NAND2_X1 U2661 ( .A1(n4163), .A2(n2930), .ZN(n3331) );
  NAND2_X1 U2662 ( .A1(n2380), .A2(n2379), .ZN(n3332) );
  NAND2_X1 U2663 ( .A1(n3329), .A2(REG2_REG_2__SCAN_IN), .ZN(n2379) );
  OR2_X1 U2664 ( .A1(n3329), .A2(REG2_REG_2__SCAN_IN), .ZN(n2380) );
  OAI21_X1 U2665 ( .B1(n3350), .B2(n2324), .A(n2322), .ZN(n3310) );
  OR2_X1 U2666 ( .A1(n3311), .A2(n4752), .ZN(n2324) );
  INV_X1 U2667 ( .A(n3311), .ZN(n2323) );
  XNOR2_X1 U2668 ( .A(n2939), .B(n3343), .ZN(n3340) );
  NAND2_X1 U2669 ( .A1(n2899), .A2(n2898), .ZN(n3535) );
  INV_X1 U2670 ( .A(n3530), .ZN(n2898) );
  XNOR2_X1 U2671 ( .A(n2308), .B(n3641), .ZN(n3638) );
  INV_X1 U2672 ( .A(n2901), .ZN(n2902) );
  NAND2_X1 U2673 ( .A1(n4186), .A2(REG2_REG_14__SCAN_IN), .ZN(n4185) );
  NOR2_X1 U2674 ( .A1(n4711), .A2(REG1_REG_16__SCAN_IN), .ZN(n4712) );
  OR2_X1 U2675 ( .A1(n3306), .A2(n4677), .ZN(n4199) );
  NAND2_X1 U2676 ( .A1(n4193), .A2(n2252), .ZN(n2251) );
  OR2_X1 U2677 ( .A1(n4192), .A2(n4194), .ZN(n2252) );
  NAND2_X1 U2678 ( .A1(n2250), .A2(n4195), .ZN(n2249) );
  NAND2_X1 U2679 ( .A1(n4709), .A2(ADDR_REG_17__SCAN_IN), .ZN(n2250) );
  NAND2_X1 U2680 ( .A1(n2330), .A2(n2329), .ZN(n2328) );
  NAND2_X1 U2681 ( .A1(n2913), .A2(n2330), .ZN(n2327) );
  INV_X1 U2682 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2329) );
  NOR2_X1 U2683 ( .A1(n2966), .A2(n2967), .ZN(n4201) );
  OR2_X1 U2684 ( .A1(n4201), .A2(n2382), .ZN(n2381) );
  AND2_X1 U2685 ( .A1(n4202), .A2(REG2_REG_18__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U2686 ( .A1(n2355), .A2(n2358), .ZN(n2877) );
  AOI21_X1 U2687 ( .B1(n2361), .B2(n2359), .A(n2371), .ZN(n2358) );
  NAND2_X1 U2688 ( .A1(n2393), .A2(n2392), .ZN(n3191) );
  AND2_X1 U2689 ( .A1(n2756), .A2(n2755), .ZN(n4229) );
  NAND2_X1 U2690 ( .A1(n2364), .A2(n2362), .ZN(n3193) );
  NAND2_X1 U2691 ( .A1(n2368), .A2(n2365), .ZN(n2364) );
  NAND2_X1 U2692 ( .A1(n4724), .A2(n2829), .ZN(n4498) );
  NAND2_X1 U2693 ( .A1(n4217), .A2(n2786), .ZN(n3230) );
  OR2_X1 U2694 ( .A1(n3209), .A2(n2785), .ZN(n2786) );
  INV_X1 U2695 ( .A(IR_REG_29__SCAN_IN), .ZN(n2288) );
  AOI21_X1 U2696 ( .B1(n2653), .B2(n2652), .A(n2651), .ZN(n2654) );
  INV_X1 U2697 ( .A(IR_REG_18__SCAN_IN), .ZN(n2652) );
  INV_X1 U2698 ( .A(n2416), .ZN(n2413) );
  INV_X1 U2699 ( .A(n2394), .ZN(n2389) );
  INV_X1 U2700 ( .A(n4055), .ZN(n2388) );
  INV_X1 U2701 ( .A(n2423), .ZN(n2422) );
  OAI21_X1 U2702 ( .B1(n2202), .B2(n2201), .A(n3892), .ZN(n2200) );
  INV_X1 U2703 ( .A(n3954), .ZN(n2201) );
  NAND2_X1 U2704 ( .A1(n2219), .A2(n2218), .ZN(n2217) );
  INV_X1 U2705 ( .A(n3768), .ZN(n2218) );
  INV_X1 U2706 ( .A(n3769), .ZN(n2219) );
  NOR2_X1 U2707 ( .A1(n3798), .A2(n2214), .ZN(n2213) );
  INV_X1 U2708 ( .A(n2216), .ZN(n2214) );
  INV_X1 U2709 ( .A(n3799), .ZN(n2210) );
  NAND2_X1 U2710 ( .A1(n3114), .A2(n2436), .ZN(n2435) );
  NAND2_X1 U2711 ( .A1(n3472), .A2(n2206), .ZN(n2205) );
  INV_X1 U2712 ( .A(n3012), .ZN(n2206) );
  NAND2_X1 U2713 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2257) );
  OR2_X1 U2714 ( .A1(n2677), .A2(n4387), .ZN(n4104) );
  NOR2_X1 U2715 ( .A1(n4290), .A2(n2269), .ZN(n2268) );
  NAND2_X1 U2716 ( .A1(n4343), .A2(n2270), .ZN(n2269) );
  NOR2_X1 U2717 ( .A1(n2248), .A2(n2245), .ZN(n2242) );
  INV_X1 U2718 ( .A(n3314), .ZN(n2230) );
  NOR2_X1 U2719 ( .A1(n2230), .A2(n2505), .ZN(n2227) );
  NOR2_X1 U2720 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2450)
         );
  NOR2_X1 U2721 ( .A1(n2316), .A2(n4968), .ZN(n2313) );
  NOR2_X1 U2722 ( .A1(n2320), .A2(n2319), .ZN(n2316) );
  NAND2_X1 U2723 ( .A1(n2318), .A2(n4685), .ZN(n2317) );
  INV_X1 U2724 ( .A(n4175), .ZN(n2378) );
  NOR2_X1 U2725 ( .A1(n2378), .A2(n3673), .ZN(n2237) );
  NAND2_X1 U2726 ( .A1(n5037), .A2(n4280), .ZN(n2874) );
  AND2_X1 U2727 ( .A1(n4261), .A2(n4280), .ZN(n4116) );
  INV_X1 U2728 ( .A(n2861), .ZN(n2339) );
  INV_X1 U2729 ( .A(n2857), .ZN(n2351) );
  AND2_X1 U2730 ( .A1(n4477), .A2(n4070), .ZN(n4038) );
  NOR2_X1 U2731 ( .A1(n3773), .A2(n2260), .ZN(n2259) );
  INV_X1 U2732 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2260) );
  INV_X1 U2733 ( .A(n3151), .ZN(n2817) );
  OR2_X1 U2734 ( .A1(n4464), .A2(n4446), .ZN(n4429) );
  OR2_X1 U2735 ( .A1(n2621), .A2(IR_REG_14__SCAN_IN), .ZN(n2622) );
  INV_X1 U2736 ( .A(IR_REG_4__SCAN_IN), .ZN(n4785) );
  INV_X1 U2737 ( .A(n3374), .ZN(n2540) );
  AND2_X1 U2738 ( .A1(n3263), .A2(n2183), .ZN(n2433) );
  NAND2_X1 U2739 ( .A1(n2433), .A2(n2435), .ZN(n2430) );
  NOR2_X1 U2740 ( .A1(n3953), .A2(n2203), .ZN(n2202) );
  INV_X1 U2741 ( .A(n2444), .ZN(n2203) );
  NAND2_X1 U2742 ( .A1(n3769), .A2(n3768), .ZN(n2216) );
  NAND2_X1 U2743 ( .A1(n3771), .A2(n2217), .ZN(n2215) );
  NOR2_X1 U2744 ( .A1(n2568), .A2(n4823), .ZN(n2579) );
  INV_X1 U2745 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4823) );
  AND2_X1 U2746 ( .A1(n3107), .A2(n3106), .ZN(n3933) );
  NAND2_X1 U2747 ( .A1(n2579), .A2(REG3_REG_10__SCAN_IN), .ZN(n2587) );
  OAI22_X1 U2748 ( .A1(n3444), .A2(n3008), .B1(n2988), .B2(n3571), .ZN(n2985)
         );
  NAND2_X1 U2749 ( .A1(n3074), .A2(n3073), .ZN(n3084) );
  INV_X1 U2750 ( .A(n3082), .ZN(n3083) );
  NOR2_X1 U2751 ( .A1(n2519), .A2(n3315), .ZN(n2529) );
  OR2_X1 U2752 ( .A1(n4540), .A2(n3156), .ZN(n3169) );
  NOR2_X1 U2753 ( .A1(n2719), .A2(n2257), .ZN(n2735) );
  NOR2_X1 U2754 ( .A1(n3177), .A2(n3176), .ZN(n4137) );
  OR2_X1 U2755 ( .A1(n3837), .A2(n3626), .ZN(n2534) );
  NAND2_X1 U2756 ( .A1(n2544), .A2(REG0_REG_1__SCAN_IN), .ZN(n2299) );
  NAND2_X1 U2757 ( .A1(n2545), .A2(REG1_REG_1__SCAN_IN), .ZN(n2298) );
  XNOR2_X1 U2758 ( .A(n2950), .B(n3641), .ZN(n3639) );
  NOR2_X1 U2759 ( .A1(n2321), .A2(n3792), .ZN(n2320) );
  INV_X1 U2760 ( .A(n2442), .ZN(n2321) );
  NAND2_X1 U2761 ( .A1(n3816), .A2(n2906), .ZN(n2907) );
  NOR2_X1 U2762 ( .A1(n4693), .A2(n2384), .ZN(n2963) );
  AND2_X1 U2763 ( .A1(n2962), .A2(REG2_REG_15__SCAN_IN), .ZN(n2384) );
  INV_X1 U2764 ( .A(n4191), .ZN(n2330) );
  NOR2_X1 U2765 ( .A1(n2360), .A2(n2357), .ZN(n2356) );
  INV_X1 U2766 ( .A(n2874), .ZN(n2357) );
  INV_X1 U2767 ( .A(n2361), .ZN(n2360) );
  INV_X1 U2768 ( .A(n2365), .ZN(n2359) );
  OR2_X1 U2769 ( .A1(n2397), .A2(n2396), .ZN(n2392) );
  AND2_X1 U2770 ( .A1(n4238), .A2(n2398), .ZN(n2397) );
  NOR2_X1 U2771 ( .A1(n2396), .A2(n2395), .ZN(n2394) );
  INV_X1 U2772 ( .A(n4121), .ZN(n2395) );
  OR2_X1 U2773 ( .A1(n2370), .A2(n2180), .ZN(n2362) );
  AND2_X1 U2774 ( .A1(n2876), .A2(n2372), .ZN(n2370) );
  INV_X1 U2775 ( .A(n4095), .ZN(n2372) );
  NOR2_X1 U2776 ( .A1(n2369), .A2(n2186), .ZN(n2367) );
  NAND2_X1 U2777 ( .A1(n4312), .A2(n4298), .ZN(n2872) );
  NAND2_X1 U2778 ( .A1(n4518), .A2(n4292), .ZN(n2871) );
  NAND2_X1 U2779 ( .A1(n2344), .A2(n2179), .ZN(n2343) );
  AOI21_X1 U2780 ( .B1(n2347), .B2(n2349), .A(n2173), .ZN(n2345) );
  NAND2_X1 U2781 ( .A1(n2664), .A2(n2154), .ZN(n2678) );
  AND2_X1 U2782 ( .A1(n2664), .A2(n2634), .ZN(n2657) );
  AND2_X1 U2783 ( .A1(n4388), .A2(n4389), .ZN(n4412) );
  NAND2_X1 U2784 ( .A1(n2140), .A2(n4454), .ZN(n4453) );
  INV_X1 U2785 ( .A(n4570), .ZN(n4446) );
  NAND2_X1 U2786 ( .A1(n2579), .A2(n2259), .ZN(n2603) );
  INV_X1 U2787 ( .A(n4014), .ZN(n2274) );
  INV_X1 U2788 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2556) );
  NAND4_X1 U2789 ( .A1(n2265), .A2(n2262), .A3(REG3_REG_5__SCAN_IN), .A4(
        REG3_REG_7__SCAN_IN), .ZN(n2568) );
  NOR2_X1 U2790 ( .A1(n2264), .A2(n2556), .ZN(n2262) );
  INV_X1 U2791 ( .A(n3585), .ZN(n3616) );
  OAI21_X1 U2792 ( .B1(n3590), .B2(n2549), .A(n4012), .ZN(n3608) );
  NAND2_X1 U2793 ( .A1(n2263), .A2(n2265), .ZN(n2542) );
  NOR2_X1 U2794 ( .A1(n3315), .A2(n2264), .ZN(n2263) );
  INV_X1 U2795 ( .A(n4007), .ZN(n2293) );
  CLKBUF_X1 U2796 ( .A(n3251), .Z(n3252) );
  NAND2_X1 U2797 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2519) );
  CLKBUF_X1 U2798 ( .A(n3539), .Z(n4087) );
  AND2_X1 U2799 ( .A1(n3432), .A2(n4154), .ZN(n3403) );
  CLKBUF_X1 U2800 ( .A(n3400), .Z(n3401) );
  AOI21_X1 U2801 ( .B1(n2817), .B2(n3287), .A(n3286), .ZN(n3213) );
  NOR2_X1 U2802 ( .A1(n4217), .A2(n4218), .ZN(n4216) );
  AND2_X1 U2803 ( .A1(n4241), .A2(n4230), .ZN(n3209) );
  NAND2_X1 U2804 ( .A1(n4316), .A2(n2156), .ZN(n4277) );
  AND2_X1 U2805 ( .A1(n4316), .A2(n4298), .ZN(n4296) );
  INV_X1 U2806 ( .A(n3886), .ZN(n4315) );
  NAND2_X1 U2807 ( .A1(n4409), .A2(n2159), .ZN(n4338) );
  NAND2_X1 U2808 ( .A1(n3832), .A2(DATAI_20_), .ZN(n4376) );
  AND2_X1 U2809 ( .A1(n4409), .A2(n2408), .ZN(n4378) );
  INV_X1 U2810 ( .A(n4393), .ZN(n4399) );
  OR2_X1 U2811 ( .A1(n4429), .A2(n4431), .ZN(n4430) );
  NAND2_X1 U2812 ( .A1(n4465), .A2(n4579), .ZN(n4464) );
  INV_X1 U2813 ( .A(n3069), .ZN(n4579) );
  AND2_X1 U2814 ( .A1(n3748), .A2(n2407), .ZN(n4465) );
  AND2_X1 U2815 ( .A1(n2151), .A2(n4588), .ZN(n2407) );
  NAND2_X1 U2816 ( .A1(n3748), .A2(n2145), .ZN(n4496) );
  NAND2_X1 U2817 ( .A1(n3748), .A2(n3774), .ZN(n3747) );
  AND2_X1 U2818 ( .A1(n3671), .A2(n3704), .ZN(n3748) );
  NOR2_X1 U2819 ( .A1(n2449), .A2(n3659), .ZN(n3671) );
  OR2_X1 U2820 ( .A1(n3617), .A2(n3616), .ZN(n2449) );
  NAND2_X1 U2821 ( .A1(n2404), .A2(n3474), .ZN(n2439) );
  NOR2_X1 U2822 ( .A1(n3399), .A2(n2784), .ZN(n3554) );
  INV_X1 U2823 ( .A(n4540), .ZN(n4603) );
  NAND2_X1 U2824 ( .A1(n3364), .A2(n3571), .ZN(n3399) );
  AND2_X1 U2825 ( .A1(n2461), .A2(n2462), .ZN(n2402) );
  NAND2_X1 U2826 ( .A1(n2795), .A2(n2789), .ZN(n2799) );
  NOR2_X1 U2827 ( .A1(IR_REG_22__SCAN_IN), .A2(n2788), .ZN(n2789) );
  NOR2_X1 U2828 ( .A1(n2575), .A2(n2647), .ZN(n2670) );
  OR2_X1 U2829 ( .A1(n2586), .A2(n2791), .ZN(n2594) );
  INV_X1 U2830 ( .A(IR_REG_7__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U2831 ( .A1(n3521), .A2(n2424), .ZN(n2419) );
  NAND2_X1 U2832 ( .A1(n3941), .A2(n2416), .ZN(n2411) );
  INV_X1 U2833 ( .A(n3701), .ZN(n3039) );
  NAND2_X1 U2834 ( .A1(n2198), .A2(n3954), .ZN(n3891) );
  NAND2_X1 U2835 ( .A1(n3087), .A2(n2202), .ZN(n2198) );
  NAND2_X1 U2836 ( .A1(n2977), .A2(n3146), .ZN(n2980) );
  NAND2_X1 U2837 ( .A1(n3832), .A2(DATAI_21_), .ZN(n4356) );
  AND2_X1 U2838 ( .A1(n2189), .A2(n2720), .ZN(n4278) );
  NAND2_X1 U2839 ( .A1(n3473), .A2(n3472), .ZN(n3471) );
  AND2_X1 U2840 ( .A1(n2711), .A2(n2719), .ZN(n4299) );
  INV_X1 U2841 ( .A(n3456), .ZN(n3009) );
  INV_X1 U2842 ( .A(n4414), .ZN(n3958) );
  INV_X1 U2843 ( .A(n3988), .ZN(n3961) );
  INV_X1 U2844 ( .A(n3984), .ZN(n3923) );
  OAI21_X1 U2845 ( .B1(n3130), .B2(n3855), .A(n3129), .ZN(n3131) );
  INV_X1 U2846 ( .A(n3993), .ZN(n3972) );
  OAI21_X1 U2847 ( .B1(n2271), .B2(n2827), .A(n2266), .ZN(n4134) );
  INV_X1 U2848 ( .A(n4229), .ZN(n4147) );
  OAI21_X1 U2849 ( .B1(n4245), .B2(n2750), .A(n2740), .ZN(n4148) );
  INV_X1 U2850 ( .A(n4332), .ZN(n4293) );
  NAND2_X1 U2851 ( .A1(n2699), .A2(n2698), .ZN(n4329) );
  NAND2_X1 U2852 ( .A1(n2684), .A2(n2683), .ZN(n4541) );
  NAND2_X1 U2853 ( .A1(n2669), .A2(n2668), .ZN(n4568) );
  OAI211_X1 U2854 ( .C1(n4447), .C2(n2750), .A(n2631), .B(n2630), .ZN(n4577)
         );
  OAI211_X1 U2855 ( .C1(n4466), .C2(n2750), .A(n2620), .B(n2619), .ZN(n4585)
         );
  OR2_X1 U2856 ( .A1(n2614), .A2(n2613), .ZN(n4576) );
  INV_X1 U2857 ( .A(n3630), .ZN(n4151) );
  NAND2_X1 U2858 ( .A1(n2491), .A2(IR_REG_2__SCAN_IN), .ZN(n2494) );
  AND2_X1 U2859 ( .A1(n2513), .A2(n2492), .ZN(n2493) );
  NAND2_X1 U2860 ( .A1(n2247), .A2(n2246), .ZN(n3290) );
  NAND2_X1 U2861 ( .A1(n2243), .A2(n2932), .ZN(n2247) );
  OR2_X1 U2862 ( .A1(n3350), .A2(n4752), .ZN(n2326) );
  INV_X1 U2863 ( .A(n2892), .ZN(n2325) );
  NAND2_X1 U2864 ( .A1(n3313), .A2(n3314), .ZN(n3312) );
  NAND2_X1 U2865 ( .A1(n2231), .A2(n2936), .ZN(n3313) );
  NAND2_X1 U2866 ( .A1(n3348), .A2(REG2_REG_4__SCAN_IN), .ZN(n2231) );
  AOI21_X1 U2867 ( .B1(n2940), .B2(n3626), .A(n2377), .ZN(n2374) );
  INV_X1 U2868 ( .A(n3377), .ZN(n2377) );
  NAND2_X1 U2869 ( .A1(n2376), .A2(n2940), .ZN(n3378) );
  NAND2_X1 U2870 ( .A1(n3340), .A2(REG2_REG_6__SCAN_IN), .ZN(n2376) );
  OR2_X1 U2871 ( .A1(n2894), .A2(n3343), .ZN(n2895) );
  NAND2_X1 U2872 ( .A1(n2308), .A2(n4687), .ZN(n2306) );
  NAND2_X1 U2873 ( .A1(n3638), .A2(REG1_REG_10__SCAN_IN), .ZN(n2307) );
  NAND2_X1 U2874 ( .A1(n2952), .A2(n2951), .ZN(n4176) );
  NAND2_X1 U2875 ( .A1(n3639), .A2(REG2_REG_10__SCAN_IN), .ZN(n2952) );
  NAND2_X1 U2876 ( .A1(n4176), .A2(n4175), .ZN(n4174) );
  OAI211_X1 U2877 ( .C1(n4168), .C2(n4685), .A(n2315), .B(n2318), .ZN(n3788)
         );
  NAND2_X1 U2878 ( .A1(n4168), .A2(n2320), .ZN(n2315) );
  NAND2_X1 U2879 ( .A1(n2905), .A2(n2904), .ZN(n3816) );
  INV_X1 U2880 ( .A(n3811), .ZN(n2904) );
  NAND2_X1 U2881 ( .A1(n2956), .A2(n2955), .ZN(n3810) );
  XNOR2_X1 U2882 ( .A(n2959), .B(n4683), .ZN(n4186) );
  INV_X1 U2883 ( .A(n2960), .ZN(n4695) );
  XNOR2_X1 U2884 ( .A(n2963), .B(n2911), .ZN(n4706) );
  NAND2_X1 U2885 ( .A1(n4706), .A2(n4704), .ZN(n4705) );
  NAND2_X1 U2886 ( .A1(n4193), .A2(n2383), .ZN(n2966) );
  OR2_X1 U2887 ( .A1(n4682), .A2(REG2_REG_17__SCAN_IN), .ZN(n2383) );
  NAND2_X1 U2888 ( .A1(n4406), .A2(n2865), .ZN(n4398) );
  OAI21_X1 U2889 ( .B1(n3754), .B2(n2400), .A(n2286), .ZN(n4442) );
  NAND2_X1 U2890 ( .A1(n2401), .A2(n4036), .ZN(n4461) );
  NAND2_X1 U2891 ( .A1(n3754), .A2(n4079), .ZN(n2401) );
  AND2_X1 U2892 ( .A1(n2353), .A2(n2163), .ZN(n3739) );
  NAND2_X1 U2893 ( .A1(n2406), .A2(n4011), .ZN(n3656) );
  NAND2_X1 U2894 ( .A1(n2276), .A2(n2281), .ZN(n2406) );
  INV_X1 U2895 ( .A(n3525), .ZN(n3632) );
  OAI21_X1 U2896 ( .B1(n4243), .B2(n4246), .A(n4242), .ZN(n4623) );
  OAI21_X1 U2897 ( .B1(n4511), .B2(n4544), .A(n4509), .ZN(n2304) );
  NAND2_X1 U2898 ( .A1(n3151), .A2(n3423), .ZN(n4728) );
  NAND2_X1 U2899 ( .A1(n3847), .A2(IR_REG_31__SCAN_IN), .ZN(n2334) );
  INV_X1 U2900 ( .A(n2975), .ZN(n4140) );
  INV_X1 U2901 ( .A(n4202), .ZN(n4732) );
  INV_X1 U2902 ( .A(n3641), .ZN(n4687) );
  XNOR2_X1 U2903 ( .A(n2566), .B(n2565), .ZN(n3533) );
  OR3_X1 U2904 ( .A1(n2563), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2564) );
  XNOR2_X1 U2905 ( .A(n2551), .B(n2550), .ZN(n3374) );
  XNOR2_X1 U2906 ( .A(n2515), .B(n2514), .ZN(n3318) );
  NAND2_X1 U2907 ( .A1(n2235), .A2(IR_REG_1__SCAN_IN), .ZN(n2232) );
  NAND2_X1 U2908 ( .A1(n2651), .A2(IR_REG_1__SCAN_IN), .ZN(n2234) );
  NAND2_X1 U2909 ( .A1(n2222), .A2(n2221), .ZN(U3232) );
  NOR3_X1 U2910 ( .A1(n3269), .A2(n3268), .A3(n3267), .ZN(n2221) );
  NAND2_X1 U2911 ( .A1(n2223), .A2(n3981), .ZN(n2222) );
  AOI21_X1 U2912 ( .B1(n2251), .B2(n4184), .A(n2249), .ZN(n4198) );
  XNOR2_X1 U2913 ( .A(n2381), .B(n4203), .ZN(n4215) );
  INV_X1 U2914 ( .A(n2883), .ZN(n2884) );
  AOI211_X1 U2915 ( .C1(n4233), .C2(n4459), .A(n4232), .B(n4231), .ZN(n4234)
         );
  OR2_X1 U2916 ( .A1(n3230), .A2(n4609), .ZN(n3224) );
  OAI21_X1 U2917 ( .B1(n4620), .B2(n4754), .A(n2301), .ZN(U3545) );
  INV_X1 U2918 ( .A(n2302), .ZN(n2301) );
  OAI22_X1 U2919 ( .A1(n4623), .A2(n4609), .B1(n4756), .B2(n4513), .ZN(n2302)
         );
  OR2_X1 U2920 ( .A1(n4225), .A2(n4674), .ZN(n3211) );
  OR2_X1 U2921 ( .A1(n3715), .A2(n4149), .ZN(n2144) );
  NOR2_X2 U2922 ( .A1(n2507), .A2(n2506), .ZN(n2836) );
  AND2_X1 U2923 ( .A1(n3774), .A2(n4602), .ZN(n2145) );
  INV_X1 U2924 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3315) );
  AND2_X1 U2925 ( .A1(n2259), .A2(n2187), .ZN(n2146) );
  AND2_X1 U2926 ( .A1(n2931), .A2(n2248), .ZN(n2147) );
  AND2_X1 U2927 ( .A1(n2857), .A2(n2144), .ZN(n2148) );
  AND2_X1 U2928 ( .A1(n2146), .A2(REG3_REG_14__SCAN_IN), .ZN(n2149) );
  NAND2_X1 U2929 ( .A1(n2343), .A2(n2182), .ZN(n2150) );
  AND2_X1 U2930 ( .A1(n2145), .A2(n3946), .ZN(n2151) );
  AND3_X1 U2931 ( .A1(n4096), .A2(n4257), .A3(n2176), .ZN(n2152) );
  INV_X1 U2932 ( .A(n2415), .ZN(n2414) );
  NOR2_X1 U2933 ( .A1(n3057), .A2(n3942), .ZN(n2415) );
  AND2_X1 U2934 ( .A1(n4325), .A2(n2182), .ZN(n2153) );
  INV_X1 U2935 ( .A(n3552), .ZN(n2404) );
  AND2_X1 U2936 ( .A1(n2634), .A2(REG3_REG_19__SCAN_IN), .ZN(n2154) );
  OR2_X1 U2937 ( .A1(n5037), .A2(n4280), .ZN(n2155) );
  AND2_X1 U2938 ( .A1(n4280), .A2(n4298), .ZN(n2156) );
  AND2_X1 U2939 ( .A1(n2154), .A2(REG3_REG_20__SCAN_IN), .ZN(n2157) );
  AND2_X1 U2940 ( .A1(n2408), .A2(n4356), .ZN(n2158) );
  AND2_X1 U2941 ( .A1(n2158), .A2(n3266), .ZN(n2159) );
  AND2_X1 U2942 ( .A1(n2404), .A2(n2193), .ZN(n2160) );
  INV_X1 U2943 ( .A(n2519), .ZN(n2265) );
  XNOR2_X1 U2944 ( .A(n2761), .B(n2760), .ZN(n2879) );
  NAND2_X1 U2945 ( .A1(n2343), .A2(n2153), .ZN(n4344) );
  INV_X1 U2946 ( .A(n2400), .ZN(n2399) );
  NAND2_X1 U2947 ( .A1(n2626), .A2(n4036), .ZN(n2400) );
  OR2_X1 U2948 ( .A1(IR_REG_10__SCAN_IN), .A2(n2642), .ZN(n2161) );
  AOI21_X1 U2949 ( .B1(n2783), .B2(n4590), .A(n2782), .ZN(n3219) );
  NAND2_X1 U2950 ( .A1(n3133), .A2(n3132), .ZN(n3964) );
  NAND2_X1 U2951 ( .A1(n3087), .A2(n2444), .ZN(n3952) );
  AND2_X1 U2952 ( .A1(n2579), .A2(n2146), .ZN(n2162) );
  INV_X1 U2953 ( .A(n3474), .ZN(n3490) );
  INV_X1 U2954 ( .A(n3046), .ZN(n4602) );
  NAND2_X1 U2955 ( .A1(n2143), .A2(n2402), .ZN(n2770) );
  NAND2_X1 U2956 ( .A1(n3715), .A2(n4149), .ZN(n2163) );
  AND3_X1 U2957 ( .A1(n2462), .A2(n2470), .A3(n2771), .ZN(n2164) );
  AND2_X1 U2958 ( .A1(n2762), .A2(n2764), .ZN(n2166) );
  NAND2_X1 U2959 ( .A1(n2143), .A2(n2461), .ZN(n2803) );
  NOR2_X1 U2960 ( .A1(n4712), .A2(n2913), .ZN(n2167) );
  AND2_X1 U2961 ( .A1(n2401), .A2(n2399), .ZN(n2168) );
  AND2_X1 U2962 ( .A1(n4568), .A2(n4431), .ZN(n2169) );
  AND2_X1 U2963 ( .A1(n3024), .A2(n3023), .ZN(n2170) );
  NOR2_X1 U2964 ( .A1(n2447), .A2(n2446), .ZN(n2171) );
  NAND2_X1 U2965 ( .A1(n2143), .A2(n2762), .ZN(n2172) );
  AND2_X1 U2966 ( .A1(n3958), .A2(n4399), .ZN(n2173) );
  INV_X1 U2967 ( .A(IR_REG_31__SCAN_IN), .ZN(n2651) );
  AND2_X1 U2968 ( .A1(n4409), .A2(n4399), .ZN(n4375) );
  OR2_X1 U2969 ( .A1(n2540), .A2(REG1_REG_7__SCAN_IN), .ZN(n2174) );
  AND2_X1 U2970 ( .A1(n3592), .A2(n3553), .ZN(n2175) );
  NOR2_X1 U2971 ( .A1(n2297), .A2(n2386), .ZN(n2296) );
  AND2_X1 U2972 ( .A1(n2268), .A2(n4074), .ZN(n2176) );
  AND2_X1 U2973 ( .A1(n3039), .A2(n3034), .ZN(n2177) );
  INV_X1 U2974 ( .A(IR_REG_26__SCAN_IN), .ZN(n2462) );
  INV_X1 U2975 ( .A(n2548), .ZN(n2333) );
  INV_X1 U2976 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3373) );
  INV_X1 U2977 ( .A(IR_REG_28__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U2978 ( .A1(n4329), .A2(n4539), .ZN(n2179) );
  AND2_X1 U2979 ( .A1(n4148), .A2(n4507), .ZN(n2180) );
  AND2_X1 U2980 ( .A1(n3748), .A2(n2151), .ZN(n2181) );
  NAND2_X1 U2981 ( .A1(n4453), .A2(n2861), .ZN(n4427) );
  OR2_X1 U2982 ( .A1(n4329), .A2(n4539), .ZN(n2182) );
  NAND2_X1 U2983 ( .A1(n3113), .A2(n3898), .ZN(n2183) );
  OAI21_X1 U2984 ( .B1(n3579), .B2(n3580), .A(n3581), .ZN(n3682) );
  AND2_X1 U2985 ( .A1(n3102), .A2(n3101), .ZN(n2184) );
  NAND2_X1 U2986 ( .A1(n2418), .A2(n2417), .ZN(n3579) );
  NAND2_X1 U2987 ( .A1(n2215), .A2(n2216), .ZN(n3797) );
  NAND2_X1 U2988 ( .A1(n2411), .A2(n2414), .ZN(n3871) );
  NAND2_X1 U2989 ( .A1(n2419), .A2(n2423), .ZN(n3560) );
  OR2_X1 U2990 ( .A1(n4148), .A2(n4246), .ZN(n2185) );
  AND2_X1 U2991 ( .A1(n4508), .A2(n4260), .ZN(n2186) );
  NAND2_X1 U2992 ( .A1(n3035), .A2(n3034), .ZN(n3700) );
  INV_X1 U2993 ( .A(n3762), .ZN(n4588) );
  INV_X1 U2994 ( .A(IR_REG_11__SCAN_IN), .ZN(n2454) );
  AND2_X1 U2995 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2187) );
  AND2_X1 U2996 ( .A1(n4355), .A2(n4336), .ZN(n2188) );
  INV_X1 U2997 ( .A(n2319), .ZN(n2318) );
  NOR2_X1 U2998 ( .A1(n2442), .A2(n4685), .ZN(n2319) );
  OR2_X1 U2999 ( .A1(n2719), .A2(n4997), .ZN(n2189) );
  AND2_X1 U3000 ( .A1(n3064), .A2(n3063), .ZN(n3872) );
  INV_X1 U3001 ( .A(n4052), .ZN(n2398) );
  NOR2_X1 U3002 ( .A1(n4511), .A2(n4230), .ZN(n2371) );
  NAND2_X1 U3003 ( .A1(n4409), .A2(n2158), .ZN(n4335) );
  NAND2_X1 U3004 ( .A1(n4488), .A2(n4487), .ZN(n2190) );
  OR2_X1 U3005 ( .A1(n2442), .A2(n3792), .ZN(n2191) );
  INV_X1 U3006 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2245) );
  AND2_X1 U3007 ( .A1(n4055), .A2(n4051), .ZN(n4068) );
  INV_X1 U3008 ( .A(n4068), .ZN(n2363) );
  INV_X1 U3009 ( .A(n2155), .ZN(n2369) );
  INV_X1 U3010 ( .A(n4756), .ZN(n4754) );
  INV_X1 U3011 ( .A(n4703), .ZN(n4184) );
  AND2_X2 U3012 ( .A1(n3214), .A2(n3207), .ZN(n4751) );
  INV_X1 U3013 ( .A(n4751), .ZN(n4749) );
  NAND2_X1 U3014 ( .A1(n2290), .A2(n4022), .ZN(n3503) );
  INV_X1 U3015 ( .A(n4246), .ZN(n4507) );
  AND2_X1 U3016 ( .A1(n3061), .A2(n3062), .ZN(n2192) );
  NAND2_X1 U3017 ( .A1(n2770), .A2(n2464), .ZN(n2775) );
  NAND2_X1 U3018 ( .A1(n2428), .A2(n3003), .ZN(n3455) );
  AND2_X1 U3019 ( .A1(n3474), .A2(n3631), .ZN(n2193) );
  INV_X1 U3020 ( .A(n4266), .ZN(n4260) );
  AND2_X1 U3021 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2194) );
  AND2_X1 U3022 ( .A1(n2409), .A2(n4246), .ZN(n2195) );
  INV_X1 U3023 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U3024 ( .A1(n2766), .A2(n2765), .ZN(n2827) );
  INV_X1 U3025 ( .A(n2932), .ZN(n2248) );
  AND2_X1 U3026 ( .A1(n2326), .A2(n2325), .ZN(n2196) );
  INV_X1 U3027 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2256) );
  NAND2_X1 U3028 ( .A1(n2340), .A2(n2341), .ZN(n4313) );
  NAND2_X1 U3029 ( .A1(n2336), .A2(n2335), .ZN(n4408) );
  AOI21_X1 U3030 ( .B1(n4512), .B2(n4607), .A(n2304), .ZN(n2303) );
  NAND2_X2 U3031 ( .A1(n2971), .A2(n2972), .ZN(n2978) );
  OR2_X1 U3032 ( .A1(n2412), .A2(n3872), .ZN(n2220) );
  NAND2_X1 U3033 ( .A1(n3348), .A2(n2227), .ZN(n2226) );
  NAND3_X2 U3034 ( .A1(n2234), .A2(n2233), .A3(n2232), .ZN(n2928) );
  NAND3_X1 U3035 ( .A1(n2236), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2233) );
  INV_X2 U3036 ( .A(IR_REG_0__SCAN_IN), .ZN(n2235) );
  NAND2_X1 U3037 ( .A1(n3639), .A2(n2237), .ZN(n2240) );
  NAND2_X1 U3038 ( .A1(n2243), .A2(n2242), .ZN(n2241) );
  NAND3_X1 U3039 ( .A1(n2934), .A2(n2244), .A3(n2241), .ZN(n2935) );
  NAND2_X1 U3040 ( .A1(n3330), .A2(n2147), .ZN(n2246) );
  NAND3_X1 U3041 ( .A1(n3330), .A2(n2147), .A3(REG2_REG_3__SCAN_IN), .ZN(n2244) );
  NAND2_X1 U3042 ( .A1(n3330), .A2(n2931), .ZN(n2933) );
  NAND2_X1 U3043 ( .A1(n2744), .A2(n2830), .ZN(n4226) );
  NAND2_X1 U3044 ( .A1(n2710), .A2(REG3_REG_24__SCAN_IN), .ZN(n2719) );
  INV_X1 U3045 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2264) );
  NAND4_X1 U3046 ( .A1(n2265), .A2(REG3_REG_6__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .A4(REG3_REG_7__SCAN_IN), .ZN(n2557) );
  NAND3_X1 U3047 ( .A1(n4073), .A2(n2757), .A3(n2152), .ZN(n2267) );
  NAND2_X1 U3048 ( .A1(n3590), .A2(n2277), .ZN(n2275) );
  NAND2_X1 U3049 ( .A1(n3754), .A2(n2286), .ZN(n2284) );
  NAND2_X1 U3050 ( .A1(n2471), .A2(n2472), .ZN(n2773) );
  NAND3_X1 U3051 ( .A1(n2472), .A2(n2471), .A3(n2288), .ZN(n3847) );
  INV_X1 U3052 ( .A(n3391), .ZN(n2289) );
  NAND2_X1 U3053 ( .A1(n2289), .A2(n2296), .ZN(n2291) );
  NAND3_X1 U3054 ( .A1(n2291), .A2(n2292), .A3(n2294), .ZN(n2290) );
  NAND3_X1 U3055 ( .A1(n2294), .A2(n4007), .A3(n2291), .ZN(n3249) );
  NOR2_X1 U3056 ( .A1(n2525), .A2(n2293), .ZN(n2292) );
  NAND2_X1 U3057 ( .A1(n2295), .A2(n2296), .ZN(n2294) );
  INV_X1 U3058 ( .A(n4077), .ZN(n2295) );
  INV_X1 U3059 ( .A(n4002), .ZN(n2297) );
  NAND2_X1 U3060 ( .A1(n3390), .A2(n4002), .ZN(n3546) );
  NAND2_X1 U3061 ( .A1(n3391), .A2(n4077), .ZN(n3390) );
  NAND4_X1 U3062 ( .A1(n2178), .A2(n2298), .A3(n2299), .A4(n3437), .ZN(n2485)
         );
  OR2_X2 U3063 ( .A1(n4273), .A2(n4116), .ZN(n4256) );
  AOI21_X2 U3065 ( .B1(n3463), .B2(REG1_REG_8__SCAN_IN), .A(n2309), .ZN(n3531)
         );
  AND2_X1 U3066 ( .A1(n2310), .A2(n2943), .ZN(n2309) );
  XNOR2_X2 U3067 ( .A(n2310), .B(n3466), .ZN(n3463) );
  NAND2_X1 U3068 ( .A1(n3372), .A2(n2174), .ZN(n2311) );
  NAND2_X1 U3069 ( .A1(n4168), .A2(n2313), .ZN(n2312) );
  OAI211_X1 U3070 ( .C1(n4168), .C2(n2314), .A(n2312), .B(n2191), .ZN(n2905)
         );
  INV_X1 U3071 ( .A(n2905), .ZN(n3812) );
  NAND2_X1 U3072 ( .A1(n2892), .A2(n2323), .ZN(n2322) );
  INV_X1 U3073 ( .A(n2326), .ZN(n3349) );
  XNOR2_X2 U3074 ( .A(n2912), .B(n2911), .ZN(n4711) );
  INV_X1 U3075 ( .A(n2331), .ZN(n2332) );
  NAND3_X1 U3076 ( .A1(n2332), .A2(n2548), .A3(n2845), .ZN(n2842) );
  NAND2_X1 U3077 ( .A1(n4455), .A2(n2337), .ZN(n2336) );
  INV_X1 U3078 ( .A(n4349), .ZN(n2344) );
  NAND2_X1 U3079 ( .A1(n4349), .A2(n2153), .ZN(n2340) );
  NAND2_X1 U3080 ( .A1(n2864), .A2(n2347), .ZN(n2346) );
  INV_X1 U3081 ( .A(n3669), .ZN(n2354) );
  AOI21_X2 U3082 ( .B1(n2354), .B2(n2148), .A(n2350), .ZN(n3757) );
  NAND2_X1 U3083 ( .A1(n2875), .A2(n2356), .ZN(n2355) );
  NAND2_X1 U3084 ( .A1(n2368), .A2(n2367), .ZN(n2373) );
  AND2_X1 U3085 ( .A1(n2368), .A2(n2155), .ZN(n4253) );
  AND2_X2 U3086 ( .A1(n2373), .A2(n2372), .ZN(n4237) );
  INV_X1 U3087 ( .A(n2940), .ZN(n2375) );
  OAI21_X1 U3088 ( .B1(n3340), .B2(n2375), .A(n2374), .ZN(n3376) );
  NAND2_X1 U3089 ( .A1(n4256), .A2(n2394), .ZN(n2393) );
  NAND2_X1 U3090 ( .A1(n2403), .A2(n3474), .ZN(n3617) );
  OAI21_X2 U3091 ( .B1(n3906), .B2(n3084), .A(n3083), .ZN(n3087) );
  NAND2_X1 U3092 ( .A1(n3521), .A2(n2420), .ZN(n2418) );
  NAND2_X1 U3093 ( .A1(n3035), .A2(n2177), .ZN(n3702) );
  NAND2_X1 U3094 ( .A1(n3929), .A2(n2433), .ZN(n2431) );
  OR2_X1 U3095 ( .A1(n3929), .A2(n2435), .ZN(n2434) );
  NOR2_X1 U3096 ( .A1(n3929), .A2(n3933), .ZN(n3897) );
  INV_X1 U3097 ( .A(n3933), .ZN(n2436) );
  OR2_X1 U3098 ( .A1(n2518), .A2(n3243), .ZN(n2487) );
  NAND2_X2 U3099 ( .A1(n2609), .A2(n4041), .ZN(n3754) );
  OAI21_X1 U3100 ( .B1(REG1_REG_2__SCAN_IN), .B2(n3329), .A(n2888), .ZN(n3335)
         );
  NAND2_X1 U3101 ( .A1(n3329), .A2(REG1_REG_2__SCAN_IN), .ZN(n2888) );
  MUX2_X1 U3102 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2516), .Z(n3432) );
  NAND2_X1 U3103 ( .A1(n2516), .A2(DATAI_1_), .ZN(n2468) );
  INV_X1 U3104 ( .A(n2819), .ZN(n4678) );
  AOI21_X1 U3105 ( .B1(n3883), .B2(n3823), .A(n3822), .ZN(n3824) );
  NAND2_X1 U3106 ( .A1(n2821), .A2(n2796), .ZN(n2797) );
  NAND2_X1 U3107 ( .A1(n2971), .A2(n4729), .ZN(n3203) );
  INV_X1 U3108 ( .A(n3824), .ZN(n3850) );
  NAND2_X1 U3109 ( .A1(n2670), .A2(n2648), .ZN(n2672) );
  INV_X1 U3110 ( .A(n3974), .ZN(n3981) );
  AND2_X1 U3111 ( .A1(n2726), .A2(n2725), .ZN(n5037) );
  INV_X1 U3112 ( .A(n4545), .ZN(n4355) );
  AND2_X1 U3113 ( .A1(n2893), .A2(REG1_REG_5__SCAN_IN), .ZN(n2437) );
  AND4_X1 U3114 ( .A1(n2460), .A2(n2764), .A3(n2822), .A4(n2794), .ZN(n2438)
         );
  AND2_X1 U3115 ( .A1(n3158), .A2(n3981), .ZN(n2440) );
  AND2_X1 U3116 ( .A1(n2448), .A2(n2844), .ZN(n2441) );
  OR2_X1 U3117 ( .A1(n4171), .A2(n4940), .ZN(n2442) );
  NOR2_X1 U3118 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2443)
         );
  OR2_X1 U3119 ( .A1(n3086), .A2(n3085), .ZN(n2444) );
  INV_X1 U3120 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3227) );
  OR2_X1 U3121 ( .A1(n4229), .A2(n4544), .ZN(n2445) );
  AND2_X1 U3122 ( .A1(n4495), .A2(n4597), .ZN(n2446) );
  NOR2_X1 U3123 ( .A1(n2856), .A2(n4489), .ZN(n2447) );
  AND2_X1 U3124 ( .A1(n2841), .A2(n3504), .ZN(n2448) );
  INV_X1 U3125 ( .A(n3266), .ZN(n4336) );
  NAND2_X1 U3126 ( .A1(n3908), .A2(n3907), .ZN(n3073) );
  INV_X1 U3127 ( .A(n4104), .ZN(n2674) );
  INV_X1 U3128 ( .A(n3943), .ZN(n3057) );
  INV_X1 U3129 ( .A(n4061), .ZN(n2757) );
  AND2_X1 U3130 ( .A1(n3596), .A2(n3595), .ZN(n2846) );
  XNOR2_X1 U3131 ( .A(n2989), .B(n3142), .ZN(n2993) );
  NAND2_X1 U3132 ( .A1(n2842), .A2(n4012), .ZN(n2844) );
  NAND2_X1 U3133 ( .A1(n4007), .A2(n4003), .ZN(n3539) );
  INV_X1 U3134 ( .A(n2142), .ZN(n3145) );
  OAI22_X1 U3135 ( .A1(n3541), .A2(n3177), .B1(n3148), .B2(n3540), .ZN(n2999)
         );
  INV_X1 U3136 ( .A(n3131), .ZN(n3132) );
  NOR2_X1 U3137 ( .A1(n2541), .A2(n2505), .ZN(n2506) );
  INV_X1 U3138 ( .A(n3271), .ZN(n2475) );
  INV_X1 U3139 ( .A(n5037), .ZN(n4261) );
  AND2_X1 U3140 ( .A1(n4140), .A2(n2878), .ZN(n3153) );
  INV_X1 U3141 ( .A(n4679), .ZN(n2801) );
  INV_X1 U3142 ( .A(n2672), .ZN(n2653) );
  INV_X1 U3143 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3987) );
  AND2_X1 U3144 ( .A1(n2693), .A2(n2692), .ZN(n4545) );
  AND2_X1 U3145 ( .A1(n2891), .A2(n4689), .ZN(n2892) );
  INV_X1 U3146 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3773) );
  INV_X1 U3147 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4855) );
  AND2_X1 U31480 ( .A1(n2717), .A2(n2716), .ZN(n4312) );
  NAND2_X1 U31490 ( .A1(n3153), .A2(n4692), .ZN(n4544) );
  INV_X1 U3150 ( .A(n4149), .ZN(n3779) );
  INV_X1 U3151 ( .A(n4480), .ZN(n4599) );
  INV_X1 U3152 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3221) );
  INV_X1 U3153 ( .A(n3693), .ZN(n3659) );
  INV_X1 U3154 ( .A(n3715), .ZN(n3704) );
  INV_X1 U3155 ( .A(n4312), .ZN(n4518) );
  AND4_X1 U3156 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n3713)
         );
  INV_X1 U3157 ( .A(n4692), .ZN(n3302) );
  INV_X1 U3158 ( .A(n4199), .ZN(n4710) );
  INV_X1 U3159 ( .A(n4456), .ZN(n4501) );
  AND2_X1 U3160 ( .A1(n4002), .A2(n3999), .ZN(n4077) );
  AND2_X1 U3161 ( .A1(n4374), .A2(n4614), .ZN(n4744) );
  AND2_X1 U3162 ( .A1(n4718), .A2(n2975), .ZN(n4742) );
  NAND2_X1 U3163 ( .A1(n2806), .A2(n4678), .ZN(n3151) );
  XNOR2_X1 U3164 ( .A(n2554), .B(n2553), .ZN(n3466) );
  AND2_X1 U3165 ( .A1(n2922), .A2(n2921), .ZN(n4709) );
  OR2_X1 U3166 ( .A1(n3183), .A2(n3157), .ZN(n3974) );
  AND2_X1 U3167 ( .A1(n3178), .A2(n3422), .ZN(n3993) );
  NAND2_X1 U3168 ( .A1(n2641), .A2(n2640), .ZN(n4414) );
  OR2_X1 U3169 ( .A1(n3306), .A2(n3302), .ZN(n4715) );
  OR2_X1 U3170 ( .A1(n3306), .A2(n4138), .ZN(n4703) );
  NAND2_X1 U3171 ( .A1(n4724), .A2(n2881), .ZN(n4456) );
  OR2_X1 U3172 ( .A1(n4225), .A2(n4609), .ZN(n3217) );
  AND2_X2 U3173 ( .A1(n3214), .A2(n3213), .ZN(n4756) );
  OR2_X1 U3174 ( .A1(n3230), .A2(n4674), .ZN(n3231) );
  INV_X1 U3175 ( .A(n4728), .ZN(n4727) );
  AND2_X1 U3176 ( .A1(n3172), .A2(STATE_REG_SCAN_IN), .ZN(n4729) );
  INV_X1 U3177 ( .A(n2911), .ZN(n4733) );
  OR2_X1 U3178 ( .A1(n2969), .A2(n2968), .ZN(U3258) );
  NAND2_X1 U3179 ( .A1(n2770), .A2(IR_REG_31__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3180 ( .A1(n2463), .A2(n2470), .ZN(n2776) );
  NAND2_X1 U3181 ( .A1(n2776), .A2(n2771), .ZN(n2466) );
  NAND2_X1 U3182 ( .A1(n2775), .A2(IR_REG_28__SCAN_IN), .ZN(n2465) );
  NAND2_X2 U3183 ( .A1(n2466), .A2(n2465), .ZN(n2516) );
  INV_X1 U3184 ( .A(n2516), .ZN(n2467) );
  NAND2_X1 U3185 ( .A1(n2467), .A2(n2928), .ZN(n2469) );
  NAND2_X2 U3186 ( .A1(n2469), .A2(n2468), .ZN(n3437) );
  XNOR2_X2 U3187 ( .A(n2473), .B(IR_REG_29__SCAN_IN), .ZN(n3271) );
  INV_X1 U3188 ( .A(n2541), .ZN(n2474) );
  NAND2_X1 U3189 ( .A1(n2474), .A2(REG2_REG_1__SCAN_IN), .ZN(n2478) );
  INV_X1 U3190 ( .A(n3278), .ZN(n2476) );
  NAND2_X1 U3191 ( .A1(n2501), .A2(REG3_REG_1__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3192 ( .A1(n3571), .A2(n4153), .ZN(n3994) );
  NAND2_X1 U3193 ( .A1(n3994), .A2(n2485), .ZN(n3400) );
  INV_X1 U3194 ( .A(n3400), .ZN(n2484) );
  INV_X1 U3195 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3434) );
  OR2_X1 U3196 ( .A1(n2518), .A2(n3434), .ZN(n2483) );
  INV_X1 U3197 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3198 ( .A1(n2544), .A2(REG0_REG_0__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3199 ( .A1(n2545), .A2(REG1_REG_0__SCAN_IN), .ZN(n2480) );
  NOR2_X2 U3200 ( .A1(n3364), .A2(n4154), .ZN(n3996) );
  NAND2_X1 U3201 ( .A1(n2484), .A2(n3996), .ZN(n3405) );
  NAND2_X1 U3202 ( .A1(n3405), .A2(n2485), .ZN(n3235) );
  NAND2_X1 U3203 ( .A1(n2545), .A2(REG1_REG_2__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3204 ( .A1(n2544), .A2(REG0_REG_2__SCAN_IN), .ZN(n2488) );
  INV_X1 U3205 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U3206 ( .A1(n2474), .A2(REG2_REG_2__SCAN_IN), .ZN(n2486) );
  INV_X1 U3207 ( .A(n3573), .ZN(n3392) );
  NOR2_X1 U3208 ( .A1(n2490), .A2(n2791), .ZN(n2491) );
  INV_X1 U3209 ( .A(DATAI_2_), .ZN(n4779) );
  MUX2_X1 U32100 ( .A(n3329), .B(n4779), .S(n2516), .Z(n2990) );
  INV_X1 U32110 ( .A(n2990), .ZN(n3446) );
  NAND2_X1 U32120 ( .A1(n3446), .A2(n3573), .ZN(n3997) );
  AND2_X2 U32130 ( .A1(n4000), .A2(n3997), .ZN(n4078) );
  NAND2_X1 U32140 ( .A1(n3235), .A2(n4078), .ZN(n3234) );
  NAND2_X1 U32150 ( .A1(n3234), .A2(n3997), .ZN(n3391) );
  NAND2_X1 U32160 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2508) );
  XNOR2_X1 U32170 ( .A(n2508), .B(n2511), .ZN(n2932) );
  INV_X1 U32180 ( .A(DATAI_3_), .ZN(n2495) );
  MUX2_X1 U32190 ( .A(n2932), .B(n2495), .S(n2516), .Z(n3540) );
  INV_X1 U32200 ( .A(n3540), .ZN(n3647) );
  NAND2_X1 U32210 ( .A1(n2544), .A2(REG0_REG_3__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U32220 ( .A1(n2545), .A2(REG1_REG_3__SCAN_IN), .ZN(n2498) );
  OR2_X1 U32230 ( .A1(n2518), .A2(REG3_REG_3__SCAN_IN), .ZN(n2497) );
  OR2_X1 U32240 ( .A1(n2541), .A2(n2245), .ZN(n2496) );
  AND4_X2 U32250 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n3541)
         );
  NAND2_X1 U32260 ( .A1(n3647), .A2(n3541), .ZN(n4002) );
  INV_X1 U32270 ( .A(n3541), .ZN(n3547) );
  NAND2_X1 U32280 ( .A1(n3540), .A2(n3547), .ZN(n3999) );
  NAND2_X1 U32290 ( .A1(n2545), .A2(REG1_REG_4__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32300 ( .A1(n2544), .A2(REG0_REG_4__SCAN_IN), .ZN(n2503) );
  OAI21_X1 U32310 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2519), .ZN(n3555) );
  INV_X1 U32320 ( .A(n3555), .ZN(n2500) );
  NAND2_X1 U32330 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NAND3_X1 U32340 ( .A1(n2504), .A2(n2503), .A3(n2502), .ZN(n2507) );
  INV_X1 U32350 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32360 ( .A1(n2508), .A2(n2511), .ZN(n2509) );
  NAND2_X1 U32370 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2510) );
  XNOR2_X1 U32380 ( .A(n2510), .B(IR_REG_4__SCAN_IN), .ZN(n4689) );
  MUX2_X1 U32390 ( .A(n4689), .B(DATAI_4_), .S(n2516), .Z(n3005) );
  NAND2_X1 U32400 ( .A1(n2836), .A2(n3005), .ZN(n4003) );
  NAND2_X2 U32410 ( .A1(n4152), .A2(n3553), .ZN(n4007) );
  NAND2_X1 U32420 ( .A1(n2511), .A2(n4785), .ZN(n2512) );
  NAND2_X1 U32430 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2515) );
  INV_X1 U32440 ( .A(DATAI_5_), .ZN(n2517) );
  MUX2_X1 U32450 ( .A(n3318), .B(n2517), .S(n2555), .Z(n3474) );
  NAND2_X1 U32460 ( .A1(n2544), .A2(REG0_REG_5__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32470 ( .A1(n3834), .A2(REG1_REG_5__SCAN_IN), .ZN(n2523) );
  AND2_X1 U32480 ( .A1(n2519), .A2(n3315), .ZN(n2520) );
  OR2_X1 U32490 ( .A1(n2520), .A2(n2529), .ZN(n3479) );
  OR2_X1 U32500 ( .A1(n2750), .A2(n3479), .ZN(n2522) );
  INV_X1 U32510 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2937) );
  OR2_X1 U32520 ( .A1(n3837), .A2(n2937), .ZN(n2521) );
  AND4_X2 U32530 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n3630)
         );
  NAND2_X1 U32540 ( .A1(n3474), .A2(n4151), .ZN(n4005) );
  INV_X1 U32550 ( .A(n4005), .ZN(n2525) );
  NAND2_X1 U32560 ( .A1(n3490), .A2(n3630), .ZN(n4022) );
  INV_X1 U32570 ( .A(n2537), .ZN(n2527) );
  NAND2_X1 U32580 ( .A1(n2527), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  XNOR2_X1 U32590 ( .A(n2528), .B(IR_REG_6__SCAN_IN), .ZN(n4688) );
  MUX2_X1 U32600 ( .A(n4688), .B(DATAI_6_), .S(n2555), .Z(n3595) );
  INV_X1 U32610 ( .A(n3595), .ZN(n3631) );
  INV_X1 U32620 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3626) );
  OR2_X1 U32630 ( .A1(n2529), .A2(REG3_REG_6__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32640 ( .A1(n2542), .A2(n2530), .ZN(n3625) );
  OR2_X1 U32650 ( .A1(n2750), .A2(n3625), .ZN(n2533) );
  NAND2_X1 U32660 ( .A1(n2544), .A2(REG0_REG_6__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32670 ( .A1(n3834), .A2(REG1_REG_6__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32680 ( .A1(n3631), .A2(n3596), .ZN(n4021) );
  NAND2_X1 U32690 ( .A1(n3503), .A2(n4021), .ZN(n2535) );
  NAND2_X1 U32700 ( .A1(n3595), .A2(n3599), .ZN(n4008) );
  NAND2_X1 U32710 ( .A1(n2535), .A2(n4008), .ZN(n3590) );
  INV_X1 U32720 ( .A(IR_REG_6__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32730 ( .A1(n2537), .A2(n2536), .ZN(n2563) );
  NAND2_X1 U32740 ( .A1(n2563), .A2(IR_REG_31__SCAN_IN), .ZN(n2551) );
  INV_X1 U32750 ( .A(DATAI_7_), .ZN(n2538) );
  INV_X1 U32760 ( .A(n3592), .ZN(n2845) );
  INV_X1 U32770 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2941) );
  OR2_X1 U32780 ( .A1(n2541), .A2(n2941), .ZN(n2548) );
  NAND2_X1 U32790 ( .A1(n2542), .A2(n3373), .ZN(n2543) );
  NAND2_X1 U32800 ( .A1(n2557), .A2(n2543), .ZN(n3603) );
  NAND2_X1 U32810 ( .A1(n2544), .A2(REG0_REG_7__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32820 ( .A1(n2545), .A2(REG1_REG_7__SCAN_IN), .ZN(n2546) );
  INV_X1 U32830 ( .A(n2842), .ZN(n2549) );
  NAND2_X1 U32840 ( .A1(n3592), .A2(n3525), .ZN(n4012) );
  NAND2_X1 U32850 ( .A1(n2551), .A2(n2550), .ZN(n2552) );
  NAND2_X1 U32860 ( .A1(n2552), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  INV_X1 U32870 ( .A(IR_REG_8__SCAN_IN), .ZN(n2553) );
  INV_X1 U32880 ( .A(DATAI_8_), .ZN(n3274) );
  MUX2_X1 U32890 ( .A(n3466), .B(n3274), .S(n3832), .Z(n3585) );
  NAND2_X1 U32900 ( .A1(n3833), .A2(REG0_REG_8__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32910 ( .A1(n3834), .A2(REG1_REG_8__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32920 ( .A1(n2557), .A2(n2556), .ZN(n2558) );
  NAND2_X1 U32930 ( .A1(n2568), .A2(n2558), .ZN(n3614) );
  OR2_X1 U32940 ( .A1(n2750), .A2(n3614), .ZN(n2560) );
  INV_X1 U32950 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3615) );
  OR2_X1 U32960 ( .A1(n3837), .A2(n3615), .ZN(n2559) );
  NAND2_X1 U32970 ( .A1(n3616), .A2(n3685), .ZN(n4013) );
  NAND2_X1 U32980 ( .A1(n3585), .A2(n3691), .ZN(n4011) );
  NAND2_X1 U32990 ( .A1(n2564), .A2(IR_REG_31__SCAN_IN), .ZN(n2566) );
  INV_X1 U33000 ( .A(IR_REG_9__SCAN_IN), .ZN(n2565) );
  INV_X1 U33010 ( .A(DATAI_9_), .ZN(n2567) );
  MUX2_X1 U33020 ( .A(n3533), .B(n2567), .S(n3832), .Z(n3693) );
  NAND2_X1 U33030 ( .A1(n3833), .A2(REG0_REG_9__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33040 ( .A1(n3834), .A2(REG1_REG_9__SCAN_IN), .ZN(n2573) );
  INV_X1 U33050 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3661) );
  OR2_X1 U33060 ( .A1(n3837), .A2(n3661), .ZN(n2572) );
  INV_X1 U33070 ( .A(n2579), .ZN(n2570) );
  NAND2_X1 U33080 ( .A1(n2568), .A2(n4823), .ZN(n2569) );
  NAND2_X1 U33090 ( .A1(n2570), .A2(n2569), .ZN(n3690) );
  OR2_X1 U33100 ( .A1(n2750), .A2(n3690), .ZN(n2571) );
  INV_X1 U33110 ( .A(n3713), .ZN(n4150) );
  NAND2_X1 U33120 ( .A1(n3693), .A2(n4150), .ZN(n4020) );
  NAND2_X1 U33130 ( .A1(n3659), .A2(n3713), .ZN(n4014) );
  NAND2_X1 U33140 ( .A1(n2575), .A2(IR_REG_31__SCAN_IN), .ZN(n2576) );
  MUX2_X1 U33150 ( .A(IR_REG_31__SCAN_IN), .B(n2576), .S(IR_REG_10__SCAN_IN), 
        .Z(n2578) );
  NOR2_X1 U33160 ( .A1(n2575), .A2(IR_REG_10__SCAN_IN), .ZN(n2586) );
  INV_X1 U33170 ( .A(n2586), .ZN(n2577) );
  NAND2_X1 U33180 ( .A1(n2578), .A2(n2577), .ZN(n3641) );
  MUX2_X1 U33190 ( .A(n4687), .B(DATAI_10_), .S(n3832), .Z(n3715) );
  OR2_X1 U33200 ( .A1(n2579), .A2(REG3_REG_10__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U33210 ( .A1(n2587), .A2(n2580), .ZN(n3709) );
  OR2_X1 U33220 ( .A1(n2750), .A2(n3709), .ZN(n2584) );
  INV_X1 U33230 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3673) );
  OR2_X1 U33240 ( .A1(n3837), .A2(n3673), .ZN(n2583) );
  NAND2_X1 U33250 ( .A1(n3833), .A2(REG0_REG_10__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33260 ( .A1(n3834), .A2(REG1_REG_10__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33270 ( .A1(n3704), .A2(n4149), .ZN(n4030) );
  NAND2_X1 U33280 ( .A1(n3668), .A2(n4030), .ZN(n2585) );
  NAND2_X1 U33290 ( .A1(n3715), .A2(n3779), .ZN(n4026) );
  NAND2_X1 U33300 ( .A1(n2585), .A2(n4026), .ZN(n3740) );
  XNOR2_X1 U33310 ( .A(n2594), .B(IR_REG_11__SCAN_IN), .ZN(n4686) );
  MUX2_X1 U33320 ( .A(n4686), .B(DATAI_11_), .S(n3832), .Z(n3043) );
  NAND2_X1 U33330 ( .A1(n3833), .A2(REG0_REG_11__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33340 ( .A1(n3834), .A2(REG1_REG_11__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U33350 ( .A1(n2587), .A2(n3773), .ZN(n2588) );
  NAND2_X1 U33360 ( .A1(n2603), .A2(n2588), .ZN(n3778) );
  OR2_X1 U33370 ( .A1(n2750), .A2(n3778), .ZN(n2590) );
  INV_X1 U33380 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3746) );
  OR2_X1 U33390 ( .A1(n3837), .A2(n3746), .ZN(n2589) );
  INV_X1 U33400 ( .A(n3732), .ZN(n4600) );
  NAND2_X1 U33410 ( .A1(n3774), .A2(n4600), .ZN(n4031) );
  NAND2_X1 U33420 ( .A1(n3740), .A2(n4031), .ZN(n2593) );
  NAND2_X1 U33430 ( .A1(n3043), .A2(n3732), .ZN(n4035) );
  NAND2_X1 U33440 ( .A1(n2593), .A2(n4035), .ZN(n3726) );
  NAND2_X1 U33450 ( .A1(n2594), .A2(n2454), .ZN(n2595) );
  NAND2_X1 U33460 ( .A1(n2595), .A2(IR_REG_31__SCAN_IN), .ZN(n2596) );
  XNOR2_X1 U33470 ( .A(n2596), .B(IR_REG_12__SCAN_IN), .ZN(n4685) );
  MUX2_X1 U33480 ( .A(n4685), .B(DATAI_12_), .S(n3832), .Z(n3046) );
  INV_X1 U33490 ( .A(REG3_REG_12__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U33500 ( .A(n2603), .B(n5035), .ZN(n3808) );
  OR2_X1 U33510 ( .A1(n3808), .A2(n2750), .ZN(n2600) );
  INV_X1 U33520 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3789) );
  OR2_X1 U3353 ( .A1(n3837), .A2(n3789), .ZN(n2599) );
  NAND2_X1 U33540 ( .A1(n3833), .A2(REG0_REG_12__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3355 ( .A1(n3834), .A2(REG1_REG_12__SCAN_IN), .ZN(n2597) );
  NAND4_X1 U3356 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n3949)
         );
  NAND2_X1 U3357 ( .A1(n4602), .A2(n3949), .ZN(n4477) );
  OR2_X1 U3358 ( .A1(n2143), .A2(n2791), .ZN(n2601) );
  XNOR2_X1 U3359 ( .A(n2601), .B(IR_REG_13__SCAN_IN), .ZN(n4684) );
  MUX2_X1 U3360 ( .A(n4684), .B(DATAI_13_), .S(n3832), .Z(n4495) );
  INV_X1 U3361 ( .A(n4495), .ZN(n3946) );
  INV_X1 U3362 ( .A(n2603), .ZN(n2602) );
  AOI21_X1 U3363 ( .B1(n2602), .B2(REG3_REG_12__SCAN_IN), .A(
        REG3_REG_13__SCAN_IN), .ZN(n2604) );
  OR2_X1 U3364 ( .A1(n2604), .A2(n2162), .ZN(n4493) );
  INV_X1 U3365 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4494) );
  OAI22_X1 U3366 ( .A1(n2750), .A2(n4493), .B1(n3837), .B2(n4494), .ZN(n2608)
         );
  NAND2_X1 U3367 ( .A1(n3833), .A2(REG0_REG_13__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U3368 ( .A1(n3834), .A2(REG1_REG_13__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U3369 ( .A1(n2606), .A2(n2605), .ZN(n2607) );
  NAND2_X1 U3370 ( .A1(n3946), .A2(n4597), .ZN(n4070) );
  NAND2_X1 U3371 ( .A1(n3726), .A2(n4038), .ZN(n2609) );
  NOR2_X1 U3372 ( .A1(n4602), .A2(n3949), .ZN(n4478) );
  NOR2_X1 U3373 ( .A1(n4597), .A2(n3946), .ZN(n4069) );
  AOI21_X1 U3374 ( .B1(n4038), .B2(n4478), .A(n4069), .ZN(n4041) );
  OR2_X1 U3375 ( .A1(n2162), .A2(REG3_REG_14__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U3376 ( .A1(n2617), .A2(n2610), .ZN(n3879) );
  INV_X1 U3377 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3759) );
  OAI22_X1 U3378 ( .A1(n3879), .A2(n2750), .B1(n3837), .B2(n3759), .ZN(n2614)
         );
  NAND2_X1 U3379 ( .A1(n3833), .A2(REG0_REG_14__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U3380 ( .A1(n3834), .A2(REG1_REG_14__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3381 ( .A1(n2612), .A2(n2611), .ZN(n2613) );
  INV_X1 U3382 ( .A(IR_REG_13__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3383 ( .A1(n2143), .A2(n2615), .ZN(n2621) );
  NAND2_X1 U3384 ( .A1(n2621), .A2(IR_REG_31__SCAN_IN), .ZN(n2616) );
  XNOR2_X1 U3385 ( .A(n2616), .B(IR_REG_14__SCAN_IN), .ZN(n4683) );
  MUX2_X1 U3386 ( .A(n4683), .B(DATAI_14_), .S(n3832), .Z(n3762) );
  NAND2_X1 U3387 ( .A1(n4482), .A2(n3762), .ZN(n4036) );
  NAND2_X1 U3388 ( .A1(n4588), .A2(n4576), .ZN(n4016) );
  NAND2_X1 U3389 ( .A1(n4036), .A2(n4016), .ZN(n3756) );
  INV_X1 U3390 ( .A(n3756), .ZN(n4079) );
  NAND2_X1 U3391 ( .A1(n2617), .A2(n3987), .ZN(n2618) );
  NAND2_X1 U3392 ( .A1(n2627), .A2(n2618), .ZN(n4466) );
  INV_X1 U3393 ( .A(n3837), .ZN(n2629) );
  AOI22_X1 U3394 ( .A1(n2629), .A2(REG2_REG_15__SCAN_IN), .B1(n3833), .B2(
        REG0_REG_15__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U3395 ( .A1(n3834), .A2(REG1_REG_15__SCAN_IN), .ZN(n2619) );
  INV_X1 U3396 ( .A(n4585), .ZN(n3875) );
  NAND2_X1 U3397 ( .A1(n2622), .A2(IR_REG_31__SCAN_IN), .ZN(n2624) );
  INV_X1 U3398 ( .A(n2624), .ZN(n2623) );
  NAND2_X1 U3399 ( .A1(n2623), .A2(IR_REG_15__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3400 ( .A1(n2624), .A2(n2643), .ZN(n2632) );
  MUX2_X1 U3401 ( .A(n2962), .B(DATAI_15_), .S(n3832), .Z(n3069) );
  NAND2_X1 U3402 ( .A1(n3875), .A2(n3069), .ZN(n4037) );
  NAND2_X1 U3403 ( .A1(n4585), .A2(n4579), .ZN(n4017) );
  NAND2_X1 U3404 ( .A1(n4037), .A2(n4017), .ZN(n4462) );
  AND2_X1 U3405 ( .A1(n2627), .A2(n4855), .ZN(n2628) );
  OR2_X1 U3406 ( .A1(n2628), .A2(n2664), .ZN(n4447) );
  AOI22_X1 U3407 ( .A1(n2629), .A2(REG2_REG_16__SCAN_IN), .B1(n3833), .B2(
        REG0_REG_16__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3408 ( .A1(n3834), .A2(REG1_REG_16__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3409 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  XNOR2_X1 U3410 ( .A(n2633), .B(IR_REG_16__SCAN_IN), .ZN(n2911) );
  INV_X1 U3411 ( .A(DATAI_16_), .ZN(n4910) );
  MUX2_X1 U3412 ( .A(n4733), .B(n4910), .S(n3832), .Z(n4570) );
  NAND2_X1 U3413 ( .A1(n4577), .A2(n4570), .ZN(n4103) );
  OR2_X1 U3414 ( .A1(n4577), .A2(n4570), .ZN(n4106) );
  NAND2_X1 U3415 ( .A1(n4103), .A2(n4106), .ZN(n4454) );
  INV_X1 U3416 ( .A(n4454), .ZN(n4441) );
  INV_X1 U3417 ( .A(n4425), .ZN(n2675) );
  AND2_X1 U3418 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2634) );
  OR2_X1 U3419 ( .A1(n2657), .A2(REG3_REG_19__SCAN_IN), .ZN(n2635) );
  AND2_X1 U3420 ( .A1(n2678), .A2(n2635), .ZN(n4401) );
  NAND2_X1 U3421 ( .A1(n4401), .A2(n2501), .ZN(n2641) );
  INV_X1 U3422 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3423 ( .A1(n3834), .A2(REG1_REG_19__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U3424 ( .A1(n3833), .A2(REG0_REG_19__SCAN_IN), .ZN(n2636) );
  OAI211_X1 U3425 ( .C1(n3837), .C2(n2638), .A(n2637), .B(n2636), .ZN(n2639)
         );
  INV_X1 U3426 ( .A(n2639), .ZN(n2640) );
  NOR2_X1 U3427 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2645)
         );
  NOR2_X1 U3428 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2644)
         );
  NAND4_X1 U3429 ( .A1(n2646), .A2(n2645), .A3(n2644), .A4(n2643), .ZN(n2647)
         );
  NOR2_X1 U3430 ( .A1(n2650), .A2(n2443), .ZN(n2759) );
  NAND2_X1 U3431 ( .A1(n2654), .A2(IR_REG_19__SCAN_IN), .ZN(n2655) );
  MUX2_X1 U3432 ( .A(n4681), .B(DATAI_19_), .S(n3832), .Z(n4393) );
  NAND2_X1 U3433 ( .A1(n4414), .A2(n4399), .ZN(n4064) );
  AOI21_X1 U3434 ( .B1(n2664), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n2656) );
  OR2_X1 U3435 ( .A1(n2657), .A2(n2656), .ZN(n4421) );
  INV_X1 U3436 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3437 ( .A1(n3833), .A2(REG0_REG_18__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3438 ( .A1(n3834), .A2(REG1_REG_18__SCAN_IN), .ZN(n2658) );
  OAI211_X1 U3439 ( .C1(n2660), .C2(n3837), .A(n2659), .B(n2658), .ZN(n2661)
         );
  INV_X1 U3440 ( .A(n2661), .ZN(n2662) );
  NAND2_X1 U3441 ( .A1(n2672), .A2(IR_REG_31__SCAN_IN), .ZN(n2663) );
  XNOR2_X1 U3442 ( .A(n2663), .B(IR_REG_18__SCAN_IN), .ZN(n4202) );
  INV_X1 U3443 ( .A(DATAI_18_), .ZN(n4731) );
  MUX2_X1 U3444 ( .A(n4732), .B(n4731), .S(n3832), .Z(n4417) );
  NAND2_X1 U3445 ( .A1(n4561), .A2(n4417), .ZN(n4389) );
  NAND2_X1 U3446 ( .A1(n4064), .A2(n4389), .ZN(n2677) );
  INV_X1 U3447 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4822) );
  XNOR2_X1 U3448 ( .A(n2664), .B(n4822), .ZN(n4432) );
  NAND2_X1 U3449 ( .A1(n4432), .A2(n2501), .ZN(n2669) );
  INV_X1 U3450 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U3451 ( .A1(n3833), .A2(REG0_REG_17__SCAN_IN), .ZN(n2666) );
  NAND2_X1 U3452 ( .A1(n3834), .A2(REG1_REG_17__SCAN_IN), .ZN(n2665) );
  OAI211_X1 U3453 ( .C1(n2965), .C2(n3837), .A(n2666), .B(n2665), .ZN(n2667)
         );
  INV_X1 U3454 ( .A(n2667), .ZN(n2668) );
  NOR2_X1 U3455 ( .A1(n2670), .A2(n2791), .ZN(n2671) );
  MUX2_X1 U3456 ( .A(n2791), .B(n2671), .S(IR_REG_17__SCAN_IN), .Z(n2673) );
  NOR2_X1 U3457 ( .A1(n2673), .A2(n2653), .ZN(n4682) );
  MUX2_X1 U34580 ( .A(n4682), .B(DATAI_17_), .S(n3832), .Z(n4431) );
  INV_X1 U34590 ( .A(n4431), .ZN(n4563) );
  AND2_X1 U3460 ( .A1(n4568), .A2(n4563), .ZN(n4387) );
  NAND2_X1 U3461 ( .A1(n2675), .A2(n2674), .ZN(n4365) );
  OR2_X1 U3462 ( .A1(n4561), .A2(n4417), .ZN(n4388) );
  OR2_X1 U3463 ( .A1(n4568), .A2(n4563), .ZN(n4386) );
  AND2_X1 U3464 ( .A1(n4388), .A2(n4386), .ZN(n2676) );
  NAND2_X1 U3465 ( .A1(n3958), .A2(n4393), .ZN(n4065) );
  OAI21_X1 U3466 ( .B1(n2677), .B2(n2676), .A(n4065), .ZN(n4363) );
  INV_X1 U34670 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3936) );
  NAND2_X1 U3468 ( .A1(n2678), .A2(n3936), .ZN(n2679) );
  NAND2_X1 U34690 ( .A1(n2694), .A2(n2679), .ZN(n4379) );
  OR2_X1 U3470 ( .A1(n4379), .A2(n2750), .ZN(n2684) );
  INV_X1 U34710 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U3472 ( .A1(n3834), .A2(REG1_REG_20__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U34730 ( .A1(n3833), .A2(REG0_REG_20__SCAN_IN), .ZN(n2680) );
  OAI211_X1 U3474 ( .C1(n3837), .C2(n4380), .A(n2681), .B(n2680), .ZN(n2682)
         );
  INV_X1 U34750 ( .A(n2682), .ZN(n2683) );
  NOR2_X1 U3476 ( .A1(n4541), .A2(n4376), .ZN(n2685) );
  INV_X1 U34770 ( .A(n4109), .ZN(n2686) );
  NAND2_X1 U3478 ( .A1(n4365), .A2(n2686), .ZN(n2687) );
  NAND2_X1 U34790 ( .A1(n4541), .A2(n4376), .ZN(n4108) );
  NAND2_X1 U3480 ( .A1(n2687), .A2(n4108), .ZN(n4304) );
  INV_X1 U34810 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3901) );
  INV_X1 U3482 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3265) );
  OAI21_X1 U34830 ( .B1(n2694), .B2(n3901), .A(n3265), .ZN(n2688) );
  AND2_X1 U3484 ( .A1(n2700), .A2(n2688), .ZN(n3264) );
  NAND2_X1 U34850 ( .A1(n3264), .A2(n2501), .ZN(n2693) );
  INV_X1 U3486 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U34870 ( .A1(n3833), .A2(REG0_REG_22__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3488 ( .A1(n3834), .A2(REG1_REG_22__SCAN_IN), .ZN(n2689) );
  OAI211_X1 U34890 ( .C1(n4340), .C2(n3837), .A(n2690), .B(n2689), .ZN(n2691)
         );
  INV_X1 U3490 ( .A(n2691), .ZN(n2692) );
  NAND2_X1 U34910 ( .A1(n3832), .A2(DATAI_22_), .ZN(n3266) );
  NAND2_X1 U3492 ( .A1(n4545), .A2(n4336), .ZN(n4306) );
  XNOR2_X1 U34930 ( .A(n2694), .B(REG3_REG_21__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U3494 ( .A1(n4351), .A2(n2501), .ZN(n2699) );
  INV_X1 U34950 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U3496 ( .A1(n3834), .A2(REG1_REG_21__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U34970 ( .A1(n3833), .A2(REG0_REG_21__SCAN_IN), .ZN(n2695) );
  OAI211_X1 U3498 ( .C1(n3837), .C2(n4353), .A(n2696), .B(n2695), .ZN(n2697)
         );
  INV_X1 U34990 ( .A(n2697), .ZN(n2698) );
  OR2_X1 U3500 ( .A1(n4329), .A2(n4356), .ZN(n4324) );
  AND2_X1 U35010 ( .A1(n4306), .A2(n4324), .ZN(n4111) );
  NAND2_X1 U3502 ( .A1(n4304), .A2(n4111), .ZN(n2709) );
  INV_X1 U35030 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3885) );
  INV_X1 U3504 ( .A(n2710), .ZN(n2702) );
  NAND2_X1 U35050 ( .A1(n2700), .A2(n3885), .ZN(n2701) );
  NAND2_X1 U35060 ( .A1(n2702), .A2(n2701), .ZN(n4319) );
  OR2_X1 U35070 ( .A1(n4319), .A2(n2750), .ZN(n2707) );
  INV_X1 U35080 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U35090 ( .A1(n3833), .A2(REG0_REG_23__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U35100 ( .A1(n3834), .A2(REG1_REG_23__SCAN_IN), .ZN(n2703) );
  OAI211_X1 U35110 ( .C1(n4318), .C2(n3837), .A(n2704), .B(n2703), .ZN(n2705)
         );
  INV_X1 U35120 ( .A(n2705), .ZN(n2706) );
  NAND2_X1 U35130 ( .A1(n3832), .A2(DATAI_23_), .ZN(n3886) );
  NAND2_X1 U35140 ( .A1(n4293), .A2(n3886), .ZN(n4063) );
  NAND2_X1 U35150 ( .A1(n4355), .A2(n3266), .ZN(n2869) );
  NAND2_X1 U35160 ( .A1(n4063), .A2(n2869), .ZN(n4113) );
  AND2_X1 U35170 ( .A1(n4329), .A2(n4356), .ZN(n4305) );
  AND2_X1 U35180 ( .A1(n4306), .A2(n4305), .ZN(n4114) );
  NOR2_X1 U35190 ( .A1(n4113), .A2(n4114), .ZN(n2708) );
  NAND2_X1 U35200 ( .A1(n2709), .A2(n2708), .ZN(n4287) );
  OR2_X1 U35210 ( .A1(n2710), .A2(REG3_REG_24__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U35220 ( .A1(n4299), .A2(n2501), .ZN(n2717) );
  INV_X1 U35230 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U35240 ( .A1(n3834), .A2(REG1_REG_24__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U35250 ( .A1(n3833), .A2(REG0_REG_24__SCAN_IN), .ZN(n2712) );
  OAI211_X1 U35260 ( .C1(n3837), .C2(n2714), .A(n2713), .B(n2712), .ZN(n2715)
         );
  INV_X1 U35270 ( .A(n2715), .ZN(n2716) );
  NAND2_X1 U35280 ( .A1(n3832), .A2(DATAI_24_), .ZN(n4298) );
  INV_X1 U35290 ( .A(n4298), .ZN(n4292) );
  NAND2_X1 U35300 ( .A1(n4312), .A2(n4292), .ZN(n4076) );
  OR2_X1 U35310 ( .A1(n4293), .A2(n3886), .ZN(n4288) );
  AND2_X1 U35320 ( .A1(n4076), .A2(n4288), .ZN(n4048) );
  NAND2_X1 U35330 ( .A1(n4287), .A2(n4048), .ZN(n2718) );
  NAND2_X1 U35340 ( .A1(n4518), .A2(n4298), .ZN(n4075) );
  NAND2_X1 U35350 ( .A1(n2718), .A2(n4075), .ZN(n4273) );
  INV_X1 U35360 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U35370 ( .A1(n2719), .A2(n4997), .ZN(n2720) );
  NAND2_X1 U35380 ( .A1(n4278), .A2(n2501), .ZN(n2726) );
  INV_X1 U35390 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U35400 ( .A1(n3833), .A2(REG0_REG_25__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U35410 ( .A1(n3834), .A2(REG1_REG_25__SCAN_IN), .ZN(n2721) );
  OAI211_X1 U35420 ( .C1(n2723), .C2(n3837), .A(n2722), .B(n2721), .ZN(n2724)
         );
  INV_X1 U35430 ( .A(n2724), .ZN(n2725) );
  NAND2_X1 U35440 ( .A1(n3832), .A2(DATAI_25_), .ZN(n4280) );
  INV_X1 U35450 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3969) );
  AND2_X1 U35460 ( .A1(n2189), .A2(n3969), .ZN(n2727) );
  NOR2_X1 U35470 ( .A1(n2735), .A2(n2727), .ZN(n4268) );
  NAND2_X1 U35480 ( .A1(n4268), .A2(n2501), .ZN(n2733) );
  INV_X1 U35490 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U35500 ( .A1(n3833), .A2(REG0_REG_26__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U35510 ( .A1(n3834), .A2(REG1_REG_26__SCAN_IN), .ZN(n2728) );
  OAI211_X1 U35520 ( .C1(n2730), .C2(n3837), .A(n2729), .B(n2728), .ZN(n2731)
         );
  INV_X1 U35530 ( .A(n2731), .ZN(n2732) );
  NAND2_X1 U35540 ( .A1(n3832), .A2(DATAI_26_), .ZN(n4266) );
  OR2_X1 U35550 ( .A1(n4508), .A2(n4266), .ZN(n2734) );
  INV_X1 U35560 ( .A(n4280), .ZN(n4517) );
  NAND2_X1 U35570 ( .A1(n5037), .A2(n4517), .ZN(n4255) );
  AND2_X1 U35580 ( .A1(n4508), .A2(n4266), .ZN(n4052) );
  NOR2_X1 U35590 ( .A1(n2735), .A2(REG3_REG_27__SCAN_IN), .ZN(n2736) );
  INV_X1 U35600 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U35610 ( .A1(n3833), .A2(REG0_REG_27__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U35620 ( .A1(n3834), .A2(REG1_REG_27__SCAN_IN), .ZN(n2737) );
  OAI211_X1 U35630 ( .C1(n4244), .C2(n3837), .A(n2738), .B(n2737), .ZN(n2739)
         );
  INV_X1 U35640 ( .A(n2739), .ZN(n2740) );
  NAND2_X1 U35650 ( .A1(n3832), .A2(DATAI_27_), .ZN(n4246) );
  XNOR2_X1 U35660 ( .A(n4148), .B(n4507), .ZN(n4238) );
  NAND2_X1 U35670 ( .A1(n2741), .A2(REG3_REG_28__SCAN_IN), .ZN(n2830) );
  INV_X1 U35680 ( .A(n2741), .ZN(n2743) );
  INV_X1 U35690 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U35700 ( .A1(n2743), .A2(n2742), .ZN(n2744) );
  INV_X1 U35710 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U35720 ( .A1(n3833), .A2(REG0_REG_28__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U35730 ( .A1(n3834), .A2(REG1_REG_28__SCAN_IN), .ZN(n2745) );
  OAI211_X1 U35740 ( .C1(n2747), .C2(n3837), .A(n2746), .B(n2745), .ZN(n2748)
         );
  INV_X1 U35750 ( .A(n2748), .ZN(n2749) );
  NAND2_X1 U35760 ( .A1(n3832), .A2(DATAI_28_), .ZN(n4230) );
  NAND2_X1 U35770 ( .A1(n3868), .A2(n4230), .ZN(n4051) );
  INV_X1 U35780 ( .A(n4230), .ZN(n3194) );
  NAND2_X1 U35790 ( .A1(n4511), .A2(n3194), .ZN(n4055) );
  OR2_X1 U35800 ( .A1(n2830), .A2(n2750), .ZN(n2756) );
  INV_X1 U35810 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U3582 ( .A1(n3834), .A2(REG1_REG_29__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U3583 ( .A1(n3833), .A2(REG0_REG_29__SCAN_IN), .ZN(n2751) );
  OAI211_X1 U3584 ( .C1(n3837), .C2(n2753), .A(n2752), .B(n2751), .ZN(n2754)
         );
  INV_X1 U3585 ( .A(n2754), .ZN(n2755) );
  NAND2_X1 U3586 ( .A1(n3832), .A2(DATAI_29_), .ZN(n2785) );
  INV_X1 U3587 ( .A(n2785), .ZN(n2780) );
  NAND2_X1 U3588 ( .A1(n4229), .A2(n2780), .ZN(n4122) );
  NAND2_X1 U3589 ( .A1(n4147), .A2(n2785), .ZN(n4050) );
  NAND2_X1 U3590 ( .A1(n4122), .A2(n4050), .ZN(n4061) );
  XNOR2_X1 U3591 ( .A(n2758), .B(n2757), .ZN(n2783) );
  INV_X1 U3592 ( .A(n2879), .ZN(n4680) );
  NAND2_X1 U3593 ( .A1(n2172), .A2(IR_REG_31__SCAN_IN), .ZN(n2763) );
  INV_X1 U3594 ( .A(n2795), .ZN(n2765) );
  NAND2_X1 U3595 ( .A1(n4680), .A2(n2878), .ZN(n2769) );
  NAND2_X1 U3596 ( .A1(n4140), .A2(n4681), .ZN(n2768) );
  OAI21_X1 U3597 ( .B1(n2770), .B2(IR_REG_27__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2772) );
  MUX2_X1 U3598 ( .A(n2772), .B(IR_REG_31__SCAN_IN), .S(n2771), .Z(n2774) );
  NAND2_X1 U3599 ( .A1(n2774), .A2(n2773), .ZN(n4692) );
  NAND2_X1 U3600 ( .A1(n3302), .A2(n3153), .ZN(n4480) );
  NAND2_X1 U3601 ( .A1(n2776), .A2(n2775), .ZN(n3300) );
  INV_X1 U3602 ( .A(B_REG_SCAN_IN), .ZN(n4987) );
  NOR2_X1 U3603 ( .A1(n3300), .A2(n4987), .ZN(n2777) );
  NOR2_X1 U3604 ( .A1(n4544), .A2(n2777), .ZN(n3838) );
  INV_X1 U3605 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U3606 ( .A1(n3834), .A2(REG1_REG_30__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U3607 ( .A1(n3833), .A2(REG0_REG_30__SCAN_IN), .ZN(n2778) );
  OAI211_X1 U3608 ( .C1(n3837), .C2(n4223), .A(n2779), .B(n2778), .ZN(n4146)
         );
  AOI22_X1 U3609 ( .A1(n3838), .A2(n4146), .B1(n4540), .B2(n2780), .ZN(n2781)
         );
  OAI21_X1 U3610 ( .B1(n4511), .B2(n4480), .A(n2781), .ZN(n2782) );
  INV_X1 U3611 ( .A(n3219), .ZN(n2832) );
  NAND2_X1 U3612 ( .A1(n2990), .A2(n3540), .ZN(n2784) );
  INV_X1 U3613 ( .A(IR_REG_24__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U3614 ( .A1(n2822), .A2(n2787), .ZN(n2788) );
  NAND2_X1 U3615 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2790) );
  AOI22_X1 U3616 ( .A1(IR_REG_24__SCAN_IN), .A2(n2791), .B1(n2790), .B2(
        IR_REG_31__SCAN_IN), .ZN(n2792) );
  INV_X1 U3617 ( .A(n2792), .ZN(n2793) );
  NAND2_X1 U3618 ( .A1(n2795), .A2(n2794), .ZN(n2821) );
  AND2_X1 U3619 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2796)
         );
  NAND2_X1 U3620 ( .A1(n2798), .A2(n2797), .ZN(n2820) );
  NAND2_X1 U3621 ( .A1(n2801), .A2(n2820), .ZN(n2802) );
  MUX2_X1 U3622 ( .A(n2820), .B(n2802), .S(B_REG_SCAN_IN), .Z(n2806) );
  NAND2_X1 U3623 ( .A1(n2803), .A2(IR_REG_31__SCAN_IN), .ZN(n2804) );
  INV_X1 U3624 ( .A(D_REG_0__SCAN_IN), .ZN(n3287) );
  AND2_X1 U3625 ( .A1(n2820), .A2(n2819), .ZN(n3286) );
  INV_X1 U3626 ( .A(n3213), .ZN(n3207) );
  INV_X1 U3627 ( .A(D_REG_13__SCAN_IN), .ZN(n4830) );
  INV_X1 U3628 ( .A(D_REG_12__SCAN_IN), .ZN(n4829) );
  INV_X1 U3629 ( .A(D_REG_14__SCAN_IN), .ZN(n4828) );
  INV_X1 U3630 ( .A(D_REG_17__SCAN_IN), .ZN(n4819) );
  NAND4_X1 U3631 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4819), .ZN(n2812)
         );
  NOR4_X1 U3632 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2810) );
  NOR4_X1 U3633 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2809) );
  NOR4_X1 U3634 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2808) );
  NOR4_X1 U3635 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2807) );
  NAND4_X1 U3636 ( .A1(n2810), .A2(n2809), .A3(n2808), .A4(n2807), .ZN(n2811)
         );
  NOR4_X1 U3637 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(n2812), 
        .A4(n2811), .ZN(n2815) );
  NOR4_X1 U3638 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2814) );
  NOR4_X1 U3639 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2813) );
  AND2_X1 U3640 ( .A1(n2814), .A2(n2813), .ZN(n4763) );
  NAND2_X1 U3641 ( .A1(n2815), .A2(n4763), .ZN(n2816) );
  NAND2_X1 U3642 ( .A1(n2817), .A2(n2816), .ZN(n3204) );
  NAND2_X1 U3643 ( .A1(n2801), .A2(n2819), .ZN(n3288) );
  NAND2_X1 U3644 ( .A1(n2879), .A2(n4211), .ZN(n2818) );
  NAND2_X1 U3645 ( .A1(n3153), .A2(n2818), .ZN(n3200) );
  AND3_X1 U3646 ( .A1(n3204), .A2(n3288), .A3(n3200), .ZN(n2826) );
  NAND2_X1 U3647 ( .A1(n2821), .A2(IR_REG_31__SCAN_IN), .ZN(n2823) );
  XNOR2_X1 U3648 ( .A(n2823), .B(n2822), .ZN(n3172) );
  INV_X1 U3649 ( .A(D_REG_1__SCAN_IN), .ZN(n2824) );
  INV_X1 U3650 ( .A(n3203), .ZN(n3423) );
  OAI21_X1 U3651 ( .B1(n3203), .B2(n2824), .A(n4728), .ZN(n2825) );
  NAND3_X1 U3652 ( .A1(n3207), .A2(n2826), .A3(n2825), .ZN(n2828) );
  AND2_X1 U3653 ( .A1(n2879), .A2(n4681), .ZN(n4718) );
  NAND2_X1 U3654 ( .A1(n4742), .A2(n2827), .ZN(n3201) );
  OR2_X2 U3655 ( .A1(n3203), .A2(n3201), .ZN(n4492) );
  AND2_X1 U3656 ( .A1(n4611), .A2(n4211), .ZN(n2829) );
  OAI22_X1 U3657 ( .A1(n3230), .A2(n4498), .B1(n2830), .B2(n4492), .ZN(n2831)
         );
  NAND2_X1 U3658 ( .A1(n3540), .A2(n3541), .ZN(n2833) );
  AND2_X1 U3659 ( .A1(n3539), .A2(n2833), .ZN(n2835) );
  NAND2_X1 U3660 ( .A1(n3400), .A2(n3403), .ZN(n3402) );
  NAND2_X1 U3661 ( .A1(n3437), .A2(n4153), .ZN(n2834) );
  NAND2_X1 U3662 ( .A1(n3402), .A2(n2834), .ZN(n3237) );
  NAND2_X1 U3663 ( .A1(n2990), .A2(n3573), .ZN(n3388) );
  NAND3_X1 U3664 ( .A1(n2835), .A2(n3237), .A3(n3388), .ZN(n2840) );
  NAND3_X1 U3665 ( .A1(n2835), .A2(n3388), .A3(n4078), .ZN(n2839) );
  NOR2_X1 U3666 ( .A1(n3541), .A2(n3540), .ZN(n2837) );
  INV_X1 U3667 ( .A(n2836), .ZN(n4152) );
  AOI22_X1 U3668 ( .A1(n3539), .A2(n2837), .B1(n3005), .B2(n4152), .ZN(n2838)
         );
  NAND3_X1 U3669 ( .A1(n2840), .A2(n2839), .A3(n2838), .ZN(n3251) );
  NAND2_X1 U3670 ( .A1(n3490), .A2(n4151), .ZN(n3505) );
  INV_X1 U3671 ( .A(n3505), .ZN(n2843) );
  OR2_X1 U3672 ( .A1(n3596), .A2(n3595), .ZN(n2841) );
  NAND2_X1 U3673 ( .A1(n3474), .A2(n3630), .ZN(n3504) );
  OAI21_X1 U3674 ( .B1(n3251), .B2(n2843), .A(n2441), .ZN(n2848) );
  AOI22_X1 U3675 ( .A1(n2844), .A2(n2846), .B1(n2845), .B2(n3525), .ZN(n2847)
         );
  NAND2_X1 U3676 ( .A1(n2848), .A2(n2847), .ZN(n3609) );
  NAND2_X1 U3677 ( .A1(n3585), .A2(n3685), .ZN(n2849) );
  NAND2_X1 U3678 ( .A1(n3609), .A2(n2849), .ZN(n2851) );
  NAND2_X1 U3679 ( .A1(n3616), .A2(n3691), .ZN(n2850) );
  NAND2_X1 U3680 ( .A1(n2851), .A2(n2850), .ZN(n3658) );
  NOR2_X1 U3681 ( .A1(n3713), .A2(n3693), .ZN(n2853) );
  NAND2_X1 U3682 ( .A1(n3693), .A2(n3713), .ZN(n2852) );
  NAND2_X1 U3683 ( .A1(n4035), .A2(n4031), .ZN(n4088) );
  NAND2_X1 U3684 ( .A1(n3774), .A2(n3732), .ZN(n3729) );
  INV_X1 U3685 ( .A(n3949), .ZN(n4481) );
  NAND2_X1 U3686 ( .A1(n4602), .A2(n4481), .ZN(n2854) );
  AND2_X1 U3687 ( .A1(n3729), .A2(n2854), .ZN(n4487) );
  NOR2_X1 U3688 ( .A1(n4597), .A2(n4495), .ZN(n2856) );
  INV_X1 U3689 ( .A(n2856), .ZN(n2855) );
  AND2_X1 U3690 ( .A1(n4487), .A2(n2855), .ZN(n2857) );
  NAND2_X1 U3691 ( .A1(n3046), .A2(n3949), .ZN(n4489) );
  NAND2_X1 U3692 ( .A1(n3757), .A2(n3756), .ZN(n3755) );
  NAND2_X1 U3693 ( .A1(n4482), .A2(n4588), .ZN(n2858) );
  NAND2_X1 U3694 ( .A1(n4585), .A2(n3069), .ZN(n2860) );
  NOR2_X1 U3695 ( .A1(n4585), .A2(n3069), .ZN(n2859) );
  NAND2_X1 U3696 ( .A1(n4577), .A2(n4446), .ZN(n2861) );
  OR2_X1 U3697 ( .A1(n4568), .A2(n4431), .ZN(n2862) );
  INV_X1 U3698 ( .A(n4408), .ZN(n2864) );
  OR2_X1 U3699 ( .A1(n4561), .A2(n3088), .ZN(n2865) );
  NAND2_X1 U3700 ( .A1(n4414), .A2(n4393), .ZN(n2866) );
  INV_X1 U3701 ( .A(n4376), .ZN(n4368) );
  NOR2_X1 U3702 ( .A1(n4541), .A2(n4368), .ZN(n2868) );
  NAND2_X1 U3703 ( .A1(n4541), .A2(n4368), .ZN(n2867) );
  INV_X1 U3704 ( .A(n4356), .ZN(n4539) );
  NAND2_X1 U3705 ( .A1(n4306), .A2(n2869), .ZN(n4325) );
  NAND2_X1 U3706 ( .A1(n4332), .A2(n3886), .ZN(n2870) );
  NAND2_X1 U3707 ( .A1(n4286), .A2(n2871), .ZN(n2873) );
  NAND2_X1 U3708 ( .A1(n2873), .A2(n2872), .ZN(n4275) );
  INV_X1 U3709 ( .A(n4275), .ZN(n2875) );
  NOR2_X1 U3710 ( .A1(n4508), .A2(n4260), .ZN(n4095) );
  INV_X1 U3711 ( .A(n4148), .ZN(n4264) );
  NAND2_X1 U3712 ( .A1(n4264), .A2(n4246), .ZN(n2876) );
  XNOR2_X1 U3713 ( .A(n2877), .B(n4061), .ZN(n3220) );
  XNOR2_X1 U3714 ( .A(n2972), .B(n4140), .ZN(n2880) );
  NAND2_X1 U3715 ( .A1(n2880), .A2(n4211), .ZN(n4374) );
  OR2_X1 U3716 ( .A1(n2972), .A2(n4211), .ZN(n3241) );
  NAND2_X1 U3717 ( .A1(n4374), .A2(n3241), .ZN(n2881) );
  NAND2_X1 U3718 ( .A1(n4726), .A2(REG2_REG_29__SCAN_IN), .ZN(n2882) );
  OAI21_X1 U3719 ( .B1(n3220), .B2(n4456), .A(n2882), .ZN(n2883) );
  NAND2_X1 U3720 ( .A1(n2885), .A2(n2884), .ZN(U3354) );
  INV_X2 U3721 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3722 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U3723 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4202), .B1(n4732), .B2(
        n4205), .ZN(n2919) );
  NOR2_X1 U3724 ( .A1(n4682), .A2(REG1_REG_17__SCAN_IN), .ZN(n2916) );
  NAND2_X1 U3725 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2962), .ZN(n2910) );
  INV_X1 U3726 ( .A(n3329), .ZN(n4690) );
  INV_X1 U3727 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2886) );
  XNOR2_X1 U3728 ( .A(n2928), .B(n2886), .ZN(n4161) );
  AND2_X1 U3729 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4160)
         );
  NAND2_X1 U3730 ( .A1(n4161), .A2(n4160), .ZN(n4159) );
  NAND2_X1 U3731 ( .A1(n2928), .A2(REG1_REG_1__SCAN_IN), .ZN(n2887) );
  NAND2_X1 U3732 ( .A1(n4159), .A2(n2887), .ZN(n3334) );
  INV_X1 U3733 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4944) );
  XNOR2_X2 U3734 ( .A(n2889), .B(n2248), .ZN(n3295) );
  INV_X1 U3735 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4983) );
  OR2_X1 U3736 ( .A1(n2889), .A2(n2932), .ZN(n2890) );
  INV_X1 U3737 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4752) );
  XOR2_X1 U3738 ( .A(REG1_REG_5__SCAN_IN), .B(n3318), .Z(n3311) );
  INV_X1 U3739 ( .A(n3318), .ZN(n2893) );
  XNOR2_X1 U3740 ( .A(n2894), .B(n4688), .ZN(n3342) );
  INV_X1 U3741 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U3742 ( .A1(n3342), .A2(REG1_REG_6__SCAN_IN), .ZN(n3341) );
  INV_X1 U3743 ( .A(n4688), .ZN(n3343) );
  NAND2_X1 U3744 ( .A1(n3341), .A2(n2895), .ZN(n3372) );
  INV_X1 U3745 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4796) );
  INV_X1 U3746 ( .A(n3466), .ZN(n2943) );
  INV_X1 U3747 ( .A(n3531), .ZN(n2899) );
  INV_X1 U3748 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2897) );
  MUX2_X1 U3749 ( .A(REG1_REG_9__SCAN_IN), .B(n2897), .S(n3533), .Z(n3530) );
  INV_X1 U3750 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4940) );
  MUX2_X1 U3751 ( .A(n4940), .B(REG1_REG_11__SCAN_IN), .S(n4686), .Z(n2901) );
  INV_X1 U3752 ( .A(n4686), .ZN(n4171) );
  INV_X1 U3753 ( .A(n4685), .ZN(n3792) );
  INV_X1 U3754 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2903) );
  MUX2_X1 U3755 ( .A(n2903), .B(REG1_REG_13__SCAN_IN), .S(n4684), .Z(n3811) );
  NAND2_X1 U3756 ( .A1(n4684), .A2(REG1_REG_13__SCAN_IN), .ZN(n2906) );
  INV_X1 U3757 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U3758 ( .A1(n2907), .A2(n4683), .ZN(n2908) );
  OAI21_X2 U3759 ( .B1(n4180), .B2(n4592), .A(n2908), .ZN(n4699) );
  INV_X1 U3760 ( .A(n2962), .ZN(n4735) );
  INV_X1 U3761 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2909) );
  AOI22_X1 U3762 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2962), .B1(n4735), .B2(
        n2909), .ZN(n4700) );
  NAND2_X1 U3763 ( .A1(n4699), .A2(n4700), .ZN(n4698) );
  NAND2_X1 U3764 ( .A1(n2910), .A2(n4698), .ZN(n2912) );
  NOR2_X1 U3765 ( .A1(n2911), .A2(n2912), .ZN(n2913) );
  INV_X1 U3766 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2915) );
  INV_X1 U3767 ( .A(n4682), .ZN(n4196) );
  INV_X1 U3768 ( .A(n2916), .ZN(n2914) );
  OAI21_X1 U3769 ( .B1(n2915), .B2(n4196), .A(n2914), .ZN(n4191) );
  OR2_X1 U3770 ( .A1(n3172), .A2(U3149), .ZN(n4143) );
  NAND2_X1 U3771 ( .A1(n3203), .A2(n4143), .ZN(n2922) );
  NAND2_X1 U3772 ( .A1(n3172), .A2(n3153), .ZN(n2917) );
  AND2_X1 U3773 ( .A1(n2917), .A2(n3832), .ZN(n2920) );
  NAND2_X1 U3774 ( .A1(n2922), .A2(n2920), .ZN(n3306) );
  INV_X1 U3775 ( .A(n3300), .ZN(n4677) );
  NAND2_X1 U3776 ( .A1(n2919), .A2(n2918), .ZN(n4204) );
  OAI211_X1 U3777 ( .C1(n2919), .C2(n2918), .A(n4710), .B(n4204), .ZN(n2926)
         );
  INV_X1 U3778 ( .A(n2920), .ZN(n2921) );
  INV_X1 U3779 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4821) );
  NOR2_X1 U3780 ( .A1(n4821), .A2(STATE_REG_SCAN_IN), .ZN(n3960) );
  AOI21_X1 U3781 ( .B1(n4709), .B2(ADDR_REG_18__SCAN_IN), .A(n3960), .ZN(n2923) );
  OAI21_X1 U3782 ( .B1(n4715), .B2(n4732), .A(n2923), .ZN(n2924) );
  INV_X1 U3783 ( .A(n2924), .ZN(n2925) );
  NAND2_X1 U3784 ( .A1(n2926), .A2(n2925), .ZN(n2969) );
  AOI22_X1 U3785 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4732), .B1(n4202), .B2(
        n2660), .ZN(n2967) );
  INV_X1 U3786 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2927) );
  INV_X1 U3787 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3568) );
  AND2_X1 U3788 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2929)
         );
  NAND2_X1 U3789 ( .A1(n4164), .A2(n2929), .ZN(n4163) );
  NAND2_X1 U3790 ( .A1(n2928), .A2(REG2_REG_1__SCAN_IN), .ZN(n2930) );
  OR2_X1 U3791 ( .A1(n3329), .A2(n2927), .ZN(n2931) );
  NAND2_X1 U3792 ( .A1(n2933), .A2(n2248), .ZN(n2934) );
  INV_X1 U3793 ( .A(n4689), .ZN(n3352) );
  XNOR2_X1 U3794 ( .A(n2935), .B(n3352), .ZN(n3348) );
  NAND2_X1 U3795 ( .A1(n2935), .A2(n4689), .ZN(n2936) );
  MUX2_X1 U3796 ( .A(n2937), .B(REG2_REG_5__SCAN_IN), .S(n3318), .Z(n3314) );
  OR2_X1 U3797 ( .A1(n3318), .A2(n2937), .ZN(n2938) );
  NAND2_X1 U3798 ( .A1(n2939), .A2(n4688), .ZN(n2940) );
  MUX2_X1 U3799 ( .A(n2941), .B(REG2_REG_7__SCAN_IN), .S(n3374), .Z(n3377) );
  OR2_X1 U3800 ( .A1(n3374), .A2(n2941), .ZN(n2942) );
  XNOR2_X1 U3801 ( .A(n2944), .B(n3466), .ZN(n3464) );
  NAND2_X1 U3802 ( .A1(n3464), .A2(REG2_REG_8__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3803 ( .A1(n2944), .A2(n2943), .ZN(n2945) );
  NAND2_X1 U3804 ( .A1(n2946), .A2(n2945), .ZN(n3529) );
  XNOR2_X1 U3805 ( .A(n3533), .B(REG2_REG_9__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U3806 ( .A1(n3529), .A2(n3528), .ZN(n2949) );
  INV_X1 U3807 ( .A(n3533), .ZN(n2947) );
  NAND2_X1 U3808 ( .A1(n2947), .A2(REG2_REG_9__SCAN_IN), .ZN(n2948) );
  NAND2_X1 U3809 ( .A1(n2950), .A2(n4687), .ZN(n2951) );
  MUX2_X1 U3810 ( .A(REG2_REG_11__SCAN_IN), .B(n3746), .S(n4686), .Z(n4175) );
  NAND2_X1 U3811 ( .A1(n4686), .A2(REG2_REG_11__SCAN_IN), .ZN(n2953) );
  NAND2_X1 U3812 ( .A1(n3790), .A2(REG2_REG_12__SCAN_IN), .ZN(n2956) );
  NAND2_X1 U3813 ( .A1(n2954), .A2(n4685), .ZN(n2955) );
  AND2_X1 U3814 ( .A1(n4684), .A2(REG2_REG_13__SCAN_IN), .ZN(n2957) );
  INV_X1 U3815 ( .A(n4684), .ZN(n3814) );
  NAND2_X1 U3816 ( .A1(n3814), .A2(n4494), .ZN(n2958) );
  INV_X1 U3817 ( .A(n4683), .ZN(n4181) );
  OAI21_X1 U3818 ( .B1(n2959), .B2(n4181), .A(n4185), .ZN(n2960) );
  NAND2_X1 U3819 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2962), .ZN(n2961) );
  OAI21_X1 U3820 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2962), .A(n2961), .ZN(n4694) );
  NAND2_X1 U3821 ( .A1(n2963), .A2(n4733), .ZN(n2964) );
  INV_X1 U3822 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4704) );
  NAND2_X1 U3823 ( .A1(n2964), .A2(n4705), .ZN(n4192) );
  XNOR2_X1 U3824 ( .A(n4682), .B(n2965), .ZN(n4194) );
  NAND2_X1 U3825 ( .A1(n4192), .A2(n4194), .ZN(n4193) );
  NAND2_X1 U3826 ( .A1(n3302), .A2(n4677), .ZN(n4138) );
  AOI211_X1 U3827 ( .C1(n2967), .C2(n2966), .A(n4201), .B(n4703), .ZN(n2968)
         );
  NAND2_X2 U3828 ( .A1(n2970), .A2(n2971), .ZN(n2988) );
  NAND2_X1 U3829 ( .A1(n2998), .A2(n4154), .ZN(n2974) );
  INV_X2 U3830 ( .A(n2978), .ZN(n3004) );
  NAND2_X1 U3831 ( .A1(n3004), .A2(n3432), .ZN(n2973) );
  AND2_X1 U3832 ( .A1(n2974), .A2(n2973), .ZN(n2977) );
  INV_X1 U3833 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3299) );
  OR2_X1 U3834 ( .A1(n2971), .A2(n3299), .ZN(n2976) );
  NAND2_X1 U3835 ( .A1(n2977), .A2(n2976), .ZN(n3323) );
  INV_X1 U3836 ( .A(n4154), .ZN(n3575) );
  INV_X1 U3837 ( .A(n2971), .ZN(n3233) );
  AOI22_X1 U3838 ( .A1(n2998), .A2(n3432), .B1(n3233), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2979) );
  OAI21_X1 U3839 ( .B1(n2142), .B2(n3575), .A(n2979), .ZN(n3322) );
  NAND2_X1 U3840 ( .A1(n3323), .A2(n3322), .ZN(n3321) );
  NAND2_X1 U3841 ( .A1(n2980), .A2(n3321), .ZN(n3439) );
  NAND2_X1 U3842 ( .A1(n4153), .A2(n2998), .ZN(n2982) );
  NAND2_X1 U3843 ( .A1(n3004), .A2(n3437), .ZN(n2981) );
  NAND2_X1 U3844 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  XNOR2_X1 U3845 ( .A(n2983), .B(n3146), .ZN(n2984) );
  INV_X1 U3846 ( .A(n4153), .ZN(n3444) );
  XNOR2_X1 U3847 ( .A(n2984), .B(n2985), .ZN(n3440) );
  NAND2_X1 U3848 ( .A1(n3439), .A2(n3440), .ZN(n3438) );
  INV_X1 U3849 ( .A(n2984), .ZN(n2986) );
  NAND2_X1 U3850 ( .A1(n2986), .A2(n2985), .ZN(n2987) );
  NAND2_X1 U3851 ( .A1(n3438), .A2(n2987), .ZN(n3420) );
  INV_X1 U3852 ( .A(n3420), .ZN(n2992) );
  OAI22_X1 U3853 ( .A1(n3573), .A2(n2988), .B1(n2978), .B2(n2990), .ZN(n2989)
         );
  OAI22_X1 U3854 ( .A1(n2142), .A2(n3573), .B1(n3177), .B2(n2990), .ZN(n2994)
         );
  XNOR2_X1 U3855 ( .A(n2993), .B(n2994), .ZN(n3417) );
  INV_X1 U3856 ( .A(n3417), .ZN(n2991) );
  NAND2_X1 U3857 ( .A1(n2992), .A2(n2991), .ZN(n3418) );
  INV_X1 U3858 ( .A(n2993), .ZN(n2996) );
  INV_X1 U3859 ( .A(n2994), .ZN(n2995) );
  NAND2_X1 U3860 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  NAND2_X1 U3861 ( .A1(n3418), .A2(n2997), .ZN(n3480) );
  INV_X4 U3862 ( .A(n2998), .ZN(n3177) );
  XNOR2_X1 U3863 ( .A(n2999), .B(n3146), .ZN(n3002) );
  OAI22_X1 U3864 ( .A1(n2142), .A2(n3541), .B1(n2988), .B2(n3540), .ZN(n3000)
         );
  XNOR2_X1 U3865 ( .A(n3002), .B(n3000), .ZN(n3481) );
  INV_X1 U3866 ( .A(n3000), .ZN(n3001) );
  NAND2_X1 U3867 ( .A1(n3002), .A2(n3001), .ZN(n3003) );
  NAND2_X1 U3868 ( .A1(n3004), .A2(n3005), .ZN(n3006) );
  OAI21_X1 U3869 ( .B1(n2836), .B2(n3177), .A(n3006), .ZN(n3007) );
  XNOR2_X1 U3870 ( .A(n3007), .B(n3142), .ZN(n3011) );
  OAI22_X1 U3871 ( .A1(n2142), .A2(n2836), .B1(n3177), .B2(n3553), .ZN(n3010)
         );
  XNOR2_X1 U3872 ( .A(n3011), .B(n3010), .ZN(n3456) );
  NAND2_X1 U3873 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  OAI22_X1 U3874 ( .A1(n3630), .A2(n3177), .B1(n3148), .B2(n3474), .ZN(n3013)
         );
  XNOR2_X1 U3875 ( .A(n3013), .B(n3146), .ZN(n3014) );
  OAI22_X1 U3876 ( .A1(n2142), .A2(n3630), .B1(n3177), .B2(n3474), .ZN(n3015)
         );
  XNOR2_X1 U3877 ( .A(n3014), .B(n3015), .ZN(n3472) );
  INV_X1 U3878 ( .A(n3014), .ZN(n3016) );
  NAND2_X1 U3879 ( .A1(n3016), .A2(n3015), .ZN(n3017) );
  OAI22_X1 U3880 ( .A1(n2142), .A2(n3599), .B1(n2988), .B2(n3631), .ZN(n3518)
         );
  NAND2_X1 U3881 ( .A1(n3004), .A2(n3595), .ZN(n3019) );
  NAND2_X1 U3882 ( .A1(n3095), .A2(n3596), .ZN(n3018) );
  NAND2_X1 U3883 ( .A1(n3019), .A2(n3018), .ZN(n3020) );
  XNOR2_X1 U3884 ( .A(n3020), .B(n3142), .ZN(n3519) );
  OAI22_X1 U3885 ( .A1(n3632), .A2(n3177), .B1(n3148), .B2(n3592), .ZN(n3021)
         );
  XNOR2_X1 U3886 ( .A(n3021), .B(n3146), .ZN(n3022) );
  OAI22_X1 U3887 ( .A1(n2142), .A2(n3632), .B1(n2988), .B2(n3592), .ZN(n3023)
         );
  XNOR2_X1 U3888 ( .A(n3022), .B(n3023), .ZN(n3561) );
  INV_X1 U3889 ( .A(n3022), .ZN(n3024) );
  OAI22_X1 U3890 ( .A1(n3685), .A2(n3177), .B1(n3148), .B2(n3585), .ZN(n3025)
         );
  XNOR2_X1 U3891 ( .A(n3025), .B(n3142), .ZN(n3026) );
  OAI22_X1 U3892 ( .A1(n2142), .A2(n3685), .B1(n3177), .B2(n3585), .ZN(n3027)
         );
  AND2_X1 U3893 ( .A1(n3026), .A2(n3027), .ZN(n3580) );
  INV_X1 U3894 ( .A(n3026), .ZN(n3029) );
  INV_X1 U3895 ( .A(n3027), .ZN(n3028) );
  NAND2_X1 U3896 ( .A1(n3029), .A2(n3028), .ZN(n3581) );
  OAI22_X1 U3897 ( .A1(n3713), .A2(n3177), .B1(n3148), .B2(n3693), .ZN(n3030)
         );
  XNOR2_X1 U3898 ( .A(n3030), .B(n3146), .ZN(n3033) );
  OAI22_X1 U3899 ( .A1(n2142), .A2(n3713), .B1(n3177), .B2(n3693), .ZN(n3031)
         );
  XNOR2_X1 U3900 ( .A(n3033), .B(n3031), .ZN(n3683) );
  NAND2_X1 U3901 ( .A1(n3682), .A2(n3683), .ZN(n3035) );
  INV_X1 U3902 ( .A(n3031), .ZN(n3032) );
  NAND2_X1 U3903 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  NAND2_X1 U3904 ( .A1(n3095), .A2(n4149), .ZN(n3037) );
  NAND2_X1 U3905 ( .A1(n3004), .A2(n3715), .ZN(n3036) );
  NAND2_X1 U3906 ( .A1(n3037), .A2(n3036), .ZN(n3038) );
  XNOR2_X1 U3907 ( .A(n3038), .B(n3142), .ZN(n3041) );
  OAI22_X1 U3908 ( .A1(n2142), .A2(n3779), .B1(n3177), .B2(n3704), .ZN(n3040)
         );
  XNOR2_X1 U3909 ( .A(n3041), .B(n3040), .ZN(n3701) );
  NAND2_X1 U3910 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  OAI22_X1 U3911 ( .A1(n2142), .A2(n3732), .B1(n3177), .B2(n3774), .ZN(n3768)
         );
  NAND2_X1 U3912 ( .A1(n3004), .A2(n3043), .ZN(n3044) );
  OAI21_X1 U3913 ( .B1(n3732), .B2(n3177), .A(n3044), .ZN(n3045) );
  XNOR2_X1 U3914 ( .A(n3045), .B(n3142), .ZN(n3769) );
  NAND2_X1 U3915 ( .A1(n3004), .A2(n3046), .ZN(n3048) );
  NAND2_X1 U3916 ( .A1(n3095), .A2(n3949), .ZN(n3047) );
  NAND2_X1 U3917 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XNOR2_X1 U3918 ( .A(n3049), .B(n3142), .ZN(n3050) );
  OAI22_X1 U3919 ( .A1(n2142), .A2(n4481), .B1(n3177), .B2(n4602), .ZN(n3051)
         );
  AND2_X1 U3920 ( .A1(n3050), .A2(n3051), .ZN(n3798) );
  INV_X1 U3921 ( .A(n3050), .ZN(n3053) );
  INV_X1 U3922 ( .A(n3051), .ZN(n3052) );
  NAND2_X1 U3923 ( .A1(n3053), .A2(n3052), .ZN(n3799) );
  NAND2_X1 U3924 ( .A1(n3095), .A2(n4597), .ZN(n3055) );
  NAND2_X1 U3925 ( .A1(n3004), .A2(n4495), .ZN(n3054) );
  NAND2_X1 U3926 ( .A1(n3055), .A2(n3054), .ZN(n3056) );
  XNOR2_X1 U3927 ( .A(n3056), .B(n3146), .ZN(n3943) );
  INV_X1 U3928 ( .A(n4597), .ZN(n3803) );
  OAI22_X1 U3929 ( .A1(n2142), .A2(n3803), .B1(n2988), .B2(n3946), .ZN(n3942)
         );
  NAND2_X1 U3930 ( .A1(n3004), .A2(n3762), .ZN(n3059) );
  NAND2_X1 U3931 ( .A1(n3095), .A2(n4576), .ZN(n3058) );
  NAND2_X1 U3932 ( .A1(n3059), .A2(n3058), .ZN(n3060) );
  XNOR2_X1 U3933 ( .A(n3060), .B(n3146), .ZN(n3063) );
  INV_X1 U3934 ( .A(n3063), .ZN(n3061) );
  OAI22_X1 U3935 ( .A1(n2142), .A2(n4482), .B1(n2988), .B2(n4588), .ZN(n3062)
         );
  INV_X1 U3936 ( .A(n3062), .ZN(n3064) );
  NAND2_X1 U3937 ( .A1(n4577), .A2(n3095), .ZN(n3066) );
  NAND2_X1 U3938 ( .A1(n4446), .A2(n3004), .ZN(n3065) );
  NAND2_X1 U3939 ( .A1(n3066), .A2(n3065), .ZN(n3067) );
  XNOR2_X1 U3940 ( .A(n3067), .B(n3146), .ZN(n3909) );
  NOR2_X1 U3941 ( .A1(n4570), .A2(n3177), .ZN(n3068) );
  AOI21_X1 U3942 ( .B1(n4577), .B2(n3145), .A(n3068), .ZN(n3910) );
  NOR2_X1 U3943 ( .A1(n3909), .A2(n3910), .ZN(n3080) );
  NAND2_X1 U3944 ( .A1(n3095), .A2(n4585), .ZN(n3071) );
  NAND2_X1 U3945 ( .A1(n3004), .A2(n3069), .ZN(n3070) );
  NAND2_X1 U3946 ( .A1(n3071), .A2(n3070), .ZN(n3072) );
  XNOR2_X1 U3947 ( .A(n3072), .B(n3142), .ZN(n3908) );
  OAI22_X1 U3948 ( .A1(n3875), .A2(n2142), .B1(n3177), .B2(n4579), .ZN(n3907)
         );
  NAND2_X1 U3949 ( .A1(n4568), .A2(n3095), .ZN(n3076) );
  NAND2_X1 U3950 ( .A1(n3004), .A2(n4431), .ZN(n3075) );
  NAND2_X1 U3951 ( .A1(n3076), .A2(n3075), .ZN(n3077) );
  XNOR2_X1 U3952 ( .A(n3077), .B(n3142), .ZN(n3920) );
  NAND2_X1 U3953 ( .A1(n4568), .A2(n3145), .ZN(n3079) );
  NAND2_X1 U3954 ( .A1(n3095), .A2(n4431), .ZN(n3078) );
  NAND2_X1 U3955 ( .A1(n3079), .A2(n3078), .ZN(n3919) );
  OR3_X1 U3956 ( .A1(n3080), .A2(n3907), .A3(n3908), .ZN(n3081) );
  NAND2_X1 U3957 ( .A1(n3909), .A2(n3910), .ZN(n3917) );
  OAI211_X1 U3958 ( .C1(n3920), .C2(n3919), .A(n3081), .B(n3917), .ZN(n3082)
         );
  INV_X1 U3959 ( .A(n3920), .ZN(n3086) );
  INV_X1 U3960 ( .A(n3919), .ZN(n3085) );
  NAND2_X1 U3961 ( .A1(n4561), .A2(n3095), .ZN(n3090) );
  NAND2_X1 U3962 ( .A1(n3004), .A2(n3088), .ZN(n3089) );
  NAND2_X1 U3963 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
  XNOR2_X1 U3964 ( .A(n3091), .B(n3146), .ZN(n3094) );
  NOR2_X1 U3965 ( .A1(n3177), .A2(n4417), .ZN(n3092) );
  AOI21_X1 U3966 ( .B1(n4561), .B2(n3145), .A(n3092), .ZN(n3093) );
  NOR2_X1 U3967 ( .A1(n3094), .A2(n3093), .ZN(n3953) );
  NAND2_X1 U3968 ( .A1(n3094), .A2(n3093), .ZN(n3954) );
  OAI22_X1 U3969 ( .A1(n3958), .A2(n2142), .B1(n2988), .B2(n4399), .ZN(n3100)
         );
  NAND2_X1 U3970 ( .A1(n4414), .A2(n3095), .ZN(n3097) );
  NAND2_X1 U3971 ( .A1(n3004), .A2(n4393), .ZN(n3096) );
  NAND2_X1 U3972 ( .A1(n3097), .A2(n3096), .ZN(n3098) );
  XNOR2_X1 U3973 ( .A(n3098), .B(n3142), .ZN(n3099) );
  XOR2_X1 U3974 ( .A(n3100), .B(n3099), .Z(n3892) );
  INV_X1 U3975 ( .A(n3099), .ZN(n3102) );
  INV_X1 U3976 ( .A(n3100), .ZN(n3101) );
  NOR2_X1 U3977 ( .A1(n3148), .A2(n4376), .ZN(n3103) );
  AOI21_X1 U3978 ( .B1(n4541), .B2(n3095), .A(n3103), .ZN(n3104) );
  XNOR2_X1 U3979 ( .A(n3104), .B(n3142), .ZN(n3107) );
  NOR2_X1 U3980 ( .A1(n3177), .A2(n4376), .ZN(n3105) );
  AOI21_X1 U3981 ( .B1(n4541), .B2(n3145), .A(n3105), .ZN(n3106) );
  NOR2_X1 U3982 ( .A1(n3107), .A2(n3106), .ZN(n3931) );
  NAND2_X1 U3983 ( .A1(n4329), .A2(n3095), .ZN(n3109) );
  OR2_X1 U3984 ( .A1(n3148), .A2(n4356), .ZN(n3108) );
  NAND2_X1 U3985 ( .A1(n3109), .A2(n3108), .ZN(n3110) );
  XNOR2_X1 U3986 ( .A(n3110), .B(n3146), .ZN(n3899) );
  NOR2_X1 U3987 ( .A1(n3177), .A2(n4356), .ZN(n3111) );
  AOI21_X1 U3988 ( .B1(n4329), .B2(n3145), .A(n3111), .ZN(n3112) );
  NAND2_X1 U3989 ( .A1(n3899), .A2(n3112), .ZN(n3114) );
  INV_X1 U3990 ( .A(n3899), .ZN(n3113) );
  INV_X1 U3991 ( .A(n3112), .ZN(n3898) );
  OAI22_X1 U3992 ( .A1(n4545), .A2(n2142), .B1(n2988), .B2(n3266), .ZN(n3117)
         );
  OAI22_X1 U3993 ( .A1(n4545), .A2(n3177), .B1(n3148), .B2(n3266), .ZN(n3115)
         );
  XNOR2_X1 U3994 ( .A(n3115), .B(n3142), .ZN(n3118) );
  XOR2_X1 U3995 ( .A(n3117), .B(n3118), .Z(n3263) );
  OAI22_X1 U3996 ( .A1(n4332), .A2(n3177), .B1(n3148), .B2(n3886), .ZN(n3116)
         );
  XNOR2_X1 U3997 ( .A(n3116), .B(n3142), .ZN(n3122) );
  OAI22_X1 U3998 ( .A1(n4332), .A2(n2142), .B1(n2988), .B2(n3886), .ZN(n3121)
         );
  XNOR2_X1 U3999 ( .A(n3122), .B(n3121), .ZN(n3880) );
  NOR2_X1 U4000 ( .A1(n3118), .A2(n3117), .ZN(n3881) );
  NOR2_X1 U4001 ( .A1(n3880), .A2(n3881), .ZN(n3119) );
  OAI22_X1 U4002 ( .A1(n5037), .A2(n3177), .B1(n3148), .B2(n4280), .ZN(n3120)
         );
  XNOR2_X1 U4003 ( .A(n3120), .B(n3142), .ZN(n3855) );
  OAI22_X1 U4004 ( .A1(n5037), .A2(n2142), .B1(n3177), .B2(n4280), .ZN(n3854)
         );
  NAND2_X1 U4005 ( .A1(n3855), .A2(n3854), .ZN(n3853) );
  NAND2_X1 U4006 ( .A1(n3122), .A2(n3121), .ZN(n3823) );
  INV_X1 U4007 ( .A(n3823), .ZN(n3125) );
  OAI22_X1 U4008 ( .A1(n4312), .A2(n3177), .B1(n3148), .B2(n4298), .ZN(n3123)
         );
  XNOR2_X1 U4009 ( .A(n3123), .B(n3142), .ZN(n3825) );
  NOR2_X1 U4010 ( .A1(n3177), .A2(n4298), .ZN(n3124) );
  AOI21_X1 U4011 ( .B1(n4518), .B2(n3145), .A(n3124), .ZN(n3822) );
  NAND2_X1 U4012 ( .A1(n3823), .A2(n3822), .ZN(n3820) );
  OAI21_X1 U4013 ( .B1(n3125), .B2(n3825), .A(n3820), .ZN(n3126) );
  NAND2_X1 U4014 ( .A1(n3883), .A2(n3127), .ZN(n3133) );
  INV_X1 U4015 ( .A(n3825), .ZN(n3851) );
  INV_X1 U4016 ( .A(n3854), .ZN(n3128) );
  AOI21_X1 U4017 ( .B1(n3851), .B2(n3822), .A(n3128), .ZN(n3130) );
  NAND3_X1 U4018 ( .A1(n3128), .A2(n3822), .A3(n3851), .ZN(n3129) );
  NAND2_X1 U4019 ( .A1(n4508), .A2(n3095), .ZN(n3135) );
  OR2_X1 U4020 ( .A1(n3148), .A2(n4266), .ZN(n3134) );
  NAND2_X1 U4021 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  XNOR2_X1 U4022 ( .A(n3136), .B(n3146), .ZN(n3139) );
  NOR2_X1 U4023 ( .A1(n3177), .A2(n4266), .ZN(n3137) );
  AOI21_X1 U4024 ( .B1(n4508), .B2(n3145), .A(n3137), .ZN(n3138) );
  OR2_X1 U4025 ( .A1(n3139), .A2(n3138), .ZN(n3966) );
  AND2_X1 U4026 ( .A1(n3139), .A2(n3138), .ZN(n3965) );
  NAND2_X1 U4027 ( .A1(n4148), .A2(n3095), .ZN(n3141) );
  OR2_X1 U4028 ( .A1(n3148), .A2(n4246), .ZN(n3140) );
  NAND2_X1 U4029 ( .A1(n3141), .A2(n3140), .ZN(n3143) );
  XNOR2_X1 U4030 ( .A(n3143), .B(n3142), .ZN(n3162) );
  NOR2_X1 U4031 ( .A1(n3177), .A2(n4246), .ZN(n3144) );
  AOI21_X1 U4032 ( .B1(n4148), .B2(n3145), .A(n3144), .ZN(n3160) );
  XNOR2_X1 U4033 ( .A(n3162), .B(n3160), .ZN(n3863) );
  NAND2_X1 U4034 ( .A1(n3864), .A2(n3863), .ZN(n3166) );
  INV_X1 U4035 ( .A(n3166), .ZN(n3159) );
  OAI22_X1 U4036 ( .A1(n4511), .A2(n2142), .B1(n2988), .B2(n4230), .ZN(n3147)
         );
  XNOR2_X1 U4037 ( .A(n3147), .B(n3146), .ZN(n3150) );
  OAI22_X1 U4038 ( .A1(n4511), .A2(n3177), .B1(n3148), .B2(n4230), .ZN(n3149)
         );
  XNOR2_X1 U4039 ( .A(n3150), .B(n3149), .ZN(n3168) );
  INV_X1 U4040 ( .A(n3168), .ZN(n3158) );
  OAI21_X1 U4041 ( .B1(n3151), .B2(D_REG_1__SCAN_IN), .A(n3288), .ZN(n3206) );
  INV_X1 U4042 ( .A(n3206), .ZN(n3152) );
  NAND3_X1 U40430 ( .A1(n3152), .A2(n3213), .A3(n3204), .ZN(n3183) );
  INV_X1 U4044 ( .A(n3153), .ZN(n3155) );
  NAND2_X1 U4045 ( .A1(n3367), .A2(n4681), .ZN(n3154) );
  NAND2_X1 U4046 ( .A1(n3155), .A2(n3154), .ZN(n3156) );
  OR2_X1 U4047 ( .A1(n3203), .A2(n3169), .ZN(n3157) );
  NAND2_X1 U4048 ( .A1(n3159), .A2(n2440), .ZN(n3190) );
  INV_X1 U4049 ( .A(n3160), .ZN(n3161) );
  NAND2_X1 U4050 ( .A1(n3162), .A2(n3161), .ZN(n3167) );
  INV_X1 U4051 ( .A(n3167), .ZN(n3163) );
  NOR2_X1 U4052 ( .A1(n3163), .A2(n3974), .ZN(n3164) );
  AND2_X1 U4053 ( .A1(n3168), .A2(n3164), .ZN(n3165) );
  NAND2_X1 U4054 ( .A1(n3166), .A2(n3165), .ZN(n3189) );
  NOR3_X1 U4055 ( .A1(n3168), .A2(n3974), .A3(n3167), .ZN(n3187) );
  NAND2_X1 U4056 ( .A1(n3169), .A2(n4603), .ZN(n3170) );
  NAND2_X1 U4057 ( .A1(n3183), .A2(n3170), .ZN(n3171) );
  NAND2_X1 U4058 ( .A1(n3171), .A2(n3200), .ZN(n3421) );
  NAND2_X1 U4059 ( .A1(n2971), .A2(n3172), .ZN(n3173) );
  OAI21_X1 U4060 ( .B1(n3421), .B2(n3173), .A(STATE_REG_SCAN_IN), .ZN(n3178)
         );
  INV_X1 U4061 ( .A(n3174), .ZN(n3175) );
  NAND2_X1 U4062 ( .A1(n4729), .A2(n3175), .ZN(n3176) );
  NAND2_X1 U4063 ( .A1(n3183), .A2(n4137), .ZN(n3422) );
  NAND2_X1 U4064 ( .A1(n4137), .A2(n4692), .ZN(n3179) );
  OR2_X1 U4065 ( .A1(n3203), .A2(n4603), .ZN(n3180) );
  OR2_X1 U4066 ( .A1(n3183), .A2(n3180), .ZN(n3181) );
  INV_X1 U4067 ( .A(n3986), .ZN(n3924) );
  AOI22_X1 U4068 ( .A1(n4147), .A2(n3923), .B1(n3194), .B2(n3924), .ZN(n3185)
         );
  NAND2_X1 U4069 ( .A1(n4137), .A2(n3302), .ZN(n3182) );
  AOI22_X1 U4070 ( .A1(n4148), .A2(n3961), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3184) );
  OAI211_X1 U4071 ( .C1(n3993), .C2(n4226), .A(n3185), .B(n3184), .ZN(n3186)
         );
  NOR2_X1 U4072 ( .A1(n3187), .A2(n3186), .ZN(n3188) );
  NAND3_X1 U4073 ( .A1(n3190), .A2(n3189), .A3(n3188), .ZN(U3217) );
  INV_X1 U4074 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3208) );
  XNOR2_X1 U4075 ( .A(n3191), .B(n2363), .ZN(n3192) );
  NAND2_X1 U4076 ( .A1(n3192), .A2(n4590), .ZN(n4236) );
  INV_X1 U4077 ( .A(n4236), .ZN(n3199) );
  XNOR2_X1 U4078 ( .A(n3193), .B(n2363), .ZN(n4224) );
  INV_X1 U4079 ( .A(n4742), .ZN(n4614) );
  AOI22_X1 U4080 ( .A1(n4148), .A2(n4599), .B1(n4540), .B2(n3194), .ZN(n3195)
         );
  AOI21_X1 U4081 ( .B1(n4224), .B2(n4607), .A(n3196), .ZN(n3197) );
  INV_X1 U4082 ( .A(n3197), .ZN(n3198) );
  NOR2_X1 U4083 ( .A1(n3199), .A2(n3198), .ZN(n3215) );
  NAND2_X1 U4084 ( .A1(n3201), .A2(n3200), .ZN(n3202) );
  NOR2_X1 U4085 ( .A1(n3203), .A2(n3202), .ZN(n3205) );
  MUX2_X1 U4086 ( .A(n3208), .B(n3215), .S(n4751), .Z(n3212) );
  INV_X1 U4087 ( .A(n3209), .ZN(n3210) );
  OAI21_X1 U4088 ( .B1(n4241), .B2(n4230), .A(n3210), .ZN(n4225) );
  NAND2_X1 U4089 ( .A1(n3212), .A2(n3211), .ZN(U3514) );
  INV_X1 U4090 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3216) );
  MUX2_X1 U4091 ( .A(n3216), .B(n3215), .S(n4756), .Z(n3218) );
  NAND2_X2 U4092 ( .A1(n4756), .A2(n4611), .ZN(n4609) );
  NAND2_X1 U4093 ( .A1(n3218), .A2(n3217), .ZN(U3546) );
  OAI21_X1 U4094 ( .B1(n3220), .B2(n4744), .A(n3219), .ZN(n3226) );
  NAND2_X1 U4095 ( .A1(n4754), .A2(n3221), .ZN(n3222) );
  NAND2_X1 U4096 ( .A1(n3223), .A2(n3222), .ZN(n3225) );
  NAND2_X1 U4097 ( .A1(n3225), .A2(n3224), .ZN(U3547) );
  NAND2_X1 U4098 ( .A1(n4749), .A2(n3227), .ZN(n3228) );
  NAND2_X1 U4099 ( .A1(n3229), .A2(n3228), .ZN(n3232) );
  NAND2_X1 U4100 ( .A1(n3232), .A2(n3231), .ZN(U3515) );
  OAI21_X1 U4101 ( .B1(n4078), .B2(n3235), .A(n3234), .ZN(n3236) );
  NAND2_X1 U4102 ( .A1(n3236), .A2(n4590), .ZN(n3240) );
  OR2_X1 U4103 ( .A1(n3237), .A2(n4078), .ZN(n3389) );
  NAND2_X1 U4104 ( .A1(n3237), .A2(n4078), .ZN(n3238) );
  NAND2_X1 U4105 ( .A1(n3389), .A2(n3238), .ZN(n3450) );
  INV_X1 U4106 ( .A(n4374), .ZN(n3742) );
  NAND2_X1 U4107 ( .A1(n3450), .A2(n3742), .ZN(n3239) );
  NAND2_X1 U4108 ( .A1(n3240), .A2(n3239), .ZN(n3448) );
  MUX2_X1 U4109 ( .A(n3448), .B(REG2_REG_2__SCAN_IN), .S(n4726), .Z(n3248) );
  NAND2_X1 U4110 ( .A1(n4724), .A2(n4599), .ZN(n4469) );
  NAND2_X1 U4111 ( .A1(n4724), .A2(n4540), .ZN(n4468) );
  OAI22_X1 U4112 ( .A1(n3444), .A2(n4469), .B1(n4468), .B2(n2990), .ZN(n3247)
         );
  INV_X1 U4113 ( .A(n3241), .ZN(n3242) );
  NAND2_X1 U4114 ( .A1(n4724), .A2(n3242), .ZN(n4385) );
  INV_X1 U4115 ( .A(n3450), .ZN(n3244) );
  OAI22_X1 U4116 ( .A1(n4385), .A2(n3244), .B1(n3243), .B2(n4492), .ZN(n3246)
         );
  NAND2_X1 U4117 ( .A1(n4724), .A2(n4598), .ZN(n4451) );
  XNOR2_X1 U4118 ( .A(n3399), .B(n3446), .ZN(n3498) );
  OAI22_X1 U4119 ( .A1(n3541), .A2(n4451), .B1(n4498), .B2(n3498), .ZN(n3245)
         );
  OR4_X1 U4120 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(U3288) );
  AND2_X1 U4121 ( .A1(n4022), .A2(n4005), .ZN(n4080) );
  XOR2_X1 U4122 ( .A(n4080), .B(n3249), .Z(n3250) );
  NAND2_X1 U4123 ( .A1(n3250), .A2(n4590), .ZN(n3492) );
  NOR2_X1 U4124 ( .A1(n3492), .A2(n4726), .ZN(n3261) );
  INV_X1 U4125 ( .A(n4080), .ZN(n3253) );
  XNOR2_X1 U4126 ( .A(n3252), .B(n3253), .ZN(n3493) );
  NOR2_X1 U4127 ( .A1(n3493), .A2(n4456), .ZN(n3260) );
  OAI22_X1 U4128 ( .A1(n4724), .A2(n2937), .B1(n3479), .B2(n4492), .ZN(n3254)
         );
  INV_X1 U4129 ( .A(n3254), .ZN(n3257) );
  NAND2_X1 U4130 ( .A1(n3552), .A2(n3490), .ZN(n3255) );
  NAND2_X1 U4131 ( .A1(n2439), .A2(n3255), .ZN(n3502) );
  OR2_X1 U4132 ( .A1(n4498), .A2(n3502), .ZN(n3256) );
  OAI211_X1 U4133 ( .C1(n4468), .C2(n3474), .A(n3257), .B(n3256), .ZN(n3259)
         );
  OAI22_X1 U4134 ( .A1(n2836), .A2(n4469), .B1(n4451), .B2(n3599), .ZN(n3258)
         );
  OR4_X1 U4135 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(U3285) );
  INV_X1 U4136 ( .A(n3264), .ZN(n4339) );
  NOR2_X1 U4137 ( .A1(n3993), .A2(n4339), .ZN(n3269) );
  OAI22_X1 U4138 ( .A1(n4332), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n3265), 
        .ZN(n3268) );
  INV_X1 U4139 ( .A(n4329), .ZN(n4370) );
  OAI22_X1 U4140 ( .A1(n3986), .A2(n3266), .B1(n4370), .B2(n3988), .ZN(n3267)
         );
  MUX2_X1 U4141 ( .A(n3318), .B(n2517), .S(U3149), .Z(n3270) );
  INV_X1 U4142 ( .A(n3270), .ZN(U3347) );
  INV_X1 U4143 ( .A(DATAI_29_), .ZN(n4871) );
  NAND2_X1 U4144 ( .A1(n3271), .A2(STATE_REG_SCAN_IN), .ZN(n3272) );
  OAI21_X1 U4145 ( .B1(STATE_REG_SCAN_IN), .B2(n4871), .A(n3272), .ZN(U3323)
         );
  MUX2_X1 U4146 ( .A(n2538), .B(n3374), .S(STATE_REG_SCAN_IN), .Z(n3273) );
  INV_X1 U4147 ( .A(n3273), .ZN(U3345) );
  MUX2_X1 U4148 ( .A(n3274), .B(n3466), .S(STATE_REG_SCAN_IN), .Z(n3275) );
  INV_X1 U4149 ( .A(n3275), .ZN(U3344) );
  INV_X1 U4150 ( .A(DATAI_21_), .ZN(n3277) );
  NAND2_X1 U4151 ( .A1(n2878), .A2(STATE_REG_SCAN_IN), .ZN(n3276) );
  OAI21_X1 U4152 ( .B1(STATE_REG_SCAN_IN), .B2(n3277), .A(n3276), .ZN(U3331)
         );
  INV_X1 U4153 ( .A(DATAI_30_), .ZN(n3280) );
  NAND2_X1 U4154 ( .A1(n2141), .A2(STATE_REG_SCAN_IN), .ZN(n3279) );
  OAI21_X1 U4155 ( .B1(STATE_REG_SCAN_IN), .B2(n3280), .A(n3279), .ZN(U3322)
         );
  MUX2_X1 U4156 ( .A(n3533), .B(n2567), .S(U3149), .Z(n3281) );
  INV_X1 U4157 ( .A(n3281), .ZN(U3343) );
  INV_X1 U4158 ( .A(DATAI_22_), .ZN(n3283) );
  NAND2_X1 U4159 ( .A1(n4140), .A2(STATE_REG_SCAN_IN), .ZN(n3282) );
  OAI21_X1 U4160 ( .B1(STATE_REG_SCAN_IN), .B2(n3283), .A(n3282), .ZN(U3330)
         );
  INV_X1 U4161 ( .A(DATAI_24_), .ZN(n3284) );
  MUX2_X1 U4162 ( .A(n2820), .B(n3284), .S(U3149), .Z(n3285) );
  INV_X1 U4163 ( .A(n3285), .ZN(U3328) );
  AOI22_X1 U4164 ( .A1(n4728), .A2(n3287), .B1(n3286), .B2(n4729), .ZN(U3458)
         );
  INV_X1 U4165 ( .A(n3288), .ZN(n3289) );
  AOI22_X1 U4166 ( .A1(n4728), .A2(n2824), .B1(n3289), .B2(n4729), .ZN(U3459)
         );
  NOR2_X1 U4167 ( .A1(n4709), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U4168 ( .A(n3290), .B(REG2_REG_3__SCAN_IN), .ZN(n3298) );
  INV_X1 U4169 ( .A(n4715), .ZN(n4158) );
  INV_X1 U4170 ( .A(n4709), .ZN(n3292) );
  INV_X1 U4171 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3291) );
  INV_X1 U4172 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3648) );
  OAI22_X1 U4173 ( .A1(n3292), .A2(n3291), .B1(STATE_REG_SCAN_IN), .B2(n3648), 
        .ZN(n3293) );
  AOI21_X1 U4174 ( .B1(n2248), .B2(n4158), .A(n3293), .ZN(n3297) );
  OAI211_X1 U4175 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3295), .A(n4710), .B(n3294), 
        .ZN(n3296) );
  OAI211_X1 U4176 ( .C1(n3298), .C2(n4703), .A(n3297), .B(n3296), .ZN(U3243)
         );
  AOI21_X1 U4177 ( .B1(n3300), .B2(n3299), .A(IR_REG_0__SCAN_IN), .ZN(n3304)
         );
  OR2_X1 U4178 ( .A1(n3300), .A2(REG2_REG_0__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4179 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  NAND2_X1 U4180 ( .A1(n3303), .A2(n2235), .ZN(n3324) );
  OAI21_X1 U4181 ( .B1(n3304), .B2(n3303), .A(n3324), .ZN(n3305) );
  OAI22_X1 U4182 ( .A1(n3306), .A2(n3305), .B1(STATE_REG_SCAN_IN), .B2(n3434), 
        .ZN(n3308) );
  NOR3_X1 U4183 ( .A1(n4199), .A2(REG1_REG_0__SCAN_IN), .A3(n2235), .ZN(n3307)
         );
  AOI211_X1 U4184 ( .C1(n4709), .C2(ADDR_REG_0__SCAN_IN), .A(n3308), .B(n3307), 
        .ZN(n3309) );
  INV_X1 U4185 ( .A(n3309), .ZN(U3240) );
  AOI211_X1 U4186 ( .C1(n2196), .C2(n3311), .A(n4199), .B(n3310), .ZN(n3320)
         );
  OAI211_X1 U4187 ( .C1(n3314), .C2(n3313), .A(n4184), .B(n3312), .ZN(n3317)
         );
  NOR2_X1 U4188 ( .A1(n3315), .A2(STATE_REG_SCAN_IN), .ZN(n3476) );
  AOI21_X1 U4189 ( .B1(n4709), .B2(ADDR_REG_5__SCAN_IN), .A(n3476), .ZN(n3316)
         );
  OAI211_X1 U4190 ( .C1(n4715), .C2(n3318), .A(n3317), .B(n3316), .ZN(n3319)
         );
  OR2_X1 U4191 ( .A1(n3320), .A2(n3319), .ZN(U3245) );
  OAI21_X1 U4192 ( .B1(n3323), .B2(n3322), .A(n3321), .ZN(n3430) );
  NOR2_X1 U4193 ( .A1(n4692), .A2(n4677), .ZN(n3326) );
  NAND2_X1 U4194 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4162) );
  OAI211_X1 U4195 ( .C1(n4162), .C2(n4138), .A(U4043), .B(n3324), .ZN(n3325)
         );
  AOI21_X1 U4196 ( .B1(n3430), .B2(n3326), .A(n3325), .ZN(n3354) );
  NAND2_X1 U4197 ( .A1(U3149), .A2(REG3_REG_2__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4198 ( .A1(n4709), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3327) );
  OAI211_X1 U4199 ( .C1(n4715), .C2(n3329), .A(n3328), .B(n3327), .ZN(n3339)
         );
  OAI21_X1 U4200 ( .B1(n3332), .B2(n3331), .A(n3330), .ZN(n3337) );
  OAI21_X1 U4201 ( .B1(n3335), .B2(n3334), .A(n3333), .ZN(n3336) );
  OAI22_X1 U4202 ( .A1(n4703), .A2(n3337), .B1(n4199), .B2(n3336), .ZN(n3338)
         );
  OR3_X1 U4203 ( .A1(n3354), .A2(n3339), .A3(n3338), .ZN(U3242) );
  XNOR2_X1 U4204 ( .A(n3340), .B(REG2_REG_6__SCAN_IN), .ZN(n3347) );
  OAI211_X1 U4205 ( .C1(n3342), .C2(REG1_REG_6__SCAN_IN), .A(n3341), .B(n4710), 
        .ZN(n3346) );
  NOR2_X1 U4206 ( .A1(STATE_REG_SCAN_IN), .A2(n2264), .ZN(n3524) );
  NOR2_X1 U4207 ( .A1(n4715), .A2(n3343), .ZN(n3344) );
  AOI211_X1 U4208 ( .C1(n4709), .C2(ADDR_REG_6__SCAN_IN), .A(n3524), .B(n3344), 
        .ZN(n3345) );
  OAI211_X1 U4209 ( .C1(n3347), .C2(n4703), .A(n3346), .B(n3345), .ZN(U3246)
         );
  XNOR2_X1 U4210 ( .A(n3348), .B(REG2_REG_4__SCAN_IN), .ZN(n3357) );
  AOI211_X1 U4211 ( .C1(n4752), .C2(n3350), .A(n4199), .B(n3349), .ZN(n3355)
         );
  AND2_X1 U4212 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3460) );
  AOI21_X1 U4213 ( .B1(n4709), .B2(ADDR_REG_4__SCAN_IN), .A(n3460), .ZN(n3351)
         );
  OAI21_X1 U4214 ( .B1(n4715), .B2(n3352), .A(n3351), .ZN(n3353) );
  NOR3_X1 U4215 ( .A1(n3355), .A2(n3354), .A3(n3353), .ZN(n3356) );
  OAI21_X1 U4216 ( .B1(n3357), .B2(n4703), .A(n3356), .ZN(U3244) );
  INV_X1 U4217 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U4218 ( .A1(n4577), .A2(U4043), .ZN(n3358) );
  OAI21_X1 U4219 ( .B1(U4043), .B2(n4873), .A(n3358), .ZN(U3566) );
  INV_X1 U4220 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U4221 ( .A1(n4329), .A2(U4043), .ZN(n3359) );
  OAI21_X1 U4222 ( .B1(U4043), .B2(n4900), .A(n3359), .ZN(U3571) );
  INV_X1 U4223 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U4224 ( .A1(U4043), .A2(n3691), .ZN(n3360) );
  OAI21_X1 U4225 ( .B1(U4043), .B2(n4865), .A(n3360), .ZN(U3558) );
  INV_X1 U4226 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U4227 ( .A1(U4043), .A2(n3547), .ZN(n3361) );
  OAI21_X1 U4228 ( .B1(U4043), .B2(n4884), .A(n3361), .ZN(U3553) );
  INV_X1 U4229 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U4230 ( .A1(U4043), .A2(n4597), .ZN(n3362) );
  OAI21_X1 U4231 ( .B1(U4043), .B2(n4894), .A(n3362), .ZN(U3563) );
  INV_X1 U4232 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4874) );
  NAND2_X1 U4233 ( .A1(U4043), .A2(n3949), .ZN(n3363) );
  OAI21_X1 U4234 ( .B1(U4043), .B2(n4874), .A(n3363), .ZN(U3562) );
  INV_X1 U4235 ( .A(n3996), .ZN(n3406) );
  NAND2_X1 U4236 ( .A1(n3364), .A2(n4154), .ZN(n3995) );
  NAND2_X1 U4237 ( .A1(n3406), .A2(n3995), .ZN(n4721) );
  NAND2_X1 U4238 ( .A1(n4374), .A2(n4485), .ZN(n3366) );
  NOR2_X1 U4239 ( .A1(n3444), .A2(n4544), .ZN(n3365) );
  AOI21_X1 U4240 ( .B1(n4721), .B2(n3366), .A(n3365), .ZN(n4716) );
  NAND2_X1 U4241 ( .A1(n3432), .A2(n3367), .ZN(n4717) );
  INV_X1 U4242 ( .A(n4717), .ZN(n3368) );
  AOI21_X1 U4243 ( .B1(n4721), .B2(n4742), .A(n3368), .ZN(n3369) );
  AND2_X1 U4244 ( .A1(n4716), .A2(n3369), .ZN(n4737) );
  NAND2_X1 U4245 ( .A1(n4754), .A2(REG1_REG_0__SCAN_IN), .ZN(n3370) );
  OAI21_X1 U4246 ( .B1(n4754), .B2(n4737), .A(n3370), .ZN(U3518) );
  MUX2_X1 U4247 ( .A(n4796), .B(REG1_REG_7__SCAN_IN), .S(n3374), .Z(n3371) );
  XNOR2_X1 U4248 ( .A(n3372), .B(n3371), .ZN(n3381) );
  NOR2_X1 U4249 ( .A1(n3373), .A2(STATE_REG_SCAN_IN), .ZN(n3564) );
  NOR2_X1 U4250 ( .A1(n4715), .A2(n3374), .ZN(n3375) );
  AOI211_X1 U4251 ( .C1(n4709), .C2(ADDR_REG_7__SCAN_IN), .A(n3564), .B(n3375), 
        .ZN(n3380) );
  OAI211_X1 U4252 ( .C1(n3378), .C2(n3377), .A(n3376), .B(n4184), .ZN(n3379)
         );
  OAI211_X1 U4253 ( .C1(n3381), .C2(n4199), .A(n3380), .B(n3379), .ZN(U3247)
         );
  INV_X1 U4254 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U4255 ( .A1(n4355), .A2(U4043), .ZN(n3382) );
  OAI21_X1 U4256 ( .B1(U4043), .B2(n4917), .A(n3382), .ZN(U3572) );
  INV_X1 U4257 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U4258 ( .A1(U4043), .A2(n3525), .ZN(n3383) );
  OAI21_X1 U4259 ( .B1(U4043), .B2(n4880), .A(n3383), .ZN(U3557) );
  INV_X1 U4260 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U4261 ( .A1(U4043), .A2(n3596), .ZN(n3384) );
  OAI21_X1 U4262 ( .B1(U4043), .B2(n4918), .A(n3384), .ZN(U3556) );
  INV_X1 U4263 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U4264 ( .A1(U4043), .A2(n4576), .ZN(n3385) );
  OAI21_X1 U4265 ( .B1(U4043), .B2(n4866), .A(n3385), .ZN(U3564) );
  INV_X1 U4266 ( .A(n3554), .ZN(n3387) );
  OAI21_X1 U4267 ( .B1(n3399), .B2(n3446), .A(n3647), .ZN(n3386) );
  NAND2_X1 U4268 ( .A1(n3387), .A2(n3386), .ZN(n3651) );
  NAND2_X1 U4269 ( .A1(n3389), .A2(n3388), .ZN(n3542) );
  XNOR2_X1 U4270 ( .A(n3542), .B(n4077), .ZN(n3655) );
  OAI21_X1 U4271 ( .B1(n4077), .B2(n3391), .A(n3390), .ZN(n3393) );
  AOI22_X1 U4272 ( .A1(n3393), .A2(n4590), .B1(n4599), .B2(n3392), .ZN(n3646)
         );
  OAI22_X1 U4273 ( .A1(n2836), .A2(n4544), .B1(n3540), .B2(n4603), .ZN(n3394)
         );
  INV_X1 U4274 ( .A(n3394), .ZN(n3395) );
  OAI211_X1 U4275 ( .C1(n4744), .C2(n3655), .A(n3646), .B(n3395), .ZN(n3486)
         );
  NAND2_X1 U4276 ( .A1(n3486), .A2(n4751), .ZN(n3397) );
  NAND2_X1 U4277 ( .A1(n4749), .A2(REG0_REG_3__SCAN_IN), .ZN(n3396) );
  OAI211_X1 U4278 ( .C1(n3651), .C2(n4674), .A(n3397), .B(n3396), .ZN(U3473)
         );
  NAND2_X1 U4279 ( .A1(n3437), .A2(n3432), .ZN(n3398) );
  NAND2_X1 U4280 ( .A1(n3399), .A2(n3398), .ZN(n3574) );
  INV_X1 U4281 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3413) );
  OAI21_X1 U4282 ( .B1(n3401), .B2(n3403), .A(n3402), .ZN(n3572) );
  INV_X1 U4283 ( .A(n3572), .ZN(n3412) );
  AOI22_X1 U4284 ( .A1(n3392), .A2(n4598), .B1(n4599), .B2(n4154), .ZN(n3404)
         );
  OAI21_X1 U4285 ( .B1(n4603), .B2(n3571), .A(n3404), .ZN(n3411) );
  OR2_X1 U4286 ( .A1(n3572), .A2(n4374), .ZN(n3410) );
  NAND2_X1 U4287 ( .A1(n3406), .A2(n3401), .ZN(n3407) );
  NAND2_X1 U4288 ( .A1(n3405), .A2(n3407), .ZN(n3408) );
  NAND2_X1 U4289 ( .A1(n3408), .A2(n4590), .ZN(n3409) );
  NAND2_X1 U4290 ( .A1(n3410), .A2(n3409), .ZN(n3567) );
  AOI211_X1 U4291 ( .C1(n4742), .C2(n3412), .A(n3411), .B(n3567), .ZN(n3415)
         );
  MUX2_X1 U4292 ( .A(n3413), .B(n3415), .S(n4751), .Z(n3414) );
  OAI21_X1 U4293 ( .B1(n4674), .B2(n3574), .A(n3414), .ZN(U3469) );
  MUX2_X1 U4294 ( .A(n2886), .B(n3415), .S(n4756), .Z(n3416) );
  OAI21_X1 U4295 ( .B1(n4609), .B2(n3574), .A(n3416), .ZN(U3519) );
  INV_X1 U4296 ( .A(n3418), .ZN(n3419) );
  AOI21_X1 U4297 ( .B1(n3417), .B2(n3420), .A(n3419), .ZN(n3428) );
  INV_X1 U4298 ( .A(n3421), .ZN(n3424) );
  NAND3_X1 U4299 ( .A1(n3424), .A2(n3423), .A3(n3422), .ZN(n3429) );
  AOI22_X1 U4300 ( .A1(n3923), .A2(n3547), .B1(n3961), .B2(n4153), .ZN(n3425)
         );
  OAI21_X1 U4301 ( .B1(n2990), .B2(n3986), .A(n3425), .ZN(n3426) );
  AOI21_X1 U4302 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3429), .A(n3426), .ZN(n3427)
         );
  OAI21_X1 U4303 ( .B1(n3428), .B2(n3974), .A(n3427), .ZN(U3234) );
  INV_X1 U4304 ( .A(n3429), .ZN(n3443) );
  OAI22_X1 U4305 ( .A1(n3444), .A2(n3984), .B1(n3974), .B2(n3430), .ZN(n3431)
         );
  AOI21_X1 U4306 ( .B1(n3432), .B2(n3924), .A(n3431), .ZN(n3433) );
  OAI21_X1 U4307 ( .B1(n3443), .B2(n3434), .A(n3433), .ZN(U3229) );
  INV_X1 U4308 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U4309 ( .A1(n4293), .A2(U4043), .ZN(n3435) );
  OAI21_X1 U4310 ( .B1(U4043), .B2(n4881), .A(n3435), .ZN(U3573) );
  INV_X1 U4311 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4155) );
  OAI22_X1 U4312 ( .A1(n3575), .A2(n3988), .B1(n3984), .B2(n3573), .ZN(n3436)
         );
  AOI21_X1 U4313 ( .B1(n3437), .B2(n3924), .A(n3436), .ZN(n3442) );
  OAI211_X1 U4314 ( .C1(n3440), .C2(n3439), .A(n3981), .B(n3438), .ZN(n3441)
         );
  OAI211_X1 U4315 ( .C1(n3443), .C2(n4155), .A(n3442), .B(n3441), .ZN(U3219)
         );
  OAI22_X1 U4316 ( .A1(n3541), .A2(n4544), .B1(n3444), .B2(n4480), .ZN(n3445)
         );
  AOI21_X1 U4317 ( .B1(n4540), .B2(n3446), .A(n3445), .ZN(n3447) );
  INV_X1 U4318 ( .A(n3447), .ZN(n3449) );
  AOI211_X1 U4319 ( .C1(n4742), .C2(n3450), .A(n3449), .B(n3448), .ZN(n3496)
         );
  INV_X1 U4320 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3451) );
  OAI22_X1 U4321 ( .A1(n4674), .A2(n3498), .B1(n4751), .B2(n3451), .ZN(n3452)
         );
  INV_X1 U4322 ( .A(n3452), .ZN(n3453) );
  OAI21_X1 U4323 ( .B1(n3496), .B2(n4749), .A(n3453), .ZN(U3471) );
  INV_X1 U4324 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U4325 ( .A1(n4518), .A2(U4043), .ZN(n3454) );
  OAI21_X1 U4326 ( .B1(U4043), .B2(n4883), .A(n3454), .ZN(U3574) );
  AOI21_X1 U4327 ( .B1(n3455), .B2(n3456), .A(n3974), .ZN(n3458) );
  NAND2_X1 U4328 ( .A1(n3458), .A2(n3457), .ZN(n3462) );
  OAI22_X1 U4329 ( .A1(n3553), .A2(n3986), .B1(n3541), .B2(n3988), .ZN(n3459)
         );
  AOI211_X1 U4330 ( .C1(n3923), .C2(n4151), .A(n3460), .B(n3459), .ZN(n3461)
         );
  OAI211_X1 U4331 ( .C1(n3993), .C2(n3555), .A(n3462), .B(n3461), .ZN(U3227)
         );
  XNOR2_X1 U4332 ( .A(n3463), .B(REG1_REG_8__SCAN_IN), .ZN(n3470) );
  XNOR2_X1 U4333 ( .A(n3464), .B(n3615), .ZN(n3468) );
  AND2_X1 U4334 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3587) );
  AOI21_X1 U4335 ( .B1(n4709), .B2(ADDR_REG_8__SCAN_IN), .A(n3587), .ZN(n3465)
         );
  OAI21_X1 U4336 ( .B1(n4715), .B2(n3466), .A(n3465), .ZN(n3467) );
  AOI21_X1 U4337 ( .B1(n3468), .B2(n4184), .A(n3467), .ZN(n3469) );
  OAI21_X1 U4338 ( .B1(n3470), .B2(n4199), .A(n3469), .ZN(U3248) );
  OAI211_X1 U4339 ( .C1(n3473), .C2(n3472), .A(n3471), .B(n3981), .ZN(n3478)
         );
  OAI22_X1 U4340 ( .A1(n3986), .A2(n3474), .B1(n2836), .B2(n3988), .ZN(n3475)
         );
  AOI211_X1 U4341 ( .C1(n3923), .C2(n3596), .A(n3476), .B(n3475), .ZN(n3477)
         );
  OAI211_X1 U4342 ( .C1(n3993), .C2(n3479), .A(n3478), .B(n3477), .ZN(U3224)
         );
  XOR2_X1 U4343 ( .A(n3481), .B(n3480), .Z(n3485) );
  OAI22_X1 U4344 ( .A1(n3573), .A2(n3988), .B1(n3984), .B2(n2836), .ZN(n3483)
         );
  MUX2_X1 U4345 ( .A(n3972), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3482) );
  AOI211_X1 U4346 ( .C1(n3647), .C2(n3924), .A(n3483), .B(n3482), .ZN(n3484)
         );
  OAI21_X1 U4347 ( .B1(n3974), .B2(n3485), .A(n3484), .ZN(U3215) );
  NAND2_X1 U4348 ( .A1(n3486), .A2(n4756), .ZN(n3488) );
  NAND2_X1 U4349 ( .A1(n4754), .A2(REG1_REG_3__SCAN_IN), .ZN(n3487) );
  OAI211_X1 U4350 ( .C1(n4609), .C2(n3651), .A(n3488), .B(n3487), .ZN(U3521)
         );
  OAI22_X1 U4351 ( .A1(n3599), .A2(n4544), .B1(n2836), .B2(n4480), .ZN(n3489)
         );
  AOI21_X1 U4352 ( .B1(n4540), .B2(n3490), .A(n3489), .ZN(n3491) );
  OAI211_X1 U4353 ( .C1(n4744), .C2(n3493), .A(n3492), .B(n3491), .ZN(n3499)
         );
  NAND2_X1 U4354 ( .A1(n3499), .A2(n4751), .ZN(n3495) );
  NAND2_X1 U4355 ( .A1(n4749), .A2(REG0_REG_5__SCAN_IN), .ZN(n3494) );
  OAI211_X1 U4356 ( .C1(n3502), .C2(n4674), .A(n3495), .B(n3494), .ZN(U3477)
         );
  MUX2_X1 U4357 ( .A(n4944), .B(n3496), .S(n4756), .Z(n3497) );
  OAI21_X1 U4358 ( .B1(n3498), .B2(n4609), .A(n3497), .ZN(U3520) );
  NAND2_X1 U4359 ( .A1(n3499), .A2(n4756), .ZN(n3501) );
  NAND2_X1 U4360 ( .A1(n4754), .A2(REG1_REG_5__SCAN_IN), .ZN(n3500) );
  OAI211_X1 U4361 ( .C1(n4609), .C2(n3502), .A(n3501), .B(n3500), .ZN(U3523)
         );
  NAND2_X1 U4362 ( .A1(n4008), .A2(n4021), .ZN(n4085) );
  XNOR2_X1 U4363 ( .A(n3503), .B(n4085), .ZN(n3623) );
  OAI22_X1 U4364 ( .A1(n3632), .A2(n4544), .B1(n3630), .B2(n4480), .ZN(n3508)
         );
  NAND2_X1 U4365 ( .A1(n3252), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U4366 ( .A1(n3506), .A2(n3505), .ZN(n3597) );
  XNOR2_X1 U4367 ( .A(n3597), .B(n4085), .ZN(n3637) );
  NOR2_X1 U4368 ( .A1(n3637), .A2(n4744), .ZN(n3507) );
  AOI211_X1 U4369 ( .C1(n3595), .C2(n4540), .A(n3508), .B(n3507), .ZN(n3509)
         );
  OAI21_X1 U4370 ( .B1(n3623), .B2(n4485), .A(n3509), .ZN(n3514) );
  INV_X1 U4371 ( .A(n3514), .ZN(n3513) );
  INV_X1 U4372 ( .A(n4674), .ZN(n3511) );
  AND2_X1 U4373 ( .A1(n2439), .A2(n3595), .ZN(n3510) );
  NOR2_X1 U4374 ( .A1(n2160), .A2(n3510), .ZN(n3624) );
  INV_X1 U4375 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U4376 ( .A1(n3511), .A2(n3624), .B1(n4749), .B2(REG0_REG_6__SCAN_IN), .ZN(n3512) );
  OAI21_X1 U4377 ( .B1(n3513), .B2(n4749), .A(n3512), .ZN(U3479) );
  NAND2_X1 U4378 ( .A1(n3514), .A2(n4756), .ZN(n3517) );
  INV_X1 U4379 ( .A(n4609), .ZN(n3515) );
  NAND2_X1 U4380 ( .A1(n3515), .A2(n3624), .ZN(n3516) );
  OAI211_X1 U4381 ( .C1(n4756), .C2(n5004), .A(n3517), .B(n3516), .ZN(U3524)
         );
  XNOR2_X1 U4382 ( .A(n3519), .B(n3518), .ZN(n3520) );
  XNOR2_X1 U4383 ( .A(n3521), .B(n3520), .ZN(n3522) );
  NAND2_X1 U4384 ( .A1(n3522), .A2(n3981), .ZN(n3527) );
  OAI22_X1 U4385 ( .A1(n3986), .A2(n3631), .B1(n3630), .B2(n3988), .ZN(n3523)
         );
  AOI211_X1 U4386 ( .C1(n3923), .C2(n3525), .A(n3524), .B(n3523), .ZN(n3526)
         );
  OAI211_X1 U4387 ( .C1(n3993), .C2(n3625), .A(n3527), .B(n3526), .ZN(U3236)
         );
  XNOR2_X1 U4388 ( .A(n3529), .B(n3528), .ZN(n3538) );
  AOI21_X1 U4389 ( .B1(n3531), .B2(n3530), .A(n4199), .ZN(n3536) );
  NOR2_X1 U4390 ( .A1(n4823), .A2(STATE_REG_SCAN_IN), .ZN(n3687) );
  AOI21_X1 U4391 ( .B1(n4709), .B2(ADDR_REG_9__SCAN_IN), .A(n3687), .ZN(n3532)
         );
  OAI21_X1 U4392 ( .B1(n4715), .B2(n3533), .A(n3532), .ZN(n3534) );
  AOI21_X1 U4393 ( .B1(n3536), .B2(n3535), .A(n3534), .ZN(n3537) );
  OAI21_X1 U4394 ( .B1(n3538), .B2(n4703), .A(n3537), .ZN(U3249) );
  INV_X1 U4395 ( .A(n3542), .ZN(n3544) );
  OAI21_X1 U4396 ( .B1(n3542), .B2(n3541), .A(n3540), .ZN(n3543) );
  OAI21_X1 U4397 ( .B1(n3544), .B2(n3547), .A(n3543), .ZN(n3545) );
  XOR2_X1 U4398 ( .A(n4087), .B(n3545), .Z(n3557) );
  XOR2_X1 U4399 ( .A(n4087), .B(n3546), .Z(n3550) );
  AOI22_X1 U4400 ( .A1(n4598), .A2(n4151), .B1(n3547), .B2(n4599), .ZN(n3548)
         );
  OAI21_X1 U4401 ( .B1(n4603), .B2(n3553), .A(n3548), .ZN(n3549) );
  AOI21_X1 U4402 ( .B1(n3550), .B2(n4590), .A(n3549), .ZN(n3551) );
  OAI21_X1 U4403 ( .B1(n3557), .B2(n4374), .A(n3551), .ZN(n4739) );
  OAI211_X1 U4404 ( .C1(n3554), .C2(n3553), .A(n3552), .B(n4611), .ZN(n4738)
         );
  OAI22_X1 U4405 ( .A1(n4738), .A2(n4681), .B1(n4492), .B2(n3555), .ZN(n3556)
         );
  OAI21_X1 U4406 ( .B1(n4739), .B2(n3556), .A(n4724), .ZN(n3559) );
  INV_X1 U4407 ( .A(n3557), .ZN(n4741) );
  INV_X1 U4408 ( .A(n4385), .ZN(n4722) );
  AOI22_X1 U4409 ( .A1(n4741), .A2(n4722), .B1(REG2_REG_4__SCAN_IN), .B2(n4726), .ZN(n3558) );
  NAND2_X1 U4410 ( .A1(n3559), .A2(n3558), .ZN(U3286) );
  XOR2_X1 U4411 ( .A(n3560), .B(n3561), .Z(n3562) );
  NAND2_X1 U4412 ( .A1(n3562), .A2(n3981), .ZN(n3566) );
  OAI22_X1 U4413 ( .A1(n3986), .A2(n3592), .B1(n3599), .B2(n3988), .ZN(n3563)
         );
  AOI211_X1 U4414 ( .C1(n3923), .C2(n3691), .A(n3564), .B(n3563), .ZN(n3565)
         );
  OAI211_X1 U4415 ( .C1(n3993), .C2(n3603), .A(n3566), .B(n3565), .ZN(U3210)
         );
  INV_X1 U4416 ( .A(n4492), .ZN(n4720) );
  AOI22_X1 U4417 ( .A1(n4724), .A2(n3567), .B1(REG3_REG_1__SCAN_IN), .B2(n4720), .ZN(n3570) );
  OR2_X1 U4418 ( .A1(n4724), .A2(n3568), .ZN(n3569) );
  OAI211_X1 U4419 ( .C1(n4468), .C2(n3571), .A(n3570), .B(n3569), .ZN(n3578)
         );
  OAI22_X1 U4420 ( .A1(n3573), .A2(n4451), .B1(n4385), .B2(n3572), .ZN(n3577)
         );
  OAI22_X1 U4421 ( .A1(n3575), .A2(n4469), .B1(n4498), .B2(n3574), .ZN(n3576)
         );
  OR3_X1 U4422 ( .A1(n3578), .A2(n3577), .A3(n3576), .ZN(U3289) );
  INV_X1 U4423 ( .A(n3580), .ZN(n3582) );
  NAND2_X1 U4424 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  XNOR2_X1 U4425 ( .A(n3579), .B(n3583), .ZN(n3584) );
  NAND2_X1 U4426 ( .A1(n3584), .A2(n3981), .ZN(n3589) );
  OAI22_X1 U4427 ( .A1(n3986), .A2(n3585), .B1(n3632), .B2(n3988), .ZN(n3586)
         );
  AOI211_X1 U4428 ( .C1(n3923), .C2(n4150), .A(n3587), .B(n3586), .ZN(n3588)
         );
  OAI211_X1 U4429 ( .C1(n3993), .C2(n3614), .A(n3589), .B(n3588), .ZN(U3218)
         );
  OAI211_X1 U4430 ( .C1(n2160), .C2(n3592), .A(n3617), .B(n4611), .ZN(n4747)
         );
  INV_X1 U4431 ( .A(n2844), .ZN(n4009) );
  XNOR2_X1 U4432 ( .A(n3590), .B(n4009), .ZN(n3594) );
  AOI22_X1 U4433 ( .A1(n3691), .A2(n4598), .B1(n4599), .B2(n3596), .ZN(n3591)
         );
  OAI21_X1 U4434 ( .B1(n4603), .B2(n3592), .A(n3591), .ZN(n3593) );
  AOI21_X1 U4435 ( .B1(n3594), .B2(n4590), .A(n3593), .ZN(n4748) );
  OAI21_X1 U4436 ( .B1(n4681), .B2(n4747), .A(n4748), .ZN(n3606) );
  INV_X1 U4437 ( .A(n3597), .ZN(n3600) );
  AOI21_X1 U4438 ( .B1(n3597), .B2(n3596), .A(n3595), .ZN(n3598) );
  AOI21_X1 U4439 ( .B1(n3600), .B2(n3599), .A(n3598), .ZN(n3601) );
  NOR2_X1 U4440 ( .A1(n3601), .A2(n2844), .ZN(n4745) );
  INV_X1 U4441 ( .A(n3601), .ZN(n3602) );
  NOR2_X1 U4442 ( .A1(n3602), .A2(n4009), .ZN(n4743) );
  NOR3_X1 U4443 ( .A1(n4745), .A2(n4743), .A3(n4456), .ZN(n3605) );
  OAI22_X1 U4444 ( .A1(n4724), .A2(n2941), .B1(n3603), .B2(n4492), .ZN(n3604)
         );
  AOI211_X1 U4445 ( .C1(n3606), .C2(n4724), .A(n3605), .B(n3604), .ZN(n3607)
         );
  INV_X1 U4446 ( .A(n3607), .ZN(U3283) );
  NAND2_X1 U4447 ( .A1(n4013), .A2(n4011), .ZN(n4086) );
  XNOR2_X1 U4448 ( .A(n3608), .B(n4086), .ZN(n3613) );
  XNOR2_X1 U4449 ( .A(n3609), .B(n4086), .ZN(n4615) );
  OAI22_X1 U4450 ( .A1(n3632), .A2(n4480), .B1(n3713), .B2(n4544), .ZN(n3610)
         );
  AOI21_X1 U4451 ( .B1(n4540), .B2(n3616), .A(n3610), .ZN(n3611) );
  OAI21_X1 U4452 ( .B1(n4615), .B2(n4374), .A(n3611), .ZN(n3612) );
  AOI21_X1 U4453 ( .B1(n3613), .B2(n4590), .A(n3612), .ZN(n4613) );
  INV_X1 U4454 ( .A(n4615), .ZN(n3620) );
  OAI22_X1 U4455 ( .A1(n4724), .A2(n3615), .B1(n3614), .B2(n4492), .ZN(n3619)
         );
  NAND2_X1 U4456 ( .A1(n3617), .A2(n3616), .ZN(n4610) );
  AND3_X1 U4457 ( .A1(n4459), .A2(n2449), .A3(n4610), .ZN(n3618) );
  AOI211_X1 U4458 ( .C1(n3620), .C2(n4722), .A(n3619), .B(n3618), .ZN(n3621)
         );
  OAI21_X1 U4459 ( .B1(n4613), .B2(n4726), .A(n3621), .ZN(U3282) );
  INV_X1 U4460 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U4461 ( .A1(n3868), .A2(U4043), .ZN(n3622) );
  OAI21_X1 U4462 ( .B1(U4043), .B2(n4869), .A(n3622), .ZN(U3578) );
  NAND2_X1 U4463 ( .A1(n4724), .A2(n4590), .ZN(n3766) );
  OR2_X1 U4464 ( .A1(n3623), .A2(n3766), .ZN(n3636) );
  NAND2_X1 U4465 ( .A1(n4459), .A2(n3624), .ZN(n3629) );
  OAI22_X1 U4466 ( .A1(n4724), .A2(n3626), .B1(n3625), .B2(n4492), .ZN(n3627)
         );
  INV_X1 U4467 ( .A(n3627), .ZN(n3628) );
  OAI211_X1 U4468 ( .C1(n3630), .C2(n4469), .A(n3629), .B(n3628), .ZN(n3634)
         );
  OAI22_X1 U4469 ( .A1(n3632), .A2(n4451), .B1(n4468), .B2(n3631), .ZN(n3633)
         );
  NOR2_X1 U4470 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  OAI211_X1 U4471 ( .C1(n4456), .C2(n3637), .A(n3636), .B(n3635), .ZN(U3284)
         );
  XNOR2_X1 U4472 ( .A(n3638), .B(REG1_REG_10__SCAN_IN), .ZN(n3645) );
  XOR2_X1 U4473 ( .A(REG2_REG_10__SCAN_IN), .B(n3639), .Z(n3643) );
  AND2_X1 U4474 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3706) );
  AOI21_X1 U4475 ( .B1(n4709), .B2(ADDR_REG_10__SCAN_IN), .A(n3706), .ZN(n3640) );
  OAI21_X1 U4476 ( .B1(n4715), .B2(n3641), .A(n3640), .ZN(n3642) );
  AOI21_X1 U4477 ( .B1(n3643), .B2(n4184), .A(n3642), .ZN(n3644) );
  OAI21_X1 U4478 ( .B1(n3645), .B2(n4199), .A(n3644), .ZN(U3250) );
  INV_X1 U4479 ( .A(n3646), .ZN(n3653) );
  INV_X1 U4480 ( .A(n4468), .ZN(n4445) );
  INV_X1 U4481 ( .A(n4451), .ZN(n4472) );
  AOI22_X1 U4482 ( .A1(n4445), .A2(n3647), .B1(n4472), .B2(n4152), .ZN(n3650)
         );
  AOI22_X1 U4483 ( .A1(n4726), .A2(REG2_REG_3__SCAN_IN), .B1(n4720), .B2(n3648), .ZN(n3649) );
  OAI211_X1 U4484 ( .C1(n4498), .C2(n3651), .A(n3650), .B(n3649), .ZN(n3652)
         );
  AOI21_X1 U4485 ( .B1(n4724), .B2(n3653), .A(n3652), .ZN(n3654) );
  OAI21_X1 U4486 ( .B1(n4456), .B2(n3655), .A(n3654), .ZN(U3287) );
  NAND2_X1 U4487 ( .A1(n4014), .A2(n4020), .ZN(n4089) );
  XOR2_X1 U4488 ( .A(n3656), .B(n4089), .Z(n3657) );
  NOR2_X1 U4489 ( .A1(n3657), .A2(n4485), .ZN(n3694) );
  INV_X1 U4490 ( .A(n3694), .ZN(n3667) );
  XOR2_X1 U4491 ( .A(n3658), .B(n4089), .Z(n3696) );
  AND2_X1 U4492 ( .A1(n2449), .A2(n3659), .ZN(n3660) );
  OR2_X1 U4493 ( .A1(n3660), .A2(n3671), .ZN(n3712) );
  OAI22_X1 U4494 ( .A1(n4724), .A2(n3661), .B1(n3690), .B2(n4492), .ZN(n3663)
         );
  OAI22_X1 U4495 ( .A1(n3685), .A2(n4469), .B1(n4468), .B2(n3693), .ZN(n3662)
         );
  AOI211_X1 U4496 ( .C1(n4472), .C2(n4149), .A(n3663), .B(n3662), .ZN(n3664)
         );
  OAI21_X1 U4497 ( .B1(n4498), .B2(n3712), .A(n3664), .ZN(n3665) );
  AOI21_X1 U4498 ( .B1(n4501), .B2(n3696), .A(n3665), .ZN(n3666) );
  OAI21_X1 U4499 ( .B1(n3667), .B2(n4726), .A(n3666), .ZN(U3281) );
  NAND2_X1 U4500 ( .A1(n4026), .A2(n4030), .ZN(n4082) );
  XOR2_X1 U4501 ( .A(n3668), .B(n4082), .Z(n3719) );
  INV_X1 U4502 ( .A(n3719), .ZN(n3681) );
  INV_X1 U4503 ( .A(n4082), .ZN(n3670) );
  XNOR2_X1 U4504 ( .A(n3669), .B(n3670), .ZN(n3717) );
  INV_X1 U4505 ( .A(n3717), .ZN(n3679) );
  NOR2_X1 U4506 ( .A1(n3671), .A2(n3704), .ZN(n3672) );
  OR2_X1 U4507 ( .A1(n3748), .A2(n3672), .ZN(n3725) );
  OAI22_X1 U4508 ( .A1(n4724), .A2(n3673), .B1(n3709), .B2(n4492), .ZN(n3674)
         );
  AOI21_X1 U4509 ( .B1(n3715), .B2(n4445), .A(n3674), .ZN(n3677) );
  OAI22_X1 U4510 ( .A1(n3713), .A2(n4469), .B1(n4451), .B2(n3732), .ZN(n3675)
         );
  INV_X1 U4511 ( .A(n3675), .ZN(n3676) );
  OAI211_X1 U4512 ( .C1(n3725), .C2(n4498), .A(n3677), .B(n3676), .ZN(n3678)
         );
  AOI21_X1 U4513 ( .B1(n4501), .B2(n3679), .A(n3678), .ZN(n3680) );
  OAI21_X1 U4514 ( .B1(n3681), .B2(n3766), .A(n3680), .ZN(U3280) );
  XNOR2_X1 U4515 ( .A(n3682), .B(n3683), .ZN(n3684) );
  NAND2_X1 U4516 ( .A1(n3684), .A2(n3981), .ZN(n3689) );
  OAI22_X1 U4517 ( .A1(n3986), .A2(n3693), .B1(n3685), .B2(n3988), .ZN(n3686)
         );
  AOI211_X1 U4518 ( .C1(n3923), .C2(n4149), .A(n3687), .B(n3686), .ZN(n3688)
         );
  OAI211_X1 U4519 ( .C1(n3993), .C2(n3690), .A(n3689), .B(n3688), .ZN(U3228)
         );
  AOI22_X1 U4520 ( .A1(n3691), .A2(n4599), .B1(n4598), .B2(n4149), .ZN(n3692)
         );
  OAI21_X1 U4521 ( .B1(n4603), .B2(n3693), .A(n3692), .ZN(n3695) );
  AOI211_X1 U4522 ( .C1(n3696), .C2(n4607), .A(n3695), .B(n3694), .ZN(n3710)
         );
  INV_X1 U4523 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3697) );
  OAI22_X1 U4524 ( .A1(n3712), .A2(n4674), .B1(n4751), .B2(n3697), .ZN(n3698)
         );
  INV_X1 U4525 ( .A(n3698), .ZN(n3699) );
  OAI21_X1 U4526 ( .B1(n3710), .B2(n4749), .A(n3699), .ZN(U3485) );
  AOI21_X1 U4527 ( .B1(n3700), .B2(n3701), .A(n3974), .ZN(n3703) );
  NAND2_X1 U4528 ( .A1(n3703), .A2(n3702), .ZN(n3708) );
  OAI22_X1 U4529 ( .A1(n3986), .A2(n3704), .B1(n3732), .B2(n3984), .ZN(n3705)
         );
  AOI211_X1 U4530 ( .C1(n3961), .C2(n4150), .A(n3706), .B(n3705), .ZN(n3707)
         );
  OAI211_X1 U4531 ( .C1(n3993), .C2(n3709), .A(n3708), .B(n3707), .ZN(U3214)
         );
  MUX2_X1 U4532 ( .A(n2897), .B(n3710), .S(n4756), .Z(n3711) );
  OAI21_X1 U4533 ( .B1(n4609), .B2(n3712), .A(n3711), .ZN(U3527) );
  INV_X1 U4534 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3720) );
  OAI22_X1 U4535 ( .A1(n3713), .A2(n4480), .B1(n3732), .B2(n4544), .ZN(n3714)
         );
  AOI21_X1 U4536 ( .B1(n4540), .B2(n3715), .A(n3714), .ZN(n3716) );
  OAI21_X1 U4537 ( .B1(n3717), .B2(n4744), .A(n3716), .ZN(n3718) );
  AOI21_X1 U4538 ( .B1(n3719), .B2(n4590), .A(n3718), .ZN(n3722) );
  MUX2_X1 U4539 ( .A(n3720), .B(n3722), .S(n4751), .Z(n3721) );
  OAI21_X1 U4540 ( .B1(n3725), .B2(n4674), .A(n3721), .ZN(U3487) );
  INV_X1 U4541 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3723) );
  MUX2_X1 U4542 ( .A(n3723), .B(n3722), .S(n4756), .Z(n3724) );
  OAI21_X1 U4543 ( .B1(n4609), .B2(n3725), .A(n3724), .ZN(U3528) );
  INV_X1 U4544 ( .A(n4477), .ZN(n3727) );
  NOR2_X1 U4545 ( .A1(n4478), .A2(n3727), .ZN(n4081) );
  XOR2_X1 U4546 ( .A(n3726), .B(n4081), .Z(n3728) );
  NOR2_X1 U4547 ( .A1(n3728), .A2(n4485), .ZN(n4604) );
  INV_X1 U4548 ( .A(n4604), .ZN(n3738) );
  NAND2_X1 U4549 ( .A1(n4488), .A2(n3729), .ZN(n3730) );
  XOR2_X1 U4550 ( .A(n3730), .B(n4081), .Z(n4606) );
  INV_X1 U4551 ( .A(n3747), .ZN(n3731) );
  OAI21_X1 U4552 ( .B1(n3731), .B2(n4602), .A(n4496), .ZN(n4675) );
  OAI22_X1 U4553 ( .A1(n4724), .A2(n3789), .B1(n3808), .B2(n4492), .ZN(n3734)
         );
  OAI22_X1 U4554 ( .A1(n3732), .A2(n4469), .B1(n4468), .B2(n4602), .ZN(n3733)
         );
  AOI211_X1 U4555 ( .C1(n4472), .C2(n4597), .A(n3734), .B(n3733), .ZN(n3735)
         );
  OAI21_X1 U4556 ( .B1(n4675), .B2(n4498), .A(n3735), .ZN(n3736) );
  AOI21_X1 U4557 ( .B1(n4606), .B2(n4501), .A(n3736), .ZN(n3737) );
  OAI21_X1 U4558 ( .B1(n3738), .B2(n4726), .A(n3737), .ZN(U3278) );
  OAI21_X1 U4559 ( .B1(n3739), .B2(n4088), .A(n4488), .ZN(n3782) );
  INV_X1 U4560 ( .A(n3782), .ZN(n3753) );
  XNOR2_X1 U4561 ( .A(n3740), .B(n4088), .ZN(n3744) );
  OAI22_X1 U4562 ( .A1(n4603), .A2(n3774), .B1(n4481), .B2(n4544), .ZN(n3741)
         );
  AOI21_X1 U4563 ( .B1(n3782), .B2(n3742), .A(n3741), .ZN(n3743) );
  OAI21_X1 U4564 ( .B1(n3744), .B2(n4485), .A(n3743), .ZN(n3780) );
  INV_X1 U4565 ( .A(n3780), .ZN(n3745) );
  MUX2_X1 U4566 ( .A(n3746), .B(n3745), .S(n4724), .Z(n3752) );
  OAI21_X1 U4567 ( .B1(n3748), .B2(n3774), .A(n3747), .ZN(n3787) );
  INV_X1 U4568 ( .A(n3787), .ZN(n3750) );
  OAI22_X1 U4569 ( .A1(n4469), .A2(n3779), .B1(n3778), .B2(n4492), .ZN(n3749)
         );
  AOI21_X1 U4570 ( .B1(n3750), .B2(n4459), .A(n3749), .ZN(n3751) );
  OAI211_X1 U4571 ( .C1(n3753), .C2(n4385), .A(n3752), .B(n3751), .ZN(U3279)
         );
  XNOR2_X1 U4572 ( .A(n3754), .B(n4079), .ZN(n4591) );
  INV_X1 U4573 ( .A(n4591), .ZN(n3767) );
  OAI21_X1 U4574 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n4584) );
  INV_X1 U4575 ( .A(n4465), .ZN(n3758) );
  OAI21_X1 U4576 ( .B1(n2181), .B2(n4588), .A(n3758), .ZN(n4666) );
  OAI22_X1 U4577 ( .A1(n4724), .A2(n3759), .B1(n3879), .B2(n4492), .ZN(n3761)
         );
  OAI22_X1 U4578 ( .A1(n3875), .A2(n4451), .B1(n4469), .B2(n3803), .ZN(n3760)
         );
  AOI211_X1 U4579 ( .C1(n3762), .C2(n4445), .A(n3761), .B(n3760), .ZN(n3763)
         );
  OAI21_X1 U4580 ( .B1(n4666), .B2(n4498), .A(n3763), .ZN(n3764) );
  AOI21_X1 U4581 ( .B1(n4584), .B2(n4501), .A(n3764), .ZN(n3765) );
  OAI21_X1 U4582 ( .B1(n3767), .B2(n3766), .A(n3765), .ZN(U3276) );
  XNOR2_X1 U4583 ( .A(n3769), .B(n3768), .ZN(n3770) );
  XNOR2_X1 U4584 ( .A(n3771), .B(n3770), .ZN(n3772) );
  NAND2_X1 U4585 ( .A1(n3772), .A2(n3981), .ZN(n3777) );
  NOR2_X1 U4586 ( .A1(n3773), .A2(STATE_REG_SCAN_IN), .ZN(n4173) );
  OAI22_X1 U4587 ( .A1(n3986), .A2(n3774), .B1(n4481), .B2(n3984), .ZN(n3775)
         );
  AOI211_X1 U4588 ( .C1(n3961), .C2(n4149), .A(n4173), .B(n3775), .ZN(n3776)
         );
  OAI211_X1 U4589 ( .C1(n3993), .C2(n3778), .A(n3777), .B(n3776), .ZN(U3233)
         );
  INV_X1 U4590 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3783) );
  NOR2_X1 U4591 ( .A1(n3779), .A2(n4480), .ZN(n3781) );
  AOI211_X1 U4592 ( .C1(n4742), .C2(n3782), .A(n3781), .B(n3780), .ZN(n3785)
         );
  MUX2_X1 U4593 ( .A(n3783), .B(n3785), .S(n4751), .Z(n3784) );
  OAI21_X1 U4594 ( .B1(n3787), .B2(n4674), .A(n3784), .ZN(U3489) );
  MUX2_X1 U4595 ( .A(n4940), .B(n3785), .S(n4756), .Z(n3786) );
  OAI21_X1 U4596 ( .B1(n4609), .B2(n3787), .A(n3786), .ZN(U3529) );
  XNOR2_X1 U4597 ( .A(n3788), .B(REG1_REG_12__SCAN_IN), .ZN(n3796) );
  XNOR2_X1 U4598 ( .A(n3790), .B(n3789), .ZN(n3794) );
  AND2_X1 U4599 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3805) );
  AOI21_X1 U4600 ( .B1(n4709), .B2(ADDR_REG_12__SCAN_IN), .A(n3805), .ZN(n3791) );
  OAI21_X1 U4601 ( .B1(n4715), .B2(n3792), .A(n3791), .ZN(n3793) );
  AOI21_X1 U4602 ( .B1(n3794), .B2(n4184), .A(n3793), .ZN(n3795) );
  OAI21_X1 U4603 ( .B1(n3796), .B2(n4199), .A(n3795), .ZN(U3252) );
  INV_X1 U4604 ( .A(n3798), .ZN(n3800) );
  NAND2_X1 U4605 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  XNOR2_X1 U4606 ( .A(n3797), .B(n3801), .ZN(n3802) );
  NAND2_X1 U4607 ( .A1(n3802), .A2(n3981), .ZN(n3807) );
  OAI22_X1 U4608 ( .A1(n3986), .A2(n4602), .B1(n3803), .B2(n3984), .ZN(n3804)
         );
  AOI211_X1 U4609 ( .C1(n3961), .C2(n4600), .A(n3805), .B(n3804), .ZN(n3806)
         );
  OAI211_X1 U4610 ( .C1(n3993), .C2(n3808), .A(n3807), .B(n3806), .ZN(U3221)
         );
  XNOR2_X1 U4611 ( .A(n4684), .B(n4494), .ZN(n3809) );
  XNOR2_X1 U4612 ( .A(n3810), .B(n3809), .ZN(n3819) );
  AOI21_X1 U4613 ( .B1(n3812), .B2(n3811), .A(n4199), .ZN(n3817) );
  AND2_X1 U4614 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3948) );
  AOI21_X1 U4615 ( .B1(n4709), .B2(ADDR_REG_13__SCAN_IN), .A(n3948), .ZN(n3813) );
  OAI21_X1 U4616 ( .B1(n4715), .B2(n3814), .A(n3813), .ZN(n3815) );
  AOI21_X1 U4617 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3818) );
  OAI21_X1 U4618 ( .B1(n4703), .B2(n3819), .A(n3818), .ZN(U3253) );
  INV_X1 U4619 ( .A(n3820), .ZN(n3821) );
  NAND2_X1 U4620 ( .A1(n3883), .A2(n3821), .ZN(n3849) );
  NAND2_X1 U4621 ( .A1(n3849), .A2(n3850), .ZN(n3826) );
  XNOR2_X1 U4622 ( .A(n3826), .B(n3825), .ZN(n3827) );
  NAND2_X1 U4623 ( .A1(n3827), .A2(n3981), .ZN(n3831) );
  OAI22_X1 U4624 ( .A1(n4332), .A2(n3988), .B1(n3986), .B2(n4298), .ZN(n3829)
         );
  OAI22_X1 U4625 ( .A1(n5037), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n2256), 
        .ZN(n3828) );
  AOI211_X1 U4626 ( .C1(n4299), .C2(n3972), .A(n3829), .B(n3828), .ZN(n3830)
         );
  NAND2_X1 U4627 ( .A1(n3831), .A2(n3830), .ZN(U3226) );
  AND2_X1 U4628 ( .A1(n3832), .A2(DATAI_30_), .ZN(n4218) );
  NAND2_X1 U4629 ( .A1(n3832), .A2(DATAI_31_), .ZN(n4132) );
  XNOR2_X1 U4630 ( .A(n4216), .B(n4132), .ZN(n3846) );
  INV_X1 U4631 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U4632 ( .A1(n3833), .A2(REG0_REG_31__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4633 ( .A1(n3834), .A2(REG1_REG_31__SCAN_IN), .ZN(n3835) );
  OAI211_X1 U4634 ( .C1(n3837), .C2(n4986), .A(n3836), .B(n3835), .ZN(n4145)
         );
  NAND2_X1 U4635 ( .A1(n3838), .A2(n4145), .ZN(n4220) );
  OAI21_X1 U4636 ( .B1(n4132), .B2(n4603), .A(n4220), .ZN(n3843) );
  NAND2_X1 U4637 ( .A1(n4751), .A2(n3843), .ZN(n3840) );
  NAND2_X1 U4638 ( .A1(n4749), .A2(REG0_REG_31__SCAN_IN), .ZN(n3839) );
  OAI211_X1 U4639 ( .C1(n3846), .C2(n4674), .A(n3840), .B(n3839), .ZN(U3517)
         );
  NAND2_X1 U4640 ( .A1(n4756), .A2(n3843), .ZN(n3842) );
  NAND2_X1 U4641 ( .A1(n4754), .A2(REG1_REG_31__SCAN_IN), .ZN(n3841) );
  OAI211_X1 U4642 ( .C1(n3846), .C2(n4609), .A(n3842), .B(n3841), .ZN(U3549)
         );
  NAND2_X1 U4643 ( .A1(n4724), .A2(n3843), .ZN(n3845) );
  NAND2_X1 U4644 ( .A1(n4726), .A2(REG2_REG_31__SCAN_IN), .ZN(n3844) );
  OAI211_X1 U4645 ( .C1(n3846), .C2(n4498), .A(n3845), .B(n3844), .ZN(U3260)
         );
  INV_X1 U4646 ( .A(IR_REG_30__SCAN_IN), .ZN(n4849) );
  NAND3_X1 U4647 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4849), 
        .ZN(n3848) );
  INV_X1 U4648 ( .A(DATAI_31_), .ZN(n5019) );
  OAI22_X1 U4649 ( .A1(n3847), .A2(n3848), .B1(STATE_REG_SCAN_IN), .B2(n5019), 
        .ZN(U3321) );
  INV_X1 U4650 ( .A(n3849), .ZN(n3852) );
  OAI21_X1 U4651 ( .B1(n3852), .B2(n3851), .A(n3850), .ZN(n3857) );
  OAI21_X1 U4652 ( .B1(n3855), .B2(n3854), .A(n3853), .ZN(n3856) );
  XNOR2_X1 U4653 ( .A(n3857), .B(n3856), .ZN(n3858) );
  NAND2_X1 U4654 ( .A1(n3858), .A2(n3981), .ZN(n3862) );
  OAI22_X1 U4655 ( .A1(n4312), .A2(n3988), .B1(n3986), .B2(n4280), .ZN(n3860)
         );
  INV_X1 U4656 ( .A(n4508), .ZN(n4521) );
  OAI22_X1 U4657 ( .A1(n4521), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n4997), 
        .ZN(n3859) );
  AOI211_X1 U4658 ( .C1(n4278), .C2(n3972), .A(n3860), .B(n3859), .ZN(n3861)
         );
  NAND2_X1 U4659 ( .A1(n3862), .A2(n3861), .ZN(U3222) );
  XNOR2_X1 U4660 ( .A(n3864), .B(n3863), .ZN(n3870) );
  NOR2_X1 U4661 ( .A1(n4245), .A2(n3993), .ZN(n3867) );
  AOI22_X1 U4662 ( .A1(n4508), .A2(n3961), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3865) );
  OAI21_X1 U4663 ( .B1(n3986), .B2(n4246), .A(n3865), .ZN(n3866) );
  AOI211_X1 U4664 ( .C1(n3923), .C2(n3868), .A(n3867), .B(n3866), .ZN(n3869)
         );
  OAI21_X1 U4665 ( .B1(n3870), .B2(n3974), .A(n3869), .ZN(U3211) );
  NOR2_X1 U4666 ( .A1(n2192), .A2(n3872), .ZN(n3873) );
  XNOR2_X1 U4667 ( .A(n3871), .B(n3873), .ZN(n3874) );
  NAND2_X1 U4668 ( .A1(n3874), .A2(n3981), .ZN(n3878) );
  AND2_X1 U4669 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4183) );
  OAI22_X1 U4670 ( .A1(n3986), .A2(n4588), .B1(n3875), .B2(n3984), .ZN(n3876)
         );
  AOI211_X1 U4671 ( .C1(n3961), .C2(n4597), .A(n4183), .B(n3876), .ZN(n3877)
         );
  OAI211_X1 U4672 ( .C1(n3993), .C2(n3879), .A(n3878), .B(n3877), .ZN(U3212)
         );
  INV_X1 U4673 ( .A(n3262), .ZN(n3882) );
  OAI21_X1 U4674 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3884) );
  NAND3_X1 U4675 ( .A1(n3884), .A2(n3981), .A3(n3883), .ZN(n3890) );
  OAI22_X1 U4676 ( .A1(n4312), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n3885), 
        .ZN(n3888) );
  OAI22_X1 U4677 ( .A1(n3986), .A2(n3886), .B1(n4545), .B2(n3988), .ZN(n3887)
         );
  NOR2_X1 U4678 ( .A1(n3888), .A2(n3887), .ZN(n3889) );
  OAI211_X1 U4679 ( .C1(n3993), .C2(n4319), .A(n3890), .B(n3889), .ZN(U3213)
         );
  XOR2_X1 U4680 ( .A(n3892), .B(n3891), .Z(n3896) );
  INV_X1 U4681 ( .A(n4541), .ZN(n4396) );
  AOI22_X1 U4682 ( .A1(n3924), .A2(n4393), .B1(n3961), .B2(n4561), .ZN(n3893)
         );
  NAND2_X1 U4683 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4210) );
  OAI211_X1 U4684 ( .C1(n4396), .C2(n3984), .A(n3893), .B(n4210), .ZN(n3894)
         );
  AOI21_X1 U4685 ( .B1(n4401), .B2(n3972), .A(n3894), .ZN(n3895) );
  OAI21_X1 U4686 ( .B1(n3896), .B2(n3974), .A(n3895), .ZN(U3216) );
  XNOR2_X1 U4687 ( .A(n3899), .B(n3898), .ZN(n3900) );
  XNOR2_X1 U4688 ( .A(n3897), .B(n3900), .ZN(n3905) );
  OAI22_X1 U4689 ( .A1(n4545), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n3901), 
        .ZN(n3903) );
  OAI22_X1 U4690 ( .A1(n3986), .A2(n4356), .B1(n4396), .B2(n3988), .ZN(n3902)
         );
  AOI211_X1 U4691 ( .C1(n3972), .C2(n4351), .A(n3903), .B(n3902), .ZN(n3904)
         );
  OAI21_X1 U4692 ( .B1(n3905), .B2(n3974), .A(n3904), .ZN(U3220) );
  NAND2_X1 U4693 ( .A1(n3906), .A2(n3908), .ZN(n3979) );
  INV_X1 U4694 ( .A(n3907), .ZN(n3978) );
  NAND2_X1 U4695 ( .A1(n3979), .A2(n3978), .ZN(n3976) );
  OR2_X1 U4696 ( .A1(n3906), .A2(n3908), .ZN(n3980) );
  NAND2_X1 U4697 ( .A1(n3976), .A2(n3980), .ZN(n3911) );
  XOR2_X1 U4698 ( .A(n3910), .B(n3909), .Z(n3916) );
  XNOR2_X1 U4699 ( .A(n3911), .B(n3916), .ZN(n3912) );
  NAND2_X1 U4700 ( .A1(n3912), .A2(n3981), .ZN(n3915) );
  NOR2_X1 U4701 ( .A1(n4855), .A2(STATE_REG_SCAN_IN), .ZN(n4708) );
  INV_X1 U4702 ( .A(n4568), .ZN(n4452) );
  OAI22_X1 U4703 ( .A1(n3986), .A2(n4570), .B1(n4452), .B2(n3984), .ZN(n3913)
         );
  AOI211_X1 U4704 ( .C1(n3961), .C2(n4585), .A(n4708), .B(n3913), .ZN(n3914)
         );
  OAI211_X1 U4705 ( .C1(n3993), .C2(n4447), .A(n3915), .B(n3914), .ZN(U3223)
         );
  INV_X1 U4706 ( .A(n3980), .ZN(n3977) );
  OAI211_X1 U4707 ( .C1(n3977), .C2(n3978), .A(n3916), .B(n3979), .ZN(n3918)
         );
  NAND2_X1 U4708 ( .A1(n3918), .A2(n3917), .ZN(n3922) );
  XNOR2_X1 U4709 ( .A(n3920), .B(n3919), .ZN(n3921) );
  XNOR2_X1 U4710 ( .A(n3922), .B(n3921), .ZN(n3928) );
  INV_X1 U4711 ( .A(n4577), .ZN(n3985) );
  AOI22_X1 U4712 ( .A1(n3924), .A2(n4431), .B1(n3923), .B2(n4561), .ZN(n3925)
         );
  NAND2_X1 U4713 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4195) );
  OAI211_X1 U4714 ( .C1(n3985), .C2(n3988), .A(n3925), .B(n4195), .ZN(n3926)
         );
  AOI21_X1 U4715 ( .B1(n4432), .B2(n3972), .A(n3926), .ZN(n3927) );
  OAI21_X1 U4716 ( .B1(n3928), .B2(n3974), .A(n3927), .ZN(U3225) );
  INV_X1 U4717 ( .A(n3929), .ZN(n3934) );
  OAI21_X1 U4718 ( .B1(n3933), .B2(n3931), .A(n3930), .ZN(n3932) );
  OAI21_X1 U4719 ( .B1(n3934), .B2(n3933), .A(n3932), .ZN(n3935) );
  NAND2_X1 U4720 ( .A1(n3935), .A2(n3981), .ZN(n3940) );
  OAI22_X1 U4721 ( .A1(n3986), .A2(n4376), .B1(n3958), .B2(n3988), .ZN(n3938)
         );
  OAI22_X1 U4722 ( .A1(n4370), .A2(n3984), .B1(STATE_REG_SCAN_IN), .B2(n3936), 
        .ZN(n3937) );
  NOR2_X1 U4723 ( .A1(n3938), .A2(n3937), .ZN(n3939) );
  OAI211_X1 U4724 ( .C1(n3993), .C2(n4379), .A(n3940), .B(n3939), .ZN(U3230)
         );
  XNOR2_X1 U4725 ( .A(n3943), .B(n3942), .ZN(n3944) );
  XNOR2_X1 U4726 ( .A(n3941), .B(n3944), .ZN(n3945) );
  NAND2_X1 U4727 ( .A1(n3945), .A2(n3981), .ZN(n3951) );
  OAI22_X1 U4728 ( .A1(n3986), .A2(n3946), .B1(n4482), .B2(n3984), .ZN(n3947)
         );
  AOI211_X1 U4729 ( .C1(n3961), .C2(n3949), .A(n3948), .B(n3947), .ZN(n3950)
         );
  OAI211_X1 U4730 ( .C1(n3993), .C2(n4493), .A(n3951), .B(n3950), .ZN(U3231)
         );
  INV_X1 U4731 ( .A(n3953), .ZN(n3955) );
  NAND2_X1 U4732 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  XNOR2_X1 U4733 ( .A(n3952), .B(n3956), .ZN(n3957) );
  NAND2_X1 U4734 ( .A1(n3957), .A2(n3981), .ZN(n3963) );
  OAI22_X1 U4735 ( .A1(n3986), .A2(n4417), .B1(n3958), .B2(n3984), .ZN(n3959)
         );
  AOI211_X1 U4736 ( .C1(n3961), .C2(n4568), .A(n3960), .B(n3959), .ZN(n3962)
         );
  OAI211_X1 U4737 ( .C1(n3993), .C2(n4421), .A(n3963), .B(n3962), .ZN(U3235)
         );
  INV_X1 U4738 ( .A(n3965), .ZN(n3967) );
  NAND2_X1 U4739 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  XNOR2_X1 U4740 ( .A(n3964), .B(n3968), .ZN(n3975) );
  OAI22_X1 U4741 ( .A1(n5037), .A2(n3988), .B1(STATE_REG_SCAN_IN), .B2(n3969), 
        .ZN(n3971) );
  OAI22_X1 U4742 ( .A1(n4264), .A2(n3984), .B1(n3986), .B2(n4266), .ZN(n3970)
         );
  AOI211_X1 U4743 ( .C1(n4268), .C2(n3972), .A(n3971), .B(n3970), .ZN(n3973)
         );
  OAI21_X1 U4744 ( .B1(n3975), .B2(n3974), .A(n3973), .ZN(U3237) );
  NOR2_X1 U4745 ( .A1(n3977), .A2(n3976), .ZN(n3983) );
  AOI21_X1 U4746 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n3982) );
  OAI21_X1 U4747 ( .B1(n3983), .B2(n3982), .A(n3981), .ZN(n3992) );
  OAI22_X1 U4748 ( .A1(n3986), .A2(n4579), .B1(n3985), .B2(n3984), .ZN(n3990)
         );
  OAI22_X1 U4749 ( .A1(n3988), .A2(n4482), .B1(STATE_REG_SCAN_IN), .B2(n3987), 
        .ZN(n3989) );
  NOR2_X1 U4750 ( .A1(n3990), .A2(n3989), .ZN(n3991) );
  OAI211_X1 U4751 ( .C1(n3993), .C2(n4466), .A(n3992), .B(n3991), .ZN(U3238)
         );
  OAI211_X1 U4752 ( .C1(n3996), .C2(n2878), .A(n3995), .B(n3994), .ZN(n3998)
         );
  NAND3_X1 U4753 ( .A1(n3998), .A2(n2485), .A3(n3997), .ZN(n4001) );
  NAND3_X1 U4754 ( .A1(n4001), .A2(n4000), .A3(n3999), .ZN(n4004) );
  NAND3_X1 U4755 ( .A1(n4004), .A2(n4003), .A3(n4002), .ZN(n4006) );
  NAND4_X1 U4756 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4021), .ZN(n4010)
         );
  AND3_X1 U4757 ( .A1(n4010), .A2(n4009), .A3(n4008), .ZN(n4015) );
  NAND2_X1 U4758 ( .A1(n4012), .A2(n4011), .ZN(n4024) );
  OAI211_X1 U4759 ( .C1(n4015), .C2(n4024), .A(n4014), .B(n4013), .ZN(n4019)
         );
  NAND2_X1 U4760 ( .A1(n4017), .A2(n4016), .ZN(n4027) );
  INV_X1 U4761 ( .A(n4027), .ZN(n4018) );
  NAND3_X1 U4762 ( .A1(n4019), .A2(n4018), .A3(n4020), .ZN(n4034) );
  INV_X1 U4763 ( .A(n4020), .ZN(n4025) );
  INV_X1 U4764 ( .A(n4021), .ZN(n4023) );
  NOR4_X1 U4765 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4029)
         );
  INV_X1 U4766 ( .A(n4026), .ZN(n4028) );
  NAND2_X1 U4767 ( .A1(n4027), .A2(n4037), .ZN(n4101) );
  OAI21_X1 U4768 ( .B1(n4029), .B2(n4028), .A(n4101), .ZN(n4033) );
  NAND3_X1 U4769 ( .A1(n4038), .A2(n4031), .A3(n4030), .ZN(n4032) );
  AOI21_X1 U4770 ( .B1(n4034), .B2(n4033), .A(n4032), .ZN(n4044) );
  INV_X1 U4771 ( .A(n4035), .ZN(n4039) );
  NAND2_X1 U4772 ( .A1(n4037), .A2(n4036), .ZN(n4102) );
  AOI21_X1 U4773 ( .B1(n4039), .B2(n4038), .A(n4102), .ZN(n4042) );
  INV_X1 U4774 ( .A(n4101), .ZN(n4040) );
  AOI21_X1 U4775 ( .B1(n4042), .B2(n4041), .A(n4040), .ZN(n4043) );
  OAI21_X1 U4776 ( .B1(n4044), .B2(n4043), .A(n4103), .ZN(n4045) );
  AOI21_X1 U4777 ( .B1(n4045), .B2(n4106), .A(n4104), .ZN(n4046) );
  INV_X1 U4778 ( .A(n4305), .ZN(n4093) );
  OAI211_X1 U4779 ( .C1(n4046), .C2(n4109), .A(n4108), .B(n4093), .ZN(n4047)
         );
  AOI21_X1 U4780 ( .B1(n4047), .B2(n4111), .A(n4113), .ZN(n4049) );
  INV_X1 U4781 ( .A(n4048), .ZN(n4118) );
  INV_X1 U4782 ( .A(n4075), .ZN(n4115) );
  NOR2_X1 U4783 ( .A1(n4116), .A2(n4115), .ZN(n4117) );
  OAI21_X1 U4784 ( .B1(n4049), .B2(n4118), .A(n4117), .ZN(n4054) );
  NAND2_X1 U4785 ( .A1(n4051), .A2(n4050), .ZN(n4056) );
  NOR2_X1 U4786 ( .A1(n4056), .A2(n4052), .ZN(n4100) );
  OAI21_X1 U4787 ( .B1(n4264), .B2(n4507), .A(n4100), .ZN(n4053) );
  AOI21_X1 U4788 ( .B1(n4121), .B2(n4054), .A(n4053), .ZN(n4060) );
  NAND2_X1 U4789 ( .A1(n4055), .A2(n2185), .ZN(n4124) );
  INV_X1 U4790 ( .A(n4124), .ZN(n4057) );
  INV_X1 U4791 ( .A(n4146), .ZN(n4058) );
  AND2_X1 U4792 ( .A1(n4145), .A2(n4132), .ZN(n4059) );
  AOI21_X1 U4793 ( .B1(n4058), .B2(n4218), .A(n4059), .ZN(n4120) );
  OAI211_X1 U4794 ( .C1(n4057), .C2(n4056), .A(n4120), .B(n4122), .ZN(n4099)
         );
  INV_X1 U4795 ( .A(n4132), .ZN(n4130) );
  INV_X1 U4796 ( .A(n4145), .ZN(n4097) );
  NOR2_X1 U4797 ( .A1(n4058), .A2(n4218), .ZN(n4098) );
  AOI21_X1 U4798 ( .B1(n4130), .B2(n4097), .A(n4098), .ZN(n4067) );
  OAI22_X1 U4799 ( .A1(n4060), .A2(n4099), .B1(n4059), .B2(n4067), .ZN(n4135)
         );
  INV_X1 U4800 ( .A(n4116), .ZN(n4062) );
  NAND2_X1 U4801 ( .A1(n4062), .A2(n4255), .ZN(n4276) );
  INV_X1 U4802 ( .A(n4276), .ZN(n4096) );
  NAND2_X1 U4803 ( .A1(n4288), .A2(n4063), .ZN(n4314) );
  INV_X1 U4804 ( .A(n4314), .ZN(n4074) );
  INV_X1 U4805 ( .A(n4325), .ZN(n4343) );
  NAND2_X1 U4806 ( .A1(n4065), .A2(n4064), .ZN(n4397) );
  INV_X1 U4807 ( .A(n4386), .ZN(n4066) );
  OR2_X1 U4808 ( .A1(n4066), .A2(n4387), .ZN(n4428) );
  NAND4_X1 U4809 ( .A1(n4068), .A2(n4238), .A3(n4067), .A4(n4120), .ZN(n4072)
         );
  INV_X1 U4810 ( .A(n4069), .ZN(n4071) );
  NAND2_X1 U4811 ( .A1(n4071), .A2(n4070), .ZN(n4490) );
  NOR4_X1 U4812 ( .A1(n4397), .A2(n4428), .A3(n4072), .A4(n4490), .ZN(n4073)
         );
  NAND2_X1 U4813 ( .A1(n4076), .A2(n4075), .ZN(n4290) );
  NAND4_X1 U4814 ( .A1(n4412), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4084)
         );
  NAND2_X1 U4815 ( .A1(n4081), .A2(n4080), .ZN(n4083) );
  NOR4_X1 U4816 ( .A1(n4084), .A2(n3401), .A3(n4083), .A4(n4082), .ZN(n4092)
         );
  XNOR2_X1 U4817 ( .A(n4541), .B(n4368), .ZN(n4366) );
  NOR4_X1 U4818 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4091)
         );
  NOR4_X1 U4819 ( .A1(n4721), .A2(n4462), .A3(n2844), .A4(n4089), .ZN(n4090)
         );
  NAND4_X1 U4820 ( .A1(n4092), .A2(n4366), .A3(n4091), .A4(n4090), .ZN(n4094)
         );
  NAND2_X1 U4821 ( .A1(n4093), .A2(n4324), .ZN(n4348) );
  NOR2_X1 U4822 ( .A1(n4095), .A2(n2186), .ZN(n4254) );
  INV_X1 U4823 ( .A(n4254), .ZN(n4257) );
  OR2_X1 U4824 ( .A1(n4098), .A2(n4097), .ZN(n4129) );
  AOI21_X1 U4825 ( .B1(n4238), .B2(n4100), .A(n4099), .ZN(n4128) );
  OAI21_X1 U4826 ( .B1(n3754), .B2(n4102), .A(n4101), .ZN(n4107) );
  INV_X1 U4827 ( .A(n4103), .ZN(n4105) );
  AOI211_X1 U4828 ( .C1(n4107), .C2(n4106), .A(n4105), .B(n4104), .ZN(n4110)
         );
  OAI21_X1 U4829 ( .B1(n4110), .B2(n4109), .A(n4108), .ZN(n4112) );
  NAND2_X1 U4830 ( .A1(n4112), .A2(n4111), .ZN(n4126) );
  NOR4_X1 U4831 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4125)
         );
  NAND2_X1 U4832 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  NAND4_X1 U4833 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  AOI211_X1 U4834 ( .C1(n4126), .C2(n4125), .A(n4124), .B(n4123), .ZN(n4127)
         );
  AOI211_X1 U4835 ( .C1(n4130), .C2(n4129), .A(n4128), .B(n4127), .ZN(n4131)
         );
  AOI21_X1 U4836 ( .B1(n4218), .B2(n4132), .A(n4131), .ZN(n4133) );
  MUX2_X1 U4837 ( .A(n4135), .B(n4134), .S(n4680), .Z(n4136) );
  XNOR2_X1 U4838 ( .A(n4136), .B(n4211), .ZN(n4144) );
  INV_X1 U4839 ( .A(n4137), .ZN(n4139) );
  NOR2_X1 U4840 ( .A1(n4139), .A2(n4138), .ZN(n4142) );
  OAI21_X1 U4841 ( .B1(n4143), .B2(n4140), .A(B_REG_SCAN_IN), .ZN(n4141) );
  OAI22_X1 U4842 ( .A1(n4144), .A2(n4143), .B1(n4142), .B2(n4141), .ZN(U3239)
         );
  MUX2_X1 U4843 ( .A(DATAO_REG_31__SCAN_IN), .B(n4145), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4844 ( .A(DATAO_REG_30__SCAN_IN), .B(n4146), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4845 ( .A(DATAO_REG_29__SCAN_IN), .B(n4147), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4846 ( .A(DATAO_REG_27__SCAN_IN), .B(n4148), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4847 ( .A(DATAO_REG_26__SCAN_IN), .B(n4508), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4848 ( .A(DATAO_REG_20__SCAN_IN), .B(n4541), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4849 ( .A(DATAO_REG_19__SCAN_IN), .B(n4414), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4850 ( .A(DATAO_REG_18__SCAN_IN), .B(n4561), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4851 ( .A(DATAO_REG_17__SCAN_IN), .B(n4568), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4852 ( .A(DATAO_REG_15__SCAN_IN), .B(n4585), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4853 ( .A(DATAO_REG_11__SCAN_IN), .B(n4600), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4854 ( .A(DATAO_REG_10__SCAN_IN), .B(n4149), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4855 ( .A(DATAO_REG_9__SCAN_IN), .B(n4150), .S(U4043), .Z(U3559) );
  MUX2_X1 U4856 ( .A(DATAO_REG_5__SCAN_IN), .B(n4151), .S(U4043), .Z(U3555) );
  MUX2_X1 U4857 ( .A(DATAO_REG_4__SCAN_IN), .B(n4152), .S(U4043), .Z(U3554) );
  MUX2_X1 U4858 ( .A(DATAO_REG_2__SCAN_IN), .B(n3392), .S(U4043), .Z(U3552) );
  MUX2_X1 U4859 ( .A(DATAO_REG_1__SCAN_IN), .B(n4153), .S(U4043), .Z(U3551) );
  MUX2_X1 U4860 ( .A(DATAO_REG_0__SCAN_IN), .B(n4154), .S(U4043), .Z(U3550) );
  AND2_X1 U4861 ( .A1(n4709), .A2(ADDR_REG_1__SCAN_IN), .ZN(n4157) );
  NOR2_X1 U4862 ( .A1(n4155), .A2(STATE_REG_SCAN_IN), .ZN(n4156) );
  AOI211_X1 U4863 ( .C1(n4158), .C2(n2928), .A(n4157), .B(n4156), .ZN(n4167)
         );
  OAI211_X1 U4864 ( .C1(n4161), .C2(n4160), .A(n4710), .B(n4159), .ZN(n4166)
         );
  OAI211_X1 U4865 ( .C1(n4164), .C2(n2929), .A(n4184), .B(n4163), .ZN(n4165)
         );
  NAND3_X1 U4866 ( .A1(n4167), .A2(n4166), .A3(n4165), .ZN(U3241) );
  MUX2_X1 U4867 ( .A(REG1_REG_11__SCAN_IN), .B(n4940), .S(n4686), .Z(n4169) );
  OAI211_X1 U4868 ( .C1(n4170), .C2(n4169), .A(n4710), .B(n4168), .ZN(n4179)
         );
  NOR2_X1 U4869 ( .A1(n4715), .A2(n4171), .ZN(n4172) );
  AOI211_X1 U4870 ( .C1(n4709), .C2(ADDR_REG_11__SCAN_IN), .A(n4173), .B(n4172), .ZN(n4178) );
  OAI211_X1 U4871 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4184), .ZN(n4177)
         );
  NAND3_X1 U4872 ( .A1(n4179), .A2(n4178), .A3(n4177), .ZN(U3251) );
  XOR2_X1 U4873 ( .A(REG1_REG_14__SCAN_IN), .B(n4180), .Z(n4189) );
  NOR2_X1 U4874 ( .A1(n4715), .A2(n4181), .ZN(n4182) );
  AOI211_X1 U4875 ( .C1(n4709), .C2(ADDR_REG_14__SCAN_IN), .A(n4183), .B(n4182), .ZN(n4188) );
  OAI211_X1 U4876 ( .C1(n4186), .C2(REG2_REG_14__SCAN_IN), .A(n4185), .B(n4184), .ZN(n4187) );
  OAI211_X1 U4877 ( .C1(n4189), .C2(n4199), .A(n4188), .B(n4187), .ZN(U3254)
         );
  AOI21_X1 U4878 ( .B1(n2167), .B2(n4191), .A(n4190), .ZN(n4200) );
  OR2_X1 U4879 ( .A1(n4715), .A2(n4196), .ZN(n4197) );
  OAI211_X1 U4880 ( .C1(n4200), .C2(n4199), .A(n4198), .B(n4197), .ZN(U3257)
         );
  MUX2_X1 U4881 ( .A(REG2_REG_19__SCAN_IN), .B(n2638), .S(n4681), .Z(n4203) );
  OAI21_X1 U4882 ( .B1(n4205), .B2(n4732), .A(n4204), .ZN(n4208) );
  INV_X1 U4883 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4206) );
  MUX2_X1 U4884 ( .A(n4206), .B(REG1_REG_19__SCAN_IN), .S(n4681), .Z(n4207) );
  XNOR2_X1 U4885 ( .A(n4208), .B(n4207), .ZN(n4213) );
  NAND2_X1 U4886 ( .A1(n4709), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4209) );
  OAI211_X1 U4887 ( .C1(n4715), .C2(n4211), .A(n4210), .B(n4209), .ZN(n4212)
         );
  AOI21_X1 U4888 ( .B1(n4213), .B2(n4710), .A(n4212), .ZN(n4214) );
  OAI21_X1 U4889 ( .B1(n4215), .B2(n4703), .A(n4214), .ZN(U3259) );
  AOI21_X1 U4890 ( .B1(n4218), .B2(n4217), .A(n4216), .ZN(n4504) );
  NAND2_X1 U4891 ( .A1(n4504), .A2(n4459), .ZN(n4222) );
  NAND2_X1 U4892 ( .A1(n4540), .A2(n4218), .ZN(n4219) );
  NAND2_X1 U4893 ( .A1(n4220), .A2(n4219), .ZN(n4616) );
  NAND2_X1 U4894 ( .A1(n4724), .A2(n4616), .ZN(n4221) );
  OAI211_X1 U4895 ( .C1(n4724), .C2(n4223), .A(n4222), .B(n4221), .ZN(U3261)
         );
  NAND2_X1 U4896 ( .A1(n4224), .A2(n4501), .ZN(n4235) );
  INV_X1 U4897 ( .A(n4225), .ZN(n4233) );
  INV_X1 U4898 ( .A(n4226), .ZN(n4227) );
  AOI22_X1 U4899 ( .A1(n4227), .A2(n4720), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4726), .ZN(n4228) );
  OAI21_X1 U4900 ( .B1(n4229), .B2(n4451), .A(n4228), .ZN(n4232) );
  OAI22_X1 U4901 ( .A1(n4264), .A2(n4469), .B1(n4468), .B2(n4230), .ZN(n4231)
         );
  OAI211_X1 U4902 ( .C1(n4726), .C2(n4236), .A(n4235), .B(n4234), .ZN(U3262)
         );
  XNOR2_X1 U4903 ( .A(n4239), .B(n4238), .ZN(n4240) );
  NAND2_X1 U4904 ( .A1(n4240), .A2(n4590), .ZN(n4510) );
  NOR2_X1 U4905 ( .A1(n4510), .A2(n4726), .ZN(n4251) );
  INV_X1 U4906 ( .A(n4265), .ZN(n4243) );
  INV_X1 U4907 ( .A(n4241), .ZN(n4242) );
  INV_X1 U4908 ( .A(n4469), .ZN(n4444) );
  OAI22_X1 U4909 ( .A1(n4245), .A2(n4492), .B1(n4244), .B2(n4724), .ZN(n4248)
         );
  OAI22_X1 U4910 ( .A1(n4511), .A2(n4451), .B1(n4246), .B2(n4468), .ZN(n4247)
         );
  AOI211_X1 U4911 ( .C1(n4444), .C2(n4508), .A(n4248), .B(n4247), .ZN(n4249)
         );
  OAI21_X1 U4912 ( .B1(n4623), .B2(n4498), .A(n4249), .ZN(n4250) );
  AOI211_X1 U4913 ( .C1(n4512), .C2(n4501), .A(n4251), .B(n4250), .ZN(n4252)
         );
  INV_X1 U4914 ( .A(n4252), .ZN(U3263) );
  XNOR2_X1 U4915 ( .A(n4253), .B(n4254), .ZN(n4515) );
  INV_X1 U4916 ( .A(n4515), .ZN(n4272) );
  NAND2_X1 U4917 ( .A1(n4256), .A2(n4255), .ZN(n4258) );
  XNOR2_X1 U4918 ( .A(n4258), .B(n4257), .ZN(n4259) );
  NAND2_X1 U4919 ( .A1(n4259), .A2(n4590), .ZN(n4263) );
  AOI22_X1 U4920 ( .A1(n4261), .A2(n4599), .B1(n4540), .B2(n4260), .ZN(n4262)
         );
  OAI211_X1 U4921 ( .C1(n4264), .C2(n4544), .A(n4263), .B(n4262), .ZN(n4514)
         );
  INV_X1 U4922 ( .A(n4277), .ZN(n4267) );
  OAI21_X1 U4923 ( .B1(n4267), .B2(n4266), .A(n4265), .ZN(n4626) );
  AOI22_X1 U4924 ( .A1(n4268), .A2(n4720), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4726), .ZN(n4269) );
  OAI21_X1 U4925 ( .B1(n4626), .B2(n4498), .A(n4269), .ZN(n4270) );
  AOI21_X1 U4926 ( .B1(n4514), .B2(n4724), .A(n4270), .ZN(n4271) );
  OAI21_X1 U4927 ( .B1(n4272), .B2(n4456), .A(n4271), .ZN(U3264) );
  XNOR2_X1 U4928 ( .A(n4273), .B(n4276), .ZN(n4274) );
  NAND2_X1 U4929 ( .A1(n4274), .A2(n4590), .ZN(n4520) );
  XNOR2_X1 U4930 ( .A(n4275), .B(n4276), .ZN(n4523) );
  NAND2_X1 U4931 ( .A1(n4523), .A2(n4501), .ZN(n4285) );
  OAI21_X1 U4932 ( .B1(n4296), .B2(n4280), .A(n4277), .ZN(n4630) );
  INV_X1 U4933 ( .A(n4630), .ZN(n4283) );
  AOI22_X1 U4934 ( .A1(n4278), .A2(n4720), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4726), .ZN(n4279) );
  OAI21_X1 U4935 ( .B1(n4521), .B2(n4451), .A(n4279), .ZN(n4282) );
  OAI22_X1 U4936 ( .A1(n4312), .A2(n4469), .B1(n4468), .B2(n4280), .ZN(n4281)
         );
  AOI211_X1 U4937 ( .C1(n4283), .C2(n4459), .A(n4282), .B(n4281), .ZN(n4284)
         );
  OAI211_X1 U4938 ( .C1(n4726), .C2(n4520), .A(n4285), .B(n4284), .ZN(U3265)
         );
  XNOR2_X1 U4939 ( .A(n2139), .B(n4290), .ZN(n4527) );
  INV_X1 U4940 ( .A(n4527), .ZN(n4303) );
  NAND2_X1 U4941 ( .A1(n4287), .A2(n4288), .ZN(n4289) );
  XOR2_X1 U4942 ( .A(n4290), .B(n4289), .Z(n4291) );
  NAND2_X1 U4943 ( .A1(n4291), .A2(n4590), .ZN(n4295) );
  AOI22_X1 U4944 ( .A1(n4293), .A2(n4599), .B1(n4540), .B2(n4292), .ZN(n4294)
         );
  OAI211_X1 U4945 ( .C1(n5037), .C2(n4544), .A(n4295), .B(n4294), .ZN(n4526)
         );
  INV_X1 U4946 ( .A(n4296), .ZN(n4297) );
  OAI21_X1 U4947 ( .B1(n4316), .B2(n4298), .A(n4297), .ZN(n4634) );
  AOI22_X1 U4948 ( .A1(n4299), .A2(n4720), .B1(n4726), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4300) );
  OAI21_X1 U4949 ( .B1(n4634), .B2(n4498), .A(n4300), .ZN(n4301) );
  AOI21_X1 U4950 ( .B1(n4526), .B2(n4724), .A(n4301), .ZN(n4302) );
  OAI21_X1 U4951 ( .B1(n4303), .B2(n4456), .A(n4302), .ZN(U3266) );
  AOI21_X1 U4952 ( .B1(n4326), .B2(n4324), .A(n4325), .ZN(n4327) );
  INV_X1 U4953 ( .A(n4306), .ZN(n4307) );
  NOR2_X1 U4954 ( .A1(n4327), .A2(n4307), .ZN(n4308) );
  XNOR2_X1 U4955 ( .A(n4308), .B(n4314), .ZN(n4309) );
  NAND2_X1 U4956 ( .A1(n4309), .A2(n4590), .ZN(n4311) );
  AOI22_X1 U4957 ( .A1(n4355), .A2(n4599), .B1(n4540), .B2(n4315), .ZN(n4310)
         );
  OAI211_X1 U4958 ( .C1(n4312), .C2(n4544), .A(n4311), .B(n4310), .ZN(n4530)
         );
  INV_X1 U4959 ( .A(n4530), .ZN(n4323) );
  XOR2_X1 U4960 ( .A(n4314), .B(n4313), .Z(n4531) );
  AND2_X1 U4961 ( .A1(n4338), .A2(n4315), .ZN(n4317) );
  OR2_X1 U4962 ( .A1(n4317), .A2(n4316), .ZN(n4638) );
  NOR2_X1 U4963 ( .A1(n4638), .A2(n4498), .ZN(n4321) );
  OAI22_X1 U4964 ( .A1(n4319), .A2(n4492), .B1(n4724), .B2(n4318), .ZN(n4320)
         );
  AOI211_X1 U4965 ( .C1(n4531), .C2(n4501), .A(n4321), .B(n4320), .ZN(n4322)
         );
  OAI21_X1 U4966 ( .B1(n4726), .B2(n4323), .A(n4322), .ZN(U3267) );
  AND3_X1 U4967 ( .A1(n4326), .A2(n4325), .A3(n4324), .ZN(n4328) );
  OR2_X1 U4968 ( .A1(n4328), .A2(n4327), .ZN(n4334) );
  NAND2_X1 U4969 ( .A1(n4540), .A2(n4336), .ZN(n4331) );
  NAND2_X1 U4970 ( .A1(n4329), .A2(n4599), .ZN(n4330) );
  OAI211_X1 U4971 ( .C1(n4332), .C2(n4544), .A(n4331), .B(n4330), .ZN(n4333)
         );
  AOI21_X1 U4972 ( .B1(n4334), .B2(n4590), .A(n4333), .ZN(n4536) );
  NAND2_X1 U4973 ( .A1(n4335), .A2(n4336), .ZN(n4337) );
  NAND2_X1 U4974 ( .A1(n4338), .A2(n4337), .ZN(n4642) );
  INV_X1 U4975 ( .A(n4642), .ZN(n4342) );
  OAI22_X1 U4976 ( .A1(n4724), .A2(n4340), .B1(n4339), .B2(n4492), .ZN(n4341)
         );
  AOI21_X1 U4977 ( .B1(n4342), .B2(n4459), .A(n4341), .ZN(n4346) );
  NAND2_X1 U4978 ( .A1(n2150), .A2(n4343), .ZN(n4534) );
  NAND3_X1 U4979 ( .A1(n4534), .A2(n4501), .A3(n4344), .ZN(n4345) );
  OAI211_X1 U4980 ( .C1(n4536), .C2(n4726), .A(n4346), .B(n4345), .ZN(U3268)
         );
  XNOR2_X1 U4981 ( .A(n4304), .B(n4348), .ZN(n4347) );
  NAND2_X1 U4982 ( .A1(n4347), .A2(n4590), .ZN(n4543) );
  XOR2_X1 U4983 ( .A(n4349), .B(n4348), .Z(n4547) );
  OR2_X1 U4984 ( .A1(n4378), .A2(n4356), .ZN(n4350) );
  NAND2_X1 U4985 ( .A1(n4335), .A2(n4350), .ZN(n4646) );
  INV_X1 U4986 ( .A(n4351), .ZN(n4352) );
  OAI22_X1 U4987 ( .A1(n4724), .A2(n4353), .B1(n4352), .B2(n4492), .ZN(n4354)
         );
  AOI21_X1 U4988 ( .B1(n4472), .B2(n4355), .A(n4354), .ZN(n4359) );
  OAI22_X1 U4989 ( .A1(n4396), .A2(n4469), .B1(n4468), .B2(n4356), .ZN(n4357)
         );
  INV_X1 U4990 ( .A(n4357), .ZN(n4358) );
  OAI211_X1 U4991 ( .C1(n4646), .C2(n4498), .A(n4359), .B(n4358), .ZN(n4360)
         );
  AOI21_X1 U4992 ( .B1(n4547), .B2(n4501), .A(n4360), .ZN(n4361) );
  OAI21_X1 U4993 ( .B1(n4726), .B2(n4543), .A(n4361), .ZN(U3269) );
  XNOR2_X1 U4994 ( .A(n4362), .B(n4366), .ZN(n4550) );
  INV_X1 U4995 ( .A(n4363), .ZN(n4364) );
  NAND2_X1 U4996 ( .A1(n4365), .A2(n4364), .ZN(n4367) );
  XNOR2_X1 U4997 ( .A(n4367), .B(n4366), .ZN(n4372) );
  AOI22_X1 U4998 ( .A1(n4414), .A2(n4599), .B1(n4540), .B2(n4368), .ZN(n4369)
         );
  OAI21_X1 U4999 ( .B1(n4370), .B2(n4544), .A(n4369), .ZN(n4371) );
  AOI21_X1 U5000 ( .B1(n4372), .B2(n4590), .A(n4371), .ZN(n4373) );
  OAI21_X1 U5001 ( .B1(n4550), .B2(n4374), .A(n4373), .ZN(n4551) );
  NAND2_X1 U5002 ( .A1(n4551), .A2(n4724), .ZN(n4384) );
  NOR2_X1 U5003 ( .A1(n4375), .A2(n4376), .ZN(n4377) );
  OR2_X1 U5004 ( .A1(n4378), .A2(n4377), .ZN(n4649) );
  INV_X1 U5005 ( .A(n4649), .ZN(n4382) );
  OAI22_X1 U5006 ( .A1(n4724), .A2(n4380), .B1(n4379), .B2(n4492), .ZN(n4381)
         );
  AOI21_X1 U5007 ( .B1(n4382), .B2(n4459), .A(n4381), .ZN(n4383) );
  OAI211_X1 U5008 ( .C1(n4550), .C2(n4385), .A(n4384), .B(n4383), .ZN(U3270)
         );
  OAI21_X1 U5009 ( .B1(n4425), .B2(n4387), .A(n4386), .ZN(n4413) );
  INV_X1 U5010 ( .A(n4388), .ZN(n4390) );
  OAI21_X1 U5011 ( .B1(n4413), .B2(n4390), .A(n4389), .ZN(n4391) );
  XNOR2_X1 U5012 ( .A(n4391), .B(n4397), .ZN(n4392) );
  NAND2_X1 U5013 ( .A1(n4392), .A2(n4590), .ZN(n4395) );
  AOI22_X1 U5014 ( .A1(n4561), .A2(n4599), .B1(n4540), .B2(n4393), .ZN(n4394)
         );
  OAI211_X1 U5015 ( .C1(n4396), .C2(n4544), .A(n4395), .B(n4394), .ZN(n4555)
         );
  INV_X1 U5016 ( .A(n4555), .ZN(n4405) );
  XNOR2_X1 U5017 ( .A(n4398), .B(n4397), .ZN(n4556) );
  NOR2_X1 U5018 ( .A1(n4409), .A2(n4399), .ZN(n4400) );
  OR2_X1 U5019 ( .A1(n4375), .A2(n4400), .ZN(n4653) );
  AOI22_X1 U5020 ( .A1(n4726), .A2(REG2_REG_19__SCAN_IN), .B1(n4401), .B2(
        n4720), .ZN(n4402) );
  OAI21_X1 U5021 ( .B1(n4653), .B2(n4498), .A(n4402), .ZN(n4403) );
  AOI21_X1 U5022 ( .B1(n4556), .B2(n4501), .A(n4403), .ZN(n4404) );
  OAI21_X1 U5023 ( .B1(n4405), .B2(n4726), .A(n4404), .ZN(U3271) );
  INV_X1 U5024 ( .A(n4406), .ZN(n4407) );
  AOI21_X1 U5025 ( .B1(n4412), .B2(n4408), .A(n4407), .ZN(n4560) );
  INV_X1 U5026 ( .A(n4430), .ZN(n4411) );
  INV_X1 U5027 ( .A(n4409), .ZN(n4410) );
  OAI211_X1 U5028 ( .C1(n4411), .C2(n4417), .A(n4410), .B(n4611), .ZN(n4558)
         );
  XNOR2_X1 U5029 ( .A(n4413), .B(n4412), .ZN(n4419) );
  NAND2_X1 U5030 ( .A1(n4414), .A2(n4598), .ZN(n4416) );
  NAND2_X1 U5031 ( .A1(n4568), .A2(n4599), .ZN(n4415) );
  OAI211_X1 U5032 ( .C1(n4417), .C2(n4603), .A(n4416), .B(n4415), .ZN(n4418)
         );
  AOI21_X1 U5033 ( .B1(n4419), .B2(n4590), .A(n4418), .ZN(n4559) );
  OAI21_X1 U5034 ( .B1(n4681), .B2(n4558), .A(n4559), .ZN(n4420) );
  NAND2_X1 U5035 ( .A1(n4420), .A2(n4724), .ZN(n4424) );
  INV_X1 U5036 ( .A(n4421), .ZN(n4422) );
  AOI22_X1 U5037 ( .A1(n4726), .A2(REG2_REG_18__SCAN_IN), .B1(n4422), .B2(
        n4720), .ZN(n4423) );
  OAI211_X1 U5038 ( .C1(n4560), .C2(n4456), .A(n4424), .B(n4423), .ZN(U3272)
         );
  XOR2_X1 U5039 ( .A(n4428), .B(n4425), .Z(n4426) );
  NOR2_X1 U5040 ( .A1(n4426), .A2(n4485), .ZN(n4564) );
  INV_X1 U5041 ( .A(n4564), .ZN(n4439) );
  XOR2_X1 U5042 ( .A(n4428), .B(n4427), .Z(n4566) );
  INV_X1 U5043 ( .A(n4429), .ZN(n4443) );
  OAI21_X1 U5044 ( .B1(n4443), .B2(n4563), .A(n4430), .ZN(n4658) );
  NOR2_X1 U5045 ( .A1(n4658), .A2(n4498), .ZN(n4437) );
  INV_X1 U5046 ( .A(n4561), .ZN(n4435) );
  AOI22_X1 U5047 ( .A1(n4445), .A2(n4431), .B1(n4444), .B2(n4577), .ZN(n4434)
         );
  AOI22_X1 U5048 ( .A1(n4726), .A2(REG2_REG_17__SCAN_IN), .B1(n4432), .B2(
        n4720), .ZN(n4433) );
  OAI211_X1 U5049 ( .C1(n4435), .C2(n4451), .A(n4434), .B(n4433), .ZN(n4436)
         );
  AOI211_X1 U5050 ( .C1(n4566), .C2(n4501), .A(n4437), .B(n4436), .ZN(n4438)
         );
  OAI21_X1 U5051 ( .B1(n4439), .B2(n4726), .A(n4438), .ZN(U3273) );
  OAI211_X1 U5052 ( .C1(n4442), .C2(n4441), .A(n4440), .B(n4590), .ZN(n4574)
         );
  AOI21_X1 U5053 ( .B1(n4446), .B2(n4464), .A(n4443), .ZN(n4572) );
  AOI22_X1 U5054 ( .A1(n4446), .A2(n4445), .B1(n4444), .B2(n4585), .ZN(n4450)
         );
  INV_X1 U5055 ( .A(n4447), .ZN(n4448) );
  AOI22_X1 U5056 ( .A1(n4726), .A2(REG2_REG_16__SCAN_IN), .B1(n4448), .B2(
        n4720), .ZN(n4449) );
  OAI211_X1 U5057 ( .C1(n4452), .C2(n4451), .A(n4450), .B(n4449), .ZN(n4458)
         );
  OAI21_X1 U5058 ( .B1(n2140), .B2(n4454), .A(n4453), .ZN(n4575) );
  NOR2_X1 U5059 ( .A1(n4575), .A2(n4456), .ZN(n4457) );
  AOI211_X1 U5060 ( .C1(n4572), .C2(n4459), .A(n4458), .B(n4457), .ZN(n4460)
         );
  OAI21_X1 U5061 ( .B1(n4726), .B2(n4574), .A(n4460), .ZN(U3274) );
  AOI211_X1 U5062 ( .C1(n4461), .C2(n4462), .A(n4485), .B(n2168), .ZN(n4580)
         );
  INV_X1 U5063 ( .A(n4580), .ZN(n4476) );
  XNOR2_X1 U5064 ( .A(n4463), .B(n4462), .ZN(n4582) );
  OAI21_X1 U5065 ( .B1(n4465), .B2(n4579), .A(n4464), .ZN(n4662) );
  INV_X1 U5066 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4467) );
  OAI22_X1 U5067 ( .A1(n4724), .A2(n4467), .B1(n4466), .B2(n4492), .ZN(n4471)
         );
  OAI22_X1 U5068 ( .A1(n4482), .A2(n4469), .B1(n4468), .B2(n4579), .ZN(n4470)
         );
  AOI211_X1 U5069 ( .C1(n4472), .C2(n4577), .A(n4471), .B(n4470), .ZN(n4473)
         );
  OAI21_X1 U5070 ( .B1(n4662), .B2(n4498), .A(n4473), .ZN(n4474) );
  AOI21_X1 U5071 ( .B1(n4582), .B2(n4501), .A(n4474), .ZN(n4475) );
  OAI21_X1 U5072 ( .B1(n4476), .B2(n4726), .A(n4475), .ZN(U3275) );
  OAI21_X1 U5073 ( .B1(n3726), .B2(n4478), .A(n4477), .ZN(n4479) );
  XOR2_X1 U5074 ( .A(n4490), .B(n4479), .Z(n4486) );
  OAI22_X1 U5075 ( .A1(n4482), .A2(n4544), .B1(n4481), .B2(n4480), .ZN(n4483)
         );
  AOI21_X1 U5076 ( .B1(n4540), .B2(n4495), .A(n4483), .ZN(n4484) );
  OAI21_X1 U5077 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4594) );
  INV_X1 U5078 ( .A(n4594), .ZN(n4503) );
  AND2_X1 U5079 ( .A1(n2190), .A2(n4489), .ZN(n4491) );
  XNOR2_X1 U5080 ( .A(n4491), .B(n4490), .ZN(n4595) );
  OAI22_X1 U5081 ( .A1(n4724), .A2(n4494), .B1(n4493), .B2(n4492), .ZN(n4500)
         );
  AND2_X1 U5082 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  OR2_X1 U5083 ( .A1(n4497), .A2(n2181), .ZN(n4670) );
  NOR2_X1 U5084 ( .A1(n4670), .A2(n4498), .ZN(n4499) );
  AOI211_X1 U5085 ( .C1(n4595), .C2(n4501), .A(n4500), .B(n4499), .ZN(n4502)
         );
  OAI21_X1 U5086 ( .B1(n4503), .B2(n4726), .A(n4502), .ZN(U3277) );
  INV_X1 U5087 ( .A(n4504), .ZN(n4619) );
  NAND2_X1 U5088 ( .A1(n4756), .A2(n4616), .ZN(n4506) );
  NAND2_X1 U5089 ( .A1(n4754), .A2(REG1_REG_30__SCAN_IN), .ZN(n4505) );
  OAI211_X1 U5090 ( .C1(n4619), .C2(n4609), .A(n4506), .B(n4505), .ZN(U3548)
         );
  INV_X1 U5091 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U5092 ( .A1(n4508), .A2(n4599), .B1(n4540), .B2(n4507), .ZN(n4509)
         );
  INV_X1 U5093 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4839) );
  AOI21_X1 U5094 ( .B1(n4515), .B2(n4607), .A(n4514), .ZN(n4624) );
  OAI21_X1 U5095 ( .B1(n4609), .B2(n4626), .A(n4516), .ZN(U3544) );
  INV_X1 U5096 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5097 ( .A1(n4518), .A2(n4599), .B1(n4540), .B2(n4517), .ZN(n4519)
         );
  OAI211_X1 U5098 ( .C1(n4521), .C2(n4544), .A(n4520), .B(n4519), .ZN(n4522)
         );
  AOI21_X1 U5099 ( .B1(n4523), .B2(n4607), .A(n4522), .ZN(n4627) );
  MUX2_X1 U5100 ( .A(n4524), .B(n4627), .S(n4756), .Z(n4525) );
  OAI21_X1 U5101 ( .B1(n4609), .B2(n4630), .A(n4525), .ZN(U3543) );
  INV_X1 U5102 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4528) );
  AOI21_X1 U5103 ( .B1(n4527), .B2(n4607), .A(n4526), .ZN(n4631) );
  MUX2_X1 U5104 ( .A(n4528), .B(n4631), .S(n4756), .Z(n4529) );
  OAI21_X1 U5105 ( .B1(n4609), .B2(n4634), .A(n4529), .ZN(U3542) );
  AOI21_X1 U5106 ( .B1(n4531), .B2(n4607), .A(n4530), .ZN(n4636) );
  INV_X1 U5107 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4532) );
  MUX2_X1 U5108 ( .A(n4636), .B(n4532), .S(n4754), .Z(n4533) );
  OAI21_X1 U5109 ( .B1(n4609), .B2(n4638), .A(n4533), .ZN(U3541) );
  NAND3_X1 U5110 ( .A1(n4534), .A2(n4607), .A3(n4344), .ZN(n4535) );
  NAND2_X1 U5111 ( .A1(n4536), .A2(n4535), .ZN(n4639) );
  MUX2_X1 U5112 ( .A(n4639), .B(REG1_REG_22__SCAN_IN), .S(n4754), .Z(n4537) );
  INV_X1 U5113 ( .A(n4537), .ZN(n4538) );
  OAI21_X1 U5114 ( .B1(n4609), .B2(n4642), .A(n4538), .ZN(U3540) );
  INV_X1 U5115 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5116 ( .A1(n4541), .A2(n4599), .B1(n4540), .B2(n4539), .ZN(n4542)
         );
  OAI211_X1 U5117 ( .C1(n4545), .C2(n4544), .A(n4543), .B(n4542), .ZN(n4546)
         );
  AOI21_X1 U5118 ( .B1(n4547), .B2(n4607), .A(n4546), .ZN(n4643) );
  MUX2_X1 U5119 ( .A(n4548), .B(n4643), .S(n4756), .Z(n4549) );
  OAI21_X1 U5120 ( .B1(n4609), .B2(n4646), .A(n4549), .ZN(U3539) );
  INV_X1 U5121 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4553) );
  INV_X1 U5122 ( .A(n4550), .ZN(n4552) );
  AOI21_X1 U5123 ( .B1(n4742), .B2(n4552), .A(n4551), .ZN(n4647) );
  MUX2_X1 U5124 ( .A(n4553), .B(n4647), .S(n4756), .Z(n4554) );
  OAI21_X1 U5125 ( .B1(n4609), .B2(n4649), .A(n4554), .ZN(U3538) );
  AOI21_X1 U5126 ( .B1(n4607), .B2(n4556), .A(n4555), .ZN(n4650) );
  MUX2_X1 U5127 ( .A(n4206), .B(n4650), .S(n4756), .Z(n4557) );
  OAI21_X1 U5128 ( .B1(n4609), .B2(n4653), .A(n4557), .ZN(U3537) );
  OAI211_X1 U5129 ( .C1(n4744), .C2(n4560), .A(n4559), .B(n4558), .ZN(n4654)
         );
  MUX2_X1 U5130 ( .A(REG1_REG_18__SCAN_IN), .B(n4654), .S(n4756), .Z(U3536) );
  AOI22_X1 U5131 ( .A1(n4561), .A2(n4598), .B1(n4599), .B2(n4577), .ZN(n4562)
         );
  OAI21_X1 U5132 ( .B1(n4603), .B2(n4563), .A(n4562), .ZN(n4565) );
  AOI211_X1 U5133 ( .C1(n4566), .C2(n4607), .A(n4565), .B(n4564), .ZN(n4655)
         );
  MUX2_X1 U5134 ( .A(n2915), .B(n4655), .S(n4756), .Z(n4567) );
  OAI21_X1 U5135 ( .B1(n4609), .B2(n4658), .A(n4567), .ZN(U3535) );
  AOI22_X1 U5136 ( .A1(n4568), .A2(n4598), .B1(n4599), .B2(n4585), .ZN(n4569)
         );
  OAI21_X1 U5137 ( .B1(n4603), .B2(n4570), .A(n4569), .ZN(n4571) );
  AOI21_X1 U5138 ( .B1(n4572), .B2(n4611), .A(n4571), .ZN(n4573) );
  OAI211_X1 U5139 ( .C1(n4744), .C2(n4575), .A(n4574), .B(n4573), .ZN(n4659)
         );
  MUX2_X1 U5140 ( .A(REG1_REG_16__SCAN_IN), .B(n4659), .S(n4756), .Z(U3534) );
  AOI22_X1 U5141 ( .A1(n4577), .A2(n4598), .B1(n4599), .B2(n4576), .ZN(n4578)
         );
  OAI21_X1 U5142 ( .B1(n4603), .B2(n4579), .A(n4578), .ZN(n4581) );
  AOI211_X1 U5143 ( .C1(n4607), .C2(n4582), .A(n4581), .B(n4580), .ZN(n4660)
         );
  MUX2_X1 U5144 ( .A(n2909), .B(n4660), .S(n4756), .Z(n4583) );
  OAI21_X1 U5145 ( .B1(n4609), .B2(n4662), .A(n4583), .ZN(U3533) );
  NAND2_X1 U5146 ( .A1(n4584), .A2(n4607), .ZN(n4587) );
  AOI22_X1 U5147 ( .A1(n4585), .A2(n4598), .B1(n4599), .B2(n4597), .ZN(n4586)
         );
  OAI211_X1 U5148 ( .C1(n4588), .C2(n4603), .A(n4587), .B(n4586), .ZN(n4589)
         );
  AOI21_X1 U5149 ( .B1(n4591), .B2(n4590), .A(n4589), .ZN(n4663) );
  MUX2_X1 U5150 ( .A(n4592), .B(n4663), .S(n4756), .Z(n4593) );
  OAI21_X1 U5151 ( .B1(n4609), .B2(n4666), .A(n4593), .ZN(U3532) );
  AOI21_X1 U5152 ( .B1(n4607), .B2(n4595), .A(n4594), .ZN(n4667) );
  MUX2_X1 U5153 ( .A(n2903), .B(n4667), .S(n4756), .Z(n4596) );
  OAI21_X1 U5154 ( .B1(n4609), .B2(n4670), .A(n4596), .ZN(U3531) );
  INV_X1 U5155 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U5156 ( .A1(n4600), .A2(n4599), .B1(n4598), .B2(n4597), .ZN(n4601)
         );
  OAI21_X1 U5157 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n4605) );
  AOI211_X1 U5158 ( .C1(n4607), .C2(n4606), .A(n4605), .B(n4604), .ZN(n4671)
         );
  MUX2_X1 U5159 ( .A(n4968), .B(n4671), .S(n4756), .Z(n4608) );
  OAI21_X1 U5160 ( .B1(n4609), .B2(n4675), .A(n4608), .ZN(U3530) );
  NAND3_X1 U5161 ( .A1(n2449), .A2(n4611), .A3(n4610), .ZN(n4612) );
  OAI211_X1 U5162 ( .C1(n4615), .C2(n4614), .A(n4613), .B(n4612), .ZN(n4676)
         );
  MUX2_X1 U5163 ( .A(REG1_REG_8__SCAN_IN), .B(n4676), .S(n4756), .Z(U3526) );
  NAND2_X1 U5164 ( .A1(n4751), .A2(n4616), .ZN(n4618) );
  NAND2_X1 U5165 ( .A1(n4749), .A2(REG0_REG_30__SCAN_IN), .ZN(n4617) );
  OAI211_X1 U5166 ( .C1(n4619), .C2(n4674), .A(n4618), .B(n4617), .ZN(U3516)
         );
  INV_X1 U5167 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4621) );
  INV_X1 U5168 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4837) );
  OAI21_X1 U5169 ( .B1(n4626), .B2(n4674), .A(n4625), .ZN(U3512) );
  INV_X1 U5170 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4628) );
  MUX2_X1 U5171 ( .A(n4628), .B(n4627), .S(n4751), .Z(n4629) );
  OAI21_X1 U5172 ( .B1(n4630), .B2(n4674), .A(n4629), .ZN(U3511) );
  INV_X1 U5173 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4632) );
  MUX2_X1 U5174 ( .A(n4632), .B(n4631), .S(n4751), .Z(n4633) );
  OAI21_X1 U5175 ( .B1(n4634), .B2(n4674), .A(n4633), .ZN(U3510) );
  INV_X1 U5176 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4635) );
  MUX2_X1 U5177 ( .A(n4636), .B(n4635), .S(n4749), .Z(n4637) );
  OAI21_X1 U5178 ( .B1(n4638), .B2(n4674), .A(n4637), .ZN(U3509) );
  MUX2_X1 U5179 ( .A(n4639), .B(REG0_REG_22__SCAN_IN), .S(n4749), .Z(n4640) );
  INV_X1 U5180 ( .A(n4640), .ZN(n4641) );
  OAI21_X1 U5181 ( .B1(n4642), .B2(n4674), .A(n4641), .ZN(U3508) );
  INV_X1 U5182 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4644) );
  MUX2_X1 U5183 ( .A(n4644), .B(n4643), .S(n4751), .Z(n4645) );
  OAI21_X1 U5184 ( .B1(n4646), .B2(n4674), .A(n4645), .ZN(U3507) );
  INV_X1 U5185 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4835) );
  MUX2_X1 U5186 ( .A(n4835), .B(n4647), .S(n4751), .Z(n4648) );
  OAI21_X1 U5187 ( .B1(n4649), .B2(n4674), .A(n4648), .ZN(U3506) );
  INV_X1 U5188 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4651) );
  MUX2_X1 U5189 ( .A(n4651), .B(n4650), .S(n4751), .Z(n4652) );
  OAI21_X1 U5190 ( .B1(n4653), .B2(n4674), .A(n4652), .ZN(U3505) );
  MUX2_X1 U5191 ( .A(REG0_REG_18__SCAN_IN), .B(n4654), .S(n4751), .Z(U3503) );
  INV_X1 U5192 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4656) );
  MUX2_X1 U5193 ( .A(n4656), .B(n4655), .S(n4751), .Z(n4657) );
  OAI21_X1 U5194 ( .B1(n4658), .B2(n4674), .A(n4657), .ZN(U3501) );
  MUX2_X1 U5195 ( .A(REG0_REG_16__SCAN_IN), .B(n4659), .S(n4751), .Z(U3499) );
  MUX2_X1 U5196 ( .A(n4931), .B(n4660), .S(n4751), .Z(n4661) );
  OAI21_X1 U5197 ( .B1(n4662), .B2(n4674), .A(n4661), .ZN(U3497) );
  INV_X1 U5198 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4664) );
  MUX2_X1 U5199 ( .A(n4664), .B(n4663), .S(n4751), .Z(n4665) );
  OAI21_X1 U5200 ( .B1(n4666), .B2(n4674), .A(n4665), .ZN(U3495) );
  INV_X1 U5201 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4668) );
  MUX2_X1 U5202 ( .A(n4668), .B(n4667), .S(n4751), .Z(n4669) );
  OAI21_X1 U5203 ( .B1(n4670), .B2(n4674), .A(n4669), .ZN(U3493) );
  INV_X1 U5204 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4672) );
  MUX2_X1 U5205 ( .A(n4672), .B(n4671), .S(n4751), .Z(n4673) );
  OAI21_X1 U5206 ( .B1(n4675), .B2(n4674), .A(n4673), .ZN(U3491) );
  MUX2_X1 U5207 ( .A(REG0_REG_8__SCAN_IN), .B(n4676), .S(n4751), .Z(U3483) );
  MUX2_X1 U5208 ( .A(DATAI_27_), .B(n4677), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5209 ( .A(n4678), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5210 ( .A(DATAI_25_), .B(n4679), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5211 ( .A(DATAI_20_), .B(n4680), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5212 ( .A(n4681), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5213 ( .A(n4682), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5214 ( .A(DATAI_14_), .B(n4683), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5215 ( .A(n4684), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5216 ( .A(n4685), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5217 ( .A(n4686), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5218 ( .A(n4687), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5219 ( .A(DATAI_6_), .B(n4688), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5220 ( .A(DATAI_4_), .B(n4689), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5221 ( .A(DATAI_3_), .B(n2248), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5222 ( .A(DATAI_2_), .B(n4690), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5223 ( .A(n2928), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5224 ( .A(DATAI_28_), .ZN(n4691) );
  AOI22_X1 U5225 ( .A1(STATE_REG_SCAN_IN), .A2(n4692), .B1(n4691), .B2(U3149), 
        .ZN(U3324) );
  AND2_X1 U5226 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4697) );
  AOI211_X1 U5227 ( .C1(n4695), .C2(n4694), .A(n4693), .B(n4703), .ZN(n4696)
         );
  AOI211_X1 U5228 ( .C1(n4709), .C2(ADDR_REG_15__SCAN_IN), .A(n4697), .B(n4696), .ZN(n4702) );
  OAI211_X1 U5229 ( .C1(n4700), .C2(n4699), .A(n4710), .B(n4698), .ZN(n4701)
         );
  OAI211_X1 U5230 ( .C1(n4715), .C2(n4735), .A(n4702), .B(n4701), .ZN(U3255)
         );
  AOI221_X1 U5231 ( .B1(n4706), .B2(n4705), .C1(n4704), .C2(n4705), .A(n4703), 
        .ZN(n4707) );
  AOI211_X1 U5232 ( .C1(n4709), .C2(ADDR_REG_16__SCAN_IN), .A(n4708), .B(n4707), .ZN(n4714) );
  OAI221_X1 U5233 ( .B1(n4712), .B2(REG1_REG_16__SCAN_IN), .C1(n4712), .C2(
        n4711), .A(n4710), .ZN(n4713) );
  OAI211_X1 U5234 ( .C1(n4715), .C2(n4733), .A(n4714), .B(n4713), .ZN(U3256)
         );
  OAI21_X1 U5235 ( .B1(n4718), .B2(n4717), .A(n4716), .ZN(n4719) );
  INV_X1 U5236 ( .A(n4719), .ZN(n4725) );
  AOI22_X1 U5237 ( .A1(n4722), .A2(n4721), .B1(REG3_REG_0__SCAN_IN), .B2(n4720), .ZN(n4723) );
  OAI221_X1 U5238 ( .B1(n4726), .B2(n4725), .C1(n4724), .C2(n2479), .A(n4723), 
        .ZN(U3290) );
  INV_X1 U5239 ( .A(D_REG_31__SCAN_IN), .ZN(n4904) );
  NOR2_X1 U5240 ( .A1(n4727), .A2(n4904), .ZN(U3291) );
  INV_X1 U5241 ( .A(D_REG_30__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U5242 ( .A1(n4727), .A2(n4898), .ZN(U3292) );
  INV_X1 U5243 ( .A(D_REG_29__SCAN_IN), .ZN(n4818) );
  NOR2_X1 U5244 ( .A1(n4727), .A2(n4818), .ZN(U3293) );
  AND2_X1 U5245 ( .A1(D_REG_28__SCAN_IN), .A2(n4728), .ZN(U3294) );
  AND2_X1 U5246 ( .A1(D_REG_27__SCAN_IN), .A2(n4728), .ZN(U3295) );
  INV_X1 U5247 ( .A(D_REG_26__SCAN_IN), .ZN(n4895) );
  NOR2_X1 U5248 ( .A1(n4727), .A2(n4895), .ZN(U3296) );
  INV_X1 U5249 ( .A(D_REG_25__SCAN_IN), .ZN(n4852) );
  NOR2_X1 U5250 ( .A1(n4727), .A2(n4852), .ZN(U3297) );
  AND2_X1 U5251 ( .A1(D_REG_24__SCAN_IN), .A2(n4728), .ZN(U3298) );
  AND2_X1 U5252 ( .A1(D_REG_23__SCAN_IN), .A2(n4728), .ZN(U3299) );
  INV_X1 U5253 ( .A(D_REG_22__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U5254 ( .A1(n4727), .A2(n4920), .ZN(U3300) );
  INV_X1 U5255 ( .A(D_REG_21__SCAN_IN), .ZN(n4853) );
  NOR2_X1 U5256 ( .A1(n4727), .A2(n4853), .ZN(U3301) );
  AND2_X1 U5257 ( .A1(D_REG_20__SCAN_IN), .A2(n4728), .ZN(U3302) );
  AND2_X1 U5258 ( .A1(D_REG_19__SCAN_IN), .A2(n4728), .ZN(U3303) );
  AND2_X1 U5259 ( .A1(D_REG_18__SCAN_IN), .A2(n4728), .ZN(U3304) );
  NOR2_X1 U5260 ( .A1(n4727), .A2(n4819), .ZN(U3305) );
  AND2_X1 U5261 ( .A1(D_REG_16__SCAN_IN), .A2(n4728), .ZN(U3306) );
  INV_X1 U5262 ( .A(D_REG_15__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U5263 ( .A1(n4727), .A2(n4912), .ZN(U3307) );
  NOR2_X1 U5264 ( .A1(n4727), .A2(n4828), .ZN(U3308) );
  NOR2_X1 U5265 ( .A1(n4727), .A2(n4830), .ZN(U3309) );
  NOR2_X1 U5266 ( .A1(n4727), .A2(n4829), .ZN(U3310) );
  AND2_X1 U5267 ( .A1(D_REG_11__SCAN_IN), .A2(n4728), .ZN(U3311) );
  AND2_X1 U5268 ( .A1(D_REG_10__SCAN_IN), .A2(n4728), .ZN(U3312) );
  AND2_X1 U5269 ( .A1(D_REG_9__SCAN_IN), .A2(n4728), .ZN(U3313) );
  AND2_X1 U5270 ( .A1(D_REG_8__SCAN_IN), .A2(n4728), .ZN(U3314) );
  INV_X1 U5271 ( .A(D_REG_7__SCAN_IN), .ZN(n4903) );
  NOR2_X1 U5272 ( .A1(n4727), .A2(n4903), .ZN(U3315) );
  AND2_X1 U5273 ( .A1(D_REG_6__SCAN_IN), .A2(n4728), .ZN(U3316) );
  AND2_X1 U5274 ( .A1(D_REG_5__SCAN_IN), .A2(n4728), .ZN(U3317) );
  AND2_X1 U5275 ( .A1(D_REG_4__SCAN_IN), .A2(n4728), .ZN(U3318) );
  AND2_X1 U5276 ( .A1(D_REG_3__SCAN_IN), .A2(n4728), .ZN(U3319) );
  AND2_X1 U5277 ( .A1(D_REG_2__SCAN_IN), .A2(n4728), .ZN(U3320) );
  INV_X1 U5278 ( .A(DATAI_23_), .ZN(n4730) );
  AOI21_X1 U5279 ( .B1(U3149), .B2(n4730), .A(n4729), .ZN(U3329) );
  AOI22_X1 U5280 ( .A1(STATE_REG_SCAN_IN), .A2(n4732), .B1(n4731), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5281 ( .A1(STATE_REG_SCAN_IN), .A2(n4733), .B1(n4910), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5282 ( .A(DATAI_15_), .ZN(n4734) );
  AOI22_X1 U5283 ( .A1(STATE_REG_SCAN_IN), .A2(n4735), .B1(n4734), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5284 ( .A(DATAI_0_), .ZN(n4736) );
  AOI22_X1 U5285 ( .A1(STATE_REG_SCAN_IN), .A2(n2235), .B1(n4736), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5286 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U5287 ( .A1(n4751), .A2(n4737), .B1(n4964), .B2(n4749), .ZN(U3467)
         );
  INV_X1 U5288 ( .A(n4738), .ZN(n4740) );
  AOI211_X1 U5289 ( .C1(n4742), .C2(n4741), .A(n4740), .B(n4739), .ZN(n4753)
         );
  INV_X1 U5290 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U5291 ( .A1(n4751), .A2(n4753), .B1(n4954), .B2(n4749), .ZN(U3475)
         );
  OR3_X1 U5292 ( .A1(n4745), .A2(n4744), .A3(n4743), .ZN(n4746) );
  AND3_X1 U5293 ( .A1(n4748), .A2(n4747), .A3(n4746), .ZN(n4755) );
  INV_X1 U5294 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5295 ( .A1(n4751), .A2(n4755), .B1(n4750), .B2(n4749), .ZN(U3481)
         );
  AOI22_X1 U5296 ( .A1(n4756), .A2(n4753), .B1(n4752), .B2(n4754), .ZN(U3522)
         );
  AOI22_X1 U5297 ( .A1(n4756), .A2(n4755), .B1(n4796), .B2(n4754), .ZN(U3525)
         );
  NAND4_X1 U5298 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .A3(
        REG2_REG_25__SCAN_IN), .A4(n2965), .ZN(n4757) );
  NOR4_X1 U5299 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_27__SCAN_IN), .A3(
        ADDR_REG_6__SCAN_IN), .A4(n4757), .ZN(n4760) );
  NAND4_X1 U5300 ( .A1(REG2_REG_21__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        DATAI_31_), .A4(n4340), .ZN(n4758) );
  NOR3_X1 U5301 ( .A1(REG2_REG_23__SCAN_IN), .A2(REG2_REG_24__SCAN_IN), .A3(
        n4758), .ZN(n4759) );
  NAND4_X1 U5302 ( .A1(REG2_REG_26__SCAN_IN), .A2(REG2_REG_31__SCAN_IN), .A3(
        n4760), .A4(n4759), .ZN(n4775) );
  NAND4_X1 U5303 ( .A1(REG2_REG_29__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(
        n4983), .A4(n2660), .ZN(n4761) );
  NOR3_X1 U5304 ( .A1(ADDR_REG_19__SCAN_IN), .A2(n4997), .A3(n4761), .ZN(n4762) );
  NAND4_X1 U5305 ( .A1(B_REG_SCAN_IN), .A2(n4763), .A3(REG3_REG_28__SCAN_IN), 
        .A4(n4762), .ZN(n4774) );
  NOR4_X1 U5306 ( .A1(ADDR_REG_15__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(DATAO_REG_13__SCAN_IN), .ZN(n4767) );
  NOR4_X1 U5307 ( .A1(IR_REG_25__SCAN_IN), .A2(DATAO_REG_3__SCAN_IN), .A3(
        DATAO_REG_24__SCAN_IN), .A4(DATAO_REG_23__SCAN_IN), .ZN(n4766) );
  NOR4_X1 U5308 ( .A1(IR_REG_29__SCAN_IN), .A2(ADDR_REG_0__SCAN_IN), .A3(n4910), .A4(n4917), .ZN(n4765) );
  INV_X1 U5309 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4897) );
  NOR4_X1 U5310 ( .A1(DATAI_13_), .A2(DATAO_REG_6__SCAN_IN), .A3(n4897), .A4(
        n4900), .ZN(n4764) );
  NAND4_X1 U5311 ( .A1(n4767), .A2(n4766), .A3(n4765), .A4(n4764), .ZN(n4773)
         );
  INV_X1 U5312 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4846) );
  NOR4_X1 U5313 ( .A1(IR_REG_30__SCAN_IN), .A2(REG1_REG_31__SCAN_IN), .A3(
        n2264), .A4(n4846), .ZN(n4771) );
  NOR4_X1 U5314 ( .A1(n4855), .A2(n3227), .A3(n4866), .A4(REG0_REG_30__SCAN_IN), .ZN(n4770) );
  NOR4_X1 U5315 ( .A1(D_REG_0__SCAN_IN), .A2(REG0_REG_25__SCAN_IN), .A3(
        DATAO_REG_12__SCAN_IN), .A4(DATAO_REG_16__SCAN_IN), .ZN(n4769) );
  INV_X1 U5316 ( .A(DATAI_20_), .ZN(n4868) );
  NOR4_X1 U5317 ( .A1(n4871), .A2(n4868), .A3(n4865), .A4(n4869), .ZN(n4768)
         );
  NAND4_X1 U5318 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4772)
         );
  NOR4_X1 U5319 ( .A1(n4775), .A2(n4774), .A3(n4773), .A4(n4772), .ZN(n4805)
         );
  NAND4_X1 U5320 ( .A1(REG0_REG_27__SCAN_IN), .A2(REG0_REG_26__SCAN_IN), .A3(
        n4513), .A4(n4839), .ZN(n4776) );
  NOR3_X1 U5321 ( .A1(REG0_REG_23__SCAN_IN), .A2(REG0_REG_21__SCAN_IN), .A3(
        n4776), .ZN(n4804) );
  NAND4_X1 U5322 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n4783) );
  INV_X1 U5323 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4778) );
  INV_X1 U5324 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4777) );
  NAND4_X1 U5325 ( .A1(n4778), .A2(n4777), .A3(DATAI_7_), .A4(
        D_REG_29__SCAN_IN), .ZN(n4782) );
  NAND4_X1 U5326 ( .A1(n4779), .A2(REG3_REG_2__SCAN_IN), .A3(
        REG0_REG_2__SCAN_IN), .A4(DATAI_1_), .ZN(n4781) );
  INV_X1 U5327 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4808) );
  OR4_X1 U5328 ( .A1(DATAI_8_), .A2(n4808), .A3(REG1_REG_8__SCAN_IN), .A4(
        REG0_REG_6__SCAN_IN), .ZN(n4780) );
  NOR4_X1 U5329 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4795)
         );
  INV_X1 U5330 ( .A(n4784), .ZN(n4791) );
  NAND4_X1 U5331 ( .A1(n4785), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_5__SCAN_IN), 
        .A4(IR_REG_11__SCAN_IN), .ZN(n4790) );
  NAND4_X1 U5332 ( .A1(IR_REG_3__SCAN_IN), .A2(DATAI_4_), .A3(DATAI_3_), .A4(
        REG0_REG_3__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U5333 ( .A1(REG0_REG_0__SCAN_IN), .A2(n4786), .ZN(n4788) );
  NOR4_X1 U5334 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_8__SCAN_IN), .A3(
        REG1_REG_6__SCAN_IN), .A4(ADDR_REG_7__SCAN_IN), .ZN(n4787) );
  NAND4_X1 U5335 ( .A1(n4788), .A2(n4954), .A3(n3697), .A4(n4787), .ZN(n4789)
         );
  NOR4_X1 U5336 ( .A1(n4791), .A2(n4790), .A3(IR_REG_12__SCAN_IN), .A4(n4789), 
        .ZN(n4794) );
  NOR4_X1 U5337 ( .A1(n4823), .A2(IR_REG_14__SCAN_IN), .A3(REG3_REG_4__SCAN_IN), .A4(REG3_REG_5__SCAN_IN), .ZN(n4793) );
  NOR4_X1 U5338 ( .A1(n4835), .A2(DATAI_26_), .A3(REG1_REG_12__SCAN_IN), .A4(
        DATAI_10_), .ZN(n4792) );
  NAND4_X1 U5339 ( .A1(n4795), .A2(n4794), .A3(n4793), .A4(n4792), .ZN(n4802)
         );
  INV_X1 U5340 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4943) );
  NOR4_X1 U5341 ( .A1(REG1_REG_11__SCAN_IN), .A2(ADDR_REG_17__SCAN_IN), .A3(
        n4796), .A4(n4943), .ZN(n4800) );
  INV_X1 U5342 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n5008) );
  NOR4_X1 U5343 ( .A1(REG3_REG_14__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        ADDR_REG_8__SCAN_IN), .A4(n5008), .ZN(n4799) );
  NOR4_X1 U5344 ( .A1(REG0_REG_15__SCAN_IN), .A2(n3759), .A3(n2937), .A4(n2941), .ZN(n4798) );
  NOR4_X1 U5345 ( .A1(REG2_REG_1__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .A3(
        n2927), .A4(n4944), .ZN(n4797) );
  NAND4_X1 U5346 ( .A1(n4800), .A2(n4799), .A3(n4798), .A4(n4797), .ZN(n4801)
         );
  NOR2_X1 U5347 ( .A1(n4802), .A2(n4801), .ZN(n4803) );
  AND3_X1 U5348 ( .A1(n4805), .A2(n4804), .A3(n4803), .ZN(n5036) );
  INV_X1 U5349 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4807) );
  AOI22_X1 U5350 ( .A1(n4808), .A2(keyinput73), .B1(n4807), .B2(keyinput16), 
        .ZN(n4806) );
  OAI221_X1 U5351 ( .B1(n4808), .B2(keyinput73), .C1(n4807), .C2(keyinput16), 
        .A(n4806), .ZN(n4816) );
  XNOR2_X1 U5352 ( .A(DATAI_8_), .B(keyinput4), .ZN(n4812) );
  XNOR2_X1 U5353 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput79), .ZN(n4811) );
  XNOR2_X1 U5354 ( .A(IR_REG_9__SCAN_IN), .B(keyinput58), .ZN(n4810) );
  XNOR2_X1 U5355 ( .A(IR_REG_8__SCAN_IN), .B(keyinput46), .ZN(n4809) );
  NAND4_X1 U5356 ( .A1(n4812), .A2(n4811), .A3(n4810), .A4(n4809), .ZN(n4815)
         );
  XNOR2_X1 U5357 ( .A(keyinput14), .B(n2514), .ZN(n4814) );
  XNOR2_X1 U5358 ( .A(keyinput117), .B(n3697), .ZN(n4813) );
  NOR4_X1 U5359 ( .A1(n4816), .A2(n4815), .A3(n4814), .A4(n4813), .ZN(n4863)
         );
  AOI22_X1 U5360 ( .A1(n4819), .A2(keyinput53), .B1(keyinput126), .B2(n4818), 
        .ZN(n4817) );
  OAI221_X1 U5361 ( .B1(n4819), .B2(keyinput53), .C1(n4818), .C2(keyinput126), 
        .A(n4817), .ZN(n4826) );
  AOI22_X1 U5362 ( .A1(n4822), .A2(keyinput19), .B1(keyinput9), .B2(n4821), 
        .ZN(n4820) );
  OAI221_X1 U5363 ( .B1(n4822), .B2(keyinput19), .C1(n4821), .C2(keyinput9), 
        .A(n4820), .ZN(n4825) );
  XNOR2_X1 U5364 ( .A(n4823), .B(keyinput90), .ZN(n4824) );
  OR3_X1 U5365 ( .A1(n4826), .A2(n4825), .A3(n4824), .ZN(n4833) );
  AOI22_X1 U5366 ( .A1(n4829), .A2(keyinput121), .B1(keyinput116), .B2(n4828), 
        .ZN(n4827) );
  OAI221_X1 U5367 ( .B1(n4829), .B2(keyinput121), .C1(n4828), .C2(keyinput116), 
        .A(n4827), .ZN(n4832) );
  XNOR2_X1 U5368 ( .A(n4830), .B(keyinput120), .ZN(n4831) );
  NOR3_X1 U5369 ( .A1(n4833), .A2(n4832), .A3(n4831), .ZN(n4862) );
  AOI22_X1 U5370 ( .A1(n4835), .A2(keyinput127), .B1(n4644), .B2(keyinput80), 
        .ZN(n4834) );
  OAI221_X1 U5371 ( .B1(n4835), .B2(keyinput127), .C1(n4644), .C2(keyinput80), 
        .A(n4834), .ZN(n4844) );
  AOI22_X1 U5372 ( .A1(n4635), .A2(keyinput50), .B1(n4837), .B2(keyinput13), 
        .ZN(n4836) );
  OAI221_X1 U5373 ( .B1(n4635), .B2(keyinput50), .C1(n4837), .C2(keyinput13), 
        .A(n4836), .ZN(n4843) );
  AOI22_X1 U5374 ( .A1(n4839), .A2(keyinput62), .B1(n4621), .B2(keyinput103), 
        .ZN(n4838) );
  OAI221_X1 U5375 ( .B1(n4839), .B2(keyinput62), .C1(n4621), .C2(keyinput103), 
        .A(n4838), .ZN(n4842) );
  AOI22_X1 U5376 ( .A1(n4513), .A2(keyinput21), .B1(n3227), .B2(keyinput111), 
        .ZN(n4840) );
  OAI221_X1 U5377 ( .B1(n4513), .B2(keyinput21), .C1(n3227), .C2(keyinput111), 
        .A(n4840), .ZN(n4841) );
  NOR4_X1 U5378 ( .A1(n4844), .A2(n4843), .A3(n4842), .A4(n4841), .ZN(n4861)
         );
  INV_X1 U5379 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4847) );
  AOI22_X1 U5380 ( .A1(n4847), .A2(keyinput10), .B1(keyinput99), .B2(n4846), 
        .ZN(n4845) );
  OAI221_X1 U5381 ( .B1(n4847), .B2(keyinput10), .C1(n4846), .C2(keyinput99), 
        .A(n4845), .ZN(n4859) );
  INV_X1 U5382 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U5383 ( .A1(n4850), .A2(keyinput1), .B1(n4849), .B2(keyinput39), 
        .ZN(n4848) );
  OAI221_X1 U5384 ( .B1(n4850), .B2(keyinput1), .C1(n4849), .C2(keyinput39), 
        .A(n4848), .ZN(n4858) );
  AOI22_X1 U5385 ( .A1(n4853), .A2(keyinput55), .B1(keyinput83), .B2(n4852), 
        .ZN(n4851) );
  OAI221_X1 U5386 ( .B1(n4853), .B2(keyinput55), .C1(n4852), .C2(keyinput83), 
        .A(n4851), .ZN(n4857) );
  AOI22_X1 U5387 ( .A1(n2264), .A2(keyinput3), .B1(n4855), .B2(keyinput7), 
        .ZN(n4854) );
  OAI221_X1 U5388 ( .B1(n2264), .B2(keyinput3), .C1(n4855), .C2(keyinput7), 
        .A(n4854), .ZN(n4856) );
  NOR4_X1 U5389 ( .A1(n4859), .A2(n4858), .A3(n4857), .A4(n4856), .ZN(n4860)
         );
  NAND4_X1 U5390 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n5033)
         );
  AOI22_X1 U5391 ( .A1(n4866), .A2(keyinput91), .B1(keyinput107), .B2(n4865), 
        .ZN(n4864) );
  OAI221_X1 U5392 ( .B1(n4866), .B2(keyinput91), .C1(n4865), .C2(keyinput107), 
        .A(n4864), .ZN(n4878) );
  AOI22_X1 U5393 ( .A1(n4869), .A2(keyinput115), .B1(n4868), .B2(keyinput59), 
        .ZN(n4867) );
  OAI221_X1 U5394 ( .B1(n4869), .B2(keyinput115), .C1(n4868), .C2(keyinput59), 
        .A(n4867), .ZN(n4877) );
  AOI22_X1 U5395 ( .A1(n4871), .A2(keyinput75), .B1(keyinput26), .B2(n4628), 
        .ZN(n4870) );
  OAI221_X1 U5396 ( .B1(n4871), .B2(keyinput75), .C1(n4628), .C2(keyinput26), 
        .A(n4870), .ZN(n4876) );
  AOI22_X1 U5397 ( .A1(n4874), .A2(keyinput22), .B1(keyinput25), .B2(n4873), 
        .ZN(n4872) );
  OAI221_X1 U5398 ( .B1(n4874), .B2(keyinput22), .C1(n4873), .C2(keyinput25), 
        .A(n4872), .ZN(n4875) );
  NOR4_X1 U5399 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4928)
         );
  AOI22_X1 U5400 ( .A1(n4881), .A2(keyinput5), .B1(keyinput122), .B2(n4880), 
        .ZN(n4879) );
  OAI221_X1 U5401 ( .B1(n4881), .B2(keyinput5), .C1(n4880), .C2(keyinput122), 
        .A(n4879), .ZN(n4892) );
  AOI22_X1 U5402 ( .A1(n4884), .A2(keyinput33), .B1(keyinput6), .B2(n4883), 
        .ZN(n4882) );
  OAI221_X1 U5403 ( .B1(n4884), .B2(keyinput33), .C1(n4883), .C2(keyinput6), 
        .A(n4882), .ZN(n4891) );
  INV_X1 U5404 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5405 ( .A1(n4886), .A2(keyinput118), .B1(keyinput106), .B2(n3291), 
        .ZN(n4885) );
  OAI221_X1 U5406 ( .B1(n4886), .B2(keyinput118), .C1(n3291), .C2(keyinput106), 
        .A(n4885), .ZN(n4890) );
  XNOR2_X1 U5407 ( .A(D_REG_0__SCAN_IN), .B(keyinput24), .ZN(n4888) );
  XNOR2_X1 U5408 ( .A(IR_REG_25__SCAN_IN), .B(keyinput36), .ZN(n4887) );
  NAND2_X1 U5409 ( .A1(n4888), .A2(n4887), .ZN(n4889) );
  NOR4_X1 U5410 ( .A1(n4892), .A2(n4891), .A3(n4890), .A4(n4889), .ZN(n4927)
         );
  AOI22_X1 U5411 ( .A1(n4895), .A2(keyinput109), .B1(keyinput104), .B2(n4894), 
        .ZN(n4893) );
  OAI221_X1 U5412 ( .B1(n4895), .B2(keyinput109), .C1(n4894), .C2(keyinput104), 
        .A(n4893), .ZN(n4908) );
  AOI22_X1 U5413 ( .A1(n4898), .A2(keyinput100), .B1(keyinput102), .B2(n4897), 
        .ZN(n4896) );
  OAI221_X1 U5414 ( .B1(n4898), .B2(keyinput100), .C1(n4897), .C2(keyinput102), 
        .A(n4896), .ZN(n4907) );
  INV_X1 U5415 ( .A(DATAI_13_), .ZN(n4901) );
  AOI22_X1 U5416 ( .A1(n4901), .A2(keyinput101), .B1(keyinput96), .B2(n4900), 
        .ZN(n4899) );
  OAI221_X1 U5417 ( .B1(n4901), .B2(keyinput101), .C1(n4900), .C2(keyinput96), 
        .A(n4899), .ZN(n4906) );
  AOI22_X1 U5418 ( .A1(n4904), .A2(keyinput92), .B1(keyinput86), .B2(n4903), 
        .ZN(n4902) );
  OAI221_X1 U5419 ( .B1(n4904), .B2(keyinput92), .C1(n4903), .C2(keyinput86), 
        .A(n4902), .ZN(n4905) );
  NOR4_X1 U5420 ( .A1(n4908), .A2(n4907), .A3(n4906), .A4(n4905), .ZN(n4926)
         );
  INV_X1 U5421 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U5422 ( .A1(n4911), .A2(keyinput77), .B1(n4910), .B2(keyinput72), 
        .ZN(n4909) );
  OAI221_X1 U5423 ( .B1(n4911), .B2(keyinput77), .C1(n4910), .C2(keyinput72), 
        .A(n4909), .ZN(n4915) );
  XNOR2_X1 U5424 ( .A(n4912), .B(keyinput64), .ZN(n4914) );
  XOR2_X1 U5425 ( .A(IR_REG_29__SCAN_IN), .B(keyinput60), .Z(n4913) );
  OR3_X1 U5426 ( .A1(n4915), .A2(n4914), .A3(n4913), .ZN(n4924) );
  AOI22_X1 U5427 ( .A1(n4918), .A2(keyinput82), .B1(keyinput81), .B2(n4917), 
        .ZN(n4916) );
  OAI221_X1 U5428 ( .B1(n4918), .B2(keyinput82), .C1(n4917), .C2(keyinput81), 
        .A(n4916), .ZN(n4923) );
  INV_X1 U5429 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4921) );
  AOI22_X1 U5430 ( .A1(n4921), .A2(keyinput52), .B1(n4920), .B2(keyinput45), 
        .ZN(n4919) );
  OAI221_X1 U5431 ( .B1(n4921), .B2(keyinput52), .C1(n4920), .C2(keyinput45), 
        .A(n4919), .ZN(n4922) );
  NOR3_X1 U5432 ( .A1(n4924), .A2(n4923), .A3(n4922), .ZN(n4925) );
  NAND4_X1 U5433 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n5032)
         );
  AOI22_X1 U5434 ( .A1(n2927), .A2(keyinput61), .B1(n2937), .B2(keyinput124), 
        .ZN(n4929) );
  OAI221_X1 U5435 ( .B1(n2927), .B2(keyinput61), .C1(n2937), .C2(keyinput124), 
        .A(n4929), .ZN(n4938) );
  AOI22_X1 U5436 ( .A1(n2941), .A2(keyinput68), .B1(n3759), .B2(keyinput31), 
        .ZN(n4930) );
  OAI221_X1 U5437 ( .B1(n2941), .B2(keyinput68), .C1(n3759), .C2(keyinput31), 
        .A(n4930), .ZN(n4937) );
  INV_X1 U5438 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4931) );
  XOR2_X1 U5439 ( .A(n4931), .B(keyinput57), .Z(n4935) );
  XNOR2_X1 U5440 ( .A(IR_REG_11__SCAN_IN), .B(keyinput38), .ZN(n4934) );
  XNOR2_X1 U5441 ( .A(IR_REG_12__SCAN_IN), .B(keyinput88), .ZN(n4933) );
  XNOR2_X1 U5442 ( .A(IR_REG_14__SCAN_IN), .B(keyinput63), .ZN(n4932) );
  NAND4_X1 U5443 ( .A1(n4935), .A2(n4934), .A3(n4933), .A4(n4932), .ZN(n4936)
         );
  NOR3_X1 U5444 ( .A1(n4938), .A2(n4937), .A3(n4936), .ZN(n4980) );
  INV_X1 U5445 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5446 ( .A1(n4941), .A2(keyinput11), .B1(n4940), .B2(keyinput112), 
        .ZN(n4939) );
  OAI221_X1 U5447 ( .B1(n4941), .B2(keyinput11), .C1(n4940), .C2(keyinput112), 
        .A(n4939), .ZN(n4951) );
  AOI22_X1 U5448 ( .A1(n2261), .A2(keyinput119), .B1(keyinput114), .B2(n4943), 
        .ZN(n4942) );
  OAI221_X1 U5449 ( .B1(n2261), .B2(keyinput119), .C1(n4943), .C2(keyinput114), 
        .A(n4942), .ZN(n4950) );
  XOR2_X1 U5450 ( .A(n4944), .B(keyinput34), .Z(n4948) );
  XNOR2_X1 U5451 ( .A(keyinput30), .B(REG1_REG_7__SCAN_IN), .ZN(n4947) );
  XNOR2_X1 U5452 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput8), .ZN(n4946) );
  XNOR2_X1 U5453 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput65), .ZN(n4945) );
  NAND4_X1 U5454 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4945), .ZN(n4949)
         );
  NOR3_X1 U5455 ( .A1(n4951), .A2(n4950), .A3(n4949), .ZN(n4979) );
  AOI22_X1 U5456 ( .A1(n3451), .A2(keyinput43), .B1(n2495), .B2(keyinput87), 
        .ZN(n4952) );
  OAI221_X1 U5457 ( .B1(n3451), .B2(keyinput43), .C1(n2495), .C2(keyinput87), 
        .A(n4952), .ZN(n4962) );
  INV_X1 U5458 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U5459 ( .A(keyinput108), .B(n4953), .ZN(n4961) );
  XNOR2_X1 U5460 ( .A(keyinput76), .B(n4954), .ZN(n4960) );
  XNOR2_X1 U5461 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput44), .ZN(n4958) );
  XNOR2_X1 U5462 ( .A(IR_REG_3__SCAN_IN), .B(keyinput71), .ZN(n4957) );
  XNOR2_X1 U5463 ( .A(IR_REG_4__SCAN_IN), .B(keyinput74), .ZN(n4956) );
  XNOR2_X1 U5464 ( .A(DATAI_4_), .B(keyinput12), .ZN(n4955) );
  NAND4_X1 U5465 ( .A1(n4958), .A2(n4957), .A3(n4956), .A4(n4955), .ZN(n4959)
         );
  NOR4_X1 U5466 ( .A1(n4962), .A2(n4961), .A3(n4960), .A4(n4959), .ZN(n4978)
         );
  AOI22_X1 U5467 ( .A1(n4965), .A2(keyinput105), .B1(keyinput2), .B2(n4964), 
        .ZN(n4963) );
  OAI221_X1 U5468 ( .B1(n4965), .B2(keyinput105), .C1(n4964), .C2(keyinput2), 
        .A(n4963), .ZN(n4976) );
  INV_X1 U5469 ( .A(DATAI_10_), .ZN(n4967) );
  AOI22_X1 U5470 ( .A1(n4968), .A2(keyinput42), .B1(keyinput89), .B2(n4967), 
        .ZN(n4966) );
  OAI221_X1 U5471 ( .B1(n4968), .B2(keyinput42), .C1(n4967), .C2(keyinput89), 
        .A(n4966), .ZN(n4975) );
  XOR2_X1 U5472 ( .A(n2538), .B(keyinput70), .Z(n4973) );
  INV_X1 U5473 ( .A(DATAI_1_), .ZN(n4969) );
  XOR2_X1 U5474 ( .A(n4969), .B(keyinput78), .Z(n4972) );
  XNOR2_X1 U5475 ( .A(IR_REG_7__SCAN_IN), .B(keyinput40), .ZN(n4971) );
  XNOR2_X1 U5476 ( .A(DATAI_2_), .B(keyinput69), .ZN(n4970) );
  NAND4_X1 U5477 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n4970), .ZN(n4974)
         );
  NOR3_X1 U5478 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n4977) );
  NAND4_X1 U5479 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n5031)
         );
  AOI22_X1 U5480 ( .A1(n2753), .A2(keyinput18), .B1(keyinput98), .B2(n2742), 
        .ZN(n4981) );
  OAI221_X1 U5481 ( .B1(n2753), .B2(keyinput18), .C1(n2742), .C2(keyinput98), 
        .A(n4981), .ZN(n4991) );
  AOI22_X1 U5482 ( .A1(U3149), .A2(keyinput37), .B1(keyinput29), .B2(n4983), 
        .ZN(n4982) );
  OAI221_X1 U5483 ( .B1(U3149), .B2(keyinput37), .C1(n4983), .C2(keyinput29), 
        .A(n4982), .ZN(n4990) );
  AOI22_X1 U5484 ( .A1(n2730), .A2(keyinput20), .B1(keyinput23), .B2(n2714), 
        .ZN(n4984) );
  OAI221_X1 U5485 ( .B1(n2730), .B2(keyinput20), .C1(n2714), .C2(keyinput23), 
        .A(n4984), .ZN(n4989) );
  AOI22_X1 U5486 ( .A1(n4987), .A2(keyinput28), .B1(keyinput67), .B2(n4986), 
        .ZN(n4985) );
  OAI221_X1 U5487 ( .B1(n4987), .B2(keyinput28), .C1(n4986), .C2(keyinput67), 
        .A(n4985), .ZN(n4988) );
  NOR4_X1 U5488 ( .A1(n4991), .A2(n4990), .A3(n4989), .A4(n4988), .ZN(n5029)
         );
  NAND2_X1 U5489 ( .A1(n2723), .A2(keyinput110), .ZN(n4992) );
  OAI221_X1 U5490 ( .B1(n5035), .B2(keyinput27), .C1(n2723), .C2(keyinput110), 
        .A(n4992), .ZN(n5001) );
  AOI22_X1 U5491 ( .A1(n2747), .A2(keyinput54), .B1(keyinput47), .B2(n4244), 
        .ZN(n4993) );
  OAI221_X1 U5492 ( .B1(n2747), .B2(keyinput54), .C1(n4244), .C2(keyinput47), 
        .A(n4993), .ZN(n5000) );
  INV_X1 U5493 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4995) );
  AOI22_X1 U5494 ( .A1(n4995), .A2(keyinput125), .B1(n2660), .B2(keyinput35), 
        .ZN(n4994) );
  OAI221_X1 U5495 ( .B1(n4995), .B2(keyinput125), .C1(n2660), .C2(keyinput35), 
        .A(n4994), .ZN(n4999) );
  AOI22_X1 U5496 ( .A1(n2965), .A2(keyinput17), .B1(n4997), .B2(keyinput15), 
        .ZN(n4996) );
  OAI221_X1 U5497 ( .B1(n2965), .B2(keyinput17), .C1(n4997), .C2(keyinput15), 
        .A(n4996), .ZN(n4998) );
  NOR4_X1 U5498 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n5028)
         );
  INV_X1 U5499 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n5003) );
  AOI22_X1 U5500 ( .A1(n5004), .A2(keyinput94), .B1(keyinput113), .B2(n5003), 
        .ZN(n5002) );
  OAI221_X1 U5501 ( .B1(n5004), .B2(keyinput94), .C1(n5003), .C2(keyinput113), 
        .A(n5002), .ZN(n5014) );
  AOI22_X1 U5502 ( .A1(n4777), .A2(keyinput0), .B1(n2235), .B2(keyinput95), 
        .ZN(n5005) );
  OAI221_X1 U5503 ( .B1(n4777), .B2(keyinput0), .C1(n2235), .C2(keyinput95), 
        .A(n5005), .ZN(n5013) );
  INV_X1 U5504 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U5505 ( .A1(n5008), .A2(keyinput49), .B1(n5007), .B2(keyinput32), 
        .ZN(n5006) );
  OAI221_X1 U5506 ( .B1(n5008), .B2(keyinput49), .C1(n5007), .C2(keyinput32), 
        .A(n5006), .ZN(n5012) );
  INV_X1 U5507 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U5508 ( .A1(n3615), .A2(keyinput84), .B1(keyinput85), .B2(n5010), 
        .ZN(n5009) );
  OAI221_X1 U5509 ( .B1(n3615), .B2(keyinput84), .C1(n5010), .C2(keyinput85), 
        .A(n5009), .ZN(n5011) );
  NOR4_X1 U5510 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n5027)
         );
  AOI22_X1 U5511 ( .A1(n4318), .A2(keyinput97), .B1(keyinput48), .B2(n4340), 
        .ZN(n5015) );
  OAI221_X1 U5512 ( .B1(n4318), .B2(keyinput97), .C1(n4340), .C2(keyinput48), 
        .A(n5015), .ZN(n5025) );
  AOI22_X1 U5513 ( .A1(n4353), .A2(keyinput123), .B1(keyinput51), .B2(n4380), 
        .ZN(n5016) );
  OAI221_X1 U5514 ( .B1(n4353), .B2(keyinput123), .C1(n4380), .C2(keyinput51), 
        .A(n5016), .ZN(n5024) );
  INV_X1 U5515 ( .A(DATAI_26_), .ZN(n5018) );
  AOI22_X1 U5516 ( .A1(n5019), .A2(keyinput66), .B1(n5018), .B2(keyinput56), 
        .ZN(n5017) );
  OAI221_X1 U5517 ( .B1(n5019), .B2(keyinput66), .C1(n5018), .C2(keyinput56), 
        .A(n5017), .ZN(n5023) );
  XOR2_X1 U5518 ( .A(n4778), .B(keyinput93), .Z(n5021) );
  XNOR2_X1 U5519 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput41), .ZN(n5020) );
  NAND2_X1 U5520 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  NOR4_X1 U5521 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5026)
         );
  NAND4_X1 U5522 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n5030)
         );
  OR4_X1 U5523 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5034) );
  AOI221_X1 U5524 ( .B1(n5036), .B2(keyinput27), .C1(n5035), .C2(keyinput27), 
        .A(n5034), .ZN(n5040) );
  NAND2_X1 U5525 ( .A1(n5037), .A2(U4043), .ZN(n5038) );
  OAI21_X1 U5526 ( .B1(U4043), .B2(DATAO_REG_25__SCAN_IN), .A(n5038), .ZN(
        n5039) );
  XNOR2_X1 U5527 ( .A(n5040), .B(n5039), .ZN(U3575) );
  INV_X1 U2384 ( .A(IR_REG_31__SCAN_IN), .ZN(n2791) );
  CLKBUF_X1 U2382 ( .A(n2998), .Z(n3095) );
  AND2_X1 U2385 ( .A1(n4510), .A2(n2303), .ZN(n4620) );
endmodule

