

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16491,
         n16492;

  AND2_X1 U7530 ( .A1(n14477), .A2(n8162), .ZN(n14431) );
  NAND2_X1 U7531 ( .A1(n9796), .A2(n14457), .ZN(n9900) );
  INV_X4 U7532 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OAI21_X1 U7533 ( .B1(n8117), .B2(n8113), .A(n8109), .ZN(n13892) );
  NAND2_X1 U7534 ( .A1(n9783), .A2(n9782), .ZN(n14664) );
  OR2_X1 U7535 ( .A1(n14554), .A2(n9718), .ZN(n9720) );
  NAND2_X1 U7536 ( .A1(n9743), .A2(n9742), .ZN(n14530) );
  NOR2_X1 U7537 ( .A1(n13119), .A2(n13120), .ZN(n13700) );
  NOR2_X1 U7538 ( .A1(n13117), .A2(n13118), .ZN(n13119) );
  INV_X2 U7539 ( .A(n14935), .ZN(n14831) );
  BUF_X1 U7541 ( .A(n11134), .Z(n15060) );
  INV_X1 U7542 ( .A(n11130), .ZN(n12183) );
  INV_X1 U7543 ( .A(n8633), .ZN(n8983) );
  NAND4_X1 U7544 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n15449) );
  CLKBUF_X2 U7546 ( .A(n8611), .Z(n8960) );
  CLKBUF_X3 U7547 ( .A(n10687), .Z(n7431) );
  CLKBUF_X2 U7548 ( .A(n11485), .Z(n7432) );
  BUF_X4 U7549 ( .A(n10831), .Z(n7434) );
  INV_X2 U7550 ( .A(n10137), .ZN(n9754) );
  INV_X1 U7551 ( .A(n9380), .ZN(n9388) );
  INV_X1 U7552 ( .A(n11067), .ZN(n9421) );
  INV_X1 U7554 ( .A(n16492), .ZN(n7430) );
  INV_X1 U7555 ( .A(n7436), .ZN(n10650) );
  INV_X4 U7556 ( .A(n10358), .ZN(n7436) );
  INV_X1 U7557 ( .A(n15236), .ZN(n15239) );
  NOR2_X1 U7558 ( .A1(n16422), .A2(n12897), .ZN(n13117) );
  NAND2_X1 U7559 ( .A1(n8825), .A2(n8824), .ZN(n14003) );
  NAND2_X1 U7560 ( .A1(n14586), .A2(n11149), .ZN(n14242) );
  OR2_X1 U7561 ( .A1(n12737), .A2(n12736), .ZN(n12740) );
  INV_X1 U7562 ( .A(n7663), .ZN(n13309) );
  NOR2_X1 U7563 ( .A1(n13466), .A2(n13608), .ZN(n13617) );
  INV_X1 U7565 ( .A(n11215), .ZN(n8304) );
  NAND2_X1 U7566 ( .A1(n14408), .A2(n14305), .ZN(n11387) );
  INV_X1 U7568 ( .A(n8611), .ZN(n8915) );
  OAI211_X1 U7569 ( .C1(n13680), .C2(n7432), .A(n8623), .B(n8622), .ZN(n12427)
         );
  OR2_X1 U7570 ( .A1(n8561), .A2(n14231), .ZN(n8563) );
  INV_X1 U7571 ( .A(n9388), .ZN(n10117) );
  CLKBUF_X3 U7573 ( .A(n14265), .Z(n14305) );
  INV_X1 U7574 ( .A(n7431), .ZN(n10714) );
  INV_X1 U7575 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n16268) );
  XNOR2_X1 U7576 ( .A(n8563), .B(n8562), .ZN(n13183) );
  NAND2_X1 U7577 ( .A1(n7492), .A2(n9426), .ZN(n14408) );
  BUF_X1 U7578 ( .A(n7725), .Z(n7660) );
  INV_X1 U7579 ( .A(n10257), .ZN(n15621) );
  INV_X1 U7580 ( .A(n10303), .ZN(n10687) );
  NAND2_X1 U7581 ( .A1(n13183), .A2(n13775), .ZN(n11485) );
  BUF_X1 U7582 ( .A(n9390), .Z(n10120) );
  NAND2_X2 U7583 ( .A1(n7743), .A2(n7742), .ZN(n10000) );
  NAND2_X2 U7584 ( .A1(n13184), .A2(n9229), .ZN(n9380) );
  OR2_X2 U7585 ( .A1(n13644), .A2(n13645), .ZN(n8239) );
  NAND2_X2 U7586 ( .A1(n9720), .A2(n9719), .ZN(n14546) );
  OAI21_X1 U7587 ( .B1(n11509), .B2(n11489), .A(n11620), .ZN(n11491) );
  NAND2_X2 U7588 ( .A1(n8573), .A2(n8572), .ZN(n11509) );
  NAND2_X2 U7589 ( .A1(n7988), .A2(n7987), .ZN(n9249) );
  INV_X1 U7590 ( .A(n11404), .ZN(n11752) );
  NOR2_X2 U7591 ( .A1(n8128), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n8341) );
  NOR2_X2 U7592 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n9673) );
  AOI211_X1 U7593 ( .C1(n14649), .C2(n14441), .A(n14692), .B(n14431), .ZN(
        n14648) );
  XNOR2_X2 U7594 ( .A(n9741), .B(n9740), .ZN(n13028) );
  NOR2_X2 U7595 ( .A1(n16202), .A2(n16201), .ZN(n16254) );
  NAND2_X4 U7596 ( .A1(n15613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10245) );
  INV_X1 U7597 ( .A(n10120), .ZN(n9906) );
  OR2_X1 U7598 ( .A1(n9230), .A2(n9229), .ZN(n9390) );
  NAND2_X2 U7599 ( .A1(n9837), .A2(n9838), .ZN(n13175) );
  XNOR2_X2 U7600 ( .A(n15489), .B(n15217), .ZN(n15236) );
  NOR4_X2 U7601 ( .A1(n15667), .A2(n15666), .A3(n15665), .A4(n15664), .ZN(
        n15671) );
  XNOR2_X2 U7602 ( .A(n8549), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8760) );
  NAND2_X2 U7603 ( .A1(n7679), .A2(n7683), .ZN(n8549) );
  INV_X1 U7604 ( .A(n15414), .ZN(n15157) );
  NOR2_X2 U7605 ( .A1(n10174), .A2(n7483), .ZN(n7614) );
  NAND2_X2 U7606 ( .A1(n14770), .A2(n9230), .ZN(n9391) );
  AOI21_X1 U7607 ( .B1(n14285), .B2(n14284), .A(n8318), .ZN(n14343) );
  OAI21_X2 U7608 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n14777), .A(n10793), 
        .ZN(n10799) );
  OAI22_X2 U7609 ( .A1(n14519), .A2(n9895), .B1(n14679), .B2(n14537), .ZN(
        n14503) );
  OAI21_X2 U7610 ( .B1(n14536), .B2(n9894), .A(n9893), .ZN(n14519) );
  OR2_X2 U7611 ( .A1(n13874), .A2(n13316), .ZN(n13596) );
  OAI22_X1 U7612 ( .A1(n14360), .A2(n14359), .B1(n14264), .B2(n16491), .ZN(
        n8320) );
  XNOR2_X2 U7613 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8569) );
  NAND2_X2 U7614 ( .A1(n10785), .A2(n13103), .ZN(n11040) );
  AND2_X2 U7615 ( .A1(n8705), .A2(n8512), .ZN(n8725) );
  NOR2_X2 U7616 ( .A1(n8619), .A2(n8511), .ZN(n8705) );
  NOR2_X2 U7617 ( .A1(n11947), .A2(n11946), .ZN(n12232) );
  NAND2_X2 U7618 ( .A1(n10623), .A2(n10622), .ZN(n15509) );
  XNOR2_X2 U7619 ( .A(n9037), .B(n9036), .ZN(n9048) );
  XNOR2_X2 U7620 ( .A(n9799), .B(n9798), .ZN(n14772) );
  MUX2_X1 U7621 ( .A(n15319), .B(n15528), .S(n10650), .Z(n10591) );
  NAND2_X2 U7622 ( .A1(n10588), .A2(n10587), .ZN(n15528) );
  INV_X1 U7623 ( .A(n10691), .ZN(n10331) );
  NAND2_X2 U7624 ( .A1(n9680), .A2(n9679), .ZN(n14704) );
  NOR2_X2 U7625 ( .A1(n13179), .A2(n12430), .ZN(n11792) );
  NOR2_X1 U7626 ( .A1(n11154), .A2(n11155), .ZN(n11156) );
  NAND2_X1 U7627 ( .A1(n10842), .A2(n10135), .ZN(n9416) );
  NAND2_X2 U7628 ( .A1(n10786), .A2(n15622), .ZN(n10892) );
  CLKBUF_X3 U7629 ( .A(n8655), .Z(n8954) );
  NAND2_X2 U7630 ( .A1(n9661), .A2(n9660), .ZN(n14709) );
  NOR2_X2 U7631 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n16268), .ZN(n9128) );
  OAI222_X1 U7632 ( .A1(n15616), .A2(P1_U3086), .B1(n15627), .B2(n15618), .C1(
        n15617), .C2(n7555), .ZN(P1_U3325) );
  XNOR2_X2 U7633 ( .A(n10245), .B(n10252), .ZN(n15616) );
  OAI21_X2 U7634 ( .B1(n9796), .B2(n14457), .A(n9900), .ZN(n14438) );
  AND2_X2 U7635 ( .A1(n9385), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8582) );
  NAND2_X2 U7636 ( .A1(n10413), .A2(n10412), .ZN(n12496) );
  XNOR2_X2 U7637 ( .A(n9228), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9229) );
  NAND2_X2 U7638 ( .A1(n9349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9228) );
  NOR2_X2 U7639 ( .A1(n12239), .A2(n8672), .ZN(n12370) );
  NAND2_X2 U7640 ( .A1(n11033), .A2(n12597), .ZN(n11053) );
  OR2_X4 U7641 ( .A1(n11058), .A2(n11033), .ZN(n16428) );
  XNOR2_X2 U7642 ( .A(n10263), .B(P1_IR_REG_21__SCAN_IN), .ZN(n11033) );
  XNOR2_X2 U7643 ( .A(n10233), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10257) );
  XNOR2_X2 U7644 ( .A(n9226), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9230) );
  NAND2_X2 U7645 ( .A1(n14765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9226) );
  NAND2_X2 U7646 ( .A1(n8551), .A2(n8550), .ZN(n8781) );
  NOR2_X4 U7647 ( .A1(n7689), .A2(n7466), .ZN(n13902) );
  AND2_X2 U7648 ( .A1(n13938), .A2(n7920), .ZN(n7466) );
  OAI222_X1 U7649 ( .A1(P3_U3151), .A2(n13183), .B1(n14237), .B2(n15637), .C1(
        n13194), .C2(n13182), .ZN(P3_U3267) );
  AND2_X2 U7650 ( .A1(n16477), .A2(n13465), .ZN(n13637) );
  NAND2_X1 U7651 ( .A1(n15495), .A2(n15243), .ZN(n15238) );
  NAND2_X2 U7652 ( .A1(n10649), .A2(n10648), .ZN(n15495) );
  OAI22_X2 U7653 ( .A1(n10984), .A2(P3_D_REG_0__SCAN_IN), .B1(n9059), .B2(
        n14239), .ZN(n13179) );
  NAND2_X2 U7654 ( .A1(n9050), .A2(n9059), .ZN(n10984) );
  AOI21_X2 U7655 ( .B1(n13610), .B2(n13609), .A(n13608), .ZN(n13615) );
  XNOR2_X2 U7656 ( .A(n10791), .B(n8953), .ZN(n13281) );
  NOR2_X2 U7657 ( .A1(n16271), .A2(n16270), .ZN(n16269) );
  NAND2_X2 U7658 ( .A1(n7967), .A2(n7965), .ZN(n16271) );
  OAI21_X2 U7659 ( .B1(n8657), .B2(n8539), .A(n8540), .ZN(n8679) );
  NAND2_X2 U7660 ( .A1(n8538), .A2(n8537), .ZN(n8657) );
  OAI22_X2 U7661 ( .A1(n8304), .A2(n8300), .B1(n11414), .B2(n8301), .ZN(n11419) );
  NAND2_X2 U7662 ( .A1(n7736), .A2(n7734), .ZN(n10791) );
  AND2_X1 U7663 ( .A1(n11160), .A2(n13175), .ZN(n7435) );
  AND2_X1 U7664 ( .A1(n11160), .A2(n13175), .ZN(n14734) );
  XNOR2_X2 U7665 ( .A(n8557), .B(n13174), .ZN(n8880) );
  NAND2_X2 U7666 ( .A1(n8187), .A2(n8185), .ZN(n8557) );
  AND3_X1 U7667 ( .A1(n8464), .A2(n8463), .A3(n8465), .ZN(n10103) );
  OAI22_X1 U7668 ( .A1(n10639), .A2(n8408), .B1(n10640), .B2(n8407), .ZN(
        n10653) );
  XNOR2_X1 U7669 ( .A(n14264), .B(n16491), .ZN(n14360) );
  NAND2_X1 U7670 ( .A1(n9336), .A2(n9335), .ZN(n9356) );
  INV_X2 U7671 ( .A(n15329), .ZN(n15522) );
  NAND2_X1 U7672 ( .A1(n13425), .A2(n13424), .ZN(n13423) );
  OAI22_X1 U7673 ( .A1(n11967), .A2(n11966), .B1(n11965), .B2(n11964), .ZN(
        n12189) );
  NAND2_X1 U7674 ( .A1(n9458), .A2(n9457), .ZN(n11979) );
  NAND2_X1 U7675 ( .A1(n11783), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11953) );
  INV_X1 U7676 ( .A(n11715), .ZN(n11696) );
  INV_X1 U7677 ( .A(n14407), .ZN(n11841) );
  NAND2_X1 U7679 ( .A1(n12210), .A2(n12146), .ZN(n13505) );
  INV_X4 U7680 ( .A(n10153), .ZN(n10176) );
  INV_X2 U7681 ( .A(n10314), .ZN(n11436) );
  INV_X1 U7682 ( .A(n14409), .ZN(n7698) );
  INV_X1 U7683 ( .A(n11249), .ZN(n11995) );
  CLKBUF_X2 U7684 ( .A(n13265), .Z(n7663) );
  INV_X4 U7685 ( .A(n13598), .ZN(n13605) );
  INV_X1 U7686 ( .A(n13665), .ZN(n12210) );
  CLKBUF_X1 U7688 ( .A(n9956), .Z(n9930) );
  INV_X1 U7689 ( .A(n12432), .ZN(n12146) );
  INV_X2 U7690 ( .A(n9956), .ZN(n10148) );
  NAND2_X1 U7691 ( .A1(n7435), .A2(n14508), .ZN(n14265) );
  NAND4_X2 U7692 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n15058) );
  OR2_X1 U7693 ( .A1(n9391), .A2(n11090), .ZN(n9371) );
  CLKBUF_X1 U7694 ( .A(n8633), .Z(n8800) );
  XNOR2_X1 U7695 ( .A(n9398), .B(n9397), .ZN(n10840) );
  INV_X1 U7696 ( .A(n10690), .ZN(n10568) );
  INV_X1 U7697 ( .A(n8523), .ZN(n8526) );
  NOR2_X1 U7698 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n9210) );
  OR2_X1 U7699 ( .A1(n10700), .A2(n10699), .ZN(n10771) );
  OAI21_X1 U7700 ( .B1(n8454), .B2(n8453), .A(n8455), .ZN(n10063) );
  OAI22_X1 U7701 ( .A1(n14304), .A2(n14303), .B1(n14302), .B2(n14301), .ZN(
        n14309) );
  NAND2_X1 U7702 ( .A1(n14981), .A2(n8256), .ZN(n14954) );
  OAI21_X1 U7703 ( .B1(n15479), .B2(n16428), .A(n8172), .ZN(n15480) );
  NAND2_X1 U7704 ( .A1(n15260), .A2(n15259), .ZN(n15258) );
  NOR2_X2 U7705 ( .A1(n13882), .A2(n13893), .ZN(n13473) );
  OR2_X1 U7706 ( .A1(n16029), .A2(n16028), .ZN(n16030) );
  XNOR2_X1 U7707 ( .A(n15204), .B(n15477), .ZN(n15479) );
  NAND2_X1 U7708 ( .A1(n9801), .A2(n9800), .ZN(n14649) );
  NAND2_X1 U7709 ( .A1(n8175), .A2(n8174), .ZN(n15276) );
  NAND2_X1 U7710 ( .A1(n15002), .A2(n15001), .ZN(n15000) );
  AOI211_X1 U7711 ( .C1(n13813), .C2(n7977), .A(n13799), .B(n13798), .ZN(
        n13800) );
  NAND2_X1 U7712 ( .A1(n8939), .A2(n7718), .ZN(n8951) );
  NAND2_X1 U7713 ( .A1(n8166), .A2(n8165), .ZN(n14540) );
  CLKBUF_X1 U7714 ( .A(n14606), .Z(n7641) );
  NAND2_X1 U7715 ( .A1(n9770), .A2(n9769), .ZN(n14671) );
  NAND2_X1 U7716 ( .A1(n9011), .A2(n9010), .ZN(n13946) );
  XNOR2_X1 U7717 ( .A(n16031), .B(n7678), .ZN(n7677) );
  XNOR2_X1 U7718 ( .A(n9174), .B(n9176), .ZN(n16031) );
  OR3_X1 U7719 ( .A1(n15782), .A2(n15781), .A3(n15780), .ZN(n15786) );
  OAI21_X1 U7720 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n16239), .A(n9173), .ZN(
        n9174) );
  CLKBUF_X1 U7721 ( .A(n13069), .Z(n7646) );
  NAND2_X1 U7722 ( .A1(n8246), .A2(n8244), .ZN(n8917) );
  NAND2_X1 U7723 ( .A1(n9709), .A2(n9708), .ZN(n14690) );
  NAND2_X1 U7724 ( .A1(n10576), .A2(n10575), .ZN(n15533) );
  NAND2_X1 U7725 ( .A1(n12740), .A2(n9879), .ZN(n12785) );
  NAND2_X1 U7726 ( .A1(n13404), .A2(n13403), .ZN(n13402) );
  NAND2_X1 U7727 ( .A1(n12945), .A2(n12944), .ZN(n12946) );
  NOR2_X1 U7728 ( .A1(n12705), .A2(n12706), .ZN(n12847) );
  NAND2_X1 U7729 ( .A1(n8190), .A2(n8188), .ZN(n8864) );
  OR2_X1 U7730 ( .A1(n12291), .A2(n12290), .ZN(n12293) );
  NAND2_X1 U7731 ( .A1(n8556), .A2(n8555), .ZN(n8846) );
  NAND2_X1 U7732 ( .A1(n10486), .A2(n10485), .ZN(n15579) );
  NAND2_X1 U7733 ( .A1(n7592), .A2(n10193), .ZN(n11844) );
  NAND2_X1 U7734 ( .A1(n8554), .A2(n8553), .ZN(n8827) );
  NAND2_X1 U7735 ( .A1(n10472), .A2(n10471), .ZN(n12967) );
  NAND2_X1 U7736 ( .A1(n7756), .A2(n7754), .ZN(n9609) );
  NAND2_X1 U7737 ( .A1(n8035), .A2(n9150), .ZN(n9153) );
  NAND2_X1 U7738 ( .A1(n8210), .A2(n8209), .ZN(n8813) );
  NAND2_X1 U7739 ( .A1(n9567), .A2(n9566), .ZN(n16462) );
  NAND2_X1 U7740 ( .A1(n11684), .A2(n8263), .ZN(n14912) );
  NAND2_X1 U7741 ( .A1(n9553), .A2(n8502), .ZN(n9283) );
  AND2_X1 U7742 ( .A1(n14914), .A2(n11683), .ZN(n8263) );
  OR2_X1 U7743 ( .A1(n11552), .A2(n11890), .ZN(n11901) );
  NAND2_X1 U7744 ( .A1(n10349), .A2(n10348), .ZN(n12029) );
  OAI21_X1 U7745 ( .B1(n11131), .B2(n11130), .A(n7617), .ZN(n11142) );
  NAND2_X1 U7746 ( .A1(n9438), .A2(n9437), .ZN(n11517) );
  AND2_X1 U7747 ( .A1(n7962), .A2(n11951), .ZN(n11783) );
  AOI21_X1 U7748 ( .B1(n16212), .B2(n9140), .A(n16209), .ZN(n9141) );
  NAND2_X1 U7749 ( .A1(n9423), .A2(n9424), .ZN(n11404) );
  INV_X1 U7750 ( .A(n14408), .ZN(n7437) );
  NAND3_X1 U7751 ( .A1(n7954), .A2(n7956), .A3(n7953), .ZN(n13484) );
  NAND2_X1 U7752 ( .A1(n8575), .A2(n8576), .ZN(n13202) );
  NOR2_X1 U7753 ( .A1(n9137), .A2(n9138), .ZN(n16207) );
  AND2_X1 U7754 ( .A1(n8574), .A2(n8500), .ZN(n8575) );
  NAND2_X2 U7755 ( .A1(n11199), .A2(n10182), .ZN(n9956) );
  OR2_X1 U7756 ( .A1(n13462), .A2(n10866), .ZN(n8576) );
  NAND2_X1 U7757 ( .A1(n11670), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n13675) );
  AND2_X1 U7758 ( .A1(n7660), .A2(n7623), .ZN(n11160) );
  OAI211_X1 U7759 ( .C1(n10309), .C2(n10840), .A(n10296), .B(n10295), .ZN(
        n11372) );
  NAND2_X2 U7760 ( .A1(n8526), .A2(n8524), .ZN(n8874) );
  AND3_X1 U7761 ( .A1(n8145), .A2(n8144), .A3(n8148), .ZN(n13685) );
  AND2_X1 U7762 ( .A1(n11669), .A2(n13673), .ZN(n11670) );
  XNOR2_X1 U7763 ( .A(n10784), .B(P1_IR_REG_25__SCAN_IN), .ZN(n13103) );
  NAND2_X1 U7764 ( .A1(n10780), .A2(n10783), .ZN(n13033) );
  NAND2_X2 U7765 ( .A1(n11485), .A2(n10838), .ZN(n13462) );
  NAND2_X1 U7766 ( .A1(n11485), .A2(n7434), .ZN(n8655) );
  AND2_X2 U7767 ( .A1(n8523), .A2(n8525), .ZN(n10810) );
  NAND2_X1 U7768 ( .A1(n10783), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10784) );
  NAND2_X2 U7769 ( .A1(n10234), .A2(n15621), .ZN(n10691) );
  XNOR2_X1 U7770 ( .A(n8522), .B(n7959), .ZN(n8525) );
  BUF_X2 U7771 ( .A(n9856), .Z(n10182) );
  CLKBUF_X1 U7772 ( .A(n10892), .Z(n7723) );
  AOI21_X1 U7773 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  AND2_X2 U7774 ( .A1(n9677), .A2(n9834), .ZN(n14444) );
  INV_X2 U7775 ( .A(n15612), .ZN(n15627) );
  NAND2_X2 U7776 ( .A1(n7434), .A2(P3_U3151), .ZN(n14237) );
  OR2_X1 U7777 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  CLKBUF_X1 U7778 ( .A(n10786), .Z(n15073) );
  INV_X1 U7779 ( .A(n10727), .ZN(n12597) );
  AND3_X2 U7780 ( .A1(n10777), .A2(n10277), .A3(n10276), .ZN(n15629) );
  XNOR2_X1 U7781 ( .A(n10279), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15414) );
  OAI21_X1 U7782 ( .B1(n9249), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7624), .ZN(
        n9239) );
  INV_X2 U7783 ( .A(n9351), .ZN(n10831) );
  OR2_X1 U7784 ( .A1(n11498), .A2(n8568), .ZN(n11626) );
  INV_X1 U7785 ( .A(n9249), .ZN(n9351) );
  NAND2_X1 U7786 ( .A1(n8642), .A2(n7787), .ZN(n11780) );
  CLKBUF_X1 U7787 ( .A(n10438), .Z(n10453) );
  NAND2_X1 U7788 ( .A1(n9084), .A2(n8032), .ZN(n9085) );
  AND2_X1 U7789 ( .A1(n9216), .A2(n8321), .ZN(n8247) );
  AND2_X1 U7790 ( .A1(n7807), .A2(n7806), .ZN(n10407) );
  AND2_X1 U7791 ( .A1(n7859), .A2(n7858), .ZN(n10408) );
  NAND4_X1 U7792 ( .A1(n8509), .A2(n8324), .A3(n8323), .A4(n8322), .ZN(n8619)
         );
  INV_X1 U7793 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n16024) );
  NOR2_X1 U7794 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7806) );
  NOR2_X1 U7795 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7807) );
  NOR2_X1 U7796 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n8510) );
  NOR2_X1 U7797 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n9219) );
  INV_X1 U7798 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8660) );
  INV_X1 U7799 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n15793) );
  INV_X1 U7800 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8322) );
  INV_X1 U7801 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9555) );
  INV_X1 U7802 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9556) );
  INV_X4 U7803 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7804 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n10222) );
  NOR2_X1 U7805 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n10223) );
  NOR2_X1 U7806 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n10224) );
  NOR3_X2 U7807 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .ZN(n10228) );
  OAI22_X2 U7808 ( .A1(n10668), .A2(n8410), .B1(n10669), .B2(n8409), .ZN(
        n10681) );
  NOR2_X2 U7809 ( .A1(n13096), .A2(n14719), .ZN(n8170) );
  AOI21_X2 U7811 ( .B1(n13965), .B2(n13962), .A(n8892), .ZN(n13948) );
  XNOR2_X2 U7812 ( .A(n11134), .B(n7438), .ZN(n11294) );
  NOR2_X2 U7813 ( .A1(n15495), .A2(n15276), .ZN(n15261) );
  NOR2_X2 U7814 ( .A1(n9819), .A2(n9818), .ZN(n9835) );
  NOR2_X2 U7815 ( .A1(n16229), .A2(n16228), .ZN(n16227) );
  AOI21_X2 U7816 ( .B1(n16225), .B2(n9158), .A(n16222), .ZN(n16229) );
  NOR2_X2 U7817 ( .A1(n14570), .A2(n14690), .ZN(n8166) );
  OR2_X2 U7818 ( .A1(n14589), .A2(n14700), .ZN(n14570) );
  NOR2_X2 U7819 ( .A1(n15522), .A2(n15336), .ZN(n15325) );
  XNOR2_X1 U7820 ( .A(n9933), .B(n12000), .ZN(n11198) );
  BUF_X2 U7821 ( .A(n9392), .Z(n9802) );
  NOR2_X2 U7822 ( .A1(n11901), .A2(n12029), .ZN(n12039) );
  OAI211_X2 U7823 ( .C1(n7723), .C2(n15098), .A(n10311), .B(n10310), .ZN(
        n10314) );
  OAI211_X1 U7824 ( .C1(n10322), .C2(n8360), .A(n8419), .B(n8418), .ZN(n15461)
         );
  AND2_X1 U7825 ( .A1(n7560), .A2(n11289), .ZN(n7559) );
  AOI21_X1 U7826 ( .B1(n13386), .B2(n13264), .A(n8350), .ZN(n8349) );
  INV_X1 U7827 ( .A(n13359), .ZN(n8350) );
  NAND2_X1 U7828 ( .A1(n14106), .A2(n13612), .ZN(n13639) );
  NAND2_X1 U7829 ( .A1(n12653), .A2(n12654), .ZN(n7846) );
  NAND2_X1 U7830 ( .A1(n8372), .A2(n7482), .ZN(n7811) );
  AOI21_X1 U7831 ( .B1(n7757), .B2(n7447), .A(n7755), .ZN(n7754) );
  INV_X1 U7832 ( .A(n9606), .ZN(n7755) );
  NAND2_X1 U7833 ( .A1(n9272), .A2(n7479), .ZN(n9539) );
  INV_X1 U7834 ( .A(n9536), .ZN(n9277) );
  INV_X1 U7835 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8969) );
  INV_X1 U7836 ( .A(n10118), .ZN(n9905) );
  NAND2_X1 U7837 ( .A1(n9230), .A2(n9229), .ZN(n9392) );
  NAND2_X1 U7838 ( .A1(n7801), .A2(n7796), .ZN(n15284) );
  NOR2_X1 U7839 ( .A1(n15288), .A2(n7797), .ZN(n7796) );
  INV_X1 U7840 ( .A(n7800), .ZN(n7797) );
  INV_X1 U7841 ( .A(n15211), .ZN(n15477) );
  XOR2_X1 U7842 ( .A(n15216), .B(n15477), .Z(n15203) );
  NAND2_X1 U7843 ( .A1(n9956), .A2(n7635), .ZN(n9936) );
  INV_X1 U7844 ( .A(n9976), .ZN(n7578) );
  AOI21_X1 U7845 ( .B1(n7868), .B2(n10345), .A(n7867), .ZN(n7866) );
  AND2_X1 U7846 ( .A1(n8383), .A2(n8381), .ZN(n10357) );
  NAND2_X1 U7847 ( .A1(n7899), .A2(n7896), .ZN(n7891) );
  OR2_X1 U7848 ( .A1(n8412), .A2(n7900), .ZN(n7899) );
  AND2_X1 U7849 ( .A1(n8395), .A2(n10458), .ZN(n8394) );
  NAND2_X1 U7850 ( .A1(n8399), .A2(n8397), .ZN(n8395) );
  AND2_X1 U7851 ( .A1(n10548), .A2(n8401), .ZN(n8400) );
  INV_X1 U7852 ( .A(n10044), .ZN(n7638) );
  INV_X1 U7853 ( .A(n10081), .ZN(n7716) );
  INV_X1 U7854 ( .A(n9318), .ZN(n8016) );
  INV_X1 U7855 ( .A(n13600), .ZN(n7659) );
  OR2_X1 U7856 ( .A1(n10281), .A2(n11033), .ZN(n10709) );
  AND2_X1 U7857 ( .A1(n8253), .A2(n13613), .ZN(n13618) );
  INV_X1 U7858 ( .A(n8525), .ZN(n8524) );
  OR2_X1 U7859 ( .A1(n12673), .A2(n16279), .ZN(n7973) );
  NAND2_X1 U7860 ( .A1(n7971), .A2(n16279), .ZN(n7970) );
  NAND2_X1 U7861 ( .A1(n12373), .A2(n7972), .ZN(n7971) );
  OAI21_X1 U7862 ( .B1(n13122), .B2(n7783), .A(n7782), .ZN(n13698) );
  NAND2_X1 U7863 ( .A1(n13124), .A2(n7784), .ZN(n7782) );
  NAND2_X1 U7864 ( .A1(n8151), .A2(n7784), .ZN(n7783) );
  NAND2_X1 U7865 ( .A1(n13701), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7784) );
  AND2_X1 U7866 ( .A1(n13188), .A2(n13860), .ZN(n13608) );
  OR2_X1 U7867 ( .A1(n13887), .A2(n13364), .ZN(n13592) );
  NOR2_X1 U7868 ( .A1(n13923), .A2(n8116), .ZN(n8115) );
  INV_X1 U7869 ( .A(n8118), .ZN(n8116) );
  OR2_X1 U7870 ( .A1(n16417), .A2(n14079), .ZN(n8097) );
  NAND2_X1 U7871 ( .A1(n11794), .A2(n13837), .ZN(n11795) );
  INV_X1 U7872 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8340) );
  NOR2_X1 U7873 ( .A1(n7449), .A2(n8200), .ZN(n8199) );
  INV_X1 U7874 ( .A(n8544), .ZN(n8200) );
  NAND2_X1 U7875 ( .A1(n9204), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9786) );
  INV_X1 U7876 ( .A(n9758), .ZN(n9204) );
  NAND2_X1 U7877 ( .A1(n14608), .A2(n14607), .ZN(n14606) );
  AOI21_X1 U7878 ( .B1(n8060), .B2(n8059), .A(n7507), .ZN(n8058) );
  INV_X1 U7879 ( .A(n7453), .ZN(n8059) );
  INV_X1 U7880 ( .A(n8207), .ZN(n8206) );
  OAI21_X1 U7881 ( .B1(n12736), .B2(n8208), .A(n9589), .ZN(n8207) );
  OAI21_X1 U7882 ( .B1(n12014), .B2(n12021), .A(n12060), .ZN(n9873) );
  AOI21_X1 U7883 ( .B1(n8073), .B2(n8072), .A(n7478), .ZN(n8071) );
  INV_X1 U7884 ( .A(n9878), .ZN(n8072) );
  NOR2_X1 U7885 ( .A1(n15187), .A2(n8443), .ZN(n8442) );
  INV_X1 U7886 ( .A(n12974), .ZN(n8443) );
  NOR2_X1 U7887 ( .A1(n12712), .A2(n12851), .ZN(n8180) );
  NAND2_X1 U7888 ( .A1(n8423), .A2(n8421), .ZN(n12033) );
  NOR2_X1 U7889 ( .A1(n7867), .A2(n8422), .ZN(n8421) );
  INV_X1 U7890 ( .A(n11892), .ZN(n8422) );
  AND2_X1 U7891 ( .A1(n10262), .A2(n16023), .ZN(n7888) );
  NAND2_X1 U7892 ( .A1(n8367), .A2(n8365), .ZN(n9644) );
  NOR2_X1 U7893 ( .A1(n9641), .A2(n8366), .ZN(n8365) );
  INV_X1 U7894 ( .A(n9297), .ZN(n8366) );
  XNOR2_X1 U7895 ( .A(n9295), .B(SI_16_), .ZN(n9629) );
  INV_X1 U7896 ( .A(n7758), .ZN(n7757) );
  OAI21_X1 U7897 ( .B1(n7761), .B2(n7447), .A(n9290), .ZN(n7758) );
  AOI21_X1 U7898 ( .B1(n7993), .B2(n7995), .A(n7499), .ZN(n7991) );
  AOI21_X1 U7899 ( .B1(n9093), .B2(n9121), .A(n9092), .ZN(n9119) );
  INV_X1 U7900 ( .A(n8347), .ZN(n8346) );
  OAI21_X1 U7901 ( .B1(n8349), .B2(n8348), .A(n13434), .ZN(n8347) );
  INV_X1 U7902 ( .A(n10810), .ZN(n8986) );
  AND2_X1 U7903 ( .A1(n8526), .A2(n8525), .ZN(n8611) );
  AOI21_X1 U7904 ( .B1(n7839), .B2(n7837), .A(n7836), .ZN(n7835) );
  INV_X1 U7905 ( .A(n7839), .ZN(n7838) );
  INV_X1 U7906 ( .A(n16274), .ZN(n7836) );
  NOR2_X1 U7907 ( .A1(n13802), .A2(n7661), .ZN(n13828) );
  AND2_X1 U7908 ( .A1(n13803), .A2(n13804), .ZN(n7661) );
  NAND2_X1 U7909 ( .A1(n13828), .A2(n13827), .ZN(n7827) );
  NOR2_X1 U7910 ( .A1(n7440), .A2(n13249), .ZN(n8119) );
  INV_X1 U7911 ( .A(n13462), .ZN(n13458) );
  INV_X1 U7912 ( .A(n14092), .ZN(n16311) );
  OR2_X1 U7913 ( .A1(n11802), .A2(n13598), .ZN(n14092) );
  AND2_X1 U7914 ( .A1(n8343), .A2(n8564), .ZN(n8342) );
  INV_X1 U7915 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U7916 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8607) );
  AOI21_X1 U7917 ( .B1(n12222), .B2(n12218), .A(n12403), .ZN(n8295) );
  NOR2_X1 U7918 ( .A1(n8296), .A2(n8294), .ZN(n8293) );
  AND2_X1 U7919 ( .A1(n14411), .A2(n14265), .ZN(n11151) );
  INV_X1 U7920 ( .A(n8305), .ZN(n8298) );
  AND2_X1 U7921 ( .A1(n14658), .A2(n14388), .ZN(n7647) );
  XNOR2_X1 U7922 ( .A(n14686), .B(n14321), .ZN(n14545) );
  NAND2_X1 U7923 ( .A1(n12319), .A2(n9552), .ZN(n12735) );
  OAI21_X1 U7924 ( .B1(n11472), .B2(n9870), .A(n9869), .ZN(n8041) );
  OR2_X1 U7925 ( .A1(n11517), .A2(n11841), .ZN(n9869) );
  AND2_X1 U7926 ( .A1(n11071), .A2(n11162), .ZN(n14600) );
  NAND2_X1 U7927 ( .A1(n9615), .A2(n9614), .ZN(n14728) );
  OR2_X1 U7928 ( .A1(n9832), .A2(n14781), .ZN(n9852) );
  NAND2_X1 U7929 ( .A1(n14892), .A2(n14893), .ZN(n14891) );
  XNOR2_X1 U7930 ( .A(n8254), .B(n12183), .ZN(n11136) );
  NAND2_X1 U7931 ( .A1(n11135), .A2(n8255), .ZN(n8254) );
  NAND2_X1 U7932 ( .A1(n11134), .A2(n11694), .ZN(n8255) );
  INV_X1 U7933 ( .A(n15370), .ZN(n15411) );
  INV_X1 U7934 ( .A(n12502), .ZN(n8269) );
  INV_X1 U7935 ( .A(n15046), .ZN(n15243) );
  NAND2_X1 U7936 ( .A1(n15517), .A2(n15320), .ZN(n7800) );
  NAND2_X1 U7937 ( .A1(n15329), .A2(n15197), .ZN(n7802) );
  NAND2_X1 U7938 ( .A1(n15423), .A2(n15424), .ZN(n8478) );
  AND2_X2 U7939 ( .A1(n12286), .A2(n12560), .ZN(n12611) );
  NAND2_X1 U7940 ( .A1(n11545), .A2(n11544), .ZN(n8426) );
  OR2_X1 U7941 ( .A1(n7771), .A2(n15236), .ZN(n7769) );
  INV_X1 U7942 ( .A(n15483), .ZN(n15227) );
  NAND2_X1 U7943 ( .A1(n8372), .A2(n8370), .ZN(n15235) );
  XNOR2_X1 U7944 ( .A(n7818), .B(n10239), .ZN(n10786) );
  OAI21_X1 U7945 ( .B1(n10240), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7818) );
  INV_X1 U7946 ( .A(n9249), .ZN(n10838) );
  NAND2_X1 U7947 ( .A1(n15793), .A2(n10293), .ZN(n10409) );
  AOI21_X1 U7948 ( .B1(n7686), .B2(n7687), .A(n7685), .ZN(n13471) );
  AND2_X1 U7949 ( .A1(n13470), .A2(n16480), .ZN(n7685) );
  OR2_X1 U7950 ( .A1(n12893), .A2(n12892), .ZN(n7853) );
  NAND2_X1 U7951 ( .A1(n9366), .A2(n9365), .ZN(n14475) );
  NAND2_X1 U7952 ( .A1(n11749), .A2(n16455), .ZN(n16458) );
  INV_X1 U7953 ( .A(n14941), .ZN(n15216) );
  NAND2_X1 U7954 ( .A1(n7774), .A2(n15568), .ZN(n7773) );
  NOR2_X1 U7955 ( .A1(n7468), .A2(n8173), .ZN(n8172) );
  INV_X1 U7956 ( .A(n15478), .ZN(n8173) );
  INV_X1 U7957 ( .A(keyinput_131), .ZN(n7606) );
  INV_X1 U7958 ( .A(n9972), .ZN(n7727) );
  INV_X1 U7959 ( .A(n9978), .ZN(n7570) );
  INV_X1 U7960 ( .A(n9982), .ZN(n7673) );
  INV_X1 U7961 ( .A(n9986), .ZN(n7580) );
  INV_X1 U7962 ( .A(n9988), .ZN(n7568) );
  AND2_X1 U7963 ( .A1(n10312), .A2(n10330), .ZN(n7560) );
  INV_X1 U7964 ( .A(n9992), .ZN(n7571) );
  NAND2_X1 U7965 ( .A1(n8470), .A2(n8471), .ZN(n8469) );
  INV_X1 U7966 ( .A(n10004), .ZN(n8470) );
  NOR2_X1 U7967 ( .A1(n10378), .A2(n10375), .ZN(n8405) );
  MUX2_X1 U7968 ( .A(n15052), .B(n12496), .S(n10358), .Z(n10415) );
  NAND2_X1 U7969 ( .A1(n10442), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U7970 ( .A1(n10473), .A2(n7911), .ZN(n7910) );
  INV_X1 U7971 ( .A(n8397), .ZN(n7558) );
  NOR2_X1 U7972 ( .A1(n7896), .A2(n7894), .ZN(n7893) );
  AND2_X1 U7973 ( .A1(n7892), .A2(n7891), .ZN(n7890) );
  AND2_X1 U7974 ( .A1(n10397), .A2(n10396), .ZN(n7889) );
  NOR2_X1 U7975 ( .A1(n8398), .A2(n10442), .ZN(n8399) );
  INV_X1 U7976 ( .A(n10028), .ZN(n7746) );
  NAND2_X1 U7977 ( .A1(n10518), .A2(n7875), .ZN(n7874) );
  NOR2_X1 U7978 ( .A1(n10532), .A2(n10529), .ZN(n8404) );
  NAND2_X1 U7979 ( .A1(n10529), .A2(n10532), .ZN(n8403) );
  NOR2_X1 U7980 ( .A1(n10503), .A2(n10506), .ZN(n8415) );
  INV_X1 U7981 ( .A(n10503), .ZN(n8414) );
  INV_X1 U7982 ( .A(n10035), .ZN(n7644) );
  INV_X1 U7983 ( .A(n10036), .ZN(n7645) );
  INV_X1 U7984 ( .A(n10041), .ZN(n7749) );
  NOR2_X1 U7985 ( .A1(n7873), .A2(n8404), .ZN(n7872) );
  INV_X1 U7986 ( .A(n7874), .ZN(n7873) );
  INV_X1 U7987 ( .A(n8403), .ZN(n7870) );
  AND2_X1 U7988 ( .A1(n10520), .A2(n7877), .ZN(n7876) );
  INV_X1 U7989 ( .A(n10518), .ZN(n7877) );
  NAND2_X1 U7990 ( .A1(n10577), .A2(n7884), .ZN(n7883) );
  NOR2_X1 U7991 ( .A1(n8387), .A2(n10589), .ZN(n8388) );
  NAND2_X1 U7992 ( .A1(n8387), .A2(n10589), .ZN(n8386) );
  NOR2_X1 U7993 ( .A1(n10566), .A2(n10563), .ZN(n8417) );
  INV_X1 U7994 ( .A(n10563), .ZN(n8416) );
  INV_X1 U7995 ( .A(n10050), .ZN(n7656) );
  NAND2_X1 U7996 ( .A1(n7612), .A2(n7611), .ZN(n7610) );
  NAND2_X1 U7997 ( .A1(n7639), .A2(n7638), .ZN(n7613) );
  INV_X1 U7998 ( .A(n10045), .ZN(n7611) );
  NAND2_X1 U7999 ( .A1(n10055), .A2(n8457), .ZN(n8456) );
  INV_X1 U8000 ( .A(n7538), .ZN(n8457) );
  NOR2_X1 U8001 ( .A1(n8388), .A2(n7882), .ZN(n7881) );
  INV_X1 U8002 ( .A(n7883), .ZN(n7882) );
  INV_X1 U8003 ( .A(n8386), .ZN(n7879) );
  AND2_X1 U8004 ( .A1(n10579), .A2(n7886), .ZN(n7885) );
  INV_X1 U8005 ( .A(n10577), .ZN(n7886) );
  AOI21_X1 U8006 ( .B1(n8392), .B2(n8393), .A(n8390), .ZN(n8389) );
  NAND2_X1 U8007 ( .A1(n7643), .A2(n7642), .ZN(n10627) );
  NOR2_X1 U8008 ( .A1(n7860), .A2(n10626), .ZN(n7642) );
  INV_X1 U8009 ( .A(n8392), .ZN(n7860) );
  NAND2_X1 U8010 ( .A1(n7502), .A2(n10078), .ZN(n8462) );
  NOR2_X1 U8011 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8129) );
  NOR2_X1 U8012 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8130) );
  INV_X1 U8013 ( .A(n10667), .ZN(n8409) );
  NOR2_X1 U8014 ( .A1(n10670), .A2(n10667), .ZN(n8410) );
  INV_X1 U8015 ( .A(n8015), .ZN(n8014) );
  OAI21_X1 U8016 ( .B1(n9316), .B2(n8016), .A(n9320), .ZN(n8015) );
  INV_X1 U8017 ( .A(n12675), .ZN(n7984) );
  NAND2_X1 U8018 ( .A1(n7776), .A2(n13739), .ZN(n13740) );
  INV_X1 U8019 ( .A(n8196), .ZN(n8195) );
  OAI21_X1 U8020 ( .B1(n14545), .B2(n8197), .A(n10205), .ZN(n8196) );
  INV_X1 U8021 ( .A(n9735), .ZN(n8197) );
  OR2_X1 U8022 ( .A1(n15629), .A2(n15414), .ZN(n10280) );
  NAND2_X1 U8023 ( .A1(n9299), .A2(n15657), .ZN(n9302) );
  OAI21_X1 U8024 ( .B1(n9259), .B2(n8358), .A(n9262), .ZN(n8357) );
  INV_X1 U8025 ( .A(n9261), .ZN(n8358) );
  OAI21_X1 U8026 ( .B1(n10831), .B2(n8010), .A(n8009), .ZN(n8008) );
  NAND2_X1 U8027 ( .A1(n10831), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U8028 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n8033), .ZN(n8032) );
  INV_X1 U8029 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8033) );
  AND2_X1 U8030 ( .A1(n13411), .A2(n13256), .ZN(n13259) );
  NAND2_X1 U8031 ( .A1(n13251), .A2(n13250), .ZN(n13254) );
  AOI21_X1 U8032 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n11780), .A(n13685), .ZN(
        n11777) );
  INV_X1 U8033 ( .A(n12673), .ZN(n7972) );
  NOR2_X1 U8034 ( .A1(n13740), .A2(n13773), .ZN(n13741) );
  NOR2_X1 U8035 ( .A1(n14175), .A2(n13364), .ZN(n8087) );
  OR2_X1 U8036 ( .A1(n13878), .A2(n8950), .ZN(n8088) );
  OAI22_X1 U8037 ( .A1(n8936), .A2(n8111), .B1(n13895), .B2(n14182), .ZN(n8110) );
  INV_X1 U8038 ( .A(n8115), .ZN(n8112) );
  NOR2_X1 U8039 ( .A1(n8808), .A2(n7931), .ZN(n7930) );
  INV_X1 U8040 ( .A(n13555), .ZN(n7931) );
  AND2_X1 U8041 ( .A1(n13561), .A2(n13560), .ZN(n13558) );
  AND2_X1 U8042 ( .A1(n12303), .A2(n8624), .ZN(n8626) );
  AND2_X1 U8043 ( .A1(n13499), .A2(n8626), .ZN(n8627) );
  NAND2_X1 U8044 ( .A1(n12331), .A2(n12476), .ZN(n13507) );
  AND2_X1 U8045 ( .A1(n13342), .A2(n13937), .ZN(n13577) );
  AND2_X1 U8046 ( .A1(n13991), .A2(n8841), .ZN(n8106) );
  OR2_X1 U8047 ( .A1(n14135), .A2(n13426), .ZN(n8497) );
  INV_X1 U8048 ( .A(n8861), .ZN(n8105) );
  NOR2_X1 U8049 ( .A1(n8746), .A2(n8099), .ZN(n8098) );
  INV_X1 U8050 ( .A(n8731), .ZN(n8099) );
  AND2_X1 U8051 ( .A1(n13630), .A2(n8684), .ZN(n8124) );
  NAND2_X1 U8052 ( .A1(n13507), .A2(n13506), .ZN(n13624) );
  OR2_X1 U8053 ( .A1(n8977), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U8054 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n8186), .ZN(n8185) );
  INV_X1 U8055 ( .A(n8213), .ZN(n8212) );
  OAI21_X1 U8056 ( .B1(n8780), .B2(n8214), .A(n8794), .ZN(n8213) );
  INV_X1 U8057 ( .A(n8552), .ZN(n8214) );
  INV_X1 U8058 ( .A(n8203), .ZN(n8202) );
  OAI21_X1 U8059 ( .B1(n8708), .B2(n7449), .A(n8722), .ZN(n8203) );
  INV_X1 U8060 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8543) );
  INV_X1 U8061 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8324) );
  INV_X1 U8062 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U8063 ( .A1(n9198), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9617) );
  INV_X1 U8064 ( .A(n9597), .ZN(n9198) );
  NAND2_X1 U8065 ( .A1(n7637), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9382) );
  AND2_X1 U8066 ( .A1(n14658), .A2(n14475), .ZN(n8238) );
  NOR2_X1 U8067 ( .A1(n14481), .A2(n8049), .ZN(n8048) );
  INV_X1 U8068 ( .A(n14487), .ZN(n8049) );
  NOR2_X1 U8069 ( .A1(n10202), .A2(n8224), .ZN(n8223) );
  INV_X1 U8070 ( .A(n9668), .ZN(n8224) );
  INV_X1 U8071 ( .A(n9640), .ZN(n8252) );
  INV_X1 U8072 ( .A(n9884), .ZN(n8061) );
  INV_X1 U8073 ( .A(n9575), .ZN(n8208) );
  NAND2_X1 U8074 ( .A1(n7599), .A2(n7598), .ZN(n12107) );
  INV_X1 U8075 ( .A(n12108), .ZN(n7599) );
  NAND2_X1 U8076 ( .A1(n11842), .A2(n9448), .ZN(n8231) );
  AND2_X1 U8077 ( .A1(n7462), .A2(n14467), .ZN(n8236) );
  AND2_X1 U8078 ( .A1(n14444), .A2(n7725), .ZN(n9938) );
  AND2_X1 U8079 ( .A1(n9216), .A2(n8249), .ZN(n8248) );
  INV_X1 U8080 ( .A(n9224), .ZN(n7730) );
  AND2_X1 U8081 ( .A1(n8321), .A2(n9342), .ZN(n8249) );
  OR2_X1 U8082 ( .A1(n9505), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U8083 ( .A1(n7509), .A2(n14826), .ZN(n8273) );
  INV_X1 U8084 ( .A(n15033), .ZN(n8278) );
  OR2_X1 U8085 ( .A1(n14972), .A2(n14816), .ZN(n8275) );
  NOR2_X1 U8086 ( .A1(n8273), .A2(n8276), .ZN(n8272) );
  NOR2_X1 U8087 ( .A1(n14964), .A2(n14818), .ZN(n8276) );
  NAND2_X1 U8088 ( .A1(n10710), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10237) );
  NOR2_X1 U8089 ( .A1(n15236), .A2(n7603), .ZN(n7602) );
  INV_X1 U8090 ( .A(n15238), .ZN(n7603) );
  NOR2_X1 U8091 ( .A1(n15274), .A2(n8376), .ZN(n8375) );
  INV_X1 U8092 ( .A(n8379), .ZN(n8376) );
  AND2_X1 U8093 ( .A1(n8180), .A2(n8179), .ZN(n8178) );
  INV_X1 U8094 ( .A(n12451), .ZN(n8446) );
  OR2_X1 U8095 ( .A1(n8447), .A2(n8446), .ZN(n8445) );
  AND2_X1 U8096 ( .A1(n12090), .A2(n10731), .ZN(n12031) );
  NAND2_X1 U8097 ( .A1(n11887), .A2(n7470), .ZN(n8483) );
  NAND2_X1 U8098 ( .A1(n12026), .A2(n12028), .ZN(n8484) );
  NAND2_X1 U8099 ( .A1(n8426), .A2(n8424), .ZN(n8423) );
  NOR2_X1 U8100 ( .A1(n11893), .A2(n8425), .ZN(n8424) );
  INV_X1 U8101 ( .A(n11546), .ZN(n8425) );
  XNOR2_X1 U8102 ( .A(n15449), .B(n11372), .ZN(n11297) );
  NAND2_X1 U8103 ( .A1(n7626), .A2(n7625), .ZN(n10778) );
  XNOR2_X1 U8104 ( .A(n9325), .B(SI_24_), .ZN(n9753) );
  XNOR2_X1 U8105 ( .A(n9304), .B(SI_18_), .ZN(n9303) );
  NAND2_X1 U8106 ( .A1(n9609), .A2(n8368), .ZN(n8367) );
  NOR2_X1 U8107 ( .A1(n9298), .A2(n8369), .ZN(n8368) );
  INV_X1 U8108 ( .A(n9629), .ZN(n9298) );
  INV_X1 U8109 ( .A(n9294), .ZN(n8369) );
  NAND2_X1 U8110 ( .A1(n7664), .A2(n9258), .ZN(n9449) );
  XNOR2_X1 U8111 ( .A(n9260), .B(n7764), .ZN(n9259) );
  INV_X1 U8112 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n9091) );
  AOI22_X1 U8113 ( .A1(n9119), .A2(n9095), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n9094), .ZN(n9096) );
  INV_X1 U8114 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n9094) );
  OAI21_X1 U8115 ( .B1(n9099), .B2(n9118), .A(n9116), .ZN(n9151) );
  NAND2_X1 U8116 ( .A1(n12866), .A2(n12865), .ZN(n13327) );
  NAND2_X2 U8117 ( .A1(n11797), .A2(n8503), .ZN(n13265) );
  NOR2_X1 U8118 ( .A1(n7481), .A2(n8337), .ZN(n8336) );
  AND2_X1 U8119 ( .A1(n13284), .A2(n8338), .ZN(n8337) );
  INV_X1 U8120 ( .A(n13224), .ZN(n8338) );
  NAND2_X1 U8121 ( .A1(n13327), .A2(n13326), .ZN(n13325) );
  NAND2_X1 U8122 ( .A1(n8330), .A2(n13256), .ZN(n13411) );
  AND2_X1 U8123 ( .A1(n8331), .A2(n13951), .ZN(n8330) );
  INV_X1 U8124 ( .A(SI_22_), .ZN(n9721) );
  INV_X1 U8125 ( .A(n13663), .ZN(n12580) );
  NAND2_X1 U8126 ( .A1(n8351), .A2(n8349), .ZN(n13357) );
  NAND2_X1 U8127 ( .A1(n7508), .A2(n13293), .ZN(n8351) );
  INV_X1 U8128 ( .A(n8598), .ZN(n13200) );
  NAND2_X1 U8129 ( .A1(n8523), .A2(n8524), .ZN(n8633) );
  XNOR2_X1 U8130 ( .A(n11664), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n11623) );
  OR2_X1 U8131 ( .A1(n11660), .A2(n11667), .ZN(n8148) );
  NAND2_X1 U8132 ( .A1(n7961), .A2(n13672), .ZN(n13677) );
  NAND2_X1 U8133 ( .A1(n13675), .A2(n13673), .ZN(n7961) );
  AND3_X1 U8134 ( .A1(n7780), .A2(n7778), .A3(P3_REG2_REG_7__SCAN_IN), .ZN(
        n12359) );
  NOR2_X1 U8135 ( .A1(n7848), .A2(n7842), .ZN(n7841) );
  INV_X1 U8136 ( .A(n7846), .ZN(n7842) );
  NAND2_X1 U8137 ( .A1(n7840), .A2(n7846), .ZN(n7839) );
  INV_X1 U8138 ( .A(n7843), .ZN(n7840) );
  INV_X1 U8139 ( .A(n12655), .ZN(n7844) );
  INV_X1 U8140 ( .A(n7973), .ZN(n7966) );
  NOR2_X1 U8141 ( .A1(n12904), .A2(n8150), .ZN(n13122) );
  NOR2_X1 U8142 ( .A1(n7448), .A2(n14068), .ZN(n8154) );
  OR2_X1 U8143 ( .A1(n13725), .A2(n13726), .ZN(n7776) );
  INV_X1 U8144 ( .A(n13774), .ZN(n13752) );
  AOI21_X1 U8145 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13797) );
  NOR2_X1 U8146 ( .A1(n13783), .A2(n7978), .ZN(n13815) );
  NOR2_X1 U8147 ( .A1(n13780), .A2(n14154), .ZN(n7978) );
  NOR2_X1 U8148 ( .A1(n8957), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8981) );
  OR2_X1 U8149 ( .A1(n8943), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8957) );
  OR2_X1 U8150 ( .A1(n8120), .A2(n7440), .ZN(n8118) );
  AND2_X1 U8151 ( .A1(n8916), .A2(n8121), .ZN(n8120) );
  AND2_X1 U8152 ( .A1(n13585), .A2(n13584), .ZN(n13923) );
  NAND2_X1 U8153 ( .A1(n13990), .A2(n8861), .ZN(n13978) );
  NAND2_X1 U8154 ( .A1(n9002), .A2(n13477), .ZN(n14000) );
  OAI21_X1 U8155 ( .B1(n14044), .B2(n8127), .A(n8125), .ZN(n8825) );
  INV_X1 U8156 ( .A(n8126), .ZN(n8125) );
  NOR2_X1 U8157 ( .A1(n9000), .A2(n7934), .ZN(n7933) );
  INV_X1 U8158 ( .A(n13552), .ZN(n7934) );
  INV_X1 U8159 ( .A(n13558), .ZN(n8808) );
  NAND2_X1 U8160 ( .A1(n14044), .A2(n7455), .ZN(n14029) );
  AND2_X1 U8161 ( .A1(n13553), .A2(n13555), .ZN(n14043) );
  NAND2_X1 U8162 ( .A1(n14055), .A2(n13542), .ZN(n8999) );
  AOI21_X1 U8163 ( .B1(n8094), .B2(n8096), .A(n7488), .ZN(n8092) );
  NAND2_X1 U8164 ( .A1(n7537), .A2(n14045), .ZN(n14044) );
  AND4_X1 U8165 ( .A1(n8753), .A2(n8752), .A3(n8751), .A4(n8750), .ZN(n14062)
         );
  AOI21_X1 U8166 ( .B1(n7941), .B2(n13534), .A(n7939), .ZN(n7938) );
  INV_X1 U8167 ( .A(n13532), .ZN(n7939) );
  INV_X1 U8168 ( .A(n13000), .ZN(n7945) );
  NAND2_X1 U8169 ( .A1(n13938), .A2(n9012), .ZN(n13926) );
  INV_X1 U8170 ( .A(n13505), .ZN(n7918) );
  INV_X1 U8171 ( .A(n13495), .ZN(n7919) );
  AND2_X1 U8172 ( .A1(n13505), .A2(n13499), .ZN(n13628) );
  NAND2_X1 U8173 ( .A1(n12153), .A2(n13489), .ZN(n13494) );
  AND3_X1 U8174 ( .A1(n8597), .A2(n8596), .A3(n8595), .ZN(n11801) );
  OAI21_X1 U8175 ( .B1(n10984), .B2(P3_D_REG_1__SCAN_IN), .A(n9056), .ZN(
        n11912) );
  AND2_X1 U8176 ( .A1(n8342), .A2(n8562), .ZN(n7960) );
  NAND2_X1 U8177 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n7735), .ZN(n7734) );
  NAND2_X1 U8178 ( .A1(n9030), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7857) );
  AND2_X1 U8179 ( .A1(n7596), .A2(n7597), .ZN(n8938) );
  INV_X1 U8180 ( .A(n8926), .ZN(n7582) );
  AND2_X2 U8181 ( .A1(n7657), .A2(n8243), .ZN(n8926) );
  NAND2_X1 U8182 ( .A1(n11511), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8243) );
  OR2_X1 U8183 ( .A1(n8917), .A2(n8918), .ZN(n7657) );
  NAND2_X1 U8184 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n12730), .ZN(n7608) );
  NAND2_X1 U8185 ( .A1(n8971), .A2(n8970), .ZN(n8973) );
  INV_X1 U8186 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8970) );
  INV_X1 U8187 ( .A(n8975), .ZN(n8971) );
  XNOR2_X1 U8188 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8826) );
  OR2_X1 U8189 ( .A1(n8783), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U8190 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8722) );
  NAND2_X1 U8191 ( .A1(n8545), .A2(n8544), .ZN(n8710) );
  XNOR2_X1 U8192 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8708) );
  INV_X1 U8193 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8618) );
  AOI21_X1 U8194 ( .B1(n8607), .B2(n8218), .A(n7505), .ZN(n8217) );
  XNOR2_X1 U8195 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8620) );
  AND2_X1 U8196 ( .A1(n7985), .A2(n8323), .ZN(n8592) );
  INV_X1 U8197 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7985) );
  NOR3_X1 U8198 ( .A1(n13035), .A2(n14781), .A3(n13105), .ZN(n10827) );
  NAND2_X1 U8199 ( .A1(n8315), .A2(n8317), .ZN(n8314) );
  NAND2_X1 U8200 ( .A1(n14368), .A2(n8316), .ZN(n8315) );
  INV_X1 U8201 ( .A(n14248), .ZN(n8316) );
  NAND2_X1 U8202 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  NAND2_X1 U8203 ( .A1(n12056), .A2(n12057), .ZN(n12220) );
  NAND2_X1 U8204 ( .A1(n9202), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9710) );
  XNOR2_X1 U8205 ( .A(n14704), .B(n14254), .ZN(n14253) );
  INV_X1 U8206 ( .A(n7452), .ZN(n8310) );
  AOI21_X1 U8207 ( .B1(n12688), .B2(n12684), .A(n12772), .ZN(n8285) );
  NOR2_X1 U8208 ( .A1(n8286), .A2(n8284), .ZN(n8283) );
  OR2_X1 U8209 ( .A1(n9710), .A2(n14319), .ZN(n9727) );
  AND2_X1 U8210 ( .A1(n14261), .A2(n14260), .ZN(n7622) );
  AND2_X1 U8211 ( .A1(n14272), .A2(n14273), .ZN(n7667) );
  NAND2_X1 U8212 ( .A1(n12946), .A2(n12947), .ZN(n13059) );
  OR2_X1 U8213 ( .A1(n8467), .A2(n7460), .ZN(n8465) );
  NOR2_X1 U8214 ( .A1(n10170), .A2(n8459), .ZN(n8458) );
  OR2_X1 U8215 ( .A1(n10173), .A2(n8460), .ZN(n8459) );
  NAND2_X1 U8216 ( .A1(n8003), .A2(n8002), .ZN(n10170) );
  NOR2_X1 U8217 ( .A1(n10171), .A2(n10172), .ZN(n8460) );
  AND2_X1 U8218 ( .A1(n8005), .A2(n8004), .ZN(n10174) );
  INV_X1 U8219 ( .A(n10173), .ZN(n8004) );
  OR2_X1 U8220 ( .A1(n9380), .A2(n7574), .ZN(n9372) );
  OR2_X1 U8221 ( .A1(n9390), .A2(n9368), .ZN(n9369) );
  INV_X1 U8222 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9675) );
  OR2_X1 U8223 ( .A1(n14482), .A2(n7527), .ZN(n8237) );
  OAI21_X1 U8224 ( .B1(n14606), .B2(n7457), .A(n8220), .ZN(n14554) );
  INV_X1 U8225 ( .A(n8221), .ZN(n8220) );
  OAI21_X1 U8226 ( .B1(n8223), .B2(n7457), .A(n8225), .ZN(n8221) );
  OR2_X1 U8227 ( .A1(n14700), .A2(n14584), .ZN(n8225) );
  NOR2_X1 U8228 ( .A1(n14566), .A2(n8069), .ZN(n8068) );
  INV_X1 U8229 ( .A(n9889), .ZN(n8069) );
  NAND2_X1 U8230 ( .A1(n14579), .A2(n10202), .ZN(n8070) );
  NAND2_X1 U8231 ( .A1(n7641), .A2(n8223), .ZN(n14580) );
  NAND2_X1 U8232 ( .A1(n8170), .A2(n8169), .ZN(n14628) );
  NAND2_X1 U8233 ( .A1(n8057), .A2(n8058), .ZN(n14620) );
  NAND2_X1 U8234 ( .A1(n7646), .A2(n8060), .ZN(n8057) );
  NAND2_X1 U8235 ( .A1(n13070), .A2(n7472), .ZN(n13088) );
  INV_X1 U8236 ( .A(n10197), .ZN(n12736) );
  NAND2_X1 U8237 ( .A1(n12735), .A2(n12736), .ZN(n12734) );
  NAND2_X1 U8238 ( .A1(n9518), .A2(n9517), .ZN(n12344) );
  NAND2_X1 U8239 ( .A1(n11844), .A2(n9871), .ZN(n12014) );
  INV_X1 U8240 ( .A(n8231), .ZN(n8230) );
  NAND2_X1 U8241 ( .A1(n9868), .A2(n9867), .ZN(n11472) );
  NAND2_X1 U8242 ( .A1(n9429), .A2(n9428), .ZN(n11471) );
  XNOR2_X1 U8243 ( .A(n11148), .B(n7660), .ZN(n9858) );
  AND2_X1 U8244 ( .A1(n14655), .A2(n14733), .ZN(n8078) );
  NAND2_X1 U8245 ( .A1(n14440), .A2(n16374), .ZN(n7731) );
  NAND2_X1 U8246 ( .A1(n9580), .A2(n9579), .ZN(n12990) );
  NAND2_X1 U8247 ( .A1(n9543), .A2(n9542), .ZN(n12487) );
  INV_X1 U8248 ( .A(n10182), .ZN(n7623) );
  NAND2_X1 U8249 ( .A1(n9421), .A2(n11079), .ZN(n7636) );
  NAND2_X1 U8250 ( .A1(n9824), .A2(n9823), .ZN(n9829) );
  XNOR2_X1 U8251 ( .A(n9849), .B(n9848), .ZN(n11171) );
  INV_X1 U8252 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9848) );
  OR2_X1 U8253 ( .A1(n9835), .A2(n9560), .ZN(n9839) );
  AND2_X1 U8254 ( .A1(n9455), .A2(n9454), .ZN(n9473) );
  INV_X1 U8255 ( .A(n12191), .ZN(n8267) );
  NAND2_X1 U8256 ( .A1(n12186), .A2(n12187), .ZN(n7648) );
  NAND2_X1 U8257 ( .A1(n11139), .A2(n11138), .ZN(n11263) );
  INV_X1 U8258 ( .A(n11142), .ZN(n11138) );
  NAND2_X1 U8259 ( .A1(n14903), .A2(n14862), .ZN(n14982) );
  OR2_X1 U8260 ( .A1(n14861), .A2(n14860), .ZN(n14862) );
  NAND2_X1 U8261 ( .A1(n14982), .A2(n14983), .ZN(n14981) );
  NOR2_X1 U8262 ( .A1(n14947), .A2(n8261), .ZN(n8260) );
  INV_X1 U8263 ( .A(n8262), .ZN(n8261) );
  NAND2_X1 U8264 ( .A1(n14891), .A2(n14812), .ZN(n14819) );
  NOR2_X1 U8265 ( .A1(n15203), .A2(n10743), .ZN(n7600) );
  AND4_X1 U8266 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n14941) );
  NAND2_X1 U8267 ( .A1(n10705), .A2(n10704), .ZN(n15165) );
  NOR2_X1 U8268 ( .A1(n15489), .A2(n15217), .ZN(n7812) );
  NAND2_X1 U8269 ( .A1(n15501), .A2(n15290), .ZN(n8377) );
  INV_X1 U8270 ( .A(n15184), .ZN(n15259) );
  NAND2_X1 U8271 ( .A1(n15284), .A2(n8375), .ZN(n8378) );
  NOR2_X1 U8272 ( .A1(n8428), .A2(n7799), .ZN(n7798) );
  INV_X1 U8273 ( .A(n7802), .ZN(n7799) );
  NAND2_X1 U8274 ( .A1(n8428), .A2(n8427), .ZN(n8430) );
  OR2_X1 U8275 ( .A1(n15317), .A2(n8433), .ZN(n8427) );
  NAND2_X1 U8276 ( .A1(n8475), .A2(n8473), .ZN(n15324) );
  NAND2_X1 U8277 ( .A1(n8181), .A2(n8474), .ZN(n8473) );
  NAND2_X1 U8278 ( .A1(n15351), .A2(n8472), .ZN(n8475) );
  NOR2_X1 U8279 ( .A1(n15340), .A2(n8477), .ZN(n8472) );
  NAND2_X1 U8280 ( .A1(n7791), .A2(n7789), .ZN(n15353) );
  OR2_X1 U8281 ( .A1(n7793), .A2(n7790), .ZN(n7789) );
  INV_X1 U8282 ( .A(n7795), .ZN(n7790) );
  NAND2_X1 U8283 ( .A1(n15353), .A2(n15352), .ZN(n15351) );
  INV_X1 U8284 ( .A(n8452), .ZN(n8449) );
  AOI21_X1 U8285 ( .B1(n8479), .B2(n12761), .A(n7485), .ZN(n7814) );
  AOI21_X1 U8286 ( .B1(n8442), .B2(n8440), .A(n7501), .ZN(n8439) );
  OR2_X1 U8287 ( .A1(n12762), .A2(n8441), .ZN(n8438) );
  INV_X1 U8288 ( .A(n8442), .ZN(n8441) );
  NOR2_X1 U8289 ( .A1(n12976), .A2(n8480), .ZN(n8479) );
  INV_X1 U8290 ( .A(n12970), .ZN(n8480) );
  INV_X1 U8291 ( .A(n12756), .ZN(n7816) );
  NAND2_X1 U8292 ( .A1(n12762), .A2(n12761), .ZN(n12975) );
  NAND2_X1 U8293 ( .A1(n12611), .A2(n8180), .ZN(n12721) );
  NOR2_X1 U8294 ( .A1(n12715), .A2(n8482), .ZN(n8481) );
  INV_X1 U8295 ( .A(n12599), .ZN(n8482) );
  NAND2_X1 U8296 ( .A1(n12457), .A2(n12456), .ZN(n7813) );
  INV_X1 U8297 ( .A(n15049), .ZN(n12722) );
  AND2_X1 U8298 ( .A1(n12294), .A2(n12292), .ZN(n8447) );
  NOR2_X2 U8299 ( .A1(n12129), .A2(n12496), .ZN(n12286) );
  NAND2_X1 U8300 ( .A1(n12115), .A2(n7474), .ZN(n12285) );
  INV_X1 U8301 ( .A(n12123), .ZN(n12116) );
  NAND2_X1 U8302 ( .A1(n7809), .A2(n7808), .ZN(n12115) );
  AND2_X1 U8303 ( .A1(n12087), .A2(n12086), .ZN(n7808) );
  NAND2_X1 U8304 ( .A1(n11440), .A2(n11439), .ZN(n11545) );
  INV_X1 U8305 ( .A(n15410), .ZN(n15448) );
  NAND2_X2 U8306 ( .A1(n7772), .A2(n10612), .ZN(n15517) );
  NAND2_X1 U8307 ( .A1(n13028), .A2(n10702), .ZN(n7772) );
  NAND2_X1 U8308 ( .A1(n10528), .A2(n10527), .ZN(n15555) );
  INV_X1 U8309 ( .A(n16437), .ZN(n16358) );
  NOR2_X1 U8310 ( .A1(n11059), .A2(n11034), .ZN(n15563) );
  OAI21_X1 U8311 ( .B1(n8020), .B2(n8019), .A(n7544), .ZN(n8018) );
  XNOR2_X1 U8312 ( .A(n10106), .B(n10105), .ZN(n14768) );
  NAND2_X1 U8313 ( .A1(n8017), .A2(n8020), .ZN(n10106) );
  AOI21_X1 U8314 ( .B1(n10778), .B2(P1_IR_REG_31__SCAN_IN), .A(n7621), .ZN(
        n7620) );
  NAND2_X1 U8315 ( .A1(n10779), .A2(n7621), .ZN(n10783) );
  INV_X1 U8316 ( .A(n10778), .ZN(n10779) );
  NAND2_X1 U8317 ( .A1(n9316), .A2(n9693), .ZN(n7753) );
  NAND2_X1 U8318 ( .A1(n7887), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10263) );
  XNOR2_X1 U8319 ( .A(n9303), .B(n8352), .ZN(n12164) );
  INV_X1 U8320 ( .A(n9655), .ZN(n8352) );
  OAI21_X1 U8321 ( .B1(n9283), .B2(n7447), .A(n7757), .ZN(n9607) );
  NAND3_X1 U8322 ( .A1(n9247), .A2(n9246), .A3(n9245), .ZN(n9397) );
  INV_X1 U8323 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7804) );
  INV_X1 U8324 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U8325 ( .A1(n16216), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n8035) );
  OAI21_X1 U8326 ( .B1(n11339), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n9103), .ZN(
        n9159) );
  OR2_X1 U8327 ( .A1(n16234), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8031) );
  OR2_X1 U8328 ( .A1(n8030), .A2(n8029), .ZN(n8028) );
  NOR2_X1 U8329 ( .A1(n16227), .A2(n16230), .ZN(n8029) );
  INV_X1 U8330 ( .A(n13274), .ZN(n7585) );
  AND2_X1 U8331 ( .A1(n8935), .A2(n8934), .ZN(n13921) );
  NAND2_X1 U8332 ( .A1(n13273), .A2(n13274), .ZN(n13323) );
  INV_X1 U8333 ( .A(n14195), .ZN(n13342) );
  AND2_X1 U8334 ( .A1(n11590), .A2(n11595), .ZN(n13442) );
  INV_X1 U8335 ( .A(n13642), .ZN(n8241) );
  NAND2_X1 U8336 ( .A1(n13644), .A2(n13643), .ZN(n8240) );
  INV_X1 U8337 ( .A(n14062), .ZN(n13658) );
  AOI21_X1 U8338 ( .B1(n12234), .B2(n12233), .A(n12232), .ZN(n12366) );
  AND2_X1 U8339 ( .A1(n12890), .A2(n12891), .ZN(n7854) );
  OR2_X1 U8340 ( .A1(n13784), .A2(n14147), .ZN(n13821) );
  AOI21_X1 U8341 ( .B1(n13821), .B2(n13820), .A(n13819), .ZN(n13843) );
  OR2_X1 U8342 ( .A1(n13810), .A2(n13808), .ZN(n8161) );
  NAND2_X1 U8343 ( .A1(n8158), .A2(n8156), .ZN(n8155) );
  INV_X1 U8344 ( .A(n8157), .ZN(n8156) );
  NAND2_X1 U8345 ( .A1(n13813), .A2(n13827), .ZN(n8158) );
  OAI21_X1 U8346 ( .B1(n16292), .B2(n13812), .A(n13811), .ZN(n8157) );
  NOR2_X1 U8347 ( .A1(n11495), .A2(n11494), .ZN(n13847) );
  NAND2_X1 U8348 ( .A1(n7786), .A2(n13840), .ZN(n7785) );
  XNOR2_X1 U8349 ( .A(n13835), .B(n13834), .ZN(n7786) );
  OR2_X1 U8350 ( .A1(n13805), .A2(n7551), .ZN(n7823) );
  NAND2_X1 U8351 ( .A1(n7824), .A2(n7821), .ZN(n7820) );
  NAND2_X1 U8352 ( .A1(n7827), .A2(n7550), .ZN(n7821) );
  AOI21_X1 U8353 ( .B1(n10818), .B2(n16309), .A(n10817), .ZN(n13185) );
  AND2_X1 U8354 ( .A1(n13862), .A2(n13861), .ZN(n14111) );
  OAI21_X1 U8355 ( .B1(n13878), .B2(n7506), .A(n8082), .ZN(n8090) );
  AND2_X1 U8356 ( .A1(n13900), .A2(n7949), .ZN(n13885) );
  AND3_X1 U8357 ( .A1(n8730), .A2(n8729), .A3(n8728), .ZN(n14101) );
  INV_X1 U8358 ( .A(n12427), .ZN(n12476) );
  INV_X1 U8359 ( .A(n16477), .ZN(n14109) );
  NAND2_X1 U8360 ( .A1(n10796), .A2(n10795), .ZN(n13866) );
  OR2_X1 U8361 ( .A1(n8954), .A2(n15637), .ZN(n10795) );
  NAND2_X1 U8362 ( .A1(n14240), .A2(n7432), .ZN(n14120) );
  NAND2_X1 U8363 ( .A1(n13460), .A2(n13459), .ZN(n16480) );
  AOI21_X1 U8364 ( .B1(n14236), .B2(n13458), .A(n10802), .ZN(n13188) );
  NAND2_X1 U8365 ( .A1(n7958), .A2(n14111), .ZN(n14168) );
  NAND2_X1 U8366 ( .A1(n14110), .A2(n10820), .ZN(n7958) );
  INV_X1 U8367 ( .A(n13874), .ZN(n13280) );
  OR2_X1 U8368 ( .A1(n13462), .A2(n10872), .ZN(n8610) );
  NAND2_X1 U8369 ( .A1(n16476), .A2(n16418), .ZN(n14221) );
  XNOR2_X1 U8370 ( .A(n8320), .B(n8319), .ZN(n14285) );
  INV_X1 U8371 ( .A(n14267), .ZN(n8319) );
  AND2_X1 U8372 ( .A1(n11150), .A2(n11151), .ZN(n7595) );
  NAND2_X1 U8373 ( .A1(n11206), .A2(n11207), .ZN(n11205) );
  NAND2_X1 U8374 ( .A1(n8307), .A2(n8306), .ZN(n8305) );
  OR2_X1 U8375 ( .A1(n8304), .A2(n8303), .ZN(n8302) );
  OR2_X1 U8376 ( .A1(n11385), .A2(n11156), .ZN(n8303) );
  AND2_X1 U8377 ( .A1(n8302), .A2(n8301), .ZN(n11415) );
  OR2_X1 U8378 ( .A1(n12844), .A2(n10113), .ZN(n9726) );
  NAND2_X1 U8379 ( .A1(n11216), .A2(n11217), .ZN(n11215) );
  INV_X1 U8380 ( .A(n14475), .ZN(n14388) );
  NAND2_X1 U8381 ( .A1(n9776), .A2(n9775), .ZN(n14474) );
  NAND4_X1 U8382 ( .A1(n9446), .A2(n9445), .A3(n9444), .A4(n9443), .ZN(n14407)
         );
  NAND2_X1 U8383 ( .A1(n10139), .A2(n10138), .ZN(n10152) );
  XNOR2_X1 U8384 ( .A(n7589), .B(n10209), .ZN(n14652) );
  NAND2_X1 U8385 ( .A1(n14437), .A2(n7590), .ZN(n7589) );
  NAND2_X1 U8386 ( .A1(n9796), .A2(n7591), .ZN(n7590) );
  INV_X1 U8387 ( .A(n14457), .ZN(n7591) );
  AOI21_X1 U8388 ( .B1(n9916), .B2(n14603), .A(n9915), .ZN(n14651) );
  NAND2_X1 U8389 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  AOI21_X1 U8390 ( .B1(n14648), .B2(n14596), .A(n9924), .ZN(n9925) );
  NAND2_X1 U8391 ( .A1(n14451), .A2(n14450), .ZN(n14653) );
  NAND2_X1 U8392 ( .A1(n9855), .A2(n16041), .ZN(n16455) );
  OAI21_X1 U8393 ( .B1(n9852), .B2(P2_D_REG_0__SCAN_IN), .A(n9851), .ZN(n16040) );
  NAND2_X1 U8394 ( .A1(n15000), .A2(n7616), .ZN(n14905) );
  NAND2_X1 U8395 ( .A1(n14854), .A2(n14855), .ZN(n7616) );
  NAND2_X1 U8396 ( .A1(n10427), .A2(n10426), .ZN(n12567) );
  OR2_X1 U8397 ( .A1(n14839), .A2(n14838), .ZN(n7703) );
  OR2_X1 U8398 ( .A1(n10892), .A2(n15067), .ZN(n8418) );
  OR2_X1 U8399 ( .A1(n10309), .A2(n10851), .ZN(n8419) );
  INV_X1 U8400 ( .A(n15369), .ZN(n15182) );
  NAND2_X1 U8401 ( .A1(n10517), .A2(n10516), .ZN(n15562) );
  NAND2_X1 U8402 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  INV_X1 U8403 ( .A(n15396), .ZN(n15545) );
  INV_X1 U8404 ( .A(n15044), .ZN(n15012) );
  INV_X1 U8405 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8565) );
  AND2_X1 U8406 ( .A1(n7515), .A2(n7605), .ZN(n15491) );
  NAND2_X1 U8407 ( .A1(n15254), .A2(n15445), .ZN(n7605) );
  NAND2_X1 U8408 ( .A1(n10455), .A2(n10454), .ZN(n12851) );
  INV_X1 U8409 ( .A(n15480), .ZN(n7819) );
  INV_X1 U8410 ( .A(n8486), .ZN(n8485) );
  XNOR2_X1 U8411 ( .A(n15202), .B(n8490), .ZN(n15481) );
  XNOR2_X1 U8412 ( .A(n8489), .B(n15203), .ZN(n15482) );
  OR2_X1 U8413 ( .A1(n16242), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8037) );
  AND2_X1 U8414 ( .A1(n16242), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8038) );
  AOI22_X1 U8415 ( .A1(n9933), .A2(n9930), .B1(n9959), .B2(n12000), .ZN(n9947)
         );
  AOI21_X1 U8416 ( .B1(n9929), .B2(n9930), .A(n9928), .ZN(n9951) );
  XNOR2_X1 U8417 ( .A(n7606), .B(SI_29_), .ZN(n15634) );
  NAND2_X1 U8418 ( .A1(n7570), .A2(n7569), .ZN(n7700) );
  INV_X1 U8419 ( .A(n9977), .ZN(n7569) );
  NAND2_X1 U8420 ( .A1(n7568), .A2(n7567), .ZN(n7691) );
  INV_X1 U8421 ( .A(n9987), .ZN(n7567) );
  INV_X1 U8422 ( .A(n9993), .ZN(n7572) );
  INV_X1 U8423 ( .A(n9999), .ZN(n7714) );
  INV_X1 U8424 ( .A(n10345), .ZN(n7864) );
  INV_X1 U8425 ( .A(n10375), .ZN(n8406) );
  INV_X1 U8426 ( .A(n10392), .ZN(n10395) );
  AOI21_X1 U8427 ( .B1(n10414), .B2(n7898), .A(n7897), .ZN(n7896) );
  INV_X1 U8428 ( .A(n10428), .ZN(n7897) );
  NOR2_X1 U8429 ( .A1(n10415), .A2(n7900), .ZN(n7898) );
  NOR2_X1 U8430 ( .A1(n7895), .A2(n10429), .ZN(n7894) );
  NOR2_X1 U8431 ( .A1(n8411), .A2(n10415), .ZN(n7895) );
  INV_X1 U8432 ( .A(n10010), .ZN(n7712) );
  OAI21_X1 U8433 ( .B1(n7910), .B2(n10489), .A(n10487), .ZN(n7907) );
  NOR2_X1 U8434 ( .A1(n7905), .A2(n10488), .ZN(n7904) );
  INV_X1 U8435 ( .A(n7910), .ZN(n7905) );
  AND2_X1 U8436 ( .A1(n10460), .A2(n10459), .ZN(n7901) );
  OAI21_X1 U8437 ( .B1(n10443), .B2(n8399), .A(n7557), .ZN(n10459) );
  NOR2_X1 U8438 ( .A1(n10458), .A2(n7558), .ZN(n7557) );
  AOI22_X1 U8439 ( .A1(n7908), .A2(n7906), .B1(n8413), .B2(n7904), .ZN(n7902)
         );
  NAND2_X1 U8440 ( .A1(n7909), .A2(n10488), .ZN(n7908) );
  INV_X1 U8441 ( .A(n8413), .ZN(n7909) );
  NOR2_X1 U8442 ( .A1(n7911), .A2(n10473), .ZN(n8413) );
  NOR2_X1 U8443 ( .A1(n7904), .A2(n7906), .ZN(n7903) );
  NAND2_X1 U8444 ( .A1(n7746), .A2(n7745), .ZN(n7744) );
  INV_X1 U8445 ( .A(n10027), .ZN(n7745) );
  NAND2_X1 U8446 ( .A1(n8404), .A2(n8403), .ZN(n8401) );
  OAI21_X1 U8447 ( .B1(n10519), .B2(n7876), .A(n7874), .ZN(n10530) );
  NAND2_X1 U8448 ( .A1(n7749), .A2(n7748), .ZN(n7747) );
  INV_X1 U8449 ( .A(n10040), .ZN(n7748) );
  AOI21_X1 U8450 ( .B1(n7872), .B2(n7876), .A(n7870), .ZN(n7869) );
  INV_X1 U8451 ( .A(n10046), .ZN(n7612) );
  NAND2_X1 U8452 ( .A1(n8388), .A2(n8386), .ZN(n8384) );
  OAI21_X1 U8453 ( .B1(n10578), .B2(n7885), .A(n7883), .ZN(n10590) );
  NAND2_X1 U8454 ( .A1(n7538), .A2(n10056), .ZN(n8455) );
  NOR2_X1 U8455 ( .A1(n10615), .A2(n10613), .ZN(n8393) );
  NAND2_X1 U8456 ( .A1(n10615), .A2(n10613), .ZN(n8392) );
  AOI21_X1 U8457 ( .B1(n7881), .B2(n7885), .A(n7879), .ZN(n7878) );
  NOR2_X1 U8458 ( .A1(n10641), .A2(n10638), .ZN(n8408) );
  NAND2_X1 U8459 ( .A1(n7777), .A2(n12902), .ZN(n12903) );
  INV_X1 U8460 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8516) );
  NOR2_X1 U8461 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8131) );
  INV_X1 U8462 ( .A(n10082), .ZN(n7709) );
  NAND2_X1 U8463 ( .A1(n7460), .A2(n8467), .ZN(n8466) );
  NOR2_X1 U8464 ( .A1(n10165), .A2(n10166), .ZN(n8006) );
  OR2_X1 U8465 ( .A1(n10151), .A2(n7531), .ZN(n7997) );
  INV_X1 U8466 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U8467 ( .A1(n9877), .A2(n9878), .ZN(n8075) );
  INV_X1 U8468 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U8469 ( .A1(n8013), .A2(n8011), .ZN(n9325) );
  AOI21_X1 U8470 ( .B1(n8014), .B2(n8016), .A(n8012), .ZN(n8011) );
  INV_X1 U8471 ( .A(n9323), .ZN(n8012) );
  INV_X1 U8472 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7750) );
  AND2_X1 U8473 ( .A1(n9669), .A2(n9309), .ZN(n9310) );
  NAND2_X1 U8474 ( .A1(n9306), .A2(n11514), .ZN(n9311) );
  NAND2_X1 U8475 ( .A1(n9644), .A2(n9302), .ZN(n9304) );
  INV_X1 U8476 ( .A(n7994), .ZN(n7993) );
  OAI21_X1 U8477 ( .B1(n9264), .B2(n7995), .A(n9267), .ZN(n7994) );
  INV_X1 U8478 ( .A(n9266), .ZN(n7995) );
  NAND2_X1 U8479 ( .A1(n9419), .A2(n9255), .ZN(n7665) );
  OAI21_X1 U8480 ( .B1(n9126), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9086), .ZN(
        n9087) );
  INV_X1 U8481 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n15806) );
  NOR2_X1 U8482 ( .A1(n13360), .A2(n8348), .ZN(n8344) );
  OR2_X1 U8483 ( .A1(n13866), .A2(n13607), .ZN(n7720) );
  NAND2_X1 U8484 ( .A1(n7563), .A2(n7561), .ZN(n13606) );
  NOR2_X1 U8485 ( .A1(n13466), .A2(n13637), .ZN(n13611) );
  NAND2_X1 U8486 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  OR2_X1 U8487 ( .A1(n12663), .A2(n12662), .ZN(n12665) );
  INV_X1 U8488 ( .A(n7968), .ZN(n7705) );
  OAI22_X1 U8489 ( .A1(n7970), .A2(n7972), .B1(n7973), .B2(n7969), .ZN(n7968)
         );
  INV_X1 U8490 ( .A(n12373), .ZN(n7969) );
  INV_X1 U8491 ( .A(n7841), .ZN(n7837) );
  OR2_X1 U8492 ( .A1(n12667), .A2(n12668), .ZN(n7777) );
  AOI21_X1 U8493 ( .B1(n7964), .B2(n7984), .A(n12894), .ZN(n7982) );
  INV_X1 U8494 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15914) );
  INV_X1 U8495 ( .A(n13856), .ZN(n8084) );
  NOR2_X1 U8496 ( .A1(n13474), .A2(n8087), .ZN(n8086) );
  OR2_X1 U8497 ( .A1(n9012), .A2(n7923), .ZN(n7922) );
  INV_X1 U8498 ( .A(n13585), .ZN(n7923) );
  NOR2_X1 U8499 ( .A1(n8928), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U8500 ( .A1(n8883), .A2(n15897), .ZN(n8910) );
  NOR2_X1 U8501 ( .A1(n8872), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8871) );
  INV_X1 U8502 ( .A(n8810), .ZN(n8127) );
  OAI21_X1 U8503 ( .B1(n7455), .B2(n8127), .A(n14017), .ZN(n8126) );
  OR2_X1 U8504 ( .A1(n14159), .A2(n14046), .ZN(n13561) );
  AND2_X1 U8505 ( .A1(n8801), .A2(n8505), .ZN(n8817) );
  NOR2_X1 U8506 ( .A1(n8802), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8801) );
  INV_X1 U8507 ( .A(n8095), .ZN(n8094) );
  OAI21_X1 U8508 ( .B1(n8098), .B2(n8096), .A(n8775), .ZN(n8095) );
  INV_X1 U8509 ( .A(n8097), .ZN(n8096) );
  NOR2_X1 U8510 ( .A1(n8748), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8747) );
  AND2_X1 U8511 ( .A1(n8669), .A2(n15892), .ZN(n8685) );
  NOR2_X1 U8512 ( .A1(n8670), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8669) );
  INV_X1 U8513 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15902) );
  NOR2_X1 U8514 ( .A1(n7918), .A2(n7919), .ZN(n7917) );
  OAI21_X1 U8515 ( .B1(n13628), .B2(n7918), .A(n13503), .ZN(n7914) );
  OR2_X1 U8516 ( .A1(n8655), .A2(n10865), .ZN(n8574) );
  AOI21_X1 U8517 ( .B1(n7949), .B2(n13893), .A(n9013), .ZN(n7947) );
  INV_X1 U8518 ( .A(n7949), .ZN(n7948) );
  NAND2_X1 U8519 ( .A1(n8341), .A2(n8726), .ZN(n8847) );
  NAND2_X1 U8520 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7684), .ZN(n7683) );
  INV_X1 U8521 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9273) );
  INV_X1 U8522 ( .A(n8534), .ZN(n8218) );
  INV_X1 U8523 ( .A(n12222), .ZN(n8296) );
  INV_X1 U8524 ( .A(n12057), .ZN(n8294) );
  NAND2_X1 U8525 ( .A1(n14250), .A2(n14251), .ZN(n8317) );
  INV_X1 U8526 ( .A(n13061), .ZN(n8291) );
  INV_X1 U8527 ( .A(n12947), .ZN(n8289) );
  INV_X1 U8528 ( .A(n12688), .ZN(n8286) );
  INV_X1 U8529 ( .A(n12486), .ZN(n8284) );
  INV_X1 U8530 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U8531 ( .A1(n9196), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9528) );
  INV_X1 U8532 ( .A(n9510), .ZN(n9196) );
  INV_X1 U8533 ( .A(n9692), .ZN(n8222) );
  NOR2_X1 U8534 ( .A1(n14628), .A2(n14709), .ZN(n8168) );
  OR2_X1 U8535 ( .A1(n9582), .A2(n9581), .ZN(n9597) );
  INV_X1 U8536 ( .A(n9447), .ZN(n8229) );
  AOI21_X1 U8537 ( .B1(n8195), .B2(n8197), .A(n8193), .ZN(n8192) );
  INV_X1 U8538 ( .A(n10204), .ZN(n8193) );
  NOR2_X2 U8539 ( .A1(n11847), .A2(n11979), .ZN(n12018) );
  INV_X1 U8540 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U8541 ( .A1(n9223), .A2(n7463), .ZN(n9224) );
  NOR2_X1 U8542 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n9820) );
  OR2_X1 U8543 ( .A1(n10281), .A2(n12597), .ZN(n10282) );
  NOR2_X1 U8544 ( .A1(n15368), .A2(n15533), .ZN(n8182) );
  AND2_X1 U8545 ( .A1(n7795), .A2(n15181), .ZN(n7792) );
  AND2_X1 U8546 ( .A1(n15365), .A2(n7461), .ZN(n7793) );
  OR2_X1 U8547 ( .A1(n15533), .A2(n15182), .ZN(n15196) );
  NAND2_X1 U8548 ( .A1(n15545), .A2(n15370), .ZN(n8452) );
  NAND2_X1 U8549 ( .A1(n10521), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10534) );
  INV_X1 U8550 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10445) );
  INV_X1 U8551 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10379) );
  OAI21_X1 U8552 ( .B1(n15239), .B2(n15238), .A(n7504), .ZN(n7771) );
  INV_X1 U8553 ( .A(n8371), .ZN(n8370) );
  OAI22_X1 U8554 ( .A1(n15259), .A2(n8377), .B1(n15267), .B2(n15243), .ZN(
        n8371) );
  NOR2_X1 U8555 ( .A1(n15259), .A2(n8374), .ZN(n8373) );
  INV_X1 U8556 ( .A(n8375), .ZN(n8374) );
  AND2_X1 U8557 ( .A1(n12597), .A2(n15157), .ZN(n11034) );
  INV_X1 U8558 ( .A(n10105), .ZN(n8019) );
  AOI21_X1 U8559 ( .B1(n8022), .B2(n9354), .A(n8021), .ZN(n8020) );
  INV_X1 U8560 ( .A(n9797), .ZN(n8021) );
  NOR2_X1 U8561 ( .A1(n9798), .A2(n8023), .ZN(n8022) );
  INV_X1 U8562 ( .A(n9338), .ZN(n8023) );
  AND2_X1 U8563 ( .A1(n9335), .A2(n9334), .ZN(n9780) );
  INV_X1 U8564 ( .A(n10261), .ZN(n10262) );
  NAND2_X1 U8565 ( .A1(n9305), .A2(SI_18_), .ZN(n9669) );
  INV_X1 U8566 ( .A(n9304), .ZN(n9305) );
  AND2_X1 U8567 ( .A1(n9294), .A2(n9293), .ZN(n9606) );
  INV_X1 U8568 ( .A(n9285), .ZN(n7759) );
  NOR2_X1 U8569 ( .A1(n9286), .A2(n7762), .ZN(n7761) );
  INV_X1 U8570 ( .A(n9282), .ZN(n7762) );
  INV_X1 U8571 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U8572 ( .A1(n8354), .A2(n8353), .ZN(n9489) );
  AOI21_X1 U8573 ( .B1(n8356), .B2(n8358), .A(n7500), .ZN(n8353) );
  OR2_X1 U8574 ( .A1(n10346), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n10370) );
  XNOR2_X1 U8575 ( .A(n9251), .B(SI_3_), .ZN(n9413) );
  NAND2_X1 U8576 ( .A1(n9249), .A2(n10847), .ZN(n7624) );
  XNOR2_X1 U8577 ( .A(n9085), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U8578 ( .A1(n9098), .A2(n9097), .ZN(n9118) );
  OR2_X1 U8579 ( .A1(n9145), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9097) );
  OAI21_X1 U8580 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9108), .A(n9107), .ZN(
        n9169) );
  NOR2_X1 U8581 ( .A1(n13303), .A2(n8326), .ZN(n8325) );
  INV_X1 U8582 ( .A(n13241), .ZN(n8326) );
  AND2_X1 U8583 ( .A1(n13269), .A2(n13268), .ZN(n13359) );
  INV_X1 U8584 ( .A(n13260), .ZN(n13387) );
  NAND2_X1 U8585 ( .A1(n13254), .A2(n7473), .ZN(n8331) );
  NAND2_X1 U8586 ( .A1(n8333), .A2(n13255), .ZN(n13256) );
  XNOR2_X1 U8587 ( .A(n13265), .B(n13202), .ZN(n11799) );
  OR2_X1 U8588 ( .A1(n12637), .A2(n12638), .ZN(n12635) );
  AND2_X1 U8589 ( .A1(n13617), .A2(n13864), .ZN(n7682) );
  NOR4_X1 U8590 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13933), .ZN(
        n13640) );
  AND2_X1 U8591 ( .A1(n7833), .A2(n7832), .ZN(n7831) );
  NAND2_X1 U8592 ( .A1(n13775), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7832) );
  OR2_X1 U8593 ( .A1(n13775), .A2(n11490), .ZN(n7833) );
  AND2_X1 U8594 ( .A1(n7831), .A2(n7830), .ZN(n11634) );
  INV_X1 U8595 ( .A(n11509), .ZN(n7830) );
  NAND2_X1 U8596 ( .A1(n11622), .A2(n11623), .ZN(n11659) );
  AND2_X1 U8597 ( .A1(n8148), .A2(n13681), .ZN(n11661) );
  NAND2_X1 U8598 ( .A1(n8148), .A2(n7553), .ZN(n13683) );
  AND2_X1 U8599 ( .A1(n11768), .A2(n13680), .ZN(n7851) );
  INV_X1 U8600 ( .A(n11782), .ZN(n7963) );
  NAND2_X1 U8601 ( .A1(n11778), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11957) );
  INV_X1 U8602 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15713) );
  OR2_X1 U8603 ( .A1(n8152), .A2(n12904), .ZN(n12905) );
  INV_X1 U8604 ( .A(n13715), .ZN(n7975) );
  NAND2_X1 U8605 ( .A1(n8139), .A2(n8138), .ZN(n13742) );
  INV_X1 U8606 ( .A(n13741), .ZN(n8139) );
  NAND2_X1 U8607 ( .A1(n13749), .A2(n7855), .ZN(n13774) );
  OR2_X1 U8608 ( .A1(n13750), .A2(n13751), .ZN(n7855) );
  NAND2_X1 U8609 ( .A1(n13766), .A2(n8140), .ZN(n8137) );
  INV_X1 U8610 ( .A(n7827), .ZN(n7826) );
  INV_X1 U8611 ( .A(n13656), .ZN(n13607) );
  INV_X1 U8612 ( .A(n8083), .ZN(n8082) );
  OAI21_X1 U8613 ( .B1(n8086), .B2(n8084), .A(n13864), .ZN(n8083) );
  OAI211_X1 U8614 ( .C1(n8089), .C2(n8081), .A(n8080), .B(n10797), .ZN(n13858)
         );
  AND2_X1 U8615 ( .A1(n13859), .A2(n13856), .ZN(n10797) );
  NAND2_X1 U8616 ( .A1(n8086), .A2(n8950), .ZN(n8080) );
  INV_X1 U8617 ( .A(n8086), .ZN(n8081) );
  INV_X1 U8618 ( .A(n8087), .ZN(n8085) );
  NAND2_X1 U8619 ( .A1(n8088), .A2(n8086), .ZN(n13857) );
  NOR2_X1 U8620 ( .A1(n13882), .A2(n7950), .ZN(n7949) );
  INV_X1 U8621 ( .A(n13590), .ZN(n7950) );
  NAND2_X1 U8622 ( .A1(n8114), .A2(n7450), .ZN(n8113) );
  INV_X1 U8623 ( .A(n8936), .ZN(n8114) );
  NAND2_X1 U8624 ( .A1(n13902), .A2(n13901), .ZN(n13900) );
  INV_X1 U8625 ( .A(n7946), .ZN(n13940) );
  OR2_X1 U8626 ( .A1(n8854), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8872) );
  INV_X1 U8627 ( .A(n13991), .ZN(n13999) );
  NAND2_X1 U8628 ( .A1(n8107), .A2(n8106), .ZN(n13990) );
  AOI21_X1 U8629 ( .B1(n7926), .B2(n7929), .A(n14017), .ZN(n7924) );
  AOI21_X1 U8630 ( .B1(n7930), .B2(n7928), .A(n7927), .ZN(n7926) );
  INV_X1 U8631 ( .A(n13561), .ZN(n7927) );
  INV_X1 U8632 ( .A(n7933), .ZN(n7928) );
  INV_X1 U8633 ( .A(n7930), .ZN(n7929) );
  NAND2_X1 U8634 ( .A1(n14029), .A2(n8810), .ZN(n14018) );
  OR2_X1 U8635 ( .A1(n8733), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8748) );
  OR2_X1 U8636 ( .A1(n8716), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8733) );
  OAI21_X1 U8637 ( .B1(n12546), .B2(n8123), .A(n8122), .ZN(n13001) );
  AOI21_X1 U8638 ( .B1(n8124), .B2(n13518), .A(n7490), .ZN(n8122) );
  INV_X1 U8639 ( .A(n8124), .ZN(n8123) );
  NAND2_X1 U8640 ( .A1(n12546), .A2(n13622), .ZN(n12545) );
  NAND2_X1 U8641 ( .A1(n12528), .A2(n8647), .ZN(n12440) );
  OR2_X1 U8642 ( .A1(n8648), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8670) );
  AND2_X1 U8643 ( .A1(n13516), .A2(n13515), .ZN(n13621) );
  OR2_X1 U8644 ( .A1(n8625), .A2(n13624), .ZN(n8629) );
  NAND2_X1 U8645 ( .A1(n13512), .A2(n13511), .ZN(n13623) );
  NAND2_X1 U8646 ( .A1(n8991), .A2(n16308), .ZN(n8585) );
  NAND2_X1 U8647 ( .A1(n8115), .A2(n8117), .ZN(n8108) );
  NAND2_X1 U8648 ( .A1(n8920), .A2(n8919), .ZN(n13257) );
  NAND2_X1 U8649 ( .A1(n8100), .A2(n8101), .ZN(n13965) );
  INV_X1 U8650 ( .A(n8102), .ZN(n8101) );
  OAI21_X1 U8651 ( .B1(n8106), .B2(n8103), .A(n8497), .ZN(n8102) );
  NAND2_X1 U8652 ( .A1(n8732), .A2(n8098), .ZN(n8093) );
  INV_X1 U8653 ( .A(n7938), .ZN(n7937) );
  AOI21_X1 U8654 ( .B1(n7938), .B2(n7940), .A(n13137), .ZN(n7936) );
  NAND2_X1 U8655 ( .A1(n12545), .A2(n8124), .ZN(n12918) );
  AND2_X1 U8656 ( .A1(n12545), .A2(n8684), .ZN(n12919) );
  AND3_X1 U8657 ( .A1(n8683), .A2(n8682), .A3(n8681), .ZN(n12586) );
  AND3_X1 U8658 ( .A1(n8646), .A2(n8645), .A3(n8644), .ZN(n12336) );
  NAND2_X1 U8659 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n7738), .ZN(n7737) );
  NAND2_X1 U8660 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n7719), .ZN(n7718) );
  AND2_X1 U8661 ( .A1(n9031), .A2(n9030), .ZN(n9059) );
  NAND2_X1 U8662 ( .A1(n9026), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U8663 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n8245), .ZN(n8244) );
  XNOR2_X1 U8664 ( .A(n8976), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12430) );
  XNOR2_X1 U8665 ( .A(n8978), .B(P3_IR_REG_20__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U8666 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n8189), .ZN(n8188) );
  INV_X1 U8667 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8189) );
  XNOR2_X1 U8668 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n8844) );
  AOI21_X1 U8669 ( .B1(n8212), .B2(n8214), .A(n7539), .ZN(n8209) );
  XNOR2_X1 U8670 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8811) );
  NOR2_X1 U8671 ( .A1(n8761), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8765) );
  XNOR2_X1 U8672 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8755) );
  NAND2_X1 U8673 ( .A1(n7688), .A2(n8547), .ZN(n8743) );
  INV_X1 U8674 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8546) );
  CLKBUF_X1 U8675 ( .A(n8725), .Z(n8726) );
  XNOR2_X1 U8676 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8695) );
  INV_X1 U8677 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8693) );
  AND2_X1 U8678 ( .A1(n10879), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U8679 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8677) );
  NOR2_X1 U8680 ( .A1(n8642), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8661) );
  XNOR2_X1 U8681 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8638) );
  INV_X1 U8682 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9493) );
  OR2_X1 U8683 ( .A1(n9494), .A2(n9493), .ZN(n9510) );
  NAND2_X1 U8684 ( .A1(n9199), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9636) );
  CLKBUF_X1 U8685 ( .A(n14334), .Z(n7666) );
  INV_X1 U8686 ( .A(n9727), .ZN(n9203) );
  NAND2_X1 U8687 ( .A1(n9197), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9569) );
  INV_X1 U8688 ( .A(n9546), .ZN(n9197) );
  AND2_X1 U8689 ( .A1(n10182), .A2(n10217), .ZN(n11162) );
  NAND2_X1 U8690 ( .A1(n9378), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8043) );
  OR2_X1 U8691 ( .A1(n9392), .A2(n11931), .ZN(n9384) );
  NAND2_X1 U8692 ( .A1(n9378), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9383) );
  NOR2_X1 U8693 ( .A1(n8164), .A2(n14658), .ZN(n8162) );
  OR2_X1 U8694 ( .A1(n14649), .A2(n14655), .ZN(n8164) );
  NAND2_X1 U8695 ( .A1(n14431), .A2(n14432), .ZN(n14430) );
  INV_X1 U8696 ( .A(n10209), .ZN(n9901) );
  OR2_X1 U8697 ( .A1(n8236), .A2(n8238), .ZN(n8234) );
  OR2_X1 U8698 ( .A1(n14482), .A2(n8235), .ZN(n8233) );
  OR2_X1 U8699 ( .A1(n8238), .A2(n7527), .ZN(n8235) );
  AOI21_X1 U8700 ( .B1(n14472), .B2(n8051), .A(n7464), .ZN(n8050) );
  INV_X1 U8701 ( .A(n9899), .ZN(n8051) );
  INV_X1 U8702 ( .A(n8166), .ZN(n14556) );
  OAI21_X1 U8703 ( .B1(n14579), .B2(n8067), .A(n8064), .ZN(n14550) );
  INV_X1 U8704 ( .A(n8068), .ZN(n8067) );
  AOI21_X1 U8705 ( .B1(n8068), .B2(n8066), .A(n8065), .ZN(n8064) );
  INV_X1 U8706 ( .A(n9891), .ZN(n8065) );
  NAND2_X1 U8707 ( .A1(n8168), .A2(n8167), .ZN(n14589) );
  INV_X1 U8708 ( .A(n8168), .ZN(n14609) );
  NOR2_X1 U8709 ( .A1(n9652), .A2(n8252), .ZN(n8251) );
  AOI21_X1 U8710 ( .B1(n8055), .B2(n8054), .A(n7487), .ZN(n8053) );
  INV_X1 U8711 ( .A(n8060), .ZN(n8054) );
  OR2_X1 U8712 ( .A1(n9636), .A2(n9635), .ZN(n9648) );
  INV_X1 U8713 ( .A(n8170), .ZN(n14630) );
  NAND2_X1 U8714 ( .A1(n8062), .A2(n9884), .ZN(n13087) );
  NAND2_X1 U8715 ( .A1(n8063), .A2(n7453), .ZN(n8062) );
  INV_X1 U8716 ( .A(n7646), .ZN(n8063) );
  OR2_X1 U8717 ( .A1(n12790), .A2(n12990), .ZN(n12880) );
  AOI21_X1 U8718 ( .B1(n8206), .B2(n8208), .A(n7465), .ZN(n8204) );
  NAND2_X1 U8719 ( .A1(n12742), .A2(n12697), .ZN(n12790) );
  NAND2_X1 U8720 ( .A1(n12321), .A2(n12320), .ZN(n12319) );
  NAND2_X1 U8721 ( .A1(n9526), .A2(n9525), .ZN(n12400) );
  INV_X1 U8722 ( .A(n14403), .ZN(n12408) );
  NAND2_X1 U8723 ( .A1(n8227), .A2(n8226), .ZN(n12012) );
  NAND2_X1 U8724 ( .A1(n8231), .A2(n9468), .ZN(n8226) );
  OR2_X1 U8725 ( .A1(n11471), .A2(n8228), .ZN(n8227) );
  NAND2_X1 U8726 ( .A1(n8229), .A2(n9468), .ZN(n8228) );
  NAND2_X1 U8727 ( .A1(n12012), .A2(n12013), .ZN(n12011) );
  INV_X1 U8728 ( .A(n8041), .ZN(n7592) );
  NAND2_X1 U8729 ( .A1(n9865), .A2(n9864), .ZN(n11397) );
  OAI21_X1 U8730 ( .B1(n11198), .B2(n11197), .A(n9387), .ZN(n11275) );
  NAND2_X1 U8731 ( .A1(n11223), .A2(n11198), .ZN(n9861) );
  AND2_X1 U8732 ( .A1(n8237), .A2(n8236), .ZN(n14662) );
  INV_X1 U8733 ( .A(n14734), .ZN(n14692) );
  NAND2_X1 U8734 ( .A1(n9595), .A2(n9594), .ZN(n14732) );
  NAND2_X1 U8735 ( .A1(n9507), .A2(n9506), .ZN(n12259) );
  INV_X1 U8736 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U8737 ( .A1(n9821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9827) );
  OR2_X1 U8738 ( .A1(n9847), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9821) );
  INV_X1 U8739 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9826) );
  INV_X1 U8740 ( .A(n9722), .ZN(n9723) );
  OR2_X1 U8741 ( .A1(n9592), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9610) );
  NOR2_X1 U8742 ( .A1(n9558), .A2(n9557), .ZN(n9562) );
  CLKBUF_X1 U8743 ( .A(n9432), .Z(n9433) );
  INV_X1 U8744 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9213) );
  AOI21_X1 U8745 ( .B1(n14803), .B2(n14802), .A(n7650), .ZN(n14892) );
  AND2_X1 U8746 ( .A1(n14800), .A2(n14801), .ZN(n7650) );
  INV_X1 U8747 ( .A(n14906), .ZN(n7629) );
  OR2_X1 U8748 ( .A1(n10553), .A2(n10552), .ZN(n10567) );
  NAND2_X1 U8749 ( .A1(n14884), .A2(n14885), .ZN(n14931) );
  INV_X1 U8750 ( .A(n8265), .ZN(n12190) );
  NAND2_X1 U8751 ( .A1(n14847), .A2(n14848), .ZN(n8262) );
  INV_X1 U8752 ( .A(n15048), .ZN(n14896) );
  INV_X1 U8753 ( .A(n10629), .ZN(n10630) );
  OR2_X1 U8754 ( .A1(n15032), .A2(n15033), .ZN(n8280) );
  NOR2_X1 U8755 ( .A1(n8272), .A2(n8271), .ZN(n8270) );
  INV_X1 U8756 ( .A(n14971), .ZN(n8271) );
  OR2_X1 U8757 ( .A1(n10380), .A2(n10379), .ZN(n10399) );
  INV_X1 U8758 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U8759 ( .A1(n10399), .A2(n10398), .ZN(n10417) );
  NAND2_X1 U8760 ( .A1(n12190), .A2(n12191), .ZN(n12503) );
  NOR2_X1 U8761 ( .A1(n10446), .A2(n10445), .ZN(n10461) );
  OR2_X1 U8762 ( .A1(n10431), .A2(n10430), .ZN(n10446) );
  NAND2_X1 U8763 ( .A1(n11703), .A2(n11704), .ZN(n11830) );
  OR2_X1 U8764 ( .A1(n10476), .A2(n10475), .ZN(n10490) );
  NOR2_X1 U8765 ( .A1(n10490), .A2(n15034), .ZN(n10507) );
  INV_X1 U8766 ( .A(n14819), .ZN(n8274) );
  NAND4_X2 U8767 ( .A1(n10237), .A2(n10235), .A3(n10236), .A4(n10238), .ZN(
        n11134) );
  OR2_X1 U8768 ( .A1(n10691), .A2(n15457), .ZN(n10235) );
  AOI21_X1 U8769 ( .B1(n15114), .B2(n15113), .A(n15112), .ZN(n15111) );
  NOR2_X1 U8770 ( .A1(n11354), .A2(n11355), .ZN(n11353) );
  AOI21_X1 U8771 ( .B1(n11347), .B2(P1_REG1_REG_10__SCAN_IN), .A(n11353), .ZN(
        n11337) );
  XNOR2_X1 U8772 ( .A(n12804), .B(n12805), .ZN(n12626) );
  NAND2_X1 U8773 ( .A1(n10718), .A2(n10717), .ZN(n15171) );
  INV_X1 U8774 ( .A(n15204), .ZN(n15226) );
  NAND2_X1 U8775 ( .A1(n15258), .A2(n7602), .ZN(n15240) );
  OAI22_X1 U8776 ( .A1(n15271), .A2(n15199), .B1(n8174), .B2(n15290), .ZN(
        n15260) );
  NAND2_X1 U8777 ( .A1(n15287), .A2(n7765), .ZN(n15271) );
  OR2_X1 U8778 ( .A1(n15509), .A2(n15198), .ZN(n7765) );
  INV_X1 U8779 ( .A(n10616), .ZN(n10617) );
  OAI21_X1 U8780 ( .B1(n15318), .B2(n8432), .A(n7766), .ZN(n15289) );
  NAND2_X1 U8781 ( .A1(n8434), .A2(n8436), .ZN(n8432) );
  NAND2_X1 U8782 ( .A1(n8430), .A2(n8434), .ZN(n7766) );
  NAND2_X1 U8783 ( .A1(n15517), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U8784 ( .A1(n15289), .A2(n15288), .ZN(n15287) );
  NAND2_X1 U8785 ( .A1(n8182), .A2(n8181), .ZN(n15336) );
  INV_X1 U8786 ( .A(n8182), .ZN(n15354) );
  NAND2_X1 U8787 ( .A1(n8184), .A2(n8183), .ZN(n15368) );
  INV_X1 U8788 ( .A(n8184), .ZN(n15392) );
  NOR2_X1 U8789 ( .A1(n15382), .A2(n8451), .ZN(n8450) );
  INV_X1 U8790 ( .A(n15192), .ZN(n8451) );
  NAND2_X1 U8791 ( .A1(n15401), .A2(n15192), .ZN(n15383) );
  NAND2_X1 U8792 ( .A1(n15190), .A2(n15189), .ZN(n15402) );
  AND2_X1 U8793 ( .A1(n8439), .A2(n15421), .ZN(n8437) );
  NAND2_X1 U8794 ( .A1(n15402), .A2(n15405), .ZN(n15401) );
  NOR2_X2 U8795 ( .A1(n15562), .A2(n15427), .ZN(n15426) );
  NOR2_X1 U8796 ( .A1(n15579), .A2(n8177), .ZN(n8176) );
  INV_X1 U8797 ( .A(n8178), .ZN(n8177) );
  AND2_X1 U8798 ( .A1(n8445), .A2(n12604), .ZN(n8444) );
  INV_X1 U8799 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10362) );
  OR2_X1 U8800 ( .A1(n10363), .A2(n10362), .ZN(n10380) );
  NAND2_X1 U8801 ( .A1(n12033), .A2(n12030), .ZN(n12091) );
  AND2_X1 U8802 ( .A1(n8483), .A2(n7458), .ZN(n12085) );
  NAND2_X1 U8803 ( .A1(n8423), .A2(n11892), .ZN(n11896) );
  NAND2_X1 U8804 ( .A1(n11887), .A2(n11886), .ZN(n12027) );
  NAND2_X1 U8805 ( .A1(n8171), .A2(n11696), .ZN(n11552) );
  INV_X1 U8806 ( .A(n11445), .ZN(n8171) );
  NAND2_X1 U8807 ( .A1(n11371), .A2(n11436), .ZN(n11445) );
  NAND2_X1 U8808 ( .A1(n11369), .A2(n11293), .ZN(n11438) );
  NAND2_X1 U8809 ( .A1(n11294), .A2(n15447), .ZN(n15446) );
  INV_X1 U8810 ( .A(n15451), .ZN(n15386) );
  INV_X1 U8811 ( .A(n11301), .ZN(n15445) );
  NAND2_X1 U8812 ( .A1(n7813), .A2(n12458), .ZN(n12459) );
  INV_X1 U8813 ( .A(n15461), .ZN(n16330) );
  INV_X1 U8814 ( .A(n15563), .ZN(n16437) );
  XNOR2_X1 U8815 ( .A(n9356), .B(n9355), .ZN(n14776) );
  XNOR2_X1 U8816 ( .A(n10264), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U8817 ( .A1(n8367), .A2(n9297), .ZN(n9642) );
  AND2_X1 U8818 ( .A1(n10470), .A2(n10483), .ZN(n12393) );
  XNOR2_X1 U8819 ( .A(n9577), .B(n9576), .ZN(n11182) );
  NAND2_X1 U8820 ( .A1(n9272), .A2(n9271), .ZN(n9537) );
  XNOR2_X1 U8821 ( .A(n9504), .B(n9503), .ZN(n10941) );
  NAND2_X1 U8822 ( .A1(n7992), .A2(n9266), .ZN(n9504) );
  NAND2_X1 U8823 ( .A1(n9489), .A2(n9264), .ZN(n7992) );
  NAND2_X1 U8824 ( .A1(n8355), .A2(n9261), .ZN(n9470) );
  NAND2_X1 U8825 ( .A1(n9449), .A2(n9259), .ZN(n8355) );
  INV_X1 U8826 ( .A(n9259), .ZN(n7763) );
  NAND2_X1 U8827 ( .A1(n9420), .A2(n9254), .ZN(n8363) );
  OR2_X1 U8828 ( .A1(n10409), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n10339) );
  XNOR2_X1 U8829 ( .A(n9420), .B(n9419), .ZN(n10837) );
  NAND2_X1 U8830 ( .A1(n9351), .A2(n9237), .ZN(n10268) );
  OAI21_X1 U8831 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n9091), .A(n9090), .ZN(
        n9121) );
  NOR2_X1 U8832 ( .A1(n9146), .A2(n9147), .ZN(n9149) );
  OAI21_X1 U8833 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n9102), .A(n9101), .ZN(
        n9112) );
  AOI22_X1 U8834 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n13127), .B1(n9159), .B2(
        n9104), .ZN(n9163) );
  AOI21_X1 U8835 ( .B1(n12638), .B2(n12585), .A(n8328), .ZN(n8327) );
  INV_X1 U8836 ( .A(n12587), .ZN(n8328) );
  NAND2_X1 U8837 ( .A1(n12635), .A2(n12585), .ZN(n12588) );
  NAND2_X1 U8838 ( .A1(n13285), .A2(n13284), .ZN(n13369) );
  NAND2_X1 U8839 ( .A1(n13402), .A2(n13224), .ZN(n13285) );
  AND2_X1 U8840 ( .A1(n13040), .A2(n13039), .ZN(n13042) );
  INV_X1 U8841 ( .A(n12145), .ZN(n12141) );
  NAND2_X1 U8842 ( .A1(n13423), .A2(n13241), .ZN(n13302) );
  AND2_X1 U8843 ( .A1(n16308), .A2(n11798), .ZN(n13197) );
  INV_X1 U8844 ( .A(n13483), .ZN(n7952) );
  AOI21_X1 U8845 ( .B1(n8336), .B2(n8339), .A(n7489), .ZN(n8335) );
  INV_X1 U8846 ( .A(n13284), .ZN(n8339) );
  CLKBUF_X1 U8847 ( .A(n12579), .Z(n12335) );
  INV_X1 U8848 ( .A(n13981), .ZN(n14007) );
  NAND2_X1 U8849 ( .A1(n12204), .A2(n12203), .ZN(n12207) );
  NAND2_X1 U8850 ( .A1(n13325), .A2(n12869), .ZN(n12872) );
  INV_X1 U8851 ( .A(n13993), .ZN(n13426) );
  AND3_X1 U8852 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n13936) );
  NAND2_X1 U8853 ( .A1(n13256), .A2(n8331), .ZN(n13413) );
  NAND2_X1 U8854 ( .A1(n8909), .A2(n8908), .ZN(n13419) );
  NAND2_X1 U8855 ( .A1(n13357), .A2(n13269), .ZN(n13433) );
  AND2_X1 U8856 ( .A1(n11805), .A2(n11804), .ZN(n13450) );
  NAND2_X1 U8857 ( .A1(n8966), .A2(n8965), .ZN(n13879) );
  NAND2_X1 U8858 ( .A1(n8949), .A2(n8948), .ZN(n13896) );
  INV_X1 U8859 ( .A(n13911), .ZN(n13880) );
  INV_X1 U8860 ( .A(n13921), .ZN(n13895) );
  NAND4_X1 U8861 ( .A1(n8617), .A2(n8616), .A3(n8615), .A4(n8614), .ZN(n13664)
         );
  NAND4_X1 U8862 ( .A1(n8604), .A2(n8603), .A3(n8602), .A4(n8601), .ZN(n13665)
         );
  NAND2_X1 U8863 ( .A1(n10810), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U8864 ( .A1(n8960), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7956) );
  NAND4_X1 U8865 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n8577), .ZN(n16312)
         );
  NOR2_X1 U8866 ( .A1(n11634), .A2(n7828), .ZN(n11487) );
  AND2_X1 U8867 ( .A1(n7829), .A2(n11509), .ZN(n7828) );
  INV_X1 U8868 ( .A(n7831), .ZN(n7829) );
  NAND2_X1 U8869 ( .A1(n14231), .A2(n8142), .ZN(n8141) );
  INV_X1 U8870 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8142) );
  INV_X1 U8871 ( .A(n13682), .ZN(n8144) );
  NAND2_X1 U8872 ( .A1(n13681), .A2(n8146), .ZN(n8145) );
  OR2_X1 U8873 ( .A1(n13682), .A2(n8147), .ZN(n8146) );
  AOI21_X1 U8874 ( .B1(n13669), .B2(n13667), .A(n13668), .ZN(n13671) );
  AND2_X1 U8875 ( .A1(n7850), .A2(n7849), .ZN(n11947) );
  INV_X1 U8876 ( .A(n11945), .ZN(n7849) );
  NAND2_X1 U8877 ( .A1(n7780), .A2(n7778), .ZN(n12248) );
  NOR2_X1 U8878 ( .A1(n12359), .A2(n7781), .ZN(n12362) );
  INV_X1 U8879 ( .A(n7780), .ZN(n7781) );
  NAND2_X1 U8880 ( .A1(n7834), .A2(n7839), .ZN(n16275) );
  NAND2_X1 U8881 ( .A1(n12366), .A2(n7841), .ZN(n7834) );
  OR2_X1 U8882 ( .A1(n12658), .A2(n12659), .ZN(n7845) );
  NOR2_X1 U8883 ( .A1(n12676), .A2(n12675), .ZN(n12895) );
  NOR2_X1 U8884 ( .A1(n16269), .A2(n7964), .ZN(n12676) );
  AND2_X1 U8885 ( .A1(n7853), .A2(n7852), .ZN(n13115) );
  NAND2_X1 U8886 ( .A1(n13110), .A2(n13111), .ZN(n7852) );
  NAND2_X1 U8887 ( .A1(n13115), .A2(n13114), .ZN(n13692) );
  INV_X1 U8888 ( .A(n16037), .ZN(n16292) );
  NOR2_X1 U8889 ( .A1(n13122), .A2(n8152), .ZN(n13123) );
  OR2_X1 U8890 ( .A1(n7448), .A2(n13724), .ZN(n13699) );
  AND2_X1 U8891 ( .A1(n8153), .A2(n8154), .ZN(n13723) );
  INV_X1 U8892 ( .A(n13724), .ZN(n8153) );
  INV_X1 U8893 ( .A(n7776), .ZN(n13738) );
  AND2_X1 U8894 ( .A1(n13720), .A2(n13719), .ZN(n7856) );
  NAND2_X1 U8895 ( .A1(n13722), .A2(n13721), .ZN(n13749) );
  OR2_X1 U8896 ( .A1(n13849), .A2(n8982), .ZN(n13867) );
  NAND2_X1 U8897 ( .A1(n8117), .A2(n8118), .ZN(n13919) );
  NAND2_X1 U8898 ( .A1(n8882), .A2(n8881), .ZN(n13972) );
  NAND2_X1 U8899 ( .A1(n7932), .A2(n13555), .ZN(n14038) );
  NAND2_X1 U8900 ( .A1(n8999), .A2(n7933), .ZN(n7932) );
  AND2_X1 U8901 ( .A1(n14044), .A2(n8793), .ZN(n14030) );
  NAND2_X1 U8902 ( .A1(n8999), .A2(n13552), .ZN(n14042) );
  NAND2_X1 U8903 ( .A1(n8768), .A2(n8767), .ZN(n16466) );
  NAND2_X1 U8904 ( .A1(n13000), .A2(n7941), .ZN(n7935) );
  NAND2_X1 U8905 ( .A1(n8732), .A2(n8731), .ZN(n13048) );
  NAND2_X1 U8906 ( .A1(n7943), .A2(n12999), .ZN(n14087) );
  NAND2_X1 U8907 ( .A1(n7945), .A2(n7944), .ZN(n7943) );
  AND2_X1 U8908 ( .A1(n16390), .A2(n16377), .ZN(n14039) );
  INV_X1 U8909 ( .A(n16348), .ZN(n16390) );
  INV_X1 U8910 ( .A(n14075), .ZN(n16384) );
  INV_X1 U8911 ( .A(n16339), .ZN(n16382) );
  INV_X1 U8912 ( .A(n16480), .ZN(n14106) );
  OAI21_X1 U8913 ( .B1(n13461), .B2(n13462), .A(n13464), .ZN(n16477) );
  INV_X1 U8914 ( .A(n13356), .ZN(n14179) );
  NAND2_X1 U8915 ( .A1(n13585), .A2(n13926), .ZN(n13908) );
  INV_X1 U8916 ( .A(n13257), .ZN(n14189) );
  AND2_X1 U8917 ( .A1(n8897), .A2(n8896), .ZN(n14195) );
  NAND2_X1 U8918 ( .A1(n8834), .A2(n8833), .ZN(n14211) );
  NAND2_X1 U8919 ( .A1(n8786), .A2(n8785), .ZN(n14219) );
  INV_X1 U8920 ( .A(n12586), .ZN(n12589) );
  AND3_X1 U8921 ( .A1(n8665), .A2(n8664), .A3(n8663), .ZN(n12646) );
  OAI21_X1 U8922 ( .B1(n13494), .B2(n7916), .A(n7915), .ZN(n12301) );
  AOI21_X1 U8923 ( .B1(n7919), .B2(n13628), .A(n7918), .ZN(n7915) );
  INV_X1 U8924 ( .A(n13628), .ZN(n7916) );
  OR2_X1 U8925 ( .A1(n8954), .A2(SI_4_), .ZN(n8622) );
  NAND2_X1 U8926 ( .A1(n12166), .A2(n13628), .ZN(n12168) );
  NAND2_X1 U8927 ( .A1(n13494), .A2(n13495), .ZN(n12166) );
  INV_X1 U8928 ( .A(n11919), .ZN(n11855) );
  INV_X1 U8929 ( .A(n13178), .ZN(n14227) );
  NAND2_X1 U8930 ( .A1(n11483), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13178) );
  NAND2_X1 U8931 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n15617), .ZN(n7681) );
  XNOR2_X1 U8932 ( .A(n13454), .B(n13455), .ZN(n13461) );
  INV_X1 U8933 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U8934 ( .A1(n14232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8520) );
  INV_X1 U8935 ( .A(SI_29_), .ZN(n15633) );
  NAND2_X1 U8936 ( .A1(n8521), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8522) );
  INV_X1 U8937 ( .A(SI_28_), .ZN(n15637) );
  INV_X1 U8938 ( .A(n9059), .ZN(n12917) );
  INV_X1 U8939 ( .A(SI_25_), .ZN(n15644) );
  XNOR2_X1 U8940 ( .A(n8938), .B(n8560), .ZN(n12750) );
  XNOR2_X1 U8941 ( .A(n9035), .B(n9034), .ZN(n12752) );
  XNOR2_X1 U8942 ( .A(n8926), .B(n7632), .ZN(n8927) );
  XNOR2_X1 U8943 ( .A(n7633), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n7632) );
  INV_X1 U8944 ( .A(n9048), .ZN(n14239) );
  NAND2_X1 U8945 ( .A1(n8974), .A2(n9024), .ZN(n12080) );
  INV_X1 U8946 ( .A(SI_20_), .ZN(n15839) );
  INV_X1 U8947 ( .A(SI_19_), .ZN(n11514) );
  XNOR2_X1 U8948 ( .A(n8866), .B(n8969), .ZN(n13837) );
  INV_X1 U8949 ( .A(SI_17_), .ZN(n15657) );
  NAND2_X1 U8950 ( .A1(n8211), .A2(n8552), .ZN(n8795) );
  NAND2_X1 U8951 ( .A1(n8781), .A2(n8780), .ZN(n8211) );
  INV_X1 U8952 ( .A(SI_14_), .ZN(n15851) );
  INV_X1 U8953 ( .A(SI_13_), .ZN(n15855) );
  INV_X1 U8954 ( .A(SI_12_), .ZN(n15856) );
  INV_X1 U8955 ( .A(SI_11_), .ZN(n15857) );
  INV_X1 U8956 ( .A(n8201), .ZN(n8724) );
  AOI21_X1 U8957 ( .B1(n8710), .B2(n8708), .A(n7449), .ZN(n8201) );
  AOI22_X1 U8958 ( .A1(n7788), .A2(n8619), .B1(n14231), .B2(n8618), .ZN(n7787)
         );
  NOR2_X1 U8959 ( .A1(n14231), .A2(n8618), .ZN(n7788) );
  NAND2_X1 U8960 ( .A1(n8219), .A2(n8534), .ZN(n8608) );
  AND2_X1 U8961 ( .A1(n11859), .A2(n11860), .ZN(n7702) );
  NAND2_X1 U8962 ( .A1(n14379), .A2(n14277), .ZN(n14304) );
  NAND2_X1 U8963 ( .A1(n8313), .A2(n8314), .ZN(n14294) );
  NAND2_X1 U8964 ( .A1(n7666), .A2(n7452), .ZN(n8313) );
  NAND2_X1 U8965 ( .A1(n12687), .A2(n12688), .ZN(n12773) );
  NAND2_X1 U8966 ( .A1(n12686), .A2(n12685), .ZN(n12687) );
  INV_X1 U8967 ( .A(n11385), .ZN(n8299) );
  NOR2_X1 U8968 ( .A1(n11156), .A2(n11414), .ZN(n8297) );
  AND2_X1 U8969 ( .A1(n7666), .A2(n14333), .ZN(n14336) );
  AND2_X1 U8970 ( .A1(n8320), .A2(n14267), .ZN(n8318) );
  NAND2_X1 U8971 ( .A1(n9756), .A2(n9755), .ZN(n14675) );
  NAND2_X1 U8972 ( .A1(n12221), .A2(n12222), .ZN(n12404) );
  NAND2_X1 U8973 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  AOI21_X1 U8974 ( .B1(n8311), .B2(n8310), .A(n7496), .ZN(n8309) );
  NAND2_X1 U8975 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  NAND2_X1 U8976 ( .A1(n12485), .A2(n12486), .ZN(n12686) );
  NAND2_X1 U8977 ( .A1(n11205), .A2(n11153), .ZN(n11216) );
  AND2_X1 U8978 ( .A1(n11166), .A2(n11165), .ZN(n14328) );
  NOR2_X1 U8979 ( .A1(n14336), .A2(n14248), .ZN(n14369) );
  NAND2_X1 U8980 ( .A1(n11203), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14373) );
  NAND2_X1 U8981 ( .A1(n11177), .A2(n16455), .ZN(n14375) );
  NAND2_X1 U8982 ( .A1(n13060), .A2(n13061), .ZN(n13151) );
  NAND2_X1 U8983 ( .A1(n13059), .A2(n13058), .ZN(n13060) );
  INV_X1 U8984 ( .A(n14377), .ZN(n14382) );
  INV_X1 U8985 ( .A(n7660), .ZN(n10217) );
  NAND2_X1 U8986 ( .A1(n9236), .A2(n9235), .ZN(n14457) );
  NAND2_X1 U8987 ( .A1(n9765), .A2(n9764), .ZN(n14523) );
  BUF_X1 U8988 ( .A(n9937), .Z(n14412) );
  NAND2_X1 U8989 ( .A1(n10115), .A2(n10114), .ZN(n14645) );
  AND2_X1 U8990 ( .A1(n8237), .A2(n7462), .ZN(n14468) );
  NAND2_X1 U8991 ( .A1(n8052), .A2(n9899), .ZN(n14473) );
  NAND2_X1 U8992 ( .A1(n14488), .A2(n14487), .ZN(n8052) );
  NAND2_X1 U8993 ( .A1(n8194), .A2(n9735), .ZN(n14521) );
  NAND2_X1 U8994 ( .A1(n14546), .A2(n14545), .ZN(n8194) );
  NAND2_X1 U8995 ( .A1(n8070), .A2(n9889), .ZN(n14565) );
  NAND2_X1 U8996 ( .A1(n14580), .A2(n9692), .ZN(n14564) );
  AND2_X1 U8997 ( .A1(n7641), .A2(n9668), .ZN(n14581) );
  NAND2_X1 U8998 ( .A1(n8057), .A2(n8055), .ZN(n14626) );
  NAND2_X1 U8999 ( .A1(n13088), .A2(n9640), .ZN(n14637) );
  NAND2_X1 U9000 ( .A1(n9634), .A2(n9633), .ZN(n14719) );
  AND2_X1 U9001 ( .A1(n13070), .A2(n9628), .ZN(n13090) );
  NAND2_X1 U9002 ( .A1(n12734), .A2(n9575), .ZN(n12782) );
  NAND2_X1 U9003 ( .A1(n8232), .A2(n8230), .ZN(n11840) );
  OR2_X1 U9004 ( .A1(n11471), .A2(n9447), .ZN(n8232) );
  NAND2_X1 U9005 ( .A1(n16458), .A2(n9919), .ZN(n14631) );
  INV_X1 U9006 ( .A(n14631), .ZN(n16463) );
  INV_X1 U9007 ( .A(n14561), .ZN(n16452) );
  INV_X1 U9008 ( .A(n14653), .ZN(n8079) );
  NOR2_X1 U9009 ( .A1(n14654), .A2(n8078), .ZN(n7732) );
  INV_X1 U9010 ( .A(n11160), .ZN(n16297) );
  AND2_X1 U9011 ( .A1(n11171), .A2(n9850), .ZN(n16041) );
  INV_X1 U9012 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9225) );
  INV_X1 U9013 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14777) );
  INV_X1 U9014 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U9015 ( .A1(n9829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U9016 ( .A1(n9829), .A2(n9825), .ZN(n13105) );
  OR2_X1 U9017 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  XNOR2_X1 U9018 ( .A(n9827), .B(n9826), .ZN(n13035) );
  NOR2_X1 U9019 ( .A1(n11171), .A2(P2_U3088), .ZN(n13024) );
  NAND2_X1 U9020 ( .A1(n9834), .A2(n7484), .ZN(n9838) );
  INV_X1 U9021 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9836) );
  INV_X1 U9022 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11825) );
  INV_X1 U9023 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11719) );
  INV_X1 U9024 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11562) );
  INV_X1 U9025 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11380) );
  INV_X1 U9026 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10990) );
  OR2_X1 U9027 ( .A1(n9475), .A2(n9474), .ZN(n16118) );
  INV_X1 U9028 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10879) );
  INV_X1 U9029 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10857) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10843) );
  INV_X1 U9031 ( .A(n8266), .ZN(n8264) );
  AOI21_X1 U9032 ( .B1(n8268), .B2(n8267), .A(n7467), .ZN(n8266) );
  AND2_X1 U9033 ( .A1(n11684), .A2(n11683), .ZN(n14913) );
  NAND2_X1 U9034 ( .A1(n10678), .A2(n10677), .ZN(n15483) );
  NAND2_X1 U9035 ( .A1(n7631), .A2(n11262), .ZN(n11141) );
  NAND2_X1 U9036 ( .A1(n7628), .A2(n7627), .ZN(n7631) );
  INV_X1 U9037 ( .A(n11137), .ZN(n7627) );
  INV_X1 U9038 ( .A(n11136), .ZN(n7628) );
  NAND2_X1 U9039 ( .A1(n11131), .A2(n11132), .ZN(n7617) );
  NAND2_X1 U9040 ( .A1(n14990), .A2(n8262), .ZN(n14946) );
  OR2_X1 U9041 ( .A1(n14864), .A2(n14865), .ZN(n8256) );
  NAND2_X1 U9042 ( .A1(n8280), .A2(n8281), .ZN(n14963) );
  INV_X1 U9043 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11736) );
  NAND2_X1 U9044 ( .A1(n14992), .A2(n14991), .ZN(n14990) );
  NAND2_X1 U9045 ( .A1(n12956), .A2(n7651), .ZN(n14803) );
  NAND2_X1 U9046 ( .A1(n7653), .A2(n7652), .ZN(n7651) );
  INV_X1 U9047 ( .A(n12958), .ZN(n7652) );
  INV_X1 U9048 ( .A(n12957), .ZN(n7653) );
  NAND2_X1 U9049 ( .A1(n8259), .A2(n7451), .ZN(n8258) );
  INV_X1 U9050 ( .A(n8260), .ZN(n8259) );
  INV_X1 U9051 ( .A(n15060), .ZN(n11291) );
  CLKBUF_X1 U9052 ( .A(n11264), .Z(n11265) );
  INV_X1 U9053 ( .A(n15042), .ZN(n15026) );
  AND2_X1 U9054 ( .A1(n11047), .A2(n11046), .ZN(n15029) );
  INV_X1 U9055 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15034) );
  NAND2_X1 U9056 ( .A1(n10502), .A2(n10501), .ZN(n15571) );
  NAND2_X1 U9057 ( .A1(n11047), .A2(n11036), .ZN(n15044) );
  NOR2_X1 U9058 ( .A1(n10767), .A2(n10770), .ZN(n10773) );
  NAND4_X1 U9059 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n15057) );
  AOI21_X1 U9060 ( .B1(n15117), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15111), .ZN(
        n10898) );
  AND2_X1 U9061 ( .A1(n11337), .A2(n11336), .ZN(n11607) );
  AND2_X1 U9062 ( .A1(n10697), .A2(n10696), .ZN(n15211) );
  NOR2_X1 U9063 ( .A1(n15234), .A2(n7812), .ZN(n15223) );
  XNOR2_X1 U9064 ( .A(n15215), .B(n15222), .ZN(n7601) );
  AND2_X1 U9065 ( .A1(n8378), .A2(n8377), .ZN(n15257) );
  NAND2_X1 U9066 ( .A1(n15284), .A2(n8379), .ZN(n15273) );
  AND2_X1 U9067 ( .A1(n7801), .A2(n7800), .ZN(n15286) );
  INV_X1 U9068 ( .A(n15517), .ZN(n15313) );
  NAND2_X1 U9069 ( .A1(n15322), .A2(n7802), .ZN(n15305) );
  INV_X1 U9070 ( .A(n7801), .ZN(n15304) );
  AOI21_X1 U9071 ( .B1(n15318), .B2(n15317), .A(n8433), .ZN(n15303) );
  NAND2_X1 U9072 ( .A1(n15630), .A2(n7723), .ZN(n15329) );
  NAND2_X1 U9073 ( .A1(n15351), .A2(n8476), .ZN(n15341) );
  AND2_X1 U9074 ( .A1(n7794), .A2(n7461), .ZN(n15366) );
  NAND2_X1 U9075 ( .A1(n15381), .A2(n15181), .ZN(n7794) );
  NAND2_X1 U9076 ( .A1(n10545), .A2(n10544), .ZN(n15396) );
  NAND2_X1 U9077 ( .A1(n8478), .A2(n7476), .ZN(n15552) );
  NAND2_X1 U9078 ( .A1(n8438), .A2(n8439), .ZN(n15422) );
  NAND2_X1 U9079 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  NAND2_X1 U9080 ( .A1(n12975), .A2(n12974), .ZN(n15188) );
  NAND2_X1 U9081 ( .A1(n12611), .A2(n16427), .ZN(n12612) );
  NAND2_X1 U9082 ( .A1(n12600), .A2(n12599), .ZN(n12602) );
  NAND2_X1 U9083 ( .A1(n12452), .A2(n12451), .ZN(n12605) );
  NAND2_X1 U9084 ( .A1(n12293), .A2(n8447), .ZN(n12452) );
  NAND2_X1 U9085 ( .A1(n12115), .A2(n12114), .ZN(n12117) );
  NAND2_X1 U9086 ( .A1(n8426), .A2(n11546), .ZN(n11894) );
  INV_X1 U9087 ( .A(n15434), .ZN(n15459) );
  INV_X1 U9088 ( .A(n15342), .ZN(n15425) );
  NAND2_X1 U9089 ( .A1(n11044), .A2(n15609), .ZN(n15428) );
  INV_X2 U9090 ( .A(n15356), .ZN(n15430) );
  NAND2_X1 U9091 ( .A1(n11055), .A2(n11056), .ZN(n15584) );
  NAND2_X1 U9092 ( .A1(n15491), .A2(n7469), .ZN(n15594) );
  OR2_X1 U9093 ( .A1(n15492), .A2(n16353), .ZN(n7604) );
  AND2_X1 U9094 ( .A1(n7513), .A2(n10231), .ZN(n8491) );
  INV_X1 U9095 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10231) );
  XNOR2_X1 U9096 ( .A(n10134), .B(n10133), .ZN(n10701) );
  XNOR2_X1 U9097 ( .A(n10782), .B(n10230), .ZN(n15628) );
  NAND2_X1 U9098 ( .A1(n7619), .A2(n7618), .ZN(n10780) );
  NAND2_X1 U9099 ( .A1(n7621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7618) );
  INV_X1 U9100 ( .A(n7620), .ZN(n7619) );
  NAND2_X1 U9101 ( .A1(n9738), .A2(n9737), .ZN(n9741) );
  XNOR2_X1 U9102 ( .A(n8380), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15630) );
  NAND2_X1 U9103 ( .A1(n10599), .A2(n10838), .ZN(n8380) );
  INV_X1 U9104 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11761) );
  INV_X1 U9105 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11564) );
  INV_X1 U9106 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11382) );
  INV_X1 U9107 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10942) );
  INV_X1 U9108 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10887) );
  INV_X1 U9109 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10881) );
  XNOR2_X1 U9110 ( .A(n10308), .B(n7858), .ZN(n15098) );
  NAND2_X1 U9111 ( .A1(n10244), .A2(n10243), .ZN(n15067) );
  NOR2_X1 U9112 ( .A1(n9132), .A2(n9131), .ZN(n16203) );
  NAND2_X1 U9113 ( .A1(n8025), .A2(n9139), .ZN(n16210) );
  AND2_X1 U9114 ( .A1(n9141), .A2(n9142), .ZN(n16250) );
  XNOR2_X1 U9115 ( .A(n9144), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n16215) );
  XNOR2_X1 U9116 ( .A(n9149), .B(n8036), .ZN(n16216) );
  INV_X1 U9117 ( .A(n9148), .ZN(n8036) );
  INV_X1 U9118 ( .A(n9154), .ZN(n8034) );
  OAI21_X1 U9119 ( .B1(n9157), .B2(n16192), .A(n16218), .ZN(n16223) );
  NOR2_X1 U9120 ( .A1(n16220), .A2(n16219), .ZN(n9157) );
  NOR2_X1 U9121 ( .A1(n16224), .A2(n16223), .ZN(n16222) );
  AND2_X1 U9122 ( .A1(n8028), .A2(n8026), .ZN(n16236) );
  AND2_X1 U9123 ( .A1(n8027), .A2(n8031), .ZN(n8026) );
  INV_X1 U9124 ( .A(n9167), .ZN(n8027) );
  NAND2_X1 U9125 ( .A1(n8028), .A2(n8031), .ZN(n9166) );
  NAND2_X1 U9126 ( .A1(n8040), .A2(n8039), .ZN(n16243) );
  NAND2_X1 U9127 ( .A1(n9175), .A2(n9176), .ZN(n8039) );
  NAND2_X1 U9128 ( .A1(n16031), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8040) );
  AND2_X1 U9129 ( .A1(n14227), .A2(n11577), .ZN(P3_U3897) );
  INV_X1 U9130 ( .A(n7669), .ZN(n7668) );
  OAI21_X1 U9131 ( .B1(n13280), .B2(n13453), .A(n13279), .ZN(n7669) );
  INV_X1 U9132 ( .A(n7853), .ZN(n13109) );
  INV_X1 U9133 ( .A(n13821), .ZN(n13814) );
  AOI21_X1 U9134 ( .B1(n8159), .B2(n13840), .A(n8155), .ZN(n13824) );
  AND2_X1 U9135 ( .A1(n7785), .A2(n7547), .ZN(n7662) );
  NAND2_X1 U9136 ( .A1(n10823), .A2(n7690), .ZN(P3_U3488) );
  NOR2_X1 U9137 ( .A1(n7443), .A2(n7542), .ZN(n7690) );
  AOI22_X1 U9138 ( .A1(n13866), .A2(n8133), .B1(P3_REG1_REG_28__SCAN_IN), .B2(
        n10822), .ZN(n8132) );
  NAND2_X1 U9139 ( .A1(n14168), .A2(n16473), .ZN(n8134) );
  OAI21_X1 U9140 ( .B1(n14171), .B2(n10822), .A(n7565), .ZN(n14114) );
  OR2_X1 U9141 ( .A1(n16473), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7565) );
  OAI21_X1 U9142 ( .B1(n14168), .B2(n16483), .A(n7957), .ZN(n14169) );
  NAND2_X1 U9143 ( .A1(n16483), .A2(n8987), .ZN(n7957) );
  NAND2_X1 U9144 ( .A1(n8302), .A2(n8305), .ZN(n11390) );
  OAI21_X1 U9145 ( .B1(n14651), .B2(n14598), .A(n9925), .ZN(n9926) );
  NAND2_X1 U9146 ( .A1(n8077), .A2(n8076), .ZN(P2_U3527) );
  NAND2_X1 U9147 ( .A1(n16412), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U9148 ( .A1(n14745), .A2(n16413), .ZN(n8077) );
  MUX2_X1 U9149 ( .A(n15159), .B(n15158), .S(n15157), .Z(n15161) );
  NAND2_X1 U9150 ( .A1(n15481), .A2(n15584), .ZN(n7775) );
  NAND2_X1 U9151 ( .A1(n16447), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8488) );
  OAI21_X1 U9152 ( .B1(n15481), .B2(n15480), .A(n8485), .ZN(n8487) );
  OAI222_X1 U9153 ( .A1(n7555), .A2(n7738), .B1(n15627), .B2(n13180), .C1(
        P1_U3086), .C2(n15073), .ZN(P1_U3327) );
  OAI222_X1 U9154 ( .A1(n7555), .A2(n15624), .B1(n15627), .B2(n15623), .C1(
        n15622), .C2(P1_U3086), .ZN(P1_U3328) );
  XNOR2_X1 U9155 ( .A(n9187), .B(n7655), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9156 ( .A(n9192), .B(n9186), .ZN(n7655) );
  NAND2_X4 U9157 ( .A1(n10720), .A2(n10282), .ZN(n10358) );
  AND2_X1 U9158 ( .A1(n8341), .A2(n8340), .ZN(n7439) );
  INV_X2 U9159 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n14231) );
  INV_X1 U9160 ( .A(n12761), .ZN(n8440) );
  INV_X1 U9161 ( .A(n11776), .ZN(n8149) );
  AOI21_X1 U9162 ( .B1(n13293), .B2(n13387), .A(n13386), .ZN(n13358) );
  OAI21_X2 U9163 ( .B1(n9421), .B2(n7554), .A(n7636), .ZN(n16298) );
  AND2_X1 U9164 ( .A1(n13419), .A2(n13657), .ZN(n7440) );
  XNOR2_X1 U9165 ( .A(n8520), .B(n8519), .ZN(n8523) );
  INV_X1 U9166 ( .A(n15528), .ZN(n8181) );
  AND4_X1 U9167 ( .A1(n15185), .A2(n10742), .A3(n15236), .A4(n15274), .ZN(
        n7441) );
  NAND2_X4 U9168 ( .A1(n11053), .A2(n11051), .ZN(n11130) );
  AND2_X1 U9169 ( .A1(n8280), .A2(n7536), .ZN(n7442) );
  NOR2_X1 U9170 ( .A1(n13188), .A2(n14164), .ZN(n7443) );
  NAND4_X1 U9171 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n15217) );
  AND3_X1 U9172 ( .A1(n7441), .A2(n7600), .A3(n10728), .ZN(n7444) );
  AND2_X1 U9173 ( .A1(n8518), .A2(n9036), .ZN(n7445) );
  NAND2_X1 U9174 ( .A1(n10003), .A2(n10004), .ZN(n7446) );
  AND2_X1 U9175 ( .A1(n13740), .A2(n13773), .ZN(n13766) );
  INV_X1 U9176 ( .A(n13766), .ZN(n8138) );
  INV_X1 U9177 ( .A(n10202), .ZN(n8066) );
  NAND2_X1 U9178 ( .A1(n8274), .A2(n14818), .ZN(n8281) );
  INV_X1 U9179 ( .A(n11694), .ZN(n11968) );
  OR2_X1 U9180 ( .A1(n9590), .A2(n7759), .ZN(n7447) );
  INV_X1 U9181 ( .A(n11888), .ZN(n7867) );
  INV_X1 U9182 ( .A(n11013), .ZN(n11695) );
  INV_X2 U9183 ( .A(n11695), .ZN(n14856) );
  AND2_X2 U9184 ( .A1(n11040), .A2(n11053), .ZN(n11013) );
  NAND2_X1 U9185 ( .A1(n13948), .A2(n8119), .ZN(n8117) );
  AND2_X1 U9186 ( .A1(n7439), .A2(n8725), .ZN(n8850) );
  AND2_X1 U9187 ( .A1(n13698), .A2(n13720), .ZN(n7448) );
  INV_X1 U9188 ( .A(n8428), .ZN(n15302) );
  XNOR2_X1 U9189 ( .A(n15517), .B(n15320), .ZN(n8428) );
  AND2_X1 U9190 ( .A1(n10942), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7449) );
  OR2_X1 U9191 ( .A1(n14189), .A2(n13936), .ZN(n7450) );
  OR2_X1 U9192 ( .A1(n14853), .A2(n14852), .ZN(n7451) );
  CLKBUF_X3 U9193 ( .A(n9959), .Z(n10153) );
  AND2_X1 U9194 ( .A1(n8317), .A2(n14333), .ZN(n7452) );
  NOR2_X1 U9195 ( .A1(n9885), .A2(n8061), .ZN(n8060) );
  NAND2_X1 U9196 ( .A1(n14728), .A2(n13157), .ZN(n7453) );
  AND2_X1 U9197 ( .A1(n13259), .A2(n13258), .ZN(n7454) );
  AND2_X1 U9198 ( .A1(n8808), .A2(n8793), .ZN(n7455) );
  OR2_X1 U9199 ( .A1(n11777), .A2(n11776), .ZN(n7456) );
  OR2_X1 U9200 ( .A1(n9705), .A2(n8222), .ZN(n7457) );
  NAND2_X1 U9201 ( .A1(n8726), .A2(n8513), .ZN(n8739) );
  INV_X1 U9202 ( .A(n9956), .ZN(n9959) );
  INV_X1 U9203 ( .A(n12999), .ZN(n7942) );
  OR2_X1 U9204 ( .A1(n12026), .A2(n12028), .ZN(n7458) );
  OR2_X1 U9205 ( .A1(n13766), .A2(n14035), .ZN(n7459) );
  OAI21_X1 U9206 ( .B1(n15309), .B2(n10690), .A(n10611), .ZN(n15320) );
  INV_X1 U9207 ( .A(n15320), .ZN(n8435) );
  NAND2_X1 U9208 ( .A1(n10562), .A2(n10561), .ZN(n15538) );
  INV_X1 U9209 ( .A(n15538), .ZN(n8183) );
  AND2_X1 U9210 ( .A1(n10094), .A2(n10093), .ZN(n7460) );
  NAND2_X1 U9211 ( .A1(n10325), .A2(n10324), .ZN(n11715) );
  XNOR2_X1 U9212 ( .A(n8008), .B(SI_4_), .ZN(n9419) );
  NAND2_X1 U9213 ( .A1(n10637), .A2(n10636), .ZN(n15501) );
  INV_X1 U9214 ( .A(n15501), .ZN(n8174) );
  INV_X1 U9215 ( .A(n14655), .ZN(n9796) );
  INV_X1 U9216 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10252) );
  INV_X1 U9217 ( .A(n10474), .ZN(n7911) );
  NAND2_X1 U9218 ( .A1(n15396), .A2(n15370), .ZN(n7461) );
  INV_X1 U9219 ( .A(n13534), .ZN(n7944) );
  INV_X1 U9220 ( .A(n10444), .ZN(n8398) );
  INV_X1 U9221 ( .A(n14964), .ZN(n8279) );
  INV_X1 U9222 ( .A(n13137), .ZN(n13632) );
  OR2_X1 U9223 ( .A1(n14664), .A2(n14395), .ZN(n7462) );
  AND3_X1 U9224 ( .A1(n9222), .A2(n9220), .A3(n9221), .ZN(n7463) );
  AND2_X1 U9225 ( .A1(n14664), .A2(n14459), .ZN(n7464) );
  NOR2_X1 U9226 ( .A1(n12505), .A2(n8269), .ZN(n8268) );
  INV_X1 U9227 ( .A(n12712), .ZN(n16427) );
  NAND2_X1 U9228 ( .A1(n10441), .A2(n10440), .ZN(n12712) );
  AND2_X1 U9229 ( .A1(n12990), .A2(n14399), .ZN(n7465) );
  AND2_X1 U9230 ( .A1(n12557), .A2(n12558), .ZN(n7467) );
  INV_X1 U9231 ( .A(n15489), .ZN(n15249) );
  AND2_X1 U9232 ( .A1(n15477), .A2(n16358), .ZN(n7468) );
  AND2_X1 U9233 ( .A1(n7604), .A2(n15490), .ZN(n7469) );
  AND2_X1 U9234 ( .A1(n11886), .A2(n8484), .ZN(n7470) );
  AND2_X1 U9235 ( .A1(n13387), .A2(n8344), .ZN(n7471) );
  AND2_X1 U9236 ( .A1(n13089), .A2(n9628), .ZN(n7472) );
  NOR2_X1 U9237 ( .A1(n14442), .A2(n14655), .ZN(n8163) );
  AND2_X1 U9238 ( .A1(n13253), .A2(n8332), .ZN(n7473) );
  AND2_X1 U9239 ( .A1(n12116), .A2(n12114), .ZN(n7474) );
  AND2_X1 U9240 ( .A1(n12205), .A2(n12203), .ZN(n7475) );
  AND2_X1 U9241 ( .A1(n15179), .A2(n15178), .ZN(n7476) );
  AND2_X1 U9242 ( .A1(n8070), .A2(n8068), .ZN(n7477) );
  AND2_X1 U9243 ( .A1(n12487), .A2(n12691), .ZN(n7478) );
  AND2_X1 U9244 ( .A1(n9277), .A2(n9271), .ZN(n7479) );
  INV_X1 U9245 ( .A(n8175), .ZN(n15294) );
  AND2_X1 U9246 ( .A1(n12461), .A2(n12458), .ZN(n7480) );
  INV_X1 U9247 ( .A(n12087), .ZN(n12119) );
  NAND2_X1 U9248 ( .A1(n13368), .A2(n13229), .ZN(n7481) );
  INV_X1 U9249 ( .A(n8477), .ZN(n8476) );
  AND2_X1 U9250 ( .A1(n8370), .A2(n15239), .ZN(n7482) );
  INV_X1 U9251 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9036) );
  INV_X1 U9252 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10241) );
  INV_X1 U9253 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7621) );
  INV_X1 U9254 ( .A(n8436), .ZN(n8433) );
  NAND2_X1 U9255 ( .A1(n15522), .A2(n15197), .ZN(n8436) );
  AND2_X1 U9256 ( .A1(n10178), .A2(n10177), .ZN(n7483) );
  NAND2_X1 U9257 ( .A1(n8008), .A2(SI_4_), .ZN(n9255) );
  AND2_X1 U9258 ( .A1(n8314), .A2(n8312), .ZN(n8311) );
  AND2_X1 U9259 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7484) );
  NOR2_X1 U9260 ( .A1(n15571), .A2(n15175), .ZN(n7485) );
  AND2_X1 U9261 ( .A1(n8429), .A2(n8431), .ZN(n7486) );
  NOR2_X1 U9262 ( .A1(n14714), .A2(n13156), .ZN(n7487) );
  NOR2_X1 U9263 ( .A1(n8779), .A2(n8778), .ZN(n7488) );
  NOR2_X1 U9264 ( .A1(n13232), .A2(n13231), .ZN(n7489) );
  INV_X1 U9265 ( .A(n12601), .ZN(n12715) );
  AND2_X1 U9266 ( .A1(n8994), .A2(n13527), .ZN(n7490) );
  INV_X1 U9267 ( .A(n10626), .ZN(n8390) );
  INV_X1 U9268 ( .A(n10429), .ZN(n7900) );
  MUX2_X1 U9269 ( .A(n15320), .B(n15517), .S(n10650), .Z(n10614) );
  AND2_X1 U9270 ( .A1(n12848), .A2(n12849), .ZN(n7491) );
  AND3_X1 U9271 ( .A1(n8043), .A2(n9425), .A3(n9427), .ZN(n7492) );
  AND2_X1 U9272 ( .A1(n7880), .A2(n7878), .ZN(n7493) );
  AND2_X1 U9273 ( .A1(n8452), .A2(n15405), .ZN(n7494) );
  AND2_X1 U9274 ( .A1(n7871), .A2(n7869), .ZN(n7495) );
  NOR2_X1 U9275 ( .A1(n14253), .A2(n14252), .ZN(n7496) );
  AND2_X1 U9276 ( .A1(n14991), .A2(n7451), .ZN(n7497) );
  AND2_X1 U9277 ( .A1(n8273), .A2(n8275), .ZN(n7498) );
  INV_X1 U9278 ( .A(n10414), .ZN(n8411) );
  AND2_X1 U9279 ( .A1(n9268), .A2(SI_9_), .ZN(n7499) );
  AND2_X1 U9280 ( .A1(n9263), .A2(SI_7_), .ZN(n7500) );
  NOR2_X1 U9281 ( .A1(n15571), .A2(n15186), .ZN(n7501) );
  INV_X1 U9282 ( .A(n13269), .ZN(n8348) );
  AND2_X1 U9283 ( .A1(n10076), .A2(n10075), .ZN(n7502) );
  OR2_X1 U9284 ( .A1(n7459), .A2(n13741), .ZN(n7503) );
  INV_X1 U9285 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U9286 ( .A1(n15489), .A2(n15200), .ZN(n7504) );
  INV_X1 U9287 ( .A(n8074), .ZN(n8073) );
  AND2_X1 U9288 ( .A1(n10843), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7505) );
  INV_X1 U9289 ( .A(n15421), .ZN(n15424) );
  OR2_X1 U9290 ( .A1(n8084), .A2(n8950), .ZN(n7506) );
  NOR2_X1 U9291 ( .A1(n13163), .A2(n14396), .ZN(n7507) );
  AND2_X1 U9292 ( .A1(n13387), .A2(n13264), .ZN(n7508) );
  INV_X1 U9293 ( .A(n8151), .ZN(n8152) );
  NAND2_X1 U9294 ( .A1(n12903), .A2(n12909), .ZN(n8151) );
  OR2_X1 U9295 ( .A1(n14964), .A2(n8278), .ZN(n7509) );
  NAND2_X1 U9296 ( .A1(n8108), .A2(n7450), .ZN(n13909) );
  INV_X1 U9297 ( .A(n15185), .ZN(n15222) );
  OR2_X1 U9298 ( .A1(n7502), .A2(n10078), .ZN(n7510) );
  OR2_X1 U9299 ( .A1(n15483), .A2(n15242), .ZN(n7511) );
  OR2_X1 U9300 ( .A1(n15227), .A2(n15242), .ZN(n7512) );
  INV_X1 U9301 ( .A(n10003), .ZN(n8471) );
  AND2_X1 U9302 ( .A1(n10239), .A2(n10241), .ZN(n7513) );
  OR2_X1 U9303 ( .A1(n15227), .A2(n15201), .ZN(n7514) );
  NOR2_X1 U9304 ( .A1(n15245), .A2(n15244), .ZN(n7515) );
  AND2_X1 U9305 ( .A1(n7503), .A2(n8138), .ZN(n7516) );
  AND2_X1 U9306 ( .A1(n8466), .A2(n10087), .ZN(n7517) );
  OR2_X1 U9307 ( .A1(n8450), .A2(n8449), .ZN(n7518) );
  AND2_X1 U9308 ( .A1(n12870), .A2(n12869), .ZN(n7519) );
  AND2_X1 U9309 ( .A1(n10602), .A2(n8384), .ZN(n7520) );
  AND2_X1 U9310 ( .A1(n12084), .A2(n7458), .ZN(n7521) );
  AND2_X1 U9311 ( .A1(n7732), .A2(n7731), .ZN(n7522) );
  AND2_X1 U9312 ( .A1(n14990), .A2(n8260), .ZN(n7523) );
  AND2_X1 U9313 ( .A1(n7819), .A2(n7773), .ZN(n7524) );
  INV_X1 U9314 ( .A(n10520), .ZN(n7875) );
  INV_X1 U9315 ( .A(n10579), .ZN(n7884) );
  INV_X1 U9316 ( .A(n8104), .ZN(n8103) );
  NOR2_X1 U9317 ( .A1(n8879), .A2(n8105), .ZN(n8104) );
  AND2_X1 U9318 ( .A1(n8466), .A2(n10091), .ZN(n7525) );
  NOR2_X1 U9319 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n8343) );
  OR2_X1 U9320 ( .A1(n8406), .A2(n10377), .ZN(n7526) );
  INV_X1 U9321 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n16023) );
  NOR2_X1 U9322 ( .A1(n10414), .A2(n10416), .ZN(n8412) );
  AND2_X1 U9323 ( .A1(n14664), .A2(n14395), .ZN(n7527) );
  NAND2_X1 U9324 ( .A1(n16234), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7528) );
  AND2_X1 U9325 ( .A1(n7960), .A2(n7959), .ZN(n7529) );
  NAND2_X1 U9326 ( .A1(n10040), .A2(n10041), .ZN(n7530) );
  NAND2_X1 U9327 ( .A1(n10171), .A2(n10172), .ZN(n7531) );
  INV_X1 U9328 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8564) );
  AND2_X1 U9329 ( .A1(n7513), .A2(n10230), .ZN(n7532) );
  NAND2_X1 U9330 ( .A1(n10027), .A2(n10028), .ZN(n7533) );
  INV_X1 U9331 ( .A(n8056), .ZN(n8055) );
  NAND2_X1 U9332 ( .A1(n8058), .A2(n9652), .ZN(n8056) );
  INV_X1 U9333 ( .A(n10356), .ZN(n7868) );
  NAND2_X1 U9334 ( .A1(n8592), .A2(n8324), .ZN(n8594) );
  INV_X1 U9335 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U9336 ( .A(n13484), .B(n7952), .ZN(n16307) );
  INV_X1 U9337 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U9338 ( .B1(n15003), .B2(n10690), .A(n10598), .ZN(n15333) );
  INV_X1 U9339 ( .A(n15333), .ZN(n15197) );
  NAND2_X1 U9340 ( .A1(n8998), .A2(n13548), .ZN(n14055) );
  NAND2_X1 U9341 ( .A1(n7815), .A2(n7814), .ZN(n15423) );
  NAND2_X1 U9342 ( .A1(n7935), .A2(n7938), .ZN(n13050) );
  INV_X1 U9343 ( .A(n14686), .ZN(n8165) );
  NAND2_X1 U9344 ( .A1(n8093), .A2(n8097), .ZN(n14056) );
  INV_X1 U9345 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8147) );
  INV_X1 U9346 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U9347 ( .A1(n8478), .A2(n15178), .ZN(n15404) );
  AND2_X1 U9348 ( .A1(n15401), .A2(n8450), .ZN(n7534) );
  NOR2_X1 U9349 ( .A1(n13347), .A2(n13348), .ZN(n7535) );
  INV_X1 U9350 ( .A(n8841), .ZN(n8842) );
  AND2_X1 U9351 ( .A1(n8281), .A2(n8279), .ZN(n7536) );
  INV_X1 U9352 ( .A(n7848), .ZN(n7847) );
  NOR2_X1 U9353 ( .A1(n12364), .A2(n12363), .ZN(n7848) );
  AND2_X1 U9354 ( .A1(n8091), .A2(n8092), .ZN(n7537) );
  AND2_X1 U9355 ( .A1(n10054), .A2(n10053), .ZN(n7538) );
  AND2_X1 U9356 ( .A1(n11564), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7539) );
  INV_X1 U9357 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n11128) );
  NOR2_X1 U9358 ( .A1(n13123), .A2(n13124), .ZN(n7540) );
  INV_X1 U9359 ( .A(n12659), .ZN(n16279) );
  INV_X1 U9360 ( .A(n9693), .ZN(n8364) );
  INV_X1 U9361 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7684) );
  INV_X1 U9362 ( .A(n16476), .ZN(n16483) );
  OAI21_X1 U9363 ( .B1(n14948), .B2(n10690), .A(n10586), .ZN(n15319) );
  INV_X1 U9364 ( .A(n12967), .ZN(n8179) );
  NAND2_X1 U9365 ( .A1(n9646), .A2(n9645), .ZN(n14714) );
  INV_X1 U9366 ( .A(n14714), .ZN(n8169) );
  NAND2_X1 U9367 ( .A1(n7813), .A2(n7480), .ZN(n12600) );
  INV_X1 U9368 ( .A(SI_6_), .ZN(n7764) );
  AND2_X1 U9369 ( .A1(n12611), .A2(n8178), .ZN(n7541) );
  AND2_X1 U9370 ( .A1(n10822), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7542) );
  INV_X1 U9371 ( .A(n13780), .ZN(n13794) );
  INV_X1 U9372 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8186) );
  INV_X1 U9373 ( .A(SI_18_), .ZN(n15843) );
  INV_X1 U9374 ( .A(n14704), .ZN(n8167) );
  NAND2_X1 U9375 ( .A1(n8850), .A2(n8518), .ZN(n9026) );
  NAND2_X1 U9376 ( .A1(n7809), .A2(n12086), .ZN(n12088) );
  AND2_X1 U9377 ( .A1(n12503), .A2(n8268), .ZN(n7543) );
  INV_X1 U9378 ( .A(n7941), .ZN(n7940) );
  NOR2_X1 U9379 ( .A1(n14088), .A2(n7942), .ZN(n7941) );
  INV_X1 U9380 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8245) );
  OR2_X1 U9381 ( .A1(n10104), .A2(SI_29_), .ZN(n7544) );
  NAND2_X1 U9382 ( .A1(n12293), .A2(n12292), .ZN(n7545) );
  INV_X1 U9383 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n12181) );
  AND2_X1 U9384 ( .A1(n8022), .A2(n10105), .ZN(n7546) );
  INV_X1 U9385 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12382) );
  INV_X1 U9386 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12733) );
  NOR2_X1 U9387 ( .A1(n13838), .A2(n13839), .ZN(n7547) );
  INV_X1 U9388 ( .A(n13767), .ZN(n8140) );
  AND2_X1 U9389 ( .A1(n8232), .A2(n9448), .ZN(n7548) );
  NAND2_X1 U9390 ( .A1(n13734), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7549) );
  INV_X1 U9391 ( .A(n13803), .ZN(n7977) );
  INV_X1 U9392 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7735) );
  INV_X1 U9393 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7719) );
  INV_X1 U9394 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7738) );
  INV_X1 U9395 ( .A(n12259), .ZN(n7598) );
  BUF_X1 U9396 ( .A(n9933), .Z(n14411) );
  INV_X1 U9397 ( .A(n14150), .ZN(n10820) );
  INV_X1 U9398 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7625) );
  AND2_X1 U9399 ( .A1(n11301), .A2(n16353), .ZN(n16425) );
  INV_X1 U9400 ( .A(n16425), .ZN(n15568) );
  OR2_X1 U9401 ( .A1(n11772), .A2(n11773), .ZN(n7850) );
  NAND2_X1 U9402 ( .A1(n13830), .A2(n13806), .ZN(n7550) );
  INV_X1 U9403 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13107) );
  INV_X1 U9404 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14782) );
  INV_X1 U9405 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12843) );
  OR2_X1 U9406 ( .A1(n13830), .A2(n13806), .ZN(n7551) );
  OR2_X1 U9407 ( .A1(n16425), .A2(n16447), .ZN(n7552) );
  INV_X1 U9408 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7633) );
  INV_X1 U9409 ( .A(n15625), .ZN(n7555) );
  INV_X1 U9410 ( .A(n13837), .ZN(n13829) );
  AND2_X1 U9411 ( .A1(n13681), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7553) );
  INV_X1 U9412 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14775) );
  XOR2_X1 U9413 ( .A(n9386), .B(n9385), .Z(n7554) );
  INV_X1 U9414 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8010) );
  INV_X1 U9415 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8359) );
  INV_X1 U9416 ( .A(n14164), .ZN(n8133) );
  AND2_X1 U9417 ( .A1(n11040), .A2(n10828), .ZN(n15609) );
  AND2_X1 U9418 ( .A1(n7434), .A2(P1_U3086), .ZN(n15625) );
  INV_X1 U9419 ( .A(n13193), .ZN(n13454) );
  NAND2_X1 U9420 ( .A1(n8533), .A2(n8532), .ZN(n8591) );
  NAND2_X1 U9421 ( .A1(n8696), .A2(n8695), .ZN(n8545) );
  NAND2_X1 U9422 ( .A1(n7739), .A2(n7737), .ZN(n13191) );
  NAND2_X1 U9423 ( .A1(n7609), .A2(n7608), .ZN(n8907) );
  OAI21_X1 U9424 ( .B1(n13615), .B2(n13614), .A(n13618), .ZN(n13616) );
  XNOR2_X1 U9425 ( .A(n7680), .B(n13457), .ZN(n14230) );
  NAND2_X1 U9426 ( .A1(n7564), .A2(n8548), .ZN(n8757) );
  INV_X1 U9427 ( .A(n10638), .ZN(n8407) );
  NAND2_X1 U9428 ( .A1(n9539), .A2(n9278), .ZN(n9553) );
  NAND2_X1 U9429 ( .A1(n7556), .A2(n8392), .ZN(n8391) );
  NAND2_X1 U9430 ( .A1(n10604), .A2(n7862), .ZN(n7556) );
  INV_X1 U9431 ( .A(P1_RD_REG_SCAN_IN), .ZN(n16294) );
  NAND2_X1 U9432 ( .A1(n9520), .A2(n9269), .ZN(n9272) );
  NAND2_X1 U9433 ( .A1(n9283), .A2(n7761), .ZN(n7760) );
  NAND2_X1 U9434 ( .A1(n7760), .A2(n9285), .ZN(n9591) );
  OAI21_X1 U9435 ( .B1(n10376), .B2(n8405), .A(n7526), .ZN(n10392) );
  NAND2_X1 U9436 ( .A1(n7588), .A2(n9248), .ZN(n9414) );
  OAI22_X1 U9437 ( .A1(n10564), .A2(n8417), .B1(n10565), .B2(n8416), .ZN(
        n10578) );
  OAI22_X1 U9438 ( .A1(n10504), .A2(n8415), .B1(n10505), .B2(n8414), .ZN(
        n10519) );
  NAND2_X1 U9439 ( .A1(n10313), .A2(n7559), .ZN(n8383) );
  INV_X2 U9440 ( .A(n10438), .ZN(n10229) );
  INV_X1 U9441 ( .A(n10438), .ZN(n10270) );
  NAND2_X1 U9442 ( .A1(n7582), .A2(n7633), .ZN(n7597) );
  OAI21_X1 U9443 ( .B1(n7889), .B2(n7893), .A(n7890), .ZN(n10443) );
  NAND2_X1 U9444 ( .A1(n7493), .A2(n10603), .ZN(n7862) );
  INV_X1 U9445 ( .A(n10591), .ZN(n8387) );
  NAND2_X1 U9446 ( .A1(n7866), .A2(n10357), .ZN(n7865) );
  NAND2_X1 U9447 ( .A1(n9314), .A2(SI_20_), .ZN(n9315) );
  NAND2_X1 U9448 ( .A1(n7990), .A2(n7991), .ZN(n9520) );
  INV_X1 U9449 ( .A(n7562), .ZN(n7561) );
  OAI21_X2 U9450 ( .B1(n13638), .B2(n13604), .A(n13603), .ZN(n7562) );
  OAI21_X1 U9451 ( .B1(n13638), .B2(n7659), .A(n7658), .ZN(n7563) );
  NAND2_X1 U9452 ( .A1(n8743), .A2(n8741), .ZN(n7564) );
  XNOR2_X1 U9453 ( .A(n8917), .B(n8918), .ZN(n12255) );
  NAND2_X1 U9454 ( .A1(n8112), .A2(n7450), .ZN(n8111) );
  INV_X1 U9455 ( .A(n8110), .ZN(n8109) );
  NAND2_X1 U9456 ( .A1(n7572), .A2(n7571), .ZN(n7742) );
  NAND2_X1 U9457 ( .A1(n7577), .A2(n7744), .ZN(n10036) );
  NAND2_X1 U9458 ( .A1(n7640), .A2(n7747), .ZN(n10046) );
  INV_X1 U9459 ( .A(n9991), .ZN(n7575) );
  NAND2_X1 U9460 ( .A1(n7566), .A2(n9942), .ZN(n9941) );
  NAND2_X1 U9461 ( .A1(n10189), .A2(n9936), .ZN(n7566) );
  NAND2_X1 U9462 ( .A1(n7711), .A2(n7708), .ZN(n10089) );
  NAND2_X1 U9463 ( .A1(n7576), .A2(n7575), .ZN(n7743) );
  NAND2_X1 U9464 ( .A1(n10046), .A2(n10045), .ZN(n7639) );
  AOI211_X1 U9465 ( .C1(n15759), .C2(n15758), .A(n15757), .B(n15756), .ZN(
        n15767) );
  OAI21_X1 U9466 ( .B1(n15660), .B2(n15659), .A(n15658), .ZN(n15663) );
  AOI21_X1 U9467 ( .B1(n15770), .B2(n15769), .A(n15768), .ZN(n7573) );
  AOI21_X1 U9468 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15739) );
  AOI211_X1 U9469 ( .C1(n15730), .C2(n15729), .A(n15728), .B(n15727), .ZN(
        n15733) );
  AOI211_X1 U9470 ( .C1(n15709), .C2(n15708), .A(n15707), .B(n15706), .ZN(
        n15712) );
  AOI211_X1 U9471 ( .C1(n15797), .C2(n15796), .A(n15795), .B(n15794), .ZN(
        n15804) );
  NOR3_X1 U9472 ( .A1(n15640), .A2(n15639), .A3(n15638), .ZN(n15643) );
  NOR3_X1 U9473 ( .A1(n15716), .A2(n15715), .A3(n15714), .ZN(n15719) );
  NOR3_X1 U9474 ( .A1(n15722), .A2(n15721), .A3(n15720), .ZN(n15726) );
  NOR3_X1 U9475 ( .A1(n15647), .A2(n15646), .A3(n15645), .ZN(n15650) );
  NOR4_X1 U9476 ( .A1(n15688), .A2(n15687), .A3(n15686), .A4(n15685), .ZN(
        n15691) );
  NOR4_X1 U9477 ( .A1(n15675), .A2(n15674), .A3(n15673), .A4(n15672), .ZN(
        n15678) );
  OAI21_X1 U9478 ( .B1(n7573), .B2(n15772), .A(n15771), .ZN(n15775) );
  NAND2_X1 U9479 ( .A1(n9993), .A2(n9992), .ZN(n7576) );
  NAND3_X1 U9480 ( .A1(n10024), .A2(n7533), .A3(n10023), .ZN(n7577) );
  NAND2_X1 U9481 ( .A1(n9937), .A2(n16298), .ZN(n10189) );
  NAND4_X1 U9482 ( .A1(n9382), .A2(n9384), .A3(n9381), .A4(n9383), .ZN(n9937)
         );
  NAND2_X1 U9483 ( .A1(n7579), .A2(n7578), .ZN(n7701) );
  NAND2_X1 U9484 ( .A1(n9978), .A2(n9977), .ZN(n7579) );
  NAND2_X1 U9485 ( .A1(n7581), .A2(n7580), .ZN(n7692) );
  NAND2_X1 U9486 ( .A1(n9988), .A2(n9987), .ZN(n7581) );
  NAND2_X1 U9487 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  INV_X1 U9488 ( .A(n13467), .ZN(n7687) );
  NAND2_X1 U9489 ( .A1(n7583), .A2(n7681), .ZN(n7680) );
  NAND2_X1 U9490 ( .A1(n13454), .A2(n13455), .ZN(n7583) );
  INV_X1 U9491 ( .A(n9391), .ZN(n7637) );
  NAND2_X1 U9492 ( .A1(n12142), .A2(n12141), .ZN(n12204) );
  AOI21_X2 U9493 ( .B1(n13221), .B2(n13220), .A(n13219), .ZN(n13404) );
  NAND2_X1 U9494 ( .A1(n8334), .A2(n8335), .ZN(n13371) );
  NAND2_X1 U9495 ( .A1(n12140), .A2(n12139), .ZN(n12144) );
  NAND2_X1 U9496 ( .A1(n13246), .A2(n13245), .ZN(n13396) );
  NAND2_X1 U9497 ( .A1(n13323), .A2(n7584), .ZN(n13275) );
  NAND2_X1 U9498 ( .A1(n7586), .A2(n7585), .ZN(n7584) );
  INV_X1 U9499 ( .A(n13273), .ZN(n7586) );
  NAND2_X1 U9500 ( .A1(n8992), .A2(n13507), .ZN(n12527) );
  OAI21_X1 U9501 ( .B1(n13946), .B2(n13577), .A(n13578), .ZN(n7946) );
  OAI21_X1 U9502 ( .B1(n13000), .B2(n7937), .A(n7936), .ZN(n8996) );
  NOR2_X1 U9503 ( .A1(n11150), .A2(n11151), .ZN(n11152) );
  NAND2_X1 U9504 ( .A1(n12774), .A2(n12775), .ZN(n12945) );
  AND2_X2 U9505 ( .A1(n13175), .A2(n9856), .ZN(n11148) );
  NOR2_X1 U9506 ( .A1(n11615), .A2(n11614), .ZN(n11862) );
  NAND2_X1 U9507 ( .A1(n7587), .A2(n9738), .ZN(n12844) );
  NAND2_X1 U9508 ( .A1(n9724), .A2(n9723), .ZN(n7587) );
  NAND2_X1 U9509 ( .A1(n9398), .A2(n9397), .ZN(n7588) );
  NAND3_X1 U9510 ( .A1(n16295), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7986) );
  OAI21_X2 U9511 ( .B1(n12343), .B2(n8074), .A(n8071), .ZN(n12737) );
  OAI21_X1 U9512 ( .B1(n13069), .B2(n8056), .A(n8053), .ZN(n14599) );
  NAND2_X1 U9513 ( .A1(n9897), .A2(n9896), .ZN(n14488) );
  NAND3_X1 U9514 ( .A1(n7593), .A2(n7825), .A3(n7662), .ZN(P3_U3201) );
  NAND2_X1 U9515 ( .A1(n13848), .A2(n13847), .ZN(n7593) );
  NAND3_X1 U9516 ( .A1(n8468), .A2(n7594), .A3(n7446), .ZN(n7733) );
  NAND2_X1 U9517 ( .A1(n7715), .A2(n7714), .ZN(n7594) );
  NOR2_X2 U9518 ( .A1(n12371), .A2(n12370), .ZN(n12374) );
  NAND2_X1 U9519 ( .A1(n8593), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n8143) );
  NOR2_X1 U9520 ( .A1(n13762), .A2(n13763), .ZN(n13765) );
  XNOR2_X1 U9521 ( .A(n13815), .B(n7977), .ZN(n13784) );
  NAND2_X1 U9522 ( .A1(n7976), .A2(n7975), .ZN(n7974) );
  NAND2_X1 U9523 ( .A1(n8047), .A2(n8050), .ZN(n14456) );
  OAI21_X1 U9524 ( .B1(n9872), .B2(n16370), .A(n14404), .ZN(n8046) );
  NAND2_X1 U9525 ( .A1(n7707), .A2(n7706), .ZN(n13703) );
  AOI21_X1 U9526 ( .B1(n10700), .B2(n10699), .A(n10698), .ZN(n10761) );
  NAND3_X1 U9527 ( .A1(n7861), .A2(n10604), .A3(n7862), .ZN(n7643) );
  OAI22_X1 U9528 ( .A1(n12878), .A2(n9883), .B1(n12955), .B2(n14398), .ZN(
        n13069) );
  OAI21_X1 U9529 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15139) );
  OAI21_X1 U9530 ( .B1(n10999), .B2(n10997), .A(n10998), .ZN(n11334) );
  NOR2_X1 U9531 ( .A1(n10928), .A2(n10929), .ZN(n10949) );
  NOR2_X1 U9532 ( .A1(n11813), .A2(n11812), .ZN(n12392) );
  NOR2_X1 U9533 ( .A1(n10967), .A2(n10966), .ZN(n10965) );
  NOR2_X1 U9534 ( .A1(n12807), .A2(n12806), .ZN(n12810) );
  OAI22_X1 U9535 ( .A1(n12625), .A2(n12624), .B1(n12623), .B2(n12622), .ZN(
        n12804) );
  INV_X2 U9536 ( .A(n14254), .ZN(n14306) );
  XNOR2_X1 U9537 ( .A(n14242), .B(n11279), .ZN(n11154) );
  NOR2_X2 U9538 ( .A1(n11419), .A2(n11418), .ZN(n11615) );
  NAND2_X1 U9539 ( .A1(n13152), .A2(n13153), .ZN(n14245) );
  NAND2_X1 U9540 ( .A1(n8287), .A2(n8290), .ZN(n13152) );
  AOI21_X1 U9541 ( .B1(n11862), .B2(n11861), .A(n7702), .ZN(n11866) );
  NOR2_X1 U9542 ( .A1(n11152), .A2(n7595), .ZN(n11206) );
  NAND2_X1 U9543 ( .A1(n8895), .A2(n8893), .ZN(n7609) );
  NAND2_X1 U9544 ( .A1(n8559), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7596) );
  NOR2_X2 U9545 ( .A1(n12107), .A2(n12400), .ZN(n12349) );
  AOI21_X1 U9547 ( .B1(n7697), .B2(n16374), .A(n7696), .ZN(n7695) );
  NAND2_X1 U9548 ( .A1(n12405), .A2(n12406), .ZN(n12484) );
  AOI21_X2 U9549 ( .B1(n7601), .B2(n15584), .A(n15220), .ZN(n15486) );
  INV_X1 U9550 ( .A(n15482), .ZN(n7774) );
  INV_X1 U9551 ( .A(n7771), .ZN(n7770) );
  NOR2_X1 U9552 ( .A1(n15185), .A2(n7812), .ZN(n7810) );
  NAND2_X1 U9553 ( .A1(n7775), .A2(n7524), .ZN(n15592) );
  AOI21_X1 U9554 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n8461) );
  NOR4_X1 U9555 ( .A1(n15743), .A2(n15742), .A3(n15741), .A4(n15740), .ZN(
        n15749) );
  NAND2_X1 U9556 ( .A1(n8438), .A2(n8437), .ZN(n15190) );
  NAND2_X1 U9557 ( .A1(n7607), .A2(n8003), .ZN(n7998) );
  NAND2_X1 U9558 ( .A1(n8000), .A2(n7999), .ZN(n7607) );
  NAND2_X1 U9559 ( .A1(n9327), .A2(n9326), .ZN(n9768) );
  INV_X1 U9560 ( .A(n8357), .ZN(n8356) );
  NAND2_X1 U9561 ( .A1(n8024), .A2(n9338), .ZN(n9799) );
  NAND2_X1 U9562 ( .A1(n10791), .A2(n10792), .ZN(n10793) );
  NAND2_X1 U9563 ( .A1(n7675), .A2(n7672), .ZN(n9988) );
  NAND2_X1 U9564 ( .A1(n7729), .A2(n7726), .ZN(n9978) );
  OAI21_X1 U9565 ( .B1(n7615), .B2(n8461), .A(n7614), .ZN(n10213) );
  NAND2_X1 U9566 ( .A1(n7613), .A2(n7610), .ZN(n10051) );
  OAI21_X1 U9567 ( .B1(n10103), .B2(n10102), .A(n8458), .ZN(n7615) );
  NAND4_X2 U9568 ( .A1(n9372), .A2(n9371), .A3(n9370), .A4(n9369), .ZN(n9933)
         );
  NAND2_X1 U9569 ( .A1(n15009), .A2(n7703), .ZN(n14924) );
  NOR2_X2 U9570 ( .A1(n12847), .A2(n7491), .ZN(n12854) );
  NAND2_X1 U9571 ( .A1(n7630), .A2(n7629), .ZN(n14903) );
  AOI21_X2 U9572 ( .B1(n14924), .B2(n14921), .A(n14920), .ZN(n14992) );
  NAND4_X2 U9573 ( .A1(n10407), .A2(n7803), .A3(n10293), .A4(n10408), .ZN(
        n10438) );
  INV_X1 U9574 ( .A(n10777), .ZN(n7626) );
  AOI21_X2 U9575 ( .B1(n14317), .B2(n14316), .A(n7622), .ZN(n14264) );
  NAND2_X1 U9576 ( .A1(n9627), .A2(n9626), .ZN(n13070) );
  NAND2_X1 U9577 ( .A1(n9779), .A2(n9778), .ZN(n14482) );
  NAND2_X1 U9578 ( .A1(n8205), .A2(n8204), .ZN(n12884) );
  INV_X1 U9579 ( .A(n7907), .ZN(n7906) );
  NAND2_X1 U9580 ( .A1(n10653), .A2(n10654), .ZN(n10652) );
  NAND2_X1 U9581 ( .A1(n10681), .A2(n10682), .ZN(n10680) );
  NAND2_X1 U9582 ( .A1(n11275), .A2(n11274), .ZN(n9405) );
  INV_X1 U9583 ( .A(n14905), .ZN(n7630) );
  NAND2_X1 U9584 ( .A1(n12854), .A2(n12853), .ZN(n12956) );
  OAI22_X2 U9585 ( .A1(n12704), .A2(n12703), .B1(n12702), .B2(n12701), .ZN(
        n12705) );
  NAND4_X2 U9586 ( .A1(n10269), .A2(n10229), .A3(n10228), .A4(n10230), .ZN(
        n10240) );
  NAND2_X1 U9587 ( .A1(n7649), .A2(n7648), .ZN(n8265) );
  INV_X1 U9588 ( .A(n11141), .ZN(n11139) );
  NAND2_X1 U9589 ( .A1(n12189), .A2(n12188), .ZN(n7649) );
  INV_X1 U9590 ( .A(n10240), .ZN(n8492) );
  AND3_X2 U9591 ( .A1(n15793), .A2(n15806), .A3(n15805), .ZN(n7803) );
  NAND2_X1 U9592 ( .A1(n13638), .A2(n13599), .ZN(n7658) );
  NAND2_X1 U9593 ( .A1(n13616), .A2(n13639), .ZN(n13644) );
  NAND2_X1 U9594 ( .A1(n7722), .A2(n8558), .ZN(n8895) );
  NAND2_X1 U9595 ( .A1(n13865), .A2(n13864), .ZN(n13863) );
  NAND2_X1 U9596 ( .A1(n13469), .A2(n13468), .ZN(n7686) );
  OAI21_X1 U9597 ( .B1(n7921), .B2(n13585), .A(n13588), .ZN(n7689) );
  NAND2_X1 U9598 ( .A1(n7634), .A2(n8536), .ZN(n8639) );
  NAND2_X1 U9599 ( .A1(n8621), .A2(n8620), .ZN(n7634) );
  NAND2_X1 U9600 ( .A1(n10013), .A2(n10012), .ZN(n10019) );
  NAND2_X1 U9601 ( .A1(n10068), .A2(n10067), .ZN(n10074) );
  OAI21_X1 U9602 ( .B1(n10051), .B2(n10052), .A(n8456), .ZN(n8454) );
  OAI21_X1 U9603 ( .B1(n7676), .B2(n10072), .A(n8462), .ZN(n10083) );
  NAND2_X1 U9604 ( .A1(n9844), .A2(n9847), .ZN(n7725) );
  INV_X1 U9605 ( .A(n16298), .ZN(n7635) );
  NAND2_X1 U9606 ( .A1(n7645), .A2(n7644), .ZN(n8501) );
  NAND3_X1 U9607 ( .A1(n10037), .A2(n8501), .A3(n7530), .ZN(n7640) );
  NAND3_X1 U9608 ( .A1(n7730), .A2(n8248), .A3(n8250), .ZN(n9344) );
  NOR2_X2 U9609 ( .A1(n9212), .A2(n9422), .ZN(n8250) );
  NAND2_X1 U9610 ( .A1(n7692), .A2(n7691), .ZN(n9993) );
  INV_X1 U9611 ( .A(n11250), .ZN(n10191) );
  INV_X1 U9612 ( .A(n14652), .ZN(n7697) );
  NAND2_X1 U9613 ( .A1(n12583), .A2(n12582), .ZN(n12637) );
  NAND2_X1 U9614 ( .A1(n8412), .A2(n7894), .ZN(n7892) );
  AOI21_X1 U9615 ( .B1(n14456), .B2(n14455), .A(n7647), .ZN(n14448) );
  NOR2_X2 U9616 ( .A1(n14412), .A2(n16298), .ZN(n11223) );
  NAND3_X1 U9617 ( .A1(n9873), .A2(n16370), .A3(n9872), .ZN(n8044) );
  NAND2_X1 U9618 ( .A1(n13423), .A2(n8325), .ZN(n13300) );
  NAND2_X1 U9619 ( .A1(n13325), .A2(n7519), .ZN(n13040) );
  NAND2_X1 U9620 ( .A1(n12204), .A2(n7475), .ZN(n12334) );
  NOR2_X2 U9621 ( .A1(n7454), .A2(n13260), .ZN(n13294) );
  NOR2_X2 U9622 ( .A1(n13259), .A2(n13258), .ZN(n13260) );
  INV_X1 U9623 ( .A(n12208), .ZN(n12205) );
  NAND2_X1 U9624 ( .A1(n8345), .A2(n8346), .ZN(n13432) );
  AOI21_X1 U9625 ( .B1(n13647), .B2(n13646), .A(n7654), .ZN(n13654) );
  OAI211_X1 U9626 ( .C1(n8242), .C2(n8241), .A(n8239), .B(n8240), .ZN(n7654)
         );
  NAND2_X2 U9627 ( .A1(n8956), .A2(n8955), .ZN(n13874) );
  XNOR2_X1 U9628 ( .A(n16030), .B(n7677), .ZN(SUB_1596_U64) );
  NOR2_X1 U9629 ( .A1(n16206), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n9137) );
  XNOR2_X1 U9630 ( .A(n9136), .B(n9135), .ZN(n16206) );
  NOR2_X2 U9631 ( .A1(n9143), .A2(n16249), .ZN(n9144) );
  XNOR2_X1 U9632 ( .A(n9153), .B(n8034), .ZN(n16217) );
  OAI21_X1 U9633 ( .B1(n16227), .B2(n9161), .A(n7528), .ZN(n8030) );
  NAND2_X1 U9634 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  NAND2_X1 U9635 ( .A1(n7733), .A2(n8469), .ZN(n10011) );
  OAI21_X1 U9636 ( .B1(n10074), .B2(n10073), .A(n7510), .ZN(n7676) );
  AOI21_X1 U9637 ( .B1(n10051), .B2(n10052), .A(n7656), .ZN(n8453) );
  OAI21_X1 U9638 ( .B1(n8045), .B2(n8046), .A(n8044), .ZN(n12101) );
  NAND2_X1 U9639 ( .A1(n9863), .A2(n9862), .ZN(n11251) );
  NAND2_X1 U9640 ( .A1(n11487), .A2(n16262), .ZN(n11641) );
  NAND2_X1 U9641 ( .A1(n7826), .A2(n13830), .ZN(n7824) );
  OAI21_X1 U9642 ( .B1(n11654), .B2(n11653), .A(n11652), .ZN(n13669) );
  NOR2_X1 U9643 ( .A1(n13671), .A2(n7851), .ZN(n11772) );
  NAND2_X1 U9644 ( .A1(n16273), .A2(n7845), .ZN(n12660) );
  NOR2_X1 U9645 ( .A1(n13718), .A2(n7856), .ZN(n13722) );
  NOR2_X1 U9646 ( .A1(n12889), .A2(n7854), .ZN(n12893) );
  NAND2_X1 U9647 ( .A1(n13196), .A2(n13197), .ZN(n13195) );
  NAND2_X1 U9648 ( .A1(n13396), .A2(n13248), .ZN(n13337) );
  NAND3_X1 U9649 ( .A1(n8362), .A2(n9256), .A3(n7665), .ZN(n7664) );
  NOR2_X2 U9650 ( .A1(n14353), .A2(n14352), .ZN(n14351) );
  INV_X1 U9651 ( .A(n14293), .ZN(n8312) );
  AOI21_X2 U9652 ( .B1(n14327), .B2(n14326), .A(n7667), .ZN(n14380) );
  NAND2_X1 U9653 ( .A1(n11401), .A2(n11752), .ZN(n11477) );
  INV_X2 U9654 ( .A(n12000), .ZN(n11211) );
  INV_X1 U9655 ( .A(n14650), .ZN(n7696) );
  NAND2_X1 U9656 ( .A1(n14651), .A2(n7695), .ZN(n14744) );
  NAND2_X1 U9657 ( .A1(n14245), .A2(n14244), .ZN(n14334) );
  INV_X1 U9658 ( .A(n14334), .ZN(n7671) );
  NAND2_X1 U9659 ( .A1(n7671), .A2(n8311), .ZN(n8308) );
  OAI22_X2 U9660 ( .A1(n14343), .A2(n14342), .B1(n14270), .B2(n14269), .ZN(
        n14327) );
  NAND2_X1 U9661 ( .A1(n7670), .A2(n7668), .ZN(P3_U3154) );
  NAND2_X1 U9662 ( .A1(n13275), .A2(n13442), .ZN(n7670) );
  NAND2_X1 U9663 ( .A1(n8329), .A2(n8327), .ZN(n12866) );
  NOR2_X1 U9664 ( .A1(n8298), .A2(n11389), .ZN(n8301) );
  OAI21_X2 U9665 ( .B1(n9386), .B2(n9385), .A(n10268), .ZN(n9373) );
  INV_X1 U9666 ( .A(n8393), .ZN(n7861) );
  INV_X1 U9667 ( .A(n10011), .ZN(n7713) );
  NAND2_X1 U9668 ( .A1(n9968), .A2(n9967), .ZN(n9973) );
  NAND2_X1 U9669 ( .A1(n7674), .A2(n7673), .ZN(n7672) );
  INV_X1 U9670 ( .A(n9983), .ZN(n7674) );
  NAND2_X1 U9671 ( .A1(n7694), .A2(n7693), .ZN(n7675) );
  INV_X1 U9672 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U9673 ( .A1(n8757), .A2(n8755), .ZN(n7679) );
  NAND2_X1 U9674 ( .A1(n10799), .A2(n10800), .ZN(n7739) );
  NAND2_X1 U9675 ( .A1(n16480), .A2(n13851), .ZN(n8253) );
  NAND2_X1 U9676 ( .A1(n8951), .A2(n8952), .ZN(n7736) );
  NAND2_X1 U9677 ( .A1(n8215), .A2(n8217), .ZN(n8621) );
  NAND4_X1 U9678 ( .A1(n13640), .A2(n13618), .A3(n13639), .A4(n7682), .ZN(
        n13641) );
  AND2_X1 U9679 ( .A1(n8607), .A2(n8590), .ZN(n8216) );
  INV_X1 U9680 ( .A(n9981), .ZN(n7693) );
  NAND2_X1 U9681 ( .A1(n8198), .A2(n8202), .ZN(n7688) );
  NAND2_X1 U9682 ( .A1(n8907), .A2(n8905), .ZN(n8246) );
  NAND2_X1 U9683 ( .A1(n8292), .A2(n8295), .ZN(n12405) );
  NAND2_X1 U9684 ( .A1(n8282), .A2(n8285), .ZN(n12774) );
  NAND2_X1 U9685 ( .A1(n13910), .A2(n7922), .ZN(n7921) );
  INV_X1 U9686 ( .A(n7921), .ZN(n7920) );
  INV_X1 U9687 ( .A(n7951), .ZN(n9014) );
  OAI21_X1 U9688 ( .B1(n10824), .B2(n16483), .A(n10825), .ZN(n10826) );
  NAND2_X1 U9689 ( .A1(n9983), .A2(n9982), .ZN(n7694) );
  NAND2_X1 U9690 ( .A1(n11251), .A2(n11250), .ZN(n9865) );
  XNOR2_X2 U9691 ( .A(n7698), .B(n11995), .ZN(n11250) );
  INV_X1 U9692 ( .A(n9239), .ZN(n9244) );
  XNOR2_X1 U9693 ( .A(n9902), .B(n9901), .ZN(n9916) );
  NAND2_X1 U9694 ( .A1(n9243), .A2(n7699), .ZN(n9238) );
  NAND2_X1 U9695 ( .A1(n9374), .A2(n9373), .ZN(n7699) );
  NAND2_X1 U9696 ( .A1(n8079), .A2(n7522), .ZN(n14745) );
  OAI21_X1 U9697 ( .B1(n12344), .B2(n9534), .A(n9535), .ZN(n12318) );
  NAND2_X1 U9698 ( .A1(n9388), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U9699 ( .A1(n7701), .A2(n7700), .ZN(n9983) );
  NAND2_X1 U9700 ( .A1(n7713), .A2(n7712), .ZN(n10012) );
  NAND2_X4 U9701 ( .A1(n10234), .A2(n10257), .ZN(n10690) );
  OAI21_X1 U9702 ( .B1(n12293), .B2(n8446), .A(n8444), .ZN(n12607) );
  NAND2_X1 U9703 ( .A1(n11264), .A2(n11266), .ZN(n11684) );
  NAND2_X1 U9704 ( .A1(n8492), .A2(n8491), .ZN(n15613) );
  AOI22_X1 U9705 ( .A1(n15364), .A2(n15194), .B1(n15193), .B2(n15538), .ZN(
        n15346) );
  INV_X1 U9706 ( .A(n8420), .ZN(n15215) );
  OAI21_X2 U9707 ( .B1(n12759), .B2(n12758), .A(n12760), .ZN(n12762) );
  NAND2_X1 U9708 ( .A1(n7963), .A2(n11776), .ZN(n7962) );
  NAND2_X1 U9709 ( .A1(n11626), .A2(n11625), .ZN(n11627) );
  INV_X1 U9710 ( .A(n7704), .ZN(n7967) );
  OAI21_X1 U9711 ( .B1(n12374), .B2(n7970), .A(n7705), .ZN(n7704) );
  NAND2_X1 U9712 ( .A1(n11953), .A2(n11951), .ZN(n11949) );
  NAND2_X1 U9713 ( .A1(n7974), .A2(n7549), .ZN(n13736) );
  NOR2_X1 U9714 ( .A1(n13703), .A2(n16472), .ZN(n13712) );
  NAND2_X1 U9715 ( .A1(n13702), .A2(n13720), .ZN(n7706) );
  INV_X1 U9716 ( .A(n13713), .ZN(n7707) );
  NAND2_X1 U9717 ( .A1(n13116), .A2(n7979), .ZN(n12897) );
  INV_X1 U9718 ( .A(n13202), .ZN(n13483) );
  NAND4_X1 U9719 ( .A1(n7439), .A2(n7445), .A3(n8725), .A4(n8343), .ZN(n9030)
         );
  NAND2_X1 U9720 ( .A1(n7710), .A2(n7709), .ZN(n7708) );
  NAND2_X1 U9721 ( .A1(n12000), .A2(n9956), .ZN(n9934) );
  INV_X1 U9722 ( .A(n10083), .ZN(n7710) );
  NAND2_X1 U9723 ( .A1(n7717), .A2(n7716), .ZN(n7711) );
  INV_X1 U9724 ( .A(n10000), .ZN(n7715) );
  NAND2_X1 U9725 ( .A1(n10083), .A2(n10082), .ZN(n7717) );
  NAND2_X1 U9726 ( .A1(n7721), .A2(n7720), .ZN(n13610) );
  XNOR2_X1 U9727 ( .A(n13606), .B(n13605), .ZN(n7721) );
  NAND2_X1 U9728 ( .A1(n8880), .A2(n12598), .ZN(n7722) );
  NAND2_X2 U9729 ( .A1(n13474), .A2(n13473), .ZN(n13638) );
  NAND2_X1 U9730 ( .A1(n15261), .A2(n15249), .ZN(n15246) );
  NOR2_X2 U9731 ( .A1(n15171), .A2(n15170), .ZN(n15169) );
  NAND2_X1 U9732 ( .A1(n8363), .A2(n9255), .ZN(n9431) );
  INV_X1 U9733 ( .A(n9971), .ZN(n7740) );
  AND2_X2 U9734 ( .A1(n9938), .A2(n13175), .ZN(n11199) );
  NAND2_X1 U9735 ( .A1(n7728), .A2(n7727), .ZN(n7726) );
  NAND2_X2 U9736 ( .A1(n8250), .A2(n8247), .ZN(n9819) );
  INV_X1 U9737 ( .A(n9973), .ZN(n7728) );
  NAND2_X1 U9738 ( .A1(n7741), .A2(n7740), .ZN(n7729) );
  OR2_X1 U9739 ( .A1(n9391), .A2(n11535), .ZN(n9394) );
  NAND2_X1 U9740 ( .A1(n14527), .A2(n14514), .ZN(n14499) );
  OR2_X1 U9741 ( .A1(n11278), .A2(n11279), .ZN(n11276) );
  AND2_X2 U9742 ( .A1(n12018), .A2(n13167), .ZN(n12020) );
  INV_X1 U9743 ( .A(n8163), .ZN(n14441) );
  NOR2_X4 U9744 ( .A1(n14491), .A2(n14664), .ZN(n14477) );
  NAND2_X1 U9745 ( .A1(n8864), .A2(n8862), .ZN(n8187) );
  NAND2_X1 U9746 ( .A1(n8846), .A2(n8844), .ZN(n8190) );
  NAND2_X1 U9747 ( .A1(n8679), .A2(n8677), .ZN(n8542) );
  XNOR2_X1 U9748 ( .A(n13641), .B(n13837), .ZN(n8242) );
  NAND2_X1 U9749 ( .A1(n10213), .A2(n10184), .ZN(n10185) );
  NAND2_X1 U9750 ( .A1(n9973), .A2(n9972), .ZN(n7741) );
  NAND3_X1 U9751 ( .A1(n8565), .A2(n7750), .A3(n16294), .ZN(n7989) );
  INV_X1 U9752 ( .A(n9315), .ZN(n7751) );
  NAND2_X1 U9753 ( .A1(n7751), .A2(n9316), .ZN(n7752) );
  OAI211_X2 U9754 ( .C1(n9694), .C2(n7753), .A(n7752), .B(n9318), .ZN(n9736)
         );
  OAI21_X2 U9755 ( .B1(n9694), .B2(n8364), .A(n9315), .ZN(n9707) );
  XNOR2_X2 U9756 ( .A(n9736), .B(n9721), .ZN(n10599) );
  NAND2_X1 U9757 ( .A1(n9283), .A2(n7757), .ZN(n7756) );
  NAND2_X1 U9758 ( .A1(n9283), .A2(n9282), .ZN(n9577) );
  XNOR2_X1 U9759 ( .A(n9449), .B(n7763), .ZN(n10878) );
  AOI21_X1 U9760 ( .B1(n15258), .B2(n15238), .A(n15239), .ZN(n15237) );
  NAND2_X1 U9761 ( .A1(n7767), .A2(n7514), .ZN(n15202) );
  NAND3_X1 U9762 ( .A1(n7769), .A2(n7511), .A3(n7768), .ZN(n7767) );
  NAND2_X1 U9763 ( .A1(n7770), .A2(n15258), .ZN(n7768) );
  OAI21_X1 U9764 ( .B1(n15258), .B2(n15239), .A(n7770), .ZN(n8420) );
  INV_X1 U9765 ( .A(n7777), .ZN(n12901) );
  NOR2_X1 U9766 ( .A1(n16276), .A2(n12666), .ZN(n12667) );
  NAND2_X1 U9767 ( .A1(n12247), .A2(n12246), .ZN(n7778) );
  NAND2_X1 U9768 ( .A1(n7779), .A2(n12363), .ZN(n7780) );
  INV_X1 U9769 ( .A(n12247), .ZN(n7779) );
  NAND2_X1 U9770 ( .A1(n15381), .A2(n7792), .ZN(n7791) );
  NAND2_X1 U9771 ( .A1(n8183), .A2(n15193), .ZN(n7795) );
  NAND2_X1 U9772 ( .A1(n15322), .A2(n7798), .ZN(n7801) );
  INV_X2 U9773 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15805) );
  AND2_X2 U9774 ( .A1(n7805), .A2(n7804), .ZN(n10293) );
  NAND2_X1 U9775 ( .A1(n8483), .A2(n7521), .ZN(n7809) );
  INV_X1 U9776 ( .A(n7811), .ZN(n15234) );
  NAND2_X1 U9777 ( .A1(n7811), .A2(n7810), .ZN(n15221) );
  NAND2_X1 U9778 ( .A1(n12756), .A2(n8479), .ZN(n7815) );
  NAND2_X1 U9779 ( .A1(n12971), .A2(n8479), .ZN(n15176) );
  NAND2_X1 U9780 ( .A1(n7816), .A2(n8440), .ZN(n12971) );
  NAND2_X2 U9781 ( .A1(n10892), .A2(n10838), .ZN(n10309) );
  XNOR2_X2 U9782 ( .A(n7817), .B(n10241), .ZN(n15622) );
  NAND2_X1 U9783 ( .A1(n10240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7817) );
  NAND3_X1 U9784 ( .A1(n13805), .A2(n7827), .A3(n13830), .ZN(n7822) );
  NOR2_X1 U9785 ( .A1(n13805), .A2(n13806), .ZN(n13826) );
  NAND4_X1 U9786 ( .A1(n7823), .A2(n7822), .A3(n7820), .A4(n16272), .ZN(n7825)
         );
  OAI21_X1 U9787 ( .B1(n12366), .B2(n7838), .A(n7835), .ZN(n16273) );
  OAI21_X1 U9788 ( .B1(n12366), .B2(n12365), .A(n7847), .ZN(n12656) );
  AOI21_X1 U9789 ( .B1(n12365), .B2(n7847), .A(n7844), .ZN(n7843) );
  XNOR2_X2 U9790 ( .A(n7857), .B(P3_IR_REG_27__SCAN_IN), .ZN(n11494) );
  INV_X2 U9791 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7858) );
  NAND3_X1 U9792 ( .A1(n7865), .A2(n10361), .A3(n7863), .ZN(n10376) );
  NAND3_X1 U9793 ( .A1(n10356), .A2(n7864), .A3(n11888), .ZN(n7863) );
  NAND2_X1 U9794 ( .A1(n10519), .A2(n7872), .ZN(n7871) );
  NAND2_X1 U9795 ( .A1(n10578), .A2(n7881), .ZN(n7880) );
  NAND2_X1 U9796 ( .A1(n7888), .A2(n10270), .ZN(n10272) );
  NAND2_X1 U9797 ( .A1(n10229), .A2(n10262), .ZN(n10278) );
  NAND3_X1 U9798 ( .A1(n7888), .A2(n10270), .A3(n16024), .ZN(n7887) );
  OAI21_X1 U9799 ( .B1(n7901), .B2(n7903), .A(n7902), .ZN(n10504) );
  NAND2_X1 U9800 ( .A1(n7917), .A2(n13494), .ZN(n7912) );
  NAND2_X1 U9801 ( .A1(n7913), .A2(n7912), .ZN(n8992) );
  INV_X1 U9802 ( .A(n7914), .ZN(n7913) );
  OAI21_X1 U9803 ( .B1(n8999), .B2(n7929), .A(n7926), .ZN(n14016) );
  NAND2_X1 U9804 ( .A1(n7925), .A2(n7924), .ZN(n9001) );
  NAND2_X1 U9805 ( .A1(n8999), .A2(n7926), .ZN(n7925) );
  OAI21_X1 U9806 ( .B1(n13902), .B2(n7948), .A(n7947), .ZN(n7951) );
  NAND2_X1 U9807 ( .A1(n13900), .A2(n13590), .ZN(n13883) );
  INV_X1 U9808 ( .A(n7955), .ZN(n7954) );
  OAI22_X1 U9809 ( .A1(n8874), .A2(n16325), .B1(n8633), .B2(n8568), .ZN(n7955)
         );
  INV_X1 U9810 ( .A(n16307), .ZN(n8991) );
  NAND2_X1 U9811 ( .A1(n9032), .A2(n7960), .ZN(n8521) );
  NAND2_X1 U9812 ( .A1(n9032), .A2(n7529), .ZN(n14232) );
  AND2_X1 U9813 ( .A1(n9032), .A2(n8342), .ZN(n8561) );
  NOR2_X1 U9814 ( .A1(n12374), .A2(n12373), .ZN(n12674) );
  AOI21_X1 U9815 ( .B1(n12374), .B2(n7972), .A(n7970), .ZN(n7964) );
  NAND2_X1 U9816 ( .A1(n12374), .A2(n7966), .ZN(n7965) );
  OR2_X2 U9817 ( .A1(n12238), .A2(n12371), .ZN(n12239) );
  AND2_X2 U9818 ( .A1(n12237), .A2(n12363), .ZN(n12371) );
  INV_X1 U9819 ( .A(n7976), .ZN(n13716) );
  INV_X1 U9820 ( .A(n7974), .ZN(n13735) );
  OR2_X1 U9821 ( .A1(n13712), .A2(n13713), .ZN(n7976) );
  NAND2_X1 U9822 ( .A1(n16269), .A2(n7984), .ZN(n7983) );
  NAND2_X1 U9823 ( .A1(n7983), .A2(n7982), .ZN(n12896) );
  NAND2_X1 U9824 ( .A1(n7983), .A2(n7980), .ZN(n7979) );
  NOR2_X1 U9825 ( .A1(n7981), .A2(n12909), .ZN(n7980) );
  INV_X1 U9826 ( .A(n7982), .ZN(n7981) );
  NAND2_X1 U9827 ( .A1(n7986), .A2(n8359), .ZN(n7987) );
  NAND2_X1 U9828 ( .A1(n7989), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9829 ( .A1(n9489), .A2(n7993), .ZN(n7990) );
  NAND2_X1 U9830 ( .A1(n7996), .A2(n8006), .ZN(n7999) );
  INV_X1 U9831 ( .A(n10146), .ZN(n7996) );
  NOR2_X1 U9832 ( .A1(n10146), .A2(n10151), .ZN(n8002) );
  OR2_X1 U9833 ( .A1(n10146), .A2(n7997), .ZN(n8000) );
  NAND3_X1 U9834 ( .A1(n8001), .A2(n8007), .A3(n7998), .ZN(n8005) );
  INV_X1 U9835 ( .A(n10186), .ZN(n8003) );
  NAND2_X1 U9836 ( .A1(n10169), .A2(n10168), .ZN(n8001) );
  INV_X1 U9837 ( .A(n10167), .ZN(n8007) );
  NAND2_X1 U9838 ( .A1(n9707), .A2(n8014), .ZN(n8013) );
  NAND2_X1 U9839 ( .A1(n9356), .A2(n8022), .ZN(n8017) );
  AOI21_X1 U9840 ( .B1(n9356), .B2(n7546), .A(n8018), .ZN(n10109) );
  OR2_X1 U9841 ( .A1(n9356), .A2(n9354), .ZN(n8024) );
  NOR2_X1 U9842 ( .A1(n16210), .A2(n16211), .ZN(n16209) );
  NAND2_X1 U9843 ( .A1(n16207), .A2(n16208), .ZN(n8025) );
  XNOR2_X1 U9844 ( .A(n9125), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n16208) );
  AOI21_X1 U9845 ( .B1(n16230), .B2(n9161), .A(n16227), .ZN(n16233) );
  NOR2_X1 U9846 ( .A1(n16233), .A2(n16234), .ZN(n16232) );
  OAI21_X2 U9847 ( .B1(n16243), .B2(n8038), .A(n8037), .ZN(n16247) );
  NAND2_X1 U9848 ( .A1(n8041), .A2(n11842), .ZN(n11843) );
  CLKBUF_X1 U9849 ( .A(n11067), .Z(n8042) );
  NAND2_X2 U9852 ( .A1(n11067), .A2(n10831), .ZN(n10113) );
  INV_X1 U9853 ( .A(n9866), .ZN(n11396) );
  XNOR2_X1 U9854 ( .A(n11752), .B(n7437), .ZN(n9866) );
  NAND2_X1 U9855 ( .A1(n9873), .A2(n9872), .ZN(n11874) );
  NOR2_X1 U9856 ( .A1(n9873), .A2(n16370), .ZN(n8045) );
  NAND2_X1 U9857 ( .A1(n14488), .A2(n8048), .ZN(n8047) );
  OAI21_X1 U9858 ( .B1(n12343), .B2(n9877), .A(n9878), .ZN(n12315) );
  NAND2_X1 U9859 ( .A1(n12314), .A2(n8075), .ZN(n8074) );
  INV_X1 U9860 ( .A(n13878), .ZN(n8089) );
  NAND2_X1 U9861 ( .A1(n8088), .A2(n8085), .ZN(n8967) );
  NAND3_X1 U9862 ( .A1(n8090), .A2(n16309), .A3(n13858), .ZN(n13862) );
  NAND2_X1 U9863 ( .A1(n8732), .A2(n8094), .ZN(n8091) );
  INV_X1 U9864 ( .A(n8843), .ZN(n8107) );
  NAND2_X1 U9865 ( .A1(n8843), .A2(n8104), .ZN(n8100) );
  NOR2_X1 U9866 ( .A1(n8843), .A2(n8842), .ZN(n13992) );
  OAI21_X1 U9867 ( .B1(n13948), .B2(n13252), .A(n8904), .ZN(n13934) );
  NAND2_X1 U9868 ( .A1(n13252), .A2(n8904), .ZN(n8121) );
  NAND4_X1 U9869 ( .A1(n8131), .A2(n8130), .A3(n8129), .A4(n8514), .ZN(n8128)
         );
  NAND2_X1 U9870 ( .A1(n8134), .A2(n8132), .ZN(P3_U3487) );
  AND2_X1 U9871 ( .A1(n8725), .A2(n7445), .ZN(n8135) );
  AND2_X2 U9872 ( .A1(n7439), .A2(n8135), .ZN(n9032) );
  OR2_X1 U9873 ( .A1(n13741), .A2(n13767), .ZN(n8136) );
  OAI21_X1 U9874 ( .B1(n7459), .B2(n8136), .A(n8137), .ZN(n13785) );
  AND3_X2 U9875 ( .A1(n8594), .A2(n8143), .A3(n8141), .ZN(n11664) );
  NAND2_X1 U9876 ( .A1(n11660), .A2(n11667), .ZN(n13681) );
  XNOR2_X1 U9877 ( .A(n11777), .B(n8149), .ZN(n11778) );
  AOI21_X1 U9878 ( .B1(n11957), .B2(n7456), .A(n11956), .ZN(n12244) );
  NAND2_X1 U9879 ( .A1(n8151), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8150) );
  NOR2_X1 U9880 ( .A1(n8154), .A2(n13724), .ZN(n13725) );
  NAND2_X1 U9881 ( .A1(n13833), .A2(n8160), .ZN(n8159) );
  OR2_X1 U9882 ( .A1(n13809), .A2(n8161), .ZN(n8160) );
  NOR2_X1 U9883 ( .A1(n12362), .A2(n12361), .ZN(n12663) );
  NAND2_X1 U9884 ( .A1(n9876), .A2(n9875), .ZN(n12343) );
  OAI211_X2 U9885 ( .C1(n8042), .C2(n16067), .A(n9416), .B(n9415), .ZN(n11249)
         );
  NOR2_X1 U9886 ( .A1(n16389), .A2(n16277), .ZN(n16276) );
  NAND2_X1 U9887 ( .A1(n12665), .A2(n16279), .ZN(n12664) );
  NOR2_X2 U9888 ( .A1(n12880), .A2(n14732), .ZN(n13077) );
  AND2_X2 U9889 ( .A1(n12349), .A2(n12324), .ZN(n12742) );
  OR2_X2 U9890 ( .A1(n11477), .A2(n11517), .ZN(n11847) );
  NOR2_X2 U9891 ( .A1(n11276), .A2(n11249), .ZN(n11401) );
  NAND2_X1 U9892 ( .A1(n14477), .A2(n14465), .ZN(n14442) );
  NOR2_X2 U9893 ( .A1(n14540), .A2(n14530), .ZN(n14527) );
  OAI21_X2 U9894 ( .B1(n9819), .B2(n9224), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9343) );
  NOR2_X2 U9895 ( .A1(n16328), .A2(n11372), .ZN(n11371) );
  NOR2_X2 U9896 ( .A1(n15306), .A2(n15509), .ZN(n8175) );
  NAND2_X1 U9897 ( .A1(n12611), .A2(n8176), .ZN(n12977) );
  NOR2_X2 U9898 ( .A1(n15406), .A2(n15396), .ZN(n8184) );
  NOR2_X2 U9899 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9399) );
  INV_X2 U9900 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U9901 ( .A1(n14546), .A2(n8195), .ZN(n8191) );
  NAND2_X1 U9902 ( .A1(n8191), .A2(n8192), .ZN(n14511) );
  NAND2_X1 U9903 ( .A1(n8545), .A2(n8199), .ZN(n8198) );
  NAND2_X1 U9904 ( .A1(n12735), .A2(n8206), .ZN(n8205) );
  NAND2_X1 U9905 ( .A1(n8781), .A2(n8212), .ZN(n8210) );
  NAND2_X1 U9906 ( .A1(n8591), .A2(n8590), .ZN(n8219) );
  NAND2_X1 U9907 ( .A1(n8591), .A2(n8216), .ZN(n8215) );
  NAND2_X1 U9908 ( .A1(n8233), .A2(n8234), .ZN(n14439) );
  NOR2_X2 U9909 ( .A1(n9344), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U9910 ( .A1(n13088), .A2(n8251), .ZN(n9654) );
  NAND2_X1 U9911 ( .A1(n14992), .A2(n7497), .ZN(n8257) );
  NAND2_X1 U9912 ( .A1(n8257), .A2(n8258), .ZN(n15002) );
  NAND2_X1 U9913 ( .A1(n14912), .A2(n11693), .ZN(n11708) );
  AOI21_X2 U9914 ( .B1(n8265), .B2(n8268), .A(n8264), .ZN(n12704) );
  OAI21_X2 U9915 ( .B1(n14819), .B2(n7498), .A(n8270), .ZN(n14970) );
  NAND2_X1 U9916 ( .A1(n8281), .A2(n8277), .ZN(n15032) );
  NAND2_X1 U9917 ( .A1(n14819), .A2(n14816), .ZN(n8277) );
  NAND4_X1 U9918 ( .A1(n10269), .A2(n10270), .A3(n10228), .A4(n7532), .ZN(
        n10232) );
  NAND3_X1 U9919 ( .A1(n10270), .A2(n10269), .A3(n10228), .ZN(n10781) );
  NAND2_X1 U9920 ( .A1(n12485), .A2(n8283), .ZN(n8282) );
  NAND2_X1 U9921 ( .A1(n12946), .A2(n8288), .ZN(n8287) );
  NOR2_X1 U9922 ( .A1(n8291), .A2(n8289), .ZN(n8288) );
  AOI21_X1 U9923 ( .B1(n13061), .B2(n13057), .A(n13150), .ZN(n8290) );
  NAND2_X1 U9924 ( .A1(n12056), .A2(n8293), .ZN(n8292) );
  NAND2_X1 U9925 ( .A1(n8299), .A2(n8297), .ZN(n8300) );
  NAND2_X1 U9926 ( .A1(n11215), .A2(n11157), .ZN(n11386) );
  INV_X1 U9927 ( .A(n11383), .ZN(n8306) );
  INV_X1 U9928 ( .A(n11384), .ZN(n8307) );
  NAND2_X1 U9929 ( .A1(n8308), .A2(n8309), .ZN(n14353) );
  NAND3_X1 U9930 ( .A1(n9218), .A2(n9216), .A3(n9217), .ZN(n9631) );
  NAND2_X1 U9931 ( .A1(n12637), .A2(n12585), .ZN(n8329) );
  NAND2_X1 U9932 ( .A1(n13254), .A2(n13253), .ZN(n8333) );
  INV_X1 U9933 ( .A(n13255), .ZN(n8332) );
  NAND2_X1 U9934 ( .A1(n13402), .A2(n8336), .ZN(n8334) );
  NAND2_X1 U9935 ( .A1(n9032), .A2(n9034), .ZN(n9028) );
  NAND2_X1 U9936 ( .A1(n13293), .A2(n7471), .ZN(n8345) );
  NAND2_X1 U9937 ( .A1(n9449), .A2(n8356), .ZN(n8354) );
  NAND2_X1 U9938 ( .A1(n9253), .A2(n8361), .ZN(n8362) );
  AND2_X1 U9939 ( .A1(n9255), .A2(n9252), .ZN(n8361) );
  NAND2_X1 U9940 ( .A1(n9253), .A2(n9252), .ZN(n9420) );
  XNOR2_X2 U9941 ( .A(n9313), .B(n15839), .ZN(n9694) );
  NAND2_X1 U9942 ( .A1(n9609), .A2(n9294), .ZN(n9630) );
  NAND2_X1 U9943 ( .A1(n15284), .A2(n8373), .ZN(n8372) );
  INV_X1 U9944 ( .A(n8378), .ZN(n15272) );
  OR2_X1 U9945 ( .A1(n15509), .A2(n15183), .ZN(n8379) );
  NAND2_X1 U9946 ( .A1(n8382), .A2(n10330), .ZN(n8381) );
  NAND2_X1 U9947 ( .A1(n10326), .A2(n11544), .ZN(n8382) );
  NAND2_X1 U9948 ( .A1(n10590), .A2(n8386), .ZN(n8385) );
  NAND2_X1 U9949 ( .A1(n8385), .A2(n7520), .ZN(n10601) );
  NAND2_X1 U9950 ( .A1(n8391), .A2(n8389), .ZN(n10625) );
  NAND2_X1 U9951 ( .A1(n10443), .A2(n8397), .ZN(n8396) );
  NAND2_X1 U9952 ( .A1(n8396), .A2(n8394), .ZN(n10457) );
  NAND2_X1 U9953 ( .A1(n10530), .A2(n8403), .ZN(n8402) );
  NAND2_X1 U9954 ( .A1(n8402), .A2(n8400), .ZN(n10547) );
  NAND2_X2 U9955 ( .A1(n10892), .A2(n7434), .ZN(n10322) );
  INV_X1 U9956 ( .A(n8430), .ZN(n8431) );
  OR2_X1 U9957 ( .A1(n15318), .A2(n8433), .ZN(n8429) );
  NAND2_X1 U9958 ( .A1(n15402), .A2(n7494), .ZN(n8448) );
  NAND2_X1 U9959 ( .A1(n8448), .A2(n7518), .ZN(n15364) );
  NAND2_X1 U9960 ( .A1(n10092), .A2(n7525), .ZN(n8463) );
  NAND2_X1 U9961 ( .A1(n10088), .A2(n7517), .ZN(n8464) );
  INV_X1 U9962 ( .A(n10095), .ZN(n8467) );
  NAND2_X1 U9963 ( .A1(n9998), .A2(n9997), .ZN(n8468) );
  NAND2_X1 U9964 ( .A1(n15324), .A2(n15323), .ZN(n15322) );
  INV_X1 U9965 ( .A(n15319), .ZN(n8474) );
  NOR2_X1 U9966 ( .A1(n15360), .A2(n15182), .ZN(n8477) );
  NAND2_X1 U9967 ( .A1(n12600), .A2(n8481), .ZN(n12720) );
  OAI21_X1 U9968 ( .B1(n15480), .B2(n15584), .A(n16338), .ZN(n8486) );
  OAI211_X1 U9969 ( .C1(n15482), .C2(n7552), .A(n8487), .B(n8488), .ZN(
        P1_U3525) );
  NAND2_X1 U9970 ( .A1(n15221), .A2(n7512), .ZN(n8489) );
  INV_X1 U9971 ( .A(n15203), .ZN(n8490) );
  AND2_X1 U9972 ( .A1(n12923), .A2(n12922), .ZN(n12930) );
  CLKBUF_X1 U9973 ( .A(n11830), .Z(n11735) );
  NAND2_X1 U9974 ( .A1(n9835), .A2(n9820), .ZN(n9847) );
  INV_X4 U9975 ( .A(n11494), .ZN(n13775) );
  INV_X1 U9976 ( .A(n13620), .ZN(n13489) );
  CLKBUF_X1 U9977 ( .A(n13221), .Z(n13136) );
  OAI21_X1 U9978 ( .B1(n10213), .B2(n10190), .A(n8495), .ZN(n10219) );
  CLKBUF_X1 U9979 ( .A(n9910), .Z(n14778) );
  CLKBUF_X1 U9980 ( .A(n9904), .Z(n11076) );
  NAND4_X2 U9981 ( .A1(n9396), .A2(n9395), .A3(n9394), .A4(n9393), .ZN(n9929)
         );
  NAND2_X2 U9982 ( .A1(n13294), .A2(n13936), .ZN(n13293) );
  NOR3_X1 U9983 ( .A1(n10761), .A2(n10726), .A3(n10769), .ZN(n10775) );
  NAND2_X1 U9984 ( .A1(n10568), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10236) );
  INV_X1 U9985 ( .A(n10019), .ZN(n10022) );
  NAND4_X1 U9986 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10261) );
  INV_X1 U9987 ( .A(n9229), .ZN(n14770) );
  NAND2_X1 U9988 ( .A1(n10837), .A2(n10702), .ZN(n10325) );
  NAND2_X1 U9989 ( .A1(n15616), .A2(n10257), .ZN(n10303) );
  NOR2_X1 U9990 ( .A1(n13214), .A2(n13213), .ZN(n8493) );
  NAND2_X1 U9991 ( .A1(n11917), .A2(n16339), .ZN(n16386) );
  INV_X2 U9992 ( .A(n16386), .ZN(n16348) );
  OR2_X1 U9993 ( .A1(n13188), .A2(n14221), .ZN(n8494) );
  AND3_X1 U9994 ( .A1(n10212), .A2(n12731), .A3(n13024), .ZN(n8495) );
  NAND2_X1 U9995 ( .A1(n11247), .A2(n16040), .ZN(n16414) );
  OR2_X1 U9996 ( .A1(n13659), .A2(n16385), .ZN(n8496) );
  AND4_X1 U9997 ( .A1(n13568), .A2(n13999), .A3(n14009), .A4(n13567), .ZN(
        n8498) );
  AND2_X1 U9998 ( .A1(n10567), .A2(n14995), .ZN(n8499) );
  NAND2_X1 U9999 ( .A1(n11455), .A2(n15428), .ZN(n15432) );
  INV_X1 U10000 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14763) );
  INV_X1 U10001 ( .A(n9230), .ZN(n13184) );
  INV_X1 U10002 ( .A(n16313), .ZN(n14090) );
  AND2_X1 U10003 ( .A1(n14097), .A2(n16468), .ZN(n14150) );
  INV_X1 U10004 ( .A(n13621), .ZN(n8666) );
  OR2_X1 U10005 ( .A1(n11485), .A2(n11509), .ZN(n8500) );
  AND2_X1 U10006 ( .A1(n9282), .A2(n9281), .ZN(n8502) );
  AND2_X1 U10007 ( .A1(n11796), .A2(n11795), .ZN(n8503) );
  OR2_X1 U10008 ( .A1(n14652), .A2(n14638), .ZN(n8504) );
  INV_X1 U10009 ( .A(n14818), .ZN(n14816) );
  AND2_X2 U10010 ( .A1(n11185), .A2(n11184), .ZN(n16446) );
  OR2_X1 U10011 ( .A1(n10302), .A2(n10301), .ZN(n10312) );
  INV_X1 U10012 ( .A(n10377), .ZN(n10378) );
  INV_X1 U10013 ( .A(n9942), .ZN(n9943) );
  NAND2_X1 U10014 ( .A1(n9943), .A2(n16298), .ZN(n9944) );
  INV_X1 U10015 ( .A(n10415), .ZN(n10416) );
  INV_X1 U10016 ( .A(n10020), .ZN(n10021) );
  INV_X1 U10017 ( .A(n10531), .ZN(n10532) );
  INV_X1 U10018 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8514) );
  INV_X1 U10019 ( .A(n11793), .ZN(n11794) );
  INV_X1 U10020 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U10021 ( .A1(n12430), .A2(n11794), .ZN(n11796) );
  OR4_X1 U10022 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9814) );
  AND2_X1 U10023 ( .A1(n13972), .A2(n13980), .ZN(n8892) );
  INV_X1 U10024 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8515) );
  INV_X1 U10025 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8512) );
  NAND2_X1 U10026 ( .A1(n9346), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9347) );
  INV_X1 U10027 ( .A(n9706), .ZN(n9316) );
  OR2_X1 U10028 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  INV_X1 U10029 ( .A(n13630), .ZN(n13523) );
  AND4_X1 U10030 ( .A1(n8517), .A2(n8969), .A3(n8516), .A4(n8515), .ZN(n8518)
         );
  INV_X1 U10031 ( .A(n9697), .ZN(n9202) );
  OR2_X1 U10032 ( .A1(n9744), .A2(n14286), .ZN(n9758) );
  INV_X1 U10033 ( .A(n9648), .ZN(n9200) );
  INV_X1 U10034 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9568) );
  INV_X1 U10035 ( .A(n13073), .ZN(n9626) );
  INV_X1 U10036 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10533) );
  INV_X1 U10037 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10430) );
  INV_X1 U10038 ( .A(n12460), .ZN(n12461) );
  INV_X1 U10039 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10230) );
  INV_X1 U10040 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n16006) );
  INV_X1 U10041 ( .A(n13217), .ZN(n13218) );
  OR2_X1 U10042 ( .A1(n8910), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8921) );
  OR2_X1 U10043 ( .A1(n8787), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8802) );
  XNOR2_X1 U10044 ( .A(n13469), .B(n13617), .ZN(n13186) );
  AND2_X1 U10045 ( .A1(n8871), .A2(n15913), .ZN(n8883) );
  NAND2_X1 U10046 ( .A1(n8817), .A2(n8506), .ZN(n8854) );
  NAND2_X1 U10047 ( .A1(n13186), .A2(n10820), .ZN(n10821) );
  NAND2_X1 U10048 ( .A1(n8667), .A2(n8666), .ZN(n12442) );
  OR2_X1 U10049 ( .A1(n8973), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U10050 ( .A1(n8827), .A2(n8826), .ZN(n8556) );
  CLKBUF_X2 U10051 ( .A(n9421), .Z(n9678) );
  NOR2_X1 U10052 ( .A1(n9787), .A2(n14278), .ZN(n9205) );
  OR3_X1 U10053 ( .A1(n9786), .A2(n9785), .A3(n9784), .ZN(n9787) );
  NAND2_X1 U10054 ( .A1(n9203), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9744) );
  INV_X1 U10055 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9635) );
  OR2_X1 U10056 ( .A1(n9528), .A2(n9527), .ZN(n9546) );
  INV_X1 U10057 ( .A(n11082), .ZN(n11077) );
  NAND2_X1 U10058 ( .A1(n9200), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9683) );
  OR2_X1 U10059 ( .A1(n9569), .A2(n9568), .ZN(n9582) );
  INV_X1 U10060 ( .A(n11191), .ZN(n9855) );
  NAND2_X1 U10061 ( .A1(n14394), .A2(n14424), .ZN(n9913) );
  NAND2_X1 U10062 ( .A1(n14734), .A2(n14444), .ZN(n11191) );
  NAND2_X1 U10063 ( .A1(n12500), .A2(n12501), .ZN(n12502) );
  INV_X1 U10064 ( .A(n10642), .ZN(n10643) );
  NOR2_X1 U10065 ( .A1(n10567), .A2(n14995), .ZN(n10580) );
  OR2_X1 U10066 ( .A1(n10534), .A2(n10533), .ZN(n10553) );
  NAND2_X1 U10067 ( .A1(n10617), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U10068 ( .A1(n9324), .A2(n9752), .ZN(n9327) );
  INV_X1 U10069 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n16007) );
  OR2_X1 U10070 ( .A1(n9113), .A2(n9112), .ZN(n9103) );
  OAI21_X1 U10071 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n9111), .A(n9110), .ZN(
        n9177) );
  OR2_X1 U10072 ( .A1(n8921), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8928) );
  INV_X1 U10073 ( .A(n13879), .ZN(n13316) );
  INV_X1 U10074 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15892) );
  INV_X1 U10075 ( .A(n13896), .ZN(n13364) );
  OR2_X1 U10076 ( .A1(n8493), .A2(n13218), .ZN(n13219) );
  INV_X1 U10077 ( .A(n13439), .ZN(n13446) );
  AND2_X1 U10078 ( .A1(n8981), .A2(n8980), .ZN(n13849) );
  INV_X1 U10079 ( .A(n8874), .ZN(n10803) );
  INV_X1 U10080 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11787) );
  INV_X1 U10081 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n12369) );
  OR2_X1 U10082 ( .A1(n8954), .A2(n13283), .ZN(n8955) );
  AND2_X1 U10083 ( .A1(n13569), .A2(n13960), .ZN(n13975) );
  OAI211_X1 U10084 ( .C1(n11913), .C2(n11912), .A(n11911), .B(n11910), .ZN(
        n11917) );
  AND2_X1 U10085 ( .A1(n11802), .A2(n13605), .ZN(n16313) );
  OR2_X1 U10086 ( .A1(n8954), .A2(n15644), .ZN(n8566) );
  INV_X1 U10087 ( .A(n13526), .ZN(n13527) );
  AND2_X1 U10088 ( .A1(n9020), .A2(n9054), .ZN(n14097) );
  INV_X1 U10089 ( .A(n11801), .ZN(n16342) );
  NAND2_X1 U10090 ( .A1(n8813), .A2(n8811), .ZN(n8554) );
  OR2_X1 U10091 ( .A1(n10137), .A2(n10843), .ZN(n9415) );
  OR2_X1 U10092 ( .A1(n9683), .A2(n9201), .ZN(n9697) );
  INV_X1 U10093 ( .A(n14401), .ZN(n12691) );
  AND2_X1 U10094 ( .A1(n11168), .A2(n16041), .ZN(n11166) );
  NAND2_X1 U10095 ( .A1(n14328), .A2(n14604), .ZN(n14387) );
  INV_X1 U10096 ( .A(n9802), .ZN(n9789) );
  AND2_X1 U10097 ( .A1(n16150), .A2(n16149), .ZN(n16151) );
  AND2_X1 U10098 ( .A1(n11077), .A2(n11072), .ZN(n11074) );
  INV_X1 U10099 ( .A(n14538), .ZN(n14569) );
  INV_X1 U10100 ( .A(n10200), .ZN(n14607) );
  INV_X1 U10101 ( .A(n12320), .ZN(n12314) );
  INV_X1 U10102 ( .A(n10194), .ZN(n12013) );
  INV_X1 U10103 ( .A(n10193), .ZN(n11842) );
  AND2_X1 U10104 ( .A1(n9903), .A2(n10125), .ZN(n14619) );
  AND2_X1 U10105 ( .A1(n16033), .A2(n11191), .ZN(n11192) );
  AND2_X1 U10106 ( .A1(n13105), .A2(n9828), .ZN(n9832) );
  NAND2_X1 U10107 ( .A1(n9822), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9824) );
  INV_X1 U10108 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U10109 ( .A1(n9399), .A2(n9213), .ZN(n9422) );
  INV_X1 U10110 ( .A(n15053), .ZN(n12508) );
  INV_X1 U10111 ( .A(n15217), .ZN(n15200) );
  NAND2_X1 U10112 ( .A1(n11710), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15036) );
  AND2_X1 U10113 ( .A1(n10592), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n10605) );
  AND2_X1 U10114 ( .A1(n10580), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n10592) );
  AND2_X1 U10115 ( .A1(n10507), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10521) );
  INV_X1 U10116 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11339) );
  INV_X1 U10117 ( .A(n15201), .ZN(n15242) );
  INV_X1 U10118 ( .A(n12031), .ZN(n12084) );
  NOR2_X1 U10119 ( .A1(n11454), .A2(n11453), .ZN(n15205) );
  OR2_X1 U10120 ( .A1(n15073), .A2(n11048), .ZN(n15451) );
  OR2_X1 U10121 ( .A1(n15608), .A2(P1_D_REG_0__SCAN_IN), .ZN(n11031) );
  OR2_X1 U10122 ( .A1(n15077), .A2(n11048), .ZN(n15410) );
  INV_X1 U10123 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10239) );
  INV_X1 U10124 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15091) );
  OAI22_X1 U10125 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n16291), .B1(n9100), .B2(
        n9151), .ZN(n9114) );
  INV_X1 U10126 ( .A(n16240), .ZN(n9173) );
  AND2_X1 U10127 ( .A1(n9038), .A2(n14239), .ZN(n9039) );
  INV_X1 U10128 ( .A(n13453), .ZN(n13418) );
  AND2_X1 U10129 ( .A1(n11593), .A2(n11804), .ZN(n13439) );
  INV_X1 U10130 ( .A(n12080), .ZN(n13651) );
  AND2_X1 U10131 ( .A1(n8531), .A2(n8530), .ZN(n13911) );
  INV_X1 U10132 ( .A(n13697), .ZN(n13720) );
  INV_X1 U10133 ( .A(n16259), .ZN(n16272) );
  INV_X1 U10134 ( .A(n16278), .ZN(n13813) );
  INV_X1 U10135 ( .A(n13645), .ZN(n12431) );
  AND2_X1 U10136 ( .A1(n9073), .A2(n9068), .ZN(n11910) );
  OR2_X1 U10137 ( .A1(n16476), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U10138 ( .A1(n12080), .A2(n13487), .ZN(n16467) );
  INV_X1 U10139 ( .A(n16467), .ZN(n16418) );
  NOR2_X1 U10140 ( .A1(n13178), .A2(n11577), .ZN(n11595) );
  INV_X1 U10141 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U10142 ( .A1(n8542), .A2(n8541), .ZN(n8696) );
  OR2_X1 U10143 ( .A1(n14443), .A2(n9802), .ZN(n9236) );
  NAND2_X1 U10144 ( .A1(n9388), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9427) );
  INV_X1 U10145 ( .A(n16168), .ZN(n16188) );
  OR2_X1 U10146 ( .A1(n16043), .A2(P2_U3088), .ZN(n16168) );
  INV_X1 U10147 ( .A(n14623), .ZN(n14604) );
  AND2_X1 U10148 ( .A1(n11162), .A2(n11076), .ZN(n14583) );
  AND2_X1 U10149 ( .A1(n9917), .A2(n14508), .ZN(n14596) );
  INV_X1 U10150 ( .A(n14638), .ZN(n14617) );
  INV_X1 U10151 ( .A(n14619), .ZN(n14603) );
  OR2_X1 U10152 ( .A1(n14641), .A2(n14692), .ZN(n14643) );
  AND2_X1 U10153 ( .A1(n14586), .A2(n16299), .ZN(n14739) );
  INV_X1 U10154 ( .A(n11199), .ZN(n16299) );
  AND2_X1 U10155 ( .A1(n11193), .A2(n11192), .ZN(n11247) );
  AND2_X1 U10156 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11170), .ZN(n9850) );
  AND2_X1 U10157 ( .A1(n9540), .A2(n9524), .ZN(n16187) );
  AND2_X1 U10158 ( .A1(n11039), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10828) );
  INV_X1 U10159 ( .A(n15036), .ZN(n15017) );
  NAND2_X1 U10160 ( .A1(n11045), .A2(n15428), .ZN(n15042) );
  AND2_X1 U10161 ( .A1(n10951), .A2(n10950), .ZN(n10999) );
  INV_X1 U10162 ( .A(n12627), .ZN(n15155) );
  OR2_X1 U10163 ( .A1(n16199), .A2(n16194), .ZN(n12627) );
  INV_X1 U10164 ( .A(n15150), .ZN(n15154) );
  INV_X1 U10165 ( .A(n16428), .ZN(n16326) );
  NAND2_X1 U10166 ( .A1(n15219), .A2(n15218), .ZN(n15220) );
  AND2_X1 U10167 ( .A1(n12115), .A2(n12089), .ZN(n16363) );
  INV_X1 U10168 ( .A(n11547), .ZN(n11550) );
  INV_X1 U10169 ( .A(n12127), .ZN(n15460) );
  INV_X1 U10170 ( .A(n11451), .ZN(n11184) );
  OR2_X1 U10171 ( .A1(n11058), .A2(n15157), .ZN(n16353) );
  INV_X1 U10172 ( .A(n15584), .ZN(n15567) );
  NAND2_X1 U10173 ( .A1(n11031), .A2(n15611), .ZN(n11451) );
  OAI21_X1 U10174 ( .B1(n13103), .B2(n11018), .A(n11017), .ZN(n15608) );
  AND2_X1 U10175 ( .A1(n10515), .A2(n10542), .ZN(n12808) );
  AND2_X1 U10176 ( .A1(n9059), .A2(n9039), .ZN(n11577) );
  AND2_X1 U10177 ( .A1(n11585), .A2(n11584), .ZN(n13447) );
  INV_X1 U10178 ( .A(n13972), .ZN(n14200) );
  NAND2_X1 U10179 ( .A1(n11596), .A2(n11914), .ZN(n13453) );
  NAND2_X1 U10180 ( .A1(n8990), .A2(n8989), .ZN(n13656) );
  INV_X1 U10181 ( .A(n13840), .ZN(n16280) );
  INV_X1 U10182 ( .A(n13847), .ZN(n16285) );
  NAND2_X1 U10183 ( .A1(n11918), .A2(n16319), .ZN(n14075) );
  INV_X1 U10184 ( .A(n14039), .ZN(n14054) );
  NAND2_X1 U10185 ( .A1(n11914), .A2(n12431), .ZN(n16339) );
  NAND2_X1 U10186 ( .A1(n16473), .A2(n16418), .ZN(n14164) );
  AND3_X2 U10187 ( .A1(n9062), .A2(n11910), .A3(n9061), .ZN(n16473) );
  INV_X1 U10188 ( .A(n13887), .ZN(n14175) );
  AND2_X2 U10189 ( .A1(n9076), .A2(n11595), .ZN(n16476) );
  NAND2_X1 U10190 ( .A1(n14227), .A2(n10984), .ZN(n10985) );
  INV_X1 U10191 ( .A(n12430), .ZN(n13487) );
  INV_X1 U10192 ( .A(SI_15_), .ZN(n15850) );
  OR2_X1 U10193 ( .A1(n11176), .A2(n11164), .ZN(n14377) );
  OR3_X1 U10194 ( .A1(n9603), .A2(n9602), .A3(n9601), .ZN(n14398) );
  INV_X1 U10195 ( .A(n16055), .ZN(n16191) );
  INV_X1 U10196 ( .A(n9926), .ZN(n9927) );
  AND2_X1 U10197 ( .A1(n14593), .A2(n9859), .ZN(n14638) );
  NAND2_X1 U10198 ( .A1(n11247), .A2(n11246), .ZN(n16412) );
  OR2_X1 U10199 ( .A1(n16038), .A2(n16035), .ZN(n16036) );
  INV_X1 U10200 ( .A(n16041), .ZN(n16038) );
  XNOR2_X1 U10201 ( .A(n9831), .B(n9830), .ZN(n14781) );
  INV_X1 U10202 ( .A(n14444), .ZN(n14508) );
  OR2_X1 U10203 ( .A1(n9564), .A2(n9563), .ZN(n11318) );
  INV_X1 U10204 ( .A(n15533), .ZN(n15360) );
  OR2_X1 U10205 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  INV_X1 U10206 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11511) );
  CLKBUF_X2 U10207 ( .A(P1_U4016), .Z(n15059) );
  OR2_X1 U10208 ( .A1(n16199), .A2(n10900), .ZN(n15150) );
  NAND2_X1 U10209 ( .A1(n15430), .A2(n11460), .ZN(n15434) );
  INV_X1 U10210 ( .A(n15269), .ZN(n15440) );
  INV_X1 U10211 ( .A(n16338), .ZN(n16447) );
  INV_X1 U10212 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11823) );
  INV_X1 U10213 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11189) );
  XNOR2_X1 U10214 ( .A(n9191), .B(n8359), .ZN(n9192) );
  NAND2_X1 U10215 ( .A1(n9067), .A2(n9066), .ZN(P3_U3486) );
  NAND2_X1 U10216 ( .A1(n9081), .A2(n9080), .ZN(P3_U3454) );
  AND2_X1 U10217 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11066), .ZN(P2_U3947) );
  NAND2_X1 U10218 ( .A1(n8504), .A2(n9927), .ZN(P2_U3236) );
  NOR2_X1 U10219 ( .A1(n11040), .A2(n10829), .ZN(P1_U4016) );
  NOR2_X1 U10220 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8612) );
  NAND2_X1 U10221 ( .A1(n8612), .A2(n15902), .ZN(n8648) );
  NAND2_X1 U10222 ( .A1(n8685), .A2(n15713), .ZN(n8716) );
  NAND2_X1 U10223 ( .A1(n8747), .A2(n15914), .ZN(n8787) );
  INV_X1 U10224 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8505) );
  INV_X1 U10225 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8506) );
  INV_X1 U10226 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15913) );
  INV_X1 U10227 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15897) );
  INV_X1 U10228 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15701) );
  NAND2_X1 U10229 ( .A1(n8507), .A2(n15701), .ZN(n8943) );
  INV_X1 U10230 ( .A(n8507), .ZN(n8930) );
  NAND2_X1 U10231 ( .A1(n8930), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10232 ( .A1(n8943), .A2(n8508), .ZN(n13903) );
  INV_X1 U10233 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8509) );
  NAND4_X1 U10234 ( .A1(n8510), .A2(n8618), .A3(n8660), .A4(n8693), .ZN(n8511)
         );
  NOR2_X1 U10235 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8517) );
  NAND2_X1 U10236 ( .A1(n13903), .A2(n10803), .ZN(n8531) );
  INV_X1 U10237 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14177) );
  NAND2_X1 U10238 ( .A1(n8983), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10239 ( .A1(n8960), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8527) );
  OAI211_X1 U10240 ( .C1(n8986), .C2(n14177), .A(n8528), .B(n8527), .ZN(n8529)
         );
  INV_X1 U10241 ( .A(n8529), .ZN(n8530) );
  INV_X1 U10242 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U10243 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11511), .B2(n13031), .ZN(n8918) );
  AOI22_X1 U10244 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n12843), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8245), .ZN(n8905) );
  INV_X1 U10245 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U10246 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n12733), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12730), .ZN(n8893) );
  AOI22_X1 U10247 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12382), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n8186), .ZN(n8862) );
  NAND2_X1 U10248 ( .A1(n8569), .A2(n8582), .ZN(n8533) );
  INV_X1 U10249 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U10250 ( .A1(n10847), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8532) );
  XNOR2_X1 U10251 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8590) );
  INV_X1 U10252 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U10253 ( .A1(n10841), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8534) );
  INV_X1 U10254 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10255 ( .A1(n8535), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10256 ( .A1(n8639), .A2(n8638), .ZN(n8538) );
  NAND2_X1 U10257 ( .A1(n10857), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10258 ( .A1(n10881), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10259 ( .A1(n10887), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10260 ( .A1(n8543), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10261 ( .A1(n8546), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8547) );
  XNOR2_X1 U10262 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8741) );
  NAND2_X1 U10263 ( .A1(n9273), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10264 ( .A1(n8760), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10265 ( .A1(n11189), .A2(n8549), .ZN(n8550) );
  XNOR2_X1 U10266 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8780) );
  NAND2_X1 U10267 ( .A1(n11382), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8552) );
  XNOR2_X1 U10268 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8794) );
  NAND2_X1 U10269 ( .A1(n11761), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10270 ( .A1(n11823), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10271 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8557), .ZN(n8558) );
  INV_X1 U10272 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13174) );
  INV_X1 U10273 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U10274 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8926), .ZN(n8559) );
  AOI22_X1 U10275 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13107), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n7719), .ZN(n8937) );
  INV_X1 U10276 ( .A(n8937), .ZN(n8560) );
  NAND2_X1 U10277 ( .A1(n12750), .A2(n13458), .ZN(n8567) );
  NAND2_X2 U10278 ( .A1(n8567), .A2(n8566), .ZN(n13356) );
  INV_X1 U10279 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n16325) );
  INV_X1 U10280 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8568) );
  INV_X1 U10281 ( .A(n8582), .ZN(n8570) );
  XNOR2_X1 U10282 ( .A(n8569), .B(n8570), .ZN(n10866) );
  INV_X1 U10283 ( .A(SI_1_), .ZN(n10865) );
  NAND2_X1 U10284 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8571) );
  MUX2_X1 U10285 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8571), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8573) );
  INV_X1 U10286 ( .A(n8592), .ZN(n8572) );
  INV_X1 U10287 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n16263) );
  OR2_X1 U10288 ( .A1(n8874), .A2(n16263), .ZN(n8580) );
  NAND2_X1 U10289 ( .A1(n10810), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8579) );
  INV_X1 U10290 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11496) );
  OR2_X1 U10291 ( .A1(n8633), .A2(n11496), .ZN(n8578) );
  INV_X1 U10292 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11915) );
  OR2_X1 U10293 ( .A1(n8915), .A2(n11915), .ZN(n8577) );
  INV_X1 U10294 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10265) );
  AND2_X1 U10295 ( .A1(n10265), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8581) );
  NOR2_X1 U10296 ( .A1(n8582), .A2(n8581), .ZN(n8583) );
  NAND2_X1 U10297 ( .A1(n9249), .A2(SI_0_), .ZN(n9386) );
  OAI21_X1 U10298 ( .B1(n7434), .B2(n8583), .A(n9386), .ZN(n14241) );
  MUX2_X1 U10299 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14241), .S(n7432), .Z(n11919)
         );
  NAND2_X1 U10300 ( .A1(n16312), .A2(n11919), .ZN(n16308) );
  INV_X1 U10301 ( .A(n13484), .ZN(n12154) );
  NAND2_X1 U10302 ( .A1(n12154), .A2(n13483), .ZN(n8584) );
  NAND2_X1 U10303 ( .A1(n8585), .A2(n8584), .ZN(n12152) );
  NAND2_X1 U10304 ( .A1(n8983), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10305 ( .A1(n10810), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8588) );
  INV_X1 U10306 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16340) );
  OR2_X1 U10307 ( .A1(n8874), .A2(n16340), .ZN(n8587) );
  INV_X1 U10308 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11657) );
  OR2_X1 U10309 ( .A1(n8915), .A2(n11657), .ZN(n8586) );
  NAND4_X1 U10310 ( .A1(n8589), .A2(n8588), .A3(n8587), .A4(n8586), .ZN(n8598)
         );
  OR2_X1 U10311 ( .A1(n8655), .A2(SI_2_), .ZN(n8597) );
  XNOR2_X1 U10312 ( .A(n8591), .B(n8590), .ZN(n10867) );
  OR2_X1 U10313 ( .A1(n13462), .A2(n10867), .ZN(n8596) );
  NOR2_X1 U10314 ( .A1(n8592), .A2(n14231), .ZN(n8593) );
  OR2_X1 U10315 ( .A1(n7432), .A2(n11664), .ZN(n8595) );
  NAND2_X1 U10316 ( .A1(n13200), .A2(n11801), .ZN(n13495) );
  NAND2_X1 U10317 ( .A1(n8598), .A2(n16342), .ZN(n13498) );
  NAND2_X1 U10318 ( .A1(n13495), .A2(n13498), .ZN(n13620) );
  NAND2_X1 U10319 ( .A1(n12152), .A2(n13620), .ZN(n8600) );
  NAND2_X1 U10320 ( .A1(n13200), .A2(n16342), .ZN(n8599) );
  NAND2_X1 U10321 ( .A1(n8600), .A2(n8599), .ZN(n12169) );
  NAND2_X1 U10322 ( .A1(n8983), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10323 ( .A1(n10810), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8603) );
  OR2_X1 U10324 ( .A1(n8874), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8602) );
  OR2_X1 U10325 ( .A1(n8915), .A2(n8147), .ZN(n8601) );
  NAND2_X1 U10326 ( .A1(n8594), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8605) );
  MUX2_X1 U10327 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8605), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n8606) );
  AND2_X1 U10328 ( .A1(n8606), .A2(n8619), .ZN(n11677) );
  XNOR2_X1 U10329 ( .A(n8608), .B(n8607), .ZN(n10872) );
  OR2_X1 U10330 ( .A1(n8655), .A2(SI_3_), .ZN(n8609) );
  OAI211_X1 U10331 ( .C1(n11677), .C2(n7432), .A(n8610), .B(n8609), .ZN(n12432) );
  NAND2_X1 U10332 ( .A1(n13665), .A2(n12146), .ZN(n12303) );
  NAND2_X1 U10333 ( .A1(n8611), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10334 ( .A1(n8983), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8616) );
  INV_X1 U10335 ( .A(n8612), .ZN(n8631) );
  NAND2_X1 U10336 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8613) );
  AND2_X1 U10337 ( .A1(n8631), .A2(n8613), .ZN(n12212) );
  OR2_X1 U10338 ( .A1(n8874), .A2(n12212), .ZN(n8615) );
  NAND2_X1 U10339 ( .A1(n10810), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8614) );
  OR2_X1 U10340 ( .A1(n8619), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8642) );
  INV_X1 U10341 ( .A(n11780), .ZN(n13680) );
  XNOR2_X1 U10342 ( .A(n8621), .B(n8620), .ZN(n10869) );
  OR2_X1 U10343 ( .A1(n13462), .A2(n10869), .ZN(n8623) );
  NAND2_X1 U10344 ( .A1(n13664), .A2(n12476), .ZN(n8624) );
  NAND2_X1 U10345 ( .A1(n12169), .A2(n8626), .ZN(n8630) );
  INV_X1 U10346 ( .A(n8624), .ZN(n8625) );
  INV_X1 U10347 ( .A(n13664), .ZN(n12331) );
  NAND2_X1 U10348 ( .A1(n13664), .A2(n12427), .ZN(n13506) );
  NAND2_X1 U10349 ( .A1(n13665), .A2(n12432), .ZN(n13499) );
  NAND2_X1 U10350 ( .A1(n8627), .A2(n13505), .ZN(n8628) );
  NAND3_X1 U10351 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n12529) );
  NAND2_X1 U10352 ( .A1(n8960), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U10353 ( .A1(n10810), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10354 ( .A1(n8631), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8632) );
  AND2_X1 U10355 ( .A1(n8648), .A2(n8632), .ZN(n12531) );
  OR2_X1 U10356 ( .A1(n8874), .A2(n12531), .ZN(n8635) );
  INV_X1 U10357 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11769) );
  OR2_X1 U10358 ( .A1(n8800), .A2(n11769), .ZN(n8634) );
  NAND4_X1 U10359 ( .A1(n8637), .A2(n8636), .A3(n8635), .A4(n8634), .ZN(n13663) );
  OR2_X1 U10360 ( .A1(n8954), .A2(SI_5_), .ZN(n8646) );
  XNOR2_X1 U10361 ( .A(n8639), .B(n8638), .ZN(n10875) );
  OR2_X1 U10362 ( .A1(n13462), .A2(n10875), .ZN(n8645) );
  NAND2_X1 U10363 ( .A1(n8642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8640) );
  MUX2_X1 U10364 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8640), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8641) );
  INV_X1 U10365 ( .A(n8641), .ZN(n8643) );
  NOR2_X1 U10366 ( .A1(n8643), .A2(n8661), .ZN(n11776) );
  OR2_X1 U10367 ( .A1(n7432), .A2(n11776), .ZN(n8644) );
  NAND2_X1 U10368 ( .A1(n12580), .A2(n12336), .ZN(n13512) );
  INV_X1 U10369 ( .A(n12336), .ZN(n12541) );
  NAND2_X1 U10370 ( .A1(n13663), .A2(n12541), .ZN(n13511) );
  NAND2_X1 U10371 ( .A1(n12529), .A2(n13623), .ZN(n12528) );
  NAND2_X1 U10372 ( .A1(n12580), .A2(n12541), .ZN(n8647) );
  INV_X1 U10373 ( .A(n12440), .ZN(n8667) );
  NAND2_X1 U10374 ( .A1(n8960), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10375 ( .A1(n8983), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U10376 ( .A1(n8648), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8649) );
  AND2_X1 U10377 ( .A1(n8670), .A2(n8649), .ZN(n12645) );
  OR2_X1 U10378 ( .A1(n8874), .A2(n12645), .ZN(n8652) );
  INV_X1 U10379 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8650) );
  OR2_X1 U10380 ( .A1(n8986), .A2(n8650), .ZN(n8651) );
  NAND4_X1 U10381 ( .A1(n8654), .A2(n8653), .A3(n8652), .A4(n8651), .ZN(n13662) );
  INV_X1 U10382 ( .A(n13662), .ZN(n12590) );
  OR2_X1 U10383 ( .A1(n8954), .A2(n7764), .ZN(n8665) );
  XNOR2_X1 U10384 ( .A(n10879), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8656) );
  XNOR2_X1 U10385 ( .A(n8657), .B(n8656), .ZN(n10832) );
  OR2_X1 U10386 ( .A1(n13462), .A2(n10832), .ZN(n8664) );
  NOR2_X1 U10387 ( .A1(n8661), .A2(n14231), .ZN(n8658) );
  MUX2_X1 U10388 ( .A(n8658), .B(n14231), .S(n8660), .Z(n8659) );
  INV_X1 U10389 ( .A(n8659), .ZN(n8662) );
  NAND2_X1 U10390 ( .A1(n8661), .A2(n8660), .ZN(n8692) );
  NAND2_X1 U10391 ( .A1(n8662), .A2(n8692), .ZN(n12245) );
  OR2_X1 U10392 ( .A1(n7432), .A2(n12245), .ZN(n8663) );
  INV_X1 U10393 ( .A(n12646), .ZN(n12639) );
  NAND2_X1 U10394 ( .A1(n12590), .A2(n12639), .ZN(n13516) );
  NAND2_X1 U10395 ( .A1(n13662), .A2(n12646), .ZN(n13515) );
  NAND2_X1 U10396 ( .A1(n13662), .A2(n12639), .ZN(n8668) );
  NAND2_X1 U10397 ( .A1(n12442), .A2(n8668), .ZN(n12546) );
  NAND2_X1 U10398 ( .A1(n8960), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U10399 ( .A1(n10810), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8675) );
  INV_X1 U10400 ( .A(n8669), .ZN(n8686) );
  NAND2_X1 U10401 ( .A1(n8670), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8671) );
  AND2_X1 U10402 ( .A1(n8686), .A2(n8671), .ZN(n12595) );
  OR2_X1 U10403 ( .A1(n8874), .A2(n12595), .ZN(n8674) );
  INV_X1 U10404 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8672) );
  OR2_X1 U10405 ( .A1(n8800), .A2(n8672), .ZN(n8673) );
  NAND4_X1 U10406 ( .A1(n8676), .A2(n8675), .A3(n8674), .A4(n8673), .ZN(n13661) );
  INV_X1 U10407 ( .A(n13661), .ZN(n12920) );
  OR2_X1 U10408 ( .A1(n8954), .A2(SI_7_), .ZN(n8683) );
  INV_X1 U10409 ( .A(n8677), .ZN(n8678) );
  XNOR2_X1 U10410 ( .A(n8679), .B(n8678), .ZN(n10860) );
  OR2_X1 U10411 ( .A1(n13462), .A2(n10860), .ZN(n8682) );
  NAND2_X1 U10412 ( .A1(n8692), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U10413 ( .A(n8680), .B(P3_IR_REG_7__SCAN_IN), .ZN(n12246) );
  OR2_X1 U10414 ( .A1(n7432), .A2(n12246), .ZN(n8681) );
  NAND2_X1 U10415 ( .A1(n12920), .A2(n12586), .ZN(n13521) );
  NAND2_X1 U10416 ( .A1(n13661), .A2(n12589), .ZN(n13520) );
  NAND2_X1 U10417 ( .A1(n13521), .A2(n13520), .ZN(n13622) );
  NAND2_X1 U10418 ( .A1(n13661), .A2(n12586), .ZN(n8684) );
  NAND2_X1 U10419 ( .A1(n8960), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U10420 ( .A1(n8983), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8690) );
  INV_X1 U10421 ( .A(n8685), .ZN(n8699) );
  NAND2_X1 U10422 ( .A1(n8686), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8687) );
  AND2_X1 U10423 ( .A1(n8699), .A2(n8687), .ZN(n13329) );
  OR2_X1 U10424 ( .A1(n8874), .A2(n13329), .ZN(n8689) );
  INV_X1 U10425 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12935) );
  OR2_X1 U10426 ( .A1(n8986), .A2(n12935), .ZN(n8688) );
  NAND4_X1 U10427 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n13660) );
  OAI21_X1 U10428 ( .B1(n8692), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8694) );
  XNOR2_X1 U10429 ( .A(n8694), .B(n8693), .ZN(n12672) );
  INV_X1 U10430 ( .A(SI_8_), .ZN(n10864) );
  OR2_X1 U10431 ( .A1(n8954), .A2(n10864), .ZN(n8698) );
  XNOR2_X1 U10432 ( .A(n8696), .B(n8695), .ZN(n10863) );
  OR2_X1 U10433 ( .A1(n13462), .A2(n10863), .ZN(n8697) );
  OAI211_X1 U10434 ( .C1(n7432), .C2(n12672), .A(n8698), .B(n8697), .ZN(n13526) );
  XNOR2_X1 U10435 ( .A(n13660), .B(n13527), .ZN(n13630) );
  INV_X1 U10436 ( .A(n13660), .ZN(n8994) );
  INV_X1 U10437 ( .A(n13001), .ZN(n8713) );
  NAND2_X1 U10438 ( .A1(n8960), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10439 ( .A1(n10810), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8703) );
  OR2_X1 U10440 ( .A1(n8800), .A2(n16270), .ZN(n8702) );
  NAND2_X1 U10441 ( .A1(n8699), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8700) );
  AND2_X1 U10442 ( .A1(n8716), .A2(n8700), .ZN(n16381) );
  OR2_X1 U10443 ( .A1(n8874), .A2(n16381), .ZN(n8701) );
  NAND4_X1 U10444 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n13659) );
  INV_X1 U10445 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U10446 ( .A1(n8706), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U10447 ( .A(n8707), .B(P3_IR_REG_9__SCAN_IN), .ZN(n12659) );
  INV_X1 U10448 ( .A(n8708), .ZN(n8709) );
  XNOR2_X1 U10449 ( .A(n8710), .B(n8709), .ZN(n10833) );
  OR2_X1 U10450 ( .A1(n13462), .A2(n10833), .ZN(n8712) );
  OR2_X1 U10451 ( .A1(n8954), .A2(SI_9_), .ZN(n8711) );
  OAI211_X1 U10452 ( .C1(n12659), .C2(n7432), .A(n8712), .B(n8711), .ZN(n13006) );
  INV_X1 U10453 ( .A(n13006), .ZN(n16385) );
  NAND2_X1 U10454 ( .A1(n8713), .A2(n8496), .ZN(n8715) );
  NAND2_X1 U10455 ( .A1(n13659), .A2(n16385), .ZN(n8714) );
  NAND2_X1 U10456 ( .A1(n8715), .A2(n8714), .ZN(n14089) );
  NAND2_X1 U10457 ( .A1(n8983), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U10458 ( .A1(n10810), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U10459 ( .A1(n8716), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8717) );
  AND2_X1 U10460 ( .A1(n8733), .A2(n8717), .ZN(n14098) );
  OR2_X1 U10461 ( .A1(n8874), .A2(n14098), .ZN(n8719) );
  INV_X1 U10462 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n14099) );
  OR2_X1 U10463 ( .A1(n8915), .A2(n14099), .ZN(n8718) );
  NAND4_X1 U10464 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n13134) );
  INV_X1 U10465 ( .A(n13134), .ZN(n13142) );
  INV_X1 U10466 ( .A(n8722), .ZN(n8723) );
  XNOR2_X1 U10467 ( .A(n8724), .B(n8723), .ZN(n10848) );
  OR2_X1 U10468 ( .A1(n13462), .A2(n10848), .ZN(n8730) );
  OR2_X1 U10469 ( .A1(n8954), .A2(SI_10_), .ZN(n8729) );
  NOR2_X1 U10470 ( .A1(n8726), .A2(n14231), .ZN(n8727) );
  XNOR2_X1 U10471 ( .A(n8727), .B(P3_IR_REG_10__SCAN_IN), .ZN(n12900) );
  INV_X1 U10472 ( .A(n12900), .ZN(n12891) );
  OR2_X1 U10473 ( .A1(n7432), .A2(n12891), .ZN(n8728) );
  NAND2_X1 U10474 ( .A1(n13142), .A2(n14101), .ZN(n13532) );
  INV_X1 U10475 ( .A(n14101), .ZN(n16399) );
  NAND2_X1 U10476 ( .A1(n13134), .A2(n16399), .ZN(n13533) );
  NAND2_X1 U10477 ( .A1(n13532), .A2(n13533), .ZN(n14088) );
  NAND2_X1 U10478 ( .A1(n14089), .A2(n14088), .ZN(n8732) );
  NAND2_X1 U10479 ( .A1(n13134), .A2(n14101), .ZN(n8731) );
  NAND2_X1 U10480 ( .A1(n8983), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U10481 ( .A1(n10810), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8737) );
  INV_X1 U10482 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13051) );
  OR2_X1 U10483 ( .A1(n8915), .A2(n13051), .ZN(n8736) );
  NAND2_X1 U10484 ( .A1(n8733), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8734) );
  AND2_X1 U10485 ( .A1(n8748), .A2(n8734), .ZN(n13139) );
  OR2_X1 U10486 ( .A1(n8874), .A2(n13139), .ZN(n8735) );
  NAND4_X1 U10487 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n14079) );
  NAND2_X1 U10488 ( .A1(n8739), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8740) );
  XNOR2_X1 U10489 ( .A(n8740), .B(P3_IR_REG_11__SCAN_IN), .ZN(n13111) );
  OR2_X1 U10490 ( .A1(n8954), .A2(SI_11_), .ZN(n8745) );
  INV_X1 U10491 ( .A(n8741), .ZN(n8742) );
  XNOR2_X1 U10492 ( .A(n8743), .B(n8742), .ZN(n10858) );
  OR2_X1 U10493 ( .A1(n13462), .A2(n10858), .ZN(n8744) );
  OAI211_X1 U10494 ( .C1(n13111), .C2(n7432), .A(n8745), .B(n8744), .ZN(n13147) );
  INV_X1 U10495 ( .A(n13147), .ZN(n16417) );
  AND2_X1 U10496 ( .A1(n14079), .A2(n16417), .ZN(n8746) );
  NAND2_X1 U10497 ( .A1(n10810), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8753) );
  INV_X1 U10498 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13691) );
  OR2_X1 U10499 ( .A1(n8915), .A2(n13691), .ZN(n8752) );
  INV_X1 U10500 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13690) );
  OR2_X1 U10501 ( .A1(n8800), .A2(n13690), .ZN(n8751) );
  INV_X1 U10502 ( .A(n8747), .ZN(n8769) );
  NAND2_X1 U10503 ( .A1(n8748), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8749) );
  AND2_X1 U10504 ( .A1(n8769), .A2(n8749), .ZN(n14074) );
  OR2_X1 U10505 ( .A1(n8874), .A2(n14074), .ZN(n8750) );
  OR2_X1 U10506 ( .A1(n8739), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U10507 ( .A1(n8761), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8754) );
  XNOR2_X1 U10508 ( .A(n8754), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13694) );
  OR2_X1 U10509 ( .A1(n8954), .A2(SI_12_), .ZN(n8759) );
  INV_X1 U10510 ( .A(n8755), .ZN(n8756) );
  XNOR2_X1 U10511 ( .A(n8757), .B(n8756), .ZN(n10882) );
  OR2_X1 U10512 ( .A1(n13462), .A2(n10882), .ZN(n8758) );
  OAI211_X1 U10513 ( .C1(n13694), .C2(n7432), .A(n8759), .B(n8758), .ZN(n14222) );
  INV_X1 U10514 ( .A(n14222), .ZN(n13353) );
  AND2_X1 U10515 ( .A1(n13658), .A2(n13353), .ZN(n13206) );
  INV_X1 U10516 ( .A(n13206), .ZN(n14057) );
  XNOR2_X1 U10517 ( .A(n8760), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U10518 ( .A1(n10938), .A2(n13458), .ZN(n8768) );
  INV_X1 U10519 ( .A(n8954), .ZN(n8868) );
  INV_X1 U10520 ( .A(n7432), .ZN(n8867) );
  NOR2_X1 U10521 ( .A1(n8765), .A2(n14231), .ZN(n8762) );
  MUX2_X1 U10522 ( .A(n14231), .B(n8762), .S(P3_IR_REG_13__SCAN_IN), .Z(n8763)
         );
  INV_X1 U10523 ( .A(n8763), .ZN(n8766) );
  INV_X1 U10524 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U10525 ( .A1(n8765), .A2(n8764), .ZN(n8783) );
  NAND2_X1 U10526 ( .A1(n8766), .A2(n8783), .ZN(n13697) );
  AOI22_X1 U10527 ( .A1(n8868), .A2(n15855), .B1(n8867), .B2(n13697), .ZN(
        n8767) );
  NAND2_X1 U10528 ( .A1(n8960), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U10529 ( .A1(n10810), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U10530 ( .A1(n8769), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8770) );
  AND2_X1 U10531 ( .A1(n8787), .A2(n8770), .ZN(n14067) );
  OR2_X1 U10532 ( .A1(n8874), .A2(n14067), .ZN(n8772) );
  OR2_X1 U10533 ( .A1(n8800), .A2(n16472), .ZN(n8771) );
  NAND4_X1 U10534 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n14078) );
  INV_X1 U10535 ( .A(n14078), .ZN(n13289) );
  OR2_X1 U10536 ( .A1(n16466), .A2(n13289), .ZN(n8776) );
  AND2_X1 U10537 ( .A1(n14057), .A2(n8776), .ZN(n8775) );
  INV_X1 U10538 ( .A(n8776), .ZN(n8779) );
  NAND2_X1 U10539 ( .A1(n14062), .A2(n14222), .ZN(n14058) );
  NAND2_X1 U10540 ( .A1(n16466), .A2(n13289), .ZN(n8777) );
  AND2_X1 U10541 ( .A1(n14058), .A2(n8777), .ZN(n8778) );
  XNOR2_X1 U10542 ( .A(n8781), .B(n8780), .ZN(n10948) );
  NAND2_X1 U10543 ( .A1(n10948), .A2(n13458), .ZN(n8786) );
  NAND2_X1 U10544 ( .A1(n8783), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8782) );
  MUX2_X1 U10545 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8782), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8784) );
  NAND2_X1 U10546 ( .A1(n8784), .A2(n8814), .ZN(n13734) );
  AOI22_X1 U10547 ( .A1(n8868), .A2(n15851), .B1(n8867), .B2(n13734), .ZN(
        n8785) );
  NAND2_X1 U10548 ( .A1(n8960), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U10549 ( .A1(n8983), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U10550 ( .A1(n8787), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8788) );
  AND2_X1 U10551 ( .A1(n8802), .A2(n8788), .ZN(n13286) );
  OR2_X1 U10552 ( .A1(n8874), .A2(n13286), .ZN(n8790) );
  INV_X1 U10553 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14217) );
  OR2_X1 U10554 ( .A1(n8986), .A2(n14217), .ZN(n8789) );
  NAND4_X1 U10555 ( .A1(n8792), .A2(n8791), .A3(n8790), .A4(n8789), .ZN(n14031) );
  OR2_X1 U10556 ( .A1(n14219), .A2(n14031), .ZN(n13553) );
  NAND2_X1 U10557 ( .A1(n14219), .A2(n14031), .ZN(n13555) );
  INV_X1 U10558 ( .A(n14031), .ZN(n14063) );
  OR2_X1 U10559 ( .A1(n14219), .A2(n14063), .ZN(n8793) );
  XNOR2_X1 U10560 ( .A(n8795), .B(n8794), .ZN(n10991) );
  NAND2_X1 U10561 ( .A1(n10991), .A2(n13458), .ZN(n8799) );
  NAND2_X1 U10562 ( .A1(n8814), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8797) );
  INV_X1 U10563 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8796) );
  XNOR2_X1 U10564 ( .A(n8797), .B(n8796), .ZN(n13773) );
  AOI22_X1 U10565 ( .A1(n8868), .A2(n15850), .B1(n8867), .B2(n13773), .ZN(
        n8798) );
  NAND2_X1 U10566 ( .A1(n8799), .A2(n8798), .ZN(n14159) );
  INV_X1 U10567 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14035) );
  OR2_X1 U10568 ( .A1(n8915), .A2(n14035), .ZN(n8807) );
  NAND2_X1 U10569 ( .A1(n10810), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8806) );
  INV_X1 U10570 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13753) );
  OR2_X1 U10571 ( .A1(n8800), .A2(n13753), .ZN(n8805) );
  INV_X1 U10572 ( .A(n8801), .ZN(n8818) );
  NAND2_X1 U10573 ( .A1(n8802), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8803) );
  AND2_X1 U10574 ( .A1(n8818), .A2(n8803), .ZN(n14034) );
  OR2_X1 U10575 ( .A1(n8874), .A2(n14034), .ZN(n8804) );
  NAND4_X1 U10576 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n14046) );
  NAND2_X1 U10577 ( .A1(n14159), .A2(n14046), .ZN(n13560) );
  INV_X1 U10578 ( .A(n14046), .ZN(n8809) );
  NAND2_X1 U10579 ( .A1(n14159), .A2(n8809), .ZN(n8810) );
  INV_X1 U10580 ( .A(n8811), .ZN(n8812) );
  XNOR2_X1 U10581 ( .A(n8813), .B(n8812), .ZN(n11087) );
  NAND2_X1 U10582 ( .A1(n11087), .A2(n13458), .ZN(n8816) );
  OAI21_X1 U10583 ( .B1(n8814), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8829) );
  XNOR2_X1 U10584 ( .A(n8829), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U10585 ( .A1(n8868), .A2(SI_16_), .B1(n8867), .B2(n13780), .ZN(
        n8815) );
  NAND2_X1 U10586 ( .A1(n8816), .A2(n8815), .ZN(n14026) );
  INV_X1 U10587 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n14154) );
  OR2_X1 U10588 ( .A1(n8800), .A2(n14154), .ZN(n8823) );
  NAND2_X1 U10589 ( .A1(n10810), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8822) );
  INV_X1 U10590 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n14024) );
  OR2_X1 U10591 ( .A1(n8915), .A2(n14024), .ZN(n8821) );
  INV_X1 U10592 ( .A(n8817), .ZN(n8835) );
  NAND2_X1 U10593 ( .A1(n8818), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8819) );
  AND2_X1 U10594 ( .A1(n8835), .A2(n8819), .ZN(n14023) );
  OR2_X1 U10595 ( .A1(n8874), .A2(n14023), .ZN(n8820) );
  NAND4_X1 U10596 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(n14032) );
  INV_X1 U10597 ( .A(n14032), .ZN(n14006) );
  OR2_X1 U10598 ( .A1(n14026), .A2(n14006), .ZN(n13566) );
  NAND2_X1 U10599 ( .A1(n14026), .A2(n14006), .ZN(n13565) );
  NAND2_X1 U10600 ( .A1(n13566), .A2(n13565), .ZN(n14017) );
  OR2_X1 U10601 ( .A1(n14026), .A2(n14032), .ZN(n8824) );
  XNOR2_X1 U10602 ( .A(n8827), .B(n8826), .ZN(n11181) );
  NAND2_X1 U10603 ( .A1(n11181), .A2(n13458), .ZN(n8834) );
  INV_X1 U10604 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U10605 ( .A1(n8829), .A2(n8828), .ZN(n8830) );
  NAND2_X1 U10606 ( .A1(n8830), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8832) );
  INV_X1 U10607 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8831) );
  XNOR2_X1 U10608 ( .A(n8832), .B(n8831), .ZN(n13803) );
  AOI22_X1 U10609 ( .A1(n8868), .A2(n15657), .B1(n8867), .B2(n13803), .ZN(
        n8833) );
  INV_X1 U10610 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14011) );
  OR2_X1 U10611 ( .A1(n8915), .A2(n14011), .ZN(n8840) );
  NAND2_X1 U10612 ( .A1(n10810), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8839) );
  INV_X1 U10613 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14147) );
  OR2_X1 U10614 ( .A1(n8800), .A2(n14147), .ZN(n8838) );
  NAND2_X1 U10615 ( .A1(n8835), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8836) );
  AND2_X1 U10616 ( .A1(n8854), .A2(n8836), .ZN(n14010) );
  OR2_X1 U10617 ( .A1(n8874), .A2(n14010), .ZN(n8837) );
  NAND4_X1 U10618 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n8837), .ZN(n14020) );
  INV_X1 U10619 ( .A(n14020), .ZN(n13374) );
  XNOR2_X1 U10620 ( .A(n14211), .B(n13374), .ZN(n14009) );
  NOR2_X1 U10621 ( .A1(n14003), .A2(n14009), .ZN(n8843) );
  OR2_X1 U10622 ( .A1(n14211), .A2(n13374), .ZN(n8841) );
  INV_X1 U10623 ( .A(n8844), .ZN(n8845) );
  XNOR2_X1 U10624 ( .A(n8846), .B(n8845), .ZN(n11287) );
  NAND2_X1 U10625 ( .A1(n11287), .A2(n13458), .ZN(n8853) );
  NAND2_X1 U10626 ( .A1(n8847), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8848) );
  MUX2_X1 U10627 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8848), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8849) );
  INV_X1 U10628 ( .A(n8849), .ZN(n8851) );
  NOR2_X1 U10629 ( .A1(n8851), .A2(n8850), .ZN(n13827) );
  AOI22_X1 U10630 ( .A1(n8868), .A2(SI_18_), .B1(n8867), .B2(n13827), .ZN(
        n8852) );
  NAND2_X1 U10631 ( .A1(n8853), .A2(n8852), .ZN(n14141) );
  NAND2_X1 U10632 ( .A1(n8960), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U10633 ( .A1(n8983), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8859) );
  NAND2_X1 U10634 ( .A1(n8854), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8855) );
  AND2_X1 U10635 ( .A1(n8872), .A2(n8855), .ZN(n13995) );
  OR2_X1 U10636 ( .A1(n8874), .A2(n13995), .ZN(n8858) );
  INV_X1 U10637 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8856) );
  OR2_X1 U10638 ( .A1(n8986), .A2(n8856), .ZN(n8857) );
  NAND4_X1 U10639 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n13981) );
  OR2_X1 U10640 ( .A1(n14141), .A2(n14007), .ZN(n13480) );
  NAND2_X1 U10641 ( .A1(n14141), .A2(n14007), .ZN(n13959) );
  NAND2_X1 U10642 ( .A1(n13480), .A2(n13959), .ZN(n13991) );
  OR2_X1 U10643 ( .A1(n14141), .A2(n13981), .ZN(n8861) );
  INV_X1 U10644 ( .A(n8862), .ZN(n8863) );
  XNOR2_X1 U10645 ( .A(n8864), .B(n8863), .ZN(n11512) );
  NAND2_X1 U10646 ( .A1(n11512), .A2(n13458), .ZN(n8870) );
  INV_X1 U10647 ( .A(n8850), .ZN(n8865) );
  NAND2_X1 U10648 ( .A1(n8865), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8866) );
  AOI22_X1 U10649 ( .A1(n8868), .A2(SI_19_), .B1(n13829), .B2(n8867), .ZN(
        n8869) );
  NAND2_X1 U10650 ( .A1(n8870), .A2(n8869), .ZN(n13987) );
  NAND2_X1 U10651 ( .A1(n8960), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U10652 ( .A1(n10810), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8877) );
  INV_X1 U10653 ( .A(n8871), .ZN(n8884) );
  NAND2_X1 U10654 ( .A1(n8872), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8873) );
  AND2_X1 U10655 ( .A1(n8884), .A2(n8873), .ZN(n13984) );
  OR2_X1 U10656 ( .A1(n8874), .A2(n13984), .ZN(n8876) );
  INV_X1 U10657 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14139) );
  OR2_X1 U10658 ( .A1(n8800), .A2(n14139), .ZN(n8875) );
  NAND4_X1 U10659 ( .A1(n8878), .A2(n8877), .A3(n8876), .A4(n8875), .ZN(n13993) );
  NOR2_X1 U10660 ( .A1(n13987), .A2(n13993), .ZN(n8879) );
  INV_X1 U10661 ( .A(n13987), .ZN(n14135) );
  XNOR2_X1 U10662 ( .A(n8880), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11826) );
  NAND2_X1 U10663 ( .A1(n11826), .A2(n13458), .ZN(n8882) );
  OR2_X1 U10664 ( .A1(n8954), .A2(n15839), .ZN(n8881) );
  NAND2_X1 U10665 ( .A1(n8960), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8891) );
  INV_X1 U10666 ( .A(n8883), .ZN(n8898) );
  NAND2_X1 U10667 ( .A1(n8884), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U10668 ( .A1(n8898), .A2(n8885), .ZN(n13971) );
  NAND2_X1 U10669 ( .A1(n10803), .A2(n13971), .ZN(n8890) );
  INV_X1 U10670 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n8886) );
  OR2_X1 U10671 ( .A1(n8800), .A2(n8886), .ZN(n8889) );
  INV_X1 U10672 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n8887) );
  OR2_X1 U10673 ( .A1(n8986), .A2(n8887), .ZN(n8888) );
  NAND4_X1 U10674 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), .ZN(n13980) );
  NAND2_X1 U10675 ( .A1(n14200), .A2(n13980), .ZN(n13574) );
  INV_X1 U10676 ( .A(n13980), .ZN(n13950) );
  NAND2_X1 U10677 ( .A1(n13972), .A2(n13950), .ZN(n13573) );
  NAND2_X1 U10678 ( .A1(n13574), .A2(n13573), .ZN(n13962) );
  INV_X1 U10679 ( .A(n8893), .ZN(n8894) );
  XNOR2_X1 U10680 ( .A(n8895), .B(n8894), .ZN(n12008) );
  NAND2_X1 U10681 ( .A1(n12008), .A2(n13458), .ZN(n8897) );
  INV_X1 U10682 ( .A(SI_21_), .ZN(n12010) );
  OR2_X1 U10683 ( .A1(n8954), .A2(n12010), .ZN(n8896) );
  NAND2_X1 U10684 ( .A1(n8898), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U10685 ( .A1(n8910), .A2(n8899), .ZN(n13338) );
  NAND2_X1 U10686 ( .A1(n13338), .A2(n10803), .ZN(n8903) );
  NAND2_X1 U10687 ( .A1(n8983), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U10688 ( .A1(n10810), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U10689 ( .A1(n8960), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8900) );
  NAND4_X1 U10690 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n13967) );
  NOR2_X1 U10691 ( .A1(n13342), .A2(n13967), .ZN(n13252) );
  AND2_X1 U10692 ( .A1(n13342), .A2(n13967), .ZN(n13249) );
  INV_X1 U10693 ( .A(n13249), .ZN(n8904) );
  INV_X1 U10694 ( .A(n8905), .ZN(n8906) );
  XNOR2_X1 U10695 ( .A(n8907), .B(n8906), .ZN(n12082) );
  NAND2_X1 U10696 ( .A1(n12082), .A2(n13458), .ZN(n8909) );
  OR2_X1 U10697 ( .A1(n8954), .A2(n9721), .ZN(n8908) );
  INV_X1 U10698 ( .A(n13419), .ZN(n14193) );
  INV_X1 U10699 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U10700 ( .A1(n8910), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U10701 ( .A1(n8921), .A2(n8911), .ZN(n13941) );
  NAND2_X1 U10702 ( .A1(n13941), .A2(n10803), .ZN(n8913) );
  AOI22_X1 U10703 ( .A1(n10810), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n8983), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n8912) );
  OAI211_X1 U10704 ( .C1(n8915), .C2(n8914), .A(n8913), .B(n8912), .ZN(n13657)
         );
  INV_X1 U10705 ( .A(n13657), .ZN(n13951) );
  NAND2_X1 U10706 ( .A1(n14193), .A2(n13951), .ZN(n8916) );
  NAND2_X1 U10707 ( .A1(n12255), .A2(n13458), .ZN(n8920) );
  INV_X1 U10708 ( .A(SI_23_), .ZN(n12258) );
  OR2_X1 U10709 ( .A1(n8954), .A2(n12258), .ZN(n8919) );
  NAND2_X1 U10710 ( .A1(n8921), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U10711 ( .A1(n8928), .A2(n8922), .ZN(n13928) );
  NAND2_X1 U10712 ( .A1(n13928), .A2(n10803), .ZN(n8925) );
  AOI22_X1 U10713 ( .A1(n10810), .A2(P3_REG0_REG_23__SCAN_IN), .B1(n8983), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U10714 ( .A1(n8960), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8923) );
  INV_X1 U10715 ( .A(n13936), .ZN(n13389) );
  NAND2_X1 U10716 ( .A1(n14189), .A2(n13389), .ZN(n13585) );
  NAND2_X1 U10717 ( .A1(n13257), .A2(n13936), .ZN(n13584) );
  MUX2_X1 U10718 ( .A(n8927), .B(SI_24_), .S(n7434), .Z(n14240) );
  NAND2_X1 U10719 ( .A1(n8928), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U10720 ( .A1(n8930), .A2(n8929), .ZN(n13916) );
  NAND2_X1 U10721 ( .A1(n13916), .A2(n10803), .ZN(n8935) );
  INV_X1 U10722 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U10723 ( .A1(n8960), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U10724 ( .A1(n8983), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8931) );
  OAI211_X1 U10725 ( .C1(n14181), .C2(n8986), .A(n8932), .B(n8931), .ZN(n8933)
         );
  INV_X1 U10726 ( .A(n8933), .ZN(n8934) );
  NOR2_X1 U10727 ( .A1(n14120), .A2(n13921), .ZN(n8936) );
  INV_X1 U10728 ( .A(n14120), .ZN(n14182) );
  XNOR2_X1 U10729 ( .A(n13356), .B(n13880), .ZN(n13901) );
  NOR2_X1 U10730 ( .A1(n13892), .A2(n13901), .ZN(n13898) );
  AOI21_X2 U10731 ( .B1(n13880), .B2(n13356), .A(n13898), .ZN(n13878) );
  AOI22_X1 U10732 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n14782), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n7735), .ZN(n8952) );
  INV_X1 U10733 ( .A(n8952), .ZN(n8940) );
  XNOR2_X1 U10734 ( .A(n8951), .B(n8940), .ZN(n12914) );
  NAND2_X1 U10735 ( .A1(n12914), .A2(n13458), .ZN(n8942) );
  INV_X1 U10736 ( .A(SI_26_), .ZN(n12916) );
  OR2_X1 U10737 ( .A1(n8954), .A2(n12916), .ZN(n8941) );
  NAND2_X2 U10738 ( .A1(n8942), .A2(n8941), .ZN(n13887) );
  NAND2_X1 U10739 ( .A1(n8943), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U10740 ( .A1(n8957), .A2(n8944), .ZN(n13886) );
  NAND2_X1 U10741 ( .A1(n13886), .A2(n10803), .ZN(n8949) );
  INV_X1 U10742 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14173) );
  NAND2_X1 U10743 ( .A1(n8983), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U10744 ( .A1(n8960), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8945) );
  OAI211_X1 U10745 ( .C1(n14173), .C2(n8986), .A(n8946), .B(n8945), .ZN(n8947)
         );
  INV_X1 U10746 ( .A(n8947), .ZN(n8948) );
  NOR2_X1 U10747 ( .A1(n13887), .A2(n13896), .ZN(n8950) );
  INV_X1 U10748 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U10749 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n14777), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n15624), .ZN(n10792) );
  INV_X1 U10750 ( .A(n10792), .ZN(n8953) );
  NAND2_X1 U10751 ( .A1(n13281), .A2(n13458), .ZN(n8956) );
  INV_X1 U10752 ( .A(SI_27_), .ZN(n13283) );
  INV_X1 U10753 ( .A(n8981), .ZN(n8959) );
  NAND2_X1 U10754 ( .A1(n8957), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U10755 ( .A1(n8959), .A2(n8958), .ZN(n13873) );
  NAND2_X1 U10756 ( .A1(n13873), .A2(n10803), .ZN(n8966) );
  INV_X1 U10757 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U10758 ( .A1(n8983), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U10759 ( .A1(n8960), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8961) );
  OAI211_X1 U10760 ( .C1(n8963), .C2(n8986), .A(n8962), .B(n8961), .ZN(n8964)
         );
  INV_X1 U10761 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U10762 ( .A1(n13874), .A2(n13316), .ZN(n13595) );
  AND2_X2 U10763 ( .A1(n13596), .A2(n13595), .ZN(n13474) );
  NAND2_X1 U10764 ( .A1(n8967), .A2(n13474), .ZN(n8968) );
  AND2_X1 U10765 ( .A1(n13857), .A2(n8968), .ZN(n9023) );
  NAND2_X1 U10766 ( .A1(n8850), .A2(n8969), .ZN(n8977) );
  NAND2_X1 U10767 ( .A1(n8973), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U10768 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8972), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8974) );
  AND2_X1 U10769 ( .A1(n13651), .A2(n13829), .ZN(n9070) );
  INV_X1 U10770 ( .A(n9070), .ZN(n8979) );
  NAND2_X1 U10771 ( .A1(n8975), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U10772 ( .A1(n8977), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10773 ( .A1(n12430), .A2(n11793), .ZN(n13472) );
  NAND2_X2 U10774 ( .A1(n8979), .A2(n13472), .ZN(n16309) );
  INV_X1 U10775 ( .A(n16309), .ZN(n14005) );
  INV_X1 U10776 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8980) );
  NOR2_X1 U10777 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  NAND2_X1 U10778 ( .A1(n13867), .A2(n10803), .ZN(n8990) );
  INV_X1 U10779 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U10780 ( .A1(n8960), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U10781 ( .A1(n8983), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8984) );
  OAI211_X1 U10782 ( .C1(n8987), .C2(n8986), .A(n8985), .B(n8984), .ZN(n8988)
         );
  INV_X1 U10783 ( .A(n8988), .ZN(n8989) );
  INV_X1 U10784 ( .A(n13183), .ZN(n13648) );
  NAND2_X1 U10785 ( .A1(n13648), .A2(n11494), .ZN(n11488) );
  NAND2_X1 U10786 ( .A1(n7432), .A2(n11488), .ZN(n11802) );
  NAND2_X1 U10787 ( .A1(n13651), .A2(n12430), .ZN(n13598) );
  AOI22_X1 U10788 ( .A1(n13656), .A2(n16313), .B1(n16311), .B2(n13896), .ZN(
        n9022) );
  NOR2_X1 U10789 ( .A1(n16312), .A2(n11855), .ZN(n16306) );
  NAND2_X1 U10790 ( .A1(n16307), .A2(n16306), .ZN(n16305) );
  NAND2_X1 U10791 ( .A1(n12154), .A2(n7952), .ZN(n13491) );
  NAND2_X1 U10792 ( .A1(n16305), .A2(n13491), .ZN(n12153) );
  INV_X1 U10793 ( .A(n13624), .ZN(n13503) );
  INV_X1 U10794 ( .A(n13623), .ZN(n13509) );
  NAND2_X1 U10795 ( .A1(n12527), .A2(n13509), .ZN(n8993) );
  NAND2_X1 U10796 ( .A1(n8993), .A2(n13512), .ZN(n12439) );
  NAND2_X1 U10797 ( .A1(n12439), .A2(n13621), .ZN(n12438) );
  NAND2_X1 U10798 ( .A1(n12438), .A2(n13516), .ZN(n12550) );
  INV_X1 U10799 ( .A(n13622), .ZN(n13518) );
  NAND2_X1 U10800 ( .A1(n12550), .A2(n13518), .ZN(n12549) );
  NAND2_X1 U10801 ( .A1(n12549), .A2(n13521), .ZN(n12921) );
  NAND2_X1 U10802 ( .A1(n12921), .A2(n13523), .ZN(n12923) );
  NAND2_X1 U10803 ( .A1(n8994), .A2(n13526), .ZN(n8995) );
  NAND2_X1 U10804 ( .A1(n12923), .A2(n8995), .ZN(n13000) );
  NOR2_X1 U10805 ( .A1(n13659), .A2(n13006), .ZN(n13534) );
  NAND2_X1 U10806 ( .A1(n13659), .A2(n13006), .ZN(n12999) );
  XNOR2_X1 U10807 ( .A(n14079), .B(n13147), .ZN(n13137) );
  INV_X1 U10808 ( .A(n14079), .ZN(n14091) );
  NAND2_X1 U10809 ( .A1(n14091), .A2(n16417), .ZN(n13540) );
  NAND2_X1 U10810 ( .A1(n8996), .A2(n13540), .ZN(n14073) );
  NAND2_X1 U10811 ( .A1(n14062), .A2(n13353), .ZN(n13548) );
  NAND2_X1 U10812 ( .A1(n13658), .A2(n14222), .ZN(n13546) );
  NAND2_X1 U10813 ( .A1(n13548), .A2(n13546), .ZN(n14076) );
  INV_X1 U10814 ( .A(n14076), .ZN(n8997) );
  NAND2_X1 U10815 ( .A1(n14073), .A2(n8997), .ZN(n8998) );
  NAND2_X1 U10816 ( .A1(n16466), .A2(n14078), .ZN(n13542) );
  OR2_X1 U10817 ( .A1(n16466), .A2(n14078), .ZN(n13552) );
  INV_X1 U10818 ( .A(n13553), .ZN(n9000) );
  INV_X1 U10819 ( .A(n14017), .ZN(n13563) );
  NAND2_X1 U10820 ( .A1(n9001), .A2(n13565), .ZN(n14008) );
  NAND2_X1 U10821 ( .A1(n14008), .A2(n14009), .ZN(n9002) );
  OR2_X1 U10822 ( .A1(n14211), .A2(n14020), .ZN(n13477) );
  NAND2_X1 U10823 ( .A1(n13987), .A2(n13426), .ZN(n13960) );
  AND2_X1 U10824 ( .A1(n13960), .A2(n13573), .ZN(n9007) );
  INV_X1 U10825 ( .A(n9007), .ZN(n9003) );
  OR2_X1 U10826 ( .A1(n13987), .A2(n13426), .ZN(n13569) );
  OR2_X1 U10827 ( .A1(n9003), .A2(n13975), .ZN(n9004) );
  AND2_X1 U10828 ( .A1(n9004), .A2(n13574), .ZN(n9006) );
  AND2_X1 U10829 ( .A1(n13999), .A2(n9006), .ZN(n9005) );
  NAND2_X1 U10830 ( .A1(n14000), .A2(n9005), .ZN(n9011) );
  INV_X1 U10831 ( .A(n9006), .ZN(n9009) );
  AND2_X1 U10832 ( .A1(n13959), .A2(n9007), .ZN(n9008) );
  INV_X1 U10833 ( .A(n13967), .ZN(n13937) );
  AND2_X1 U10834 ( .A1(n14195), .A2(n13967), .ZN(n13476) );
  INV_X1 U10835 ( .A(n13476), .ZN(n13578) );
  OR2_X1 U10836 ( .A1(n13419), .A2(n13951), .ZN(n13475) );
  NAND2_X1 U10837 ( .A1(n13419), .A2(n13951), .ZN(n13922) );
  NAND2_X1 U10838 ( .A1(n13475), .A2(n13922), .ZN(n13933) );
  NAND2_X1 U10839 ( .A1(n13940), .A2(n13939), .ZN(n13938) );
  AND2_X1 U10840 ( .A1(n13923), .A2(n13922), .ZN(n9012) );
  XNOR2_X1 U10841 ( .A(n14120), .B(n13921), .ZN(n13910) );
  NAND2_X1 U10842 ( .A1(n14120), .A2(n13895), .ZN(n13588) );
  INV_X1 U10843 ( .A(n13901), .ZN(n13893) );
  NAND2_X1 U10844 ( .A1(n13356), .A2(n13911), .ZN(n13590) );
  NAND2_X1 U10845 ( .A1(n13887), .A2(n13364), .ZN(n13591) );
  NAND2_X1 U10846 ( .A1(n13592), .A2(n13591), .ZN(n13882) );
  INV_X1 U10847 ( .A(n13592), .ZN(n9013) );
  NAND2_X1 U10848 ( .A1(n9014), .A2(n13474), .ZN(n10819) );
  OAI21_X1 U10849 ( .B1(n9014), .B2(n13474), .A(n10819), .ZN(n9064) );
  AND2_X1 U10850 ( .A1(n13487), .A2(n11794), .ZN(n9015) );
  XNOR2_X1 U10851 ( .A(n12080), .B(n9015), .ZN(n9017) );
  NAND2_X1 U10852 ( .A1(n13487), .A2(n13837), .ZN(n9016) );
  NAND2_X1 U10853 ( .A1(n9017), .A2(n9016), .ZN(n11587) );
  INV_X1 U10854 ( .A(n11795), .ZN(n13643) );
  AND2_X1 U10855 ( .A1(n16467), .A2(n13643), .ZN(n9018) );
  NAND2_X1 U10856 ( .A1(n11587), .A2(n9018), .ZN(n9020) );
  AND2_X1 U10857 ( .A1(n11795), .A2(n13837), .ZN(n9019) );
  NAND2_X1 U10858 ( .A1(n13651), .A2(n9019), .ZN(n9054) );
  INV_X1 U10859 ( .A(n14097), .ZN(n12302) );
  NAND2_X1 U10860 ( .A1(n9064), .A2(n12302), .ZN(n9021) );
  OAI211_X1 U10861 ( .C1(n9023), .C2(n14005), .A(n9022), .B(n9021), .ZN(n13871) );
  NAND2_X1 U10862 ( .A1(n9024), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9025) );
  MUX2_X1 U10863 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9025), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n9027) );
  NAND2_X1 U10864 ( .A1(n9027), .A2(n9026), .ZN(n11483) );
  NAND2_X1 U10865 ( .A1(n9028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9029) );
  MUX2_X1 U10866 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9029), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9031) );
  INV_X1 U10867 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U10868 ( .A1(n9033), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9035) );
  INV_X1 U10869 ( .A(n12752), .ZN(n9038) );
  NOR2_X1 U10870 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9043) );
  NOR4_X1 U10871 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9042) );
  NOR4_X1 U10872 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9041) );
  NOR4_X1 U10873 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9040) );
  NAND4_X1 U10874 ( .A1(n9043), .A2(n9042), .A3(n9041), .A4(n9040), .ZN(n9053)
         );
  NOR4_X1 U10875 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9047) );
  NOR4_X1 U10876 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9046) );
  NOR4_X1 U10877 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9045) );
  NOR4_X1 U10878 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9044) );
  NAND4_X1 U10879 ( .A1(n9047), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(n9052)
         );
  XNOR2_X1 U10880 ( .A(n9048), .B(P3_B_REG_SCAN_IN), .ZN(n9049) );
  NAND2_X1 U10881 ( .A1(n9049), .A2(n12752), .ZN(n9050) );
  INV_X1 U10882 ( .A(n10984), .ZN(n9051) );
  OAI21_X1 U10883 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9071) );
  NAND2_X1 U10884 ( .A1(n11595), .A2(n9071), .ZN(n11909) );
  AND2_X1 U10885 ( .A1(n9054), .A2(n13598), .ZN(n11913) );
  NAND3_X1 U10886 ( .A1(n16418), .A2(n11794), .A3(n11795), .ZN(n9055) );
  NAND2_X1 U10887 ( .A1(n11913), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U10888 ( .A1(n12917), .A2(n12752), .ZN(n9056) );
  AND2_X1 U10889 ( .A1(n9057), .A2(n11912), .ZN(n9058) );
  NOR2_X1 U10890 ( .A1(n11909), .A2(n9058), .ZN(n9062) );
  NAND2_X1 U10891 ( .A1(n13179), .A2(n11912), .ZN(n9073) );
  OR2_X1 U10892 ( .A1(n13179), .A2(n11912), .ZN(n9068) );
  INV_X1 U10893 ( .A(n11912), .ZN(n14228) );
  NAND2_X1 U10894 ( .A1(n13605), .A2(n11795), .ZN(n11579) );
  INV_X1 U10895 ( .A(n11913), .ZN(n9060) );
  NAND2_X1 U10896 ( .A1(n11579), .A2(n9060), .ZN(n11907) );
  NAND2_X1 U10897 ( .A1(n14228), .A2(n11907), .ZN(n9061) );
  MUX2_X1 U10898 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13871), .S(n16473), .Z(
        n9063) );
  INV_X1 U10899 ( .A(n9063), .ZN(n9067) );
  INV_X1 U10900 ( .A(n9064), .ZN(n13877) );
  NAND2_X1 U10901 ( .A1(n11794), .A2(n13829), .ZN(n13645) );
  NAND2_X1 U10902 ( .A1(n12080), .A2(n12431), .ZN(n16468) );
  INV_X1 U10903 ( .A(n16468), .ZN(n9078) );
  NAND2_X1 U10904 ( .A1(n16473), .A2(n9078), .ZN(n14165) );
  OAI22_X1 U10905 ( .A1(n13877), .A2(n14165), .B1(n13280), .B2(n14164), .ZN(
        n9065) );
  INV_X1 U10906 ( .A(n9065), .ZN(n9066) );
  INV_X1 U10907 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U10908 ( .A1(n9069), .A2(n9071), .ZN(n11594) );
  AND2_X1 U10909 ( .A1(n13487), .A2(n11793), .ZN(n13642) );
  NAND2_X1 U10910 ( .A1(n9070), .A2(n13642), .ZN(n11588) );
  INV_X1 U10911 ( .A(n11588), .ZN(n11578) );
  NOR2_X1 U10912 ( .A1(n13598), .A2(n11795), .ZN(n11762) );
  NOR2_X1 U10913 ( .A1(n11578), .A2(n11762), .ZN(n9075) );
  INV_X1 U10914 ( .A(n9071), .ZN(n9072) );
  OR2_X1 U10915 ( .A1(n9073), .A2(n9072), .ZN(n11592) );
  INV_X1 U10916 ( .A(n11587), .ZN(n9074) );
  OAI22_X1 U10917 ( .A1(n11594), .A2(n9075), .B1(n11592), .B2(n9074), .ZN(
        n9076) );
  MUX2_X1 U10918 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13871), .S(n16476), .Z(
        n9077) );
  INV_X1 U10919 ( .A(n9077), .ZN(n9081) );
  NAND2_X1 U10920 ( .A1(n16476), .A2(n9078), .ZN(n14223) );
  OAI22_X1 U10921 ( .A1(n13877), .A2(n14223), .B1(n13280), .B2(n14221), .ZN(
        n9079) );
  INV_X1 U10922 ( .A(n9079), .ZN(n9080) );
  INV_X1 U10923 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9111) );
  INV_X1 U10924 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13747) );
  XNOR2_X1 U10925 ( .A(n13747), .B(n9111), .ZN(n9170) );
  INV_X1 U10926 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U10927 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9165) );
  INV_X1 U10928 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9106) );
  INV_X1 U10929 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13127) );
  INV_X1 U10930 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9082) );
  XOR2_X1 U10931 ( .A(n9082), .B(n11339), .Z(n9113) );
  INV_X1 U10932 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U10933 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9115) );
  INV_X1 U10934 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n16291) );
  AND2_X1 U10935 ( .A1(n16291), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n9100) );
  NOR2_X1 U10936 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n12369), .ZN(n9099) );
  NAND2_X1 U10937 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n11787), .ZN(n9093) );
  NOR2_X1 U10938 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n9091), .ZN(n9083) );
  AOI21_X1 U10939 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n9091), .A(n9083), .ZN(
        n9123) );
  XNOR2_X1 U10940 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n9127) );
  NAND2_X1 U10941 ( .A1(n9128), .A2(n9127), .ZN(n9084) );
  NAND2_X1 U10942 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n9085), .ZN(n9086) );
  NAND2_X1 U10943 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n9087), .ZN(n9089) );
  XOR2_X1 U10944 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(n9087), .Z(n9134) );
  NAND2_X1 U10945 ( .A1(n9134), .A2(n15091), .ZN(n9088) );
  NAND2_X1 U10946 ( .A1(n9089), .A2(n9088), .ZN(n9124) );
  NAND2_X1 U10947 ( .A1(n9123), .A2(n9124), .ZN(n9090) );
  NOR2_X1 U10948 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n11787), .ZN(n9092) );
  OR2_X1 U10949 ( .A1(n9094), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U10950 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n9096), .ZN(n9098) );
  XNOR2_X1 U10951 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n9096), .ZN(n9145) );
  NAND2_X1 U10952 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n12369), .ZN(n9116) );
  NAND2_X1 U10953 ( .A1(n9115), .A2(n9114), .ZN(n9101) );
  INV_X1 U10954 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U10955 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n11603), .ZN(n9104) );
  XNOR2_X1 U10956 ( .A(n9106), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n9162) );
  NOR2_X1 U10957 ( .A1(n9163), .A2(n9162), .ZN(n9105) );
  AOI21_X1 U10958 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n9106), .A(n9105), .ZN(
        n9164) );
  NAND2_X1 U10959 ( .A1(n9165), .A2(n9164), .ZN(n9107) );
  INV_X1 U10960 ( .A(n9169), .ZN(n9109) );
  NAND2_X1 U10961 ( .A1(n9170), .A2(n9109), .ZN(n9110) );
  XNOR2_X1 U10962 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9177), .ZN(n9178) );
  XOR2_X1 U10963 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9178), .Z(n9176) );
  INV_X1 U10964 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n16230) );
  INV_X1 U10965 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n16225) );
  XOR2_X1 U10966 ( .A(n9113), .B(n9112), .Z(n16224) );
  XNOR2_X1 U10967 ( .A(n9115), .B(n9114), .ZN(n16220) );
  OAI21_X1 U10968 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n12369), .A(n9116), .ZN(
        n9117) );
  XOR2_X1 U10969 ( .A(n9118), .B(n9117), .Z(n9148) );
  XNOR2_X1 U10970 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9120) );
  XOR2_X1 U10971 ( .A(n9120), .B(n9119), .Z(n9142) );
  INV_X1 U10972 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n16212) );
  XNOR2_X1 U10973 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9122) );
  XNOR2_X1 U10974 ( .A(n9122), .B(n9121), .ZN(n16211) );
  INV_X1 U10975 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n16085) );
  XOR2_X1 U10976 ( .A(n9124), .B(n9123), .Z(n9125) );
  OR2_X1 U10977 ( .A1(n16085), .A2(n9125), .ZN(n9139) );
  XOR2_X1 U10978 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n9126), .Z(n9132) );
  AOI21_X1 U10979 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n16268), .A(n9128), .ZN(
        n16202) );
  INV_X1 U10980 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n16201) );
  XNOR2_X1 U10981 ( .A(n9128), .B(n9127), .ZN(n16255) );
  OR2_X1 U10982 ( .A1(n16254), .A2(n16255), .ZN(n9130) );
  NAND2_X1 U10983 ( .A1(n16254), .A2(n16255), .ZN(n16253) );
  INV_X1 U10984 ( .A(n16253), .ZN(n9129) );
  AOI21_X1 U10985 ( .B1(n9130), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9129), .ZN(
        n9131) );
  AND2_X1 U10986 ( .A1(n9132), .A2(n9131), .ZN(n16204) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n16203), .ZN(n9133) );
  NOR2_X1 U10988 ( .A1(n16204), .A2(n9133), .ZN(n9136) );
  XNOR2_X1 U10989 ( .A(n15091), .B(n9134), .ZN(n9135) );
  NOR2_X1 U10990 ( .A1(n9136), .A2(n9135), .ZN(n9138) );
  NAND2_X1 U10991 ( .A1(n16211), .A2(n16210), .ZN(n9140) );
  NOR2_X1 U10992 ( .A1(n9142), .A2(n9141), .ZN(n16249) );
  NOR2_X1 U10993 ( .A1(n16250), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9143) );
  NOR2_X1 U10994 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9144), .ZN(n9147) );
  XNOR2_X1 U10995 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9145), .ZN(n16214) );
  NOR2_X1 U10996 ( .A1(n16215), .A2(n16214), .ZN(n9146) );
  NAND2_X1 U10997 ( .A1(n9148), .A2(n9149), .ZN(n9150) );
  XNOR2_X1 U10998 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9152) );
  XOR2_X1 U10999 ( .A(n9152), .B(n9151), .Z(n9154) );
  NAND2_X1 U11000 ( .A1(n9153), .A2(n9154), .ZN(n9156) );
  NAND2_X1 U11001 ( .A1(n16217), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U11002 ( .A1(n9156), .A2(n9155), .ZN(n16219) );
  INV_X1 U11003 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n16192) );
  NAND2_X1 U11004 ( .A1(n16220), .A2(n16219), .ZN(n16218) );
  NAND2_X1 U11005 ( .A1(n16224), .A2(n16223), .ZN(n9158) );
  XNOR2_X1 U11006 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9160) );
  XOR2_X1 U11007 ( .A(n9160), .B(n9159), .Z(n16228) );
  NAND2_X1 U11008 ( .A1(n16229), .A2(n16228), .ZN(n9161) );
  XOR2_X1 U11009 ( .A(n9163), .B(n9162), .Z(n16234) );
  XOR2_X1 U11010 ( .A(n9165), .B(n9164), .Z(n9167) );
  AND2_X1 U11011 ( .A1(n9166), .A2(n9167), .ZN(n16237) );
  NOR2_X1 U11012 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n16236), .ZN(n9168) );
  NOR2_X1 U11013 ( .A1(n16237), .A2(n9168), .ZN(n9172) );
  XNOR2_X1 U11014 ( .A(n9170), .B(n9169), .ZN(n9171) );
  AND2_X1 U11015 ( .A1(n9172), .A2(n9171), .ZN(n16239) );
  NOR2_X1 U11016 ( .A1(n9172), .A2(n9171), .ZN(n16240) );
  INV_X1 U11017 ( .A(n9174), .ZN(n9175) );
  INV_X1 U11018 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13792) );
  INV_X1 U11019 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U11020 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n9178), .B1(n13771), 
        .B2(n9177), .ZN(n9181) );
  XNOR2_X1 U11021 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n9181), .ZN(n9182) );
  XOR2_X1 U11022 ( .A(n13792), .B(n9182), .Z(n16242) );
  INV_X1 U11023 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13812) );
  NAND2_X1 U11024 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n13812), .ZN(n9179) );
  OAI21_X1 U11025 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13812), .A(n9179), .ZN(
        n9189) );
  INV_X1 U11026 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11027 ( .A1(n9181), .A2(n9180), .ZN(n9184) );
  NAND2_X1 U11028 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9182), .ZN(n9183) );
  NAND2_X1 U11029 ( .A1(n9184), .A2(n9183), .ZN(n9188) );
  XNOR2_X1 U11030 ( .A(n9189), .B(n9188), .ZN(n16246) );
  NAND2_X1 U11031 ( .A1(n16247), .A2(n16246), .ZN(n9185) );
  NOR2_X1 U11032 ( .A1(n16247), .A2(n16246), .ZN(n16245) );
  AOI21_X1 U11033 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9185), .A(n16245), .ZN(
        n9187) );
  XNOR2_X1 U11034 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9186) );
  NOR2_X1 U11035 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  AOI21_X1 U11036 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13812), .A(n9190), .ZN(
        n9191) );
  NAND2_X1 U11037 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9441) );
  INV_X1 U11038 ( .A(n9441), .ZN(n9193) );
  NAND2_X1 U11039 ( .A1(n9193), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9461) );
  INV_X1 U11040 ( .A(n9461), .ZN(n9194) );
  NAND2_X1 U11041 ( .A1(n9194), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9480) );
  INV_X1 U11042 ( .A(n9480), .ZN(n9195) );
  NAND2_X1 U11043 ( .A1(n9195), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9494) );
  INV_X1 U11044 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9581) );
  INV_X1 U11045 ( .A(n9617), .ZN(n9199) );
  NAND2_X1 U11046 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9201) );
  INV_X1 U11047 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14319) );
  INV_X1 U11048 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14286) );
  INV_X1 U11049 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9785) );
  INV_X1 U11050 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9784) );
  INV_X1 U11051 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14278) );
  NAND2_X1 U11052 ( .A1(n9205), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9920) );
  INV_X1 U11053 ( .A(n9205), .ZN(n9360) );
  INV_X1 U11054 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U11055 ( .A1(n9360), .A2(n14310), .ZN(n9206) );
  NAND2_X1 U11056 ( .A1(n9920), .A2(n9206), .ZN(n14443) );
  INV_X2 U11057 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9432) );
  INV_X1 U11058 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11059 ( .A1(n9432), .A2(n9207), .ZN(n9450) );
  INV_X1 U11060 ( .A(n9450), .ZN(n9211) );
  NOR2_X1 U11061 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n9209) );
  NOR2_X1 U11062 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n9208) );
  NAND4_X1 U11063 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n9212)
         );
  INV_X1 U11064 ( .A(n9212), .ZN(n9218) );
  INV_X1 U11065 ( .A(n9422), .ZN(n9217) );
  NOR2_X1 U11066 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9215) );
  AND4_X2 U11067 ( .A1(n9215), .A2(n9214), .A3(n9556), .A4(n9555), .ZN(n9216)
         );
  NAND2_X1 U11068 ( .A1(n9673), .A2(n9219), .ZN(n9818) );
  INV_X1 U11069 ( .A(n9818), .ZN(n9223) );
  NOR2_X1 U11070 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9222) );
  NOR2_X1 U11071 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n9221) );
  NOR2_X1 U11072 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9220) );
  NAND2_X1 U11073 ( .A1(n9227), .A2(n9225), .ZN(n14765) );
  INV_X1 U11074 ( .A(n9227), .ZN(n9349) );
  INV_X1 U11075 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11076 ( .A1(n9905), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11077 ( .A1(n9906), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9231) );
  OAI211_X1 U11078 ( .C1(n10117), .C2(n9233), .A(n9232), .B(n9231), .ZN(n9234)
         );
  INV_X1 U11079 ( .A(n9234), .ZN(n9235) );
  XNOR2_X1 U11080 ( .A(n9239), .B(SI_1_), .ZN(n9374) );
  AND2_X1 U11081 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n9237) );
  NAND2_X1 U11082 ( .A1(n9244), .A2(SI_1_), .ZN(n9243) );
  NAND2_X1 U11083 ( .A1(n9238), .A2(SI_2_), .ZN(n9248) );
  INV_X1 U11084 ( .A(SI_2_), .ZN(n15873) );
  OAI21_X1 U11085 ( .B1(SI_1_), .B2(n15873), .A(n9239), .ZN(n9241) );
  OAI21_X1 U11086 ( .B1(SI_2_), .B2(n10865), .A(n9244), .ZN(n9240) );
  NAND2_X1 U11087 ( .A1(n9241), .A2(n9240), .ZN(n9247) );
  NOR2_X1 U11088 ( .A1(n9373), .A2(n15873), .ZN(n9242) );
  NAND2_X1 U11089 ( .A1(n9243), .A2(n9242), .ZN(n9246) );
  OAI211_X1 U11090 ( .C1(n9244), .C2(SI_1_), .A(n9373), .B(n15873), .ZN(n9245)
         );
  MUX2_X1 U11091 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n10831), .Z(n9398) );
  MUX2_X1 U11092 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9249), .Z(n9251) );
  INV_X1 U11093 ( .A(n9413), .ZN(n9250) );
  NAND2_X1 U11094 ( .A1(n9414), .A2(n9250), .ZN(n9253) );
  NAND2_X1 U11095 ( .A1(n9251), .A2(SI_3_), .ZN(n9252) );
  INV_X1 U11096 ( .A(n9419), .ZN(n9254) );
  MUX2_X1 U11097 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10831), .Z(n9257) );
  XNOR2_X1 U11098 ( .A(n9257), .B(SI_5_), .ZN(n9430) );
  INV_X1 U11099 ( .A(n9430), .ZN(n9256) );
  NAND2_X1 U11100 ( .A1(n9257), .A2(SI_5_), .ZN(n9258) );
  MUX2_X1 U11101 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10831), .Z(n9260) );
  NAND2_X1 U11102 ( .A1(n9260), .A2(SI_6_), .ZN(n9261) );
  MUX2_X1 U11103 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10831), .Z(n9263) );
  XNOR2_X1 U11104 ( .A(n9263), .B(SI_7_), .ZN(n9469) );
  INV_X1 U11105 ( .A(n9469), .ZN(n9262) );
  MUX2_X1 U11106 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10831), .Z(n9265) );
  XNOR2_X1 U11107 ( .A(n9265), .B(SI_8_), .ZN(n9488) );
  INV_X1 U11108 ( .A(n9488), .ZN(n9264) );
  NAND2_X1 U11109 ( .A1(n9265), .A2(SI_8_), .ZN(n9266) );
  MUX2_X1 U11110 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10831), .Z(n9268) );
  XNOR2_X1 U11111 ( .A(n9268), .B(SI_9_), .ZN(n9503) );
  INV_X1 U11112 ( .A(n9503), .ZN(n9267) );
  MUX2_X1 U11113 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10831), .Z(n9270) );
  XNOR2_X1 U11114 ( .A(n9270), .B(SI_10_), .ZN(n9519) );
  INV_X1 U11115 ( .A(n9519), .ZN(n9269) );
  NAND2_X1 U11116 ( .A1(n9270), .A2(SI_10_), .ZN(n9271) );
  MUX2_X1 U11117 ( .A(n9273), .B(n10990), .S(n10831), .Z(n9274) );
  NAND2_X1 U11118 ( .A1(n9274), .A2(n15857), .ZN(n9278) );
  INV_X1 U11119 ( .A(n9274), .ZN(n9275) );
  NAND2_X1 U11120 ( .A1(n9275), .A2(SI_11_), .ZN(n9276) );
  NAND2_X1 U11121 ( .A1(n9278), .A2(n9276), .ZN(n9536) );
  MUX2_X1 U11122 ( .A(n7684), .B(n11128), .S(n10831), .Z(n9279) );
  NAND2_X1 U11123 ( .A1(n9279), .A2(n15856), .ZN(n9282) );
  INV_X1 U11124 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U11125 ( .A1(n9280), .A2(SI_12_), .ZN(n9281) );
  MUX2_X1 U11126 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10831), .Z(n9284) );
  XNOR2_X1 U11127 ( .A(n9284), .B(n15855), .ZN(n9576) );
  INV_X1 U11128 ( .A(n9576), .ZN(n9286) );
  NAND2_X1 U11129 ( .A1(n9284), .A2(SI_13_), .ZN(n9285) );
  MUX2_X1 U11130 ( .A(n11382), .B(n11380), .S(n7434), .Z(n9287) );
  NAND2_X1 U11131 ( .A1(n9287), .A2(n15851), .ZN(n9290) );
  INV_X1 U11132 ( .A(n9287), .ZN(n9288) );
  NAND2_X1 U11133 ( .A1(n9288), .A2(SI_14_), .ZN(n9289) );
  NAND2_X1 U11134 ( .A1(n9290), .A2(n9289), .ZN(n9590) );
  MUX2_X1 U11135 ( .A(n11564), .B(n11562), .S(n7434), .Z(n9291) );
  NAND2_X1 U11136 ( .A1(n9291), .A2(n15850), .ZN(n9294) );
  INV_X1 U11137 ( .A(n9291), .ZN(n9292) );
  NAND2_X1 U11138 ( .A1(n9292), .A2(SI_15_), .ZN(n9293) );
  MUX2_X1 U11139 ( .A(n11761), .B(n11719), .S(n7434), .Z(n9295) );
  INV_X1 U11140 ( .A(n9295), .ZN(n9296) );
  NAND2_X1 U11141 ( .A1(n9296), .A2(SI_16_), .ZN(n9297) );
  MUX2_X1 U11142 ( .A(n11823), .B(n11825), .S(n7434), .Z(n9299) );
  INV_X1 U11143 ( .A(n9299), .ZN(n9300) );
  NAND2_X1 U11144 ( .A1(n9300), .A2(SI_17_), .ZN(n9301) );
  NAND2_X1 U11145 ( .A1(n9302), .A2(n9301), .ZN(n9641) );
  MUX2_X1 U11146 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7434), .Z(n9655) );
  NAND2_X1 U11147 ( .A1(n9303), .A2(n9655), .ZN(n9670) );
  MUX2_X1 U11148 ( .A(n8186), .B(n12382), .S(n7434), .Z(n9306) );
  INV_X1 U11149 ( .A(n9306), .ZN(n9307) );
  NAND2_X1 U11150 ( .A1(n9307), .A2(SI_19_), .ZN(n9308) );
  NAND2_X1 U11151 ( .A1(n9311), .A2(n9308), .ZN(n9671) );
  INV_X1 U11152 ( .A(n9671), .ZN(n9309) );
  NAND2_X1 U11153 ( .A1(n9670), .A2(n9310), .ZN(n9312) );
  NAND2_X1 U11154 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  MUX2_X1 U11155 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n7434), .Z(n9693) );
  INV_X1 U11156 ( .A(n9313), .ZN(n9314) );
  MUX2_X1 U11157 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7434), .Z(n9317) );
  XNOR2_X1 U11158 ( .A(n9317), .B(SI_21_), .ZN(n9706) );
  NAND2_X1 U11159 ( .A1(n9317), .A2(SI_21_), .ZN(n9318) );
  MUX2_X1 U11160 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7434), .Z(n9722) );
  MUX2_X1 U11161 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7434), .Z(n9739) );
  INV_X1 U11162 ( .A(n9739), .ZN(n9319) );
  AOI22_X1 U11163 ( .A1(n9721), .A2(n9723), .B1(n9319), .B2(n12258), .ZN(n9320) );
  OAI21_X1 U11164 ( .B1(n9723), .B2(n9721), .A(n12258), .ZN(n9322) );
  AND2_X1 U11165 ( .A1(SI_22_), .A2(SI_23_), .ZN(n9321) );
  AOI22_X1 U11166 ( .A1(n9322), .A2(n9739), .B1(n9722), .B2(n9321), .ZN(n9323)
         );
  INV_X1 U11167 ( .A(n9753), .ZN(n9324) );
  MUX2_X1 U11168 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7434), .Z(n9752) );
  NAND2_X1 U11169 ( .A1(n9325), .A2(SI_24_), .ZN(n9326) );
  MUX2_X1 U11170 ( .A(n7719), .B(n13107), .S(n7434), .Z(n9328) );
  NAND2_X1 U11171 ( .A1(n9328), .A2(n15644), .ZN(n9331) );
  INV_X1 U11172 ( .A(n9328), .ZN(n9329) );
  NAND2_X1 U11173 ( .A1(n9329), .A2(SI_25_), .ZN(n9330) );
  NAND2_X1 U11174 ( .A1(n9331), .A2(n9330), .ZN(n9767) );
  OAI21_X2 U11175 ( .B1(n9768), .B2(n9767), .A(n9331), .ZN(n9781) );
  MUX2_X1 U11176 ( .A(n7735), .B(n14782), .S(n7434), .Z(n9332) );
  NAND2_X1 U11177 ( .A1(n9332), .A2(n12916), .ZN(n9335) );
  INV_X1 U11178 ( .A(n9332), .ZN(n9333) );
  NAND2_X1 U11179 ( .A1(n9333), .A2(SI_26_), .ZN(n9334) );
  NAND2_X1 U11180 ( .A1(n9781), .A2(n9780), .ZN(n9336) );
  MUX2_X1 U11181 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7434), .Z(n9337) );
  XNOR2_X1 U11182 ( .A(n9337), .B(SI_27_), .ZN(n9354) );
  NAND2_X1 U11183 ( .A1(n9337), .A2(SI_27_), .ZN(n9338) );
  MUX2_X1 U11184 ( .A(n7738), .B(n14775), .S(n7434), .Z(n9339) );
  NAND2_X1 U11185 ( .A1(n9339), .A2(n15637), .ZN(n9797) );
  INV_X1 U11186 ( .A(n9339), .ZN(n9340) );
  NAND2_X1 U11187 ( .A1(n9340), .A2(SI_28_), .ZN(n9341) );
  NAND2_X1 U11188 ( .A1(n9797), .A2(n9341), .ZN(n9798) );
  NAND2_X1 U11189 ( .A1(n9344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U11190 ( .A1(n9345), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11191 ( .A1(n9348), .A2(n9347), .ZN(n9350) );
  NAND2_X1 U11192 ( .A1(n9350), .A2(n9349), .ZN(n9904) );
  INV_X4 U11193 ( .A(n10113), .ZN(n10135) );
  NAND2_X1 U11194 ( .A1(n14772), .A2(n10135), .ZN(n9353) );
  OR2_X1 U11195 ( .A1(n10137), .A2(n14775), .ZN(n9352) );
  NAND2_X2 U11196 ( .A1(n9353), .A2(n9352), .ZN(n14655) );
  INV_X1 U11197 ( .A(n9354), .ZN(n9355) );
  NAND2_X1 U11198 ( .A1(n14776), .A2(n10135), .ZN(n9358) );
  OR2_X1 U11199 ( .A1(n10137), .A2(n14777), .ZN(n9357) );
  NAND2_X2 U11200 ( .A1(n9358), .A2(n9357), .ZN(n14658) );
  NAND2_X1 U11201 ( .A1(n9787), .A2(n14278), .ZN(n9359) );
  NAND2_X1 U11202 ( .A1(n9360), .A2(n9359), .ZN(n14462) );
  OR2_X1 U11203 ( .A1(n14462), .A2(n9802), .ZN(n9366) );
  INV_X1 U11204 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11205 ( .A1(n9906), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11206 ( .A1(n9905), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U11207 ( .C1(n10117), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9364)
         );
  INV_X1 U11208 ( .A(n9364), .ZN(n9365) );
  INV_X1 U11209 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11090) );
  INV_X1 U11210 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9367) );
  OR2_X1 U11211 ( .A1(n9392), .A2(n9367), .ZN(n9370) );
  INV_X1 U11212 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9368) );
  XNOR2_X1 U11213 ( .A(n9373), .B(n9374), .ZN(n10851) );
  NAND2_X1 U11215 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9375) );
  XNOR2_X1 U11216 ( .A(n9375), .B(P2_IR_REG_1__SCAN_IN), .ZN(n14419) );
  NAND2_X1 U11217 ( .A1(n9421), .A2(n14419), .ZN(n9376) );
  OAI211_X2 U11218 ( .C1(n10113), .C2(n10851), .A(n9377), .B(n9376), .ZN(
        n12000) );
  INV_X1 U11219 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11931) );
  INV_X1 U11220 ( .A(n9390), .ZN(n9378) );
  INV_X1 U11221 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9379) );
  INV_X1 U11222 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11075) );
  OR2_X1 U11223 ( .A1(n9380), .A2(n11075), .ZN(n9381) );
  INV_X1 U11224 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n11079) );
  AND2_X1 U11225 ( .A1(n7635), .A2(n14412), .ZN(n11197) );
  OR2_X1 U11226 ( .A1(n14411), .A2(n12000), .ZN(n9387) );
  INV_X1 U11227 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9389) );
  OR2_X1 U11228 ( .A1(n9390), .A2(n9389), .ZN(n9395) );
  INV_X1 U11229 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11535) );
  INV_X1 U11230 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11534) );
  OR2_X1 U11231 ( .A1(n9392), .A2(n11534), .ZN(n9393) );
  OR2_X1 U11232 ( .A1(n9399), .A2(n9560), .ZN(n9400) );
  XNOR2_X1 U11233 ( .A(n9400), .B(P2_IR_REG_2__SCAN_IN), .ZN(n11106) );
  NAND2_X1 U11234 ( .A1(n9421), .A2(n11106), .ZN(n9403) );
  OR2_X1 U11235 ( .A1(n9401), .A2(n10841), .ZN(n9402) );
  OAI211_X2 U11236 ( .C1(n10113), .C2(n10840), .A(n9403), .B(n9402), .ZN(
        n11279) );
  XNOR2_X1 U11237 ( .A(n9929), .B(n11279), .ZN(n11280) );
  INV_X1 U11238 ( .A(n11280), .ZN(n11274) );
  OR2_X1 U11239 ( .A1(n9929), .A2(n11279), .ZN(n9404) );
  NAND2_X1 U11240 ( .A1(n9405), .A2(n9404), .ZN(n11248) );
  NAND2_X1 U11241 ( .A1(n9388), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9410) );
  INV_X1 U11242 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9406) );
  OR2_X1 U11243 ( .A1(n9390), .A2(n9406), .ZN(n9409) );
  INV_X1 U11244 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11093) );
  OR2_X1 U11245 ( .A1(n9391), .A2(n11093), .ZN(n9408) );
  OR2_X1 U11246 ( .A1(n9802), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9407) );
  NAND4_X2 U11247 ( .A1(n9407), .A2(n9409), .A3(n9408), .A4(n9410), .ZN(n14409) );
  NAND2_X1 U11248 ( .A1(n9422), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9412) );
  INV_X1 U11249 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9411) );
  XNOR2_X1 U11250 ( .A(n9412), .B(n9411), .ZN(n16067) );
  XNOR2_X1 U11251 ( .A(n9414), .B(n9413), .ZN(n10842) );
  NAND2_X1 U11252 ( .A1(n11248), .A2(n10191), .ZN(n9418) );
  OR2_X1 U11253 ( .A1(n14409), .A2(n11249), .ZN(n9417) );
  NAND2_X1 U11254 ( .A1(n9418), .A2(n9417), .ZN(n11395) );
  NAND2_X1 U11255 ( .A1(n10837), .A2(n10135), .ZN(n9424) );
  OR2_X1 U11256 ( .A1(n9422), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U11257 ( .A1(n9452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9434) );
  XNOR2_X1 U11258 ( .A(n9434), .B(P2_IR_REG_4__SCAN_IN), .ZN(n16078) );
  AOI22_X1 U11259 ( .A1(n9754), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9678), .B2(
        n16078), .ZN(n9423) );
  OAI21_X1 U11260 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9441), .ZN(n11750) );
  OR2_X1 U11261 ( .A1(n9802), .A2(n11750), .ZN(n9426) );
  INV_X1 U11262 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11751) );
  OR2_X1 U11263 ( .A1(n9391), .A2(n11751), .ZN(n9425) );
  NAND2_X1 U11264 ( .A1(n11395), .A2(n11396), .ZN(n9429) );
  OR2_X1 U11265 ( .A1(n14408), .A2(n11404), .ZN(n9428) );
  XNOR2_X1 U11266 ( .A(n9431), .B(n9430), .ZN(n10854) );
  NAND2_X1 U11267 ( .A1(n10854), .A2(n10135), .ZN(n9438) );
  NAND2_X1 U11268 ( .A1(n9434), .A2(n9433), .ZN(n9435) );
  NAND2_X1 U11269 ( .A1(n9435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9436) );
  XNOR2_X1 U11270 ( .A(n9436), .B(P2_IR_REG_5__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U11271 ( .A1(n9754), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9678), .B2(
        n11112), .ZN(n9437) );
  NAND2_X1 U11272 ( .A1(n9378), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9446) );
  INV_X1 U11273 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9439) );
  OR2_X1 U11274 ( .A1(n10117), .A2(n9439), .ZN(n9445) );
  INV_X1 U11275 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11276 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  NAND2_X1 U11277 ( .A1(n9461), .A2(n9442), .ZN(n11518) );
  OR2_X1 U11278 ( .A1(n9802), .A2(n11518), .ZN(n9444) );
  INV_X1 U11279 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11516) );
  OR2_X1 U11280 ( .A1(n10118), .A2(n11516), .ZN(n9443) );
  NOR2_X1 U11281 ( .A1(n11517), .A2(n14407), .ZN(n9447) );
  NAND2_X1 U11282 ( .A1(n11517), .A2(n14407), .ZN(n9448) );
  NAND2_X1 U11283 ( .A1(n10878), .A2(n10135), .ZN(n9458) );
  CLKBUF_X1 U11284 ( .A(n9450), .Z(n9451) );
  NOR2_X1 U11285 ( .A1(n9452), .A2(n9451), .ZN(n9455) );
  NOR2_X1 U11286 ( .A1(n9455), .A2(n9560), .ZN(n9453) );
  MUX2_X1 U11287 ( .A(n9560), .B(n9453), .S(P2_IR_REG_6__SCAN_IN), .Z(n9456)
         );
  INV_X1 U11288 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9454) );
  OR2_X1 U11289 ( .A1(n9456), .A2(n9473), .ZN(n16106) );
  INV_X1 U11290 ( .A(n16106), .ZN(n11114) );
  AOI22_X1 U11291 ( .A1(n9754), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9678), .B2(
        n11114), .ZN(n9457) );
  NAND2_X1 U11292 ( .A1(n9685), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9467) );
  INV_X1 U11293 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9459) );
  OR2_X1 U11294 ( .A1(n10118), .A2(n9459), .ZN(n9466) );
  INV_X1 U11295 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U11296 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  NAND2_X1 U11297 ( .A1(n9480), .A2(n9462), .ZN(n11980) );
  OR2_X1 U11298 ( .A1(n9802), .A2(n11980), .ZN(n9465) );
  INV_X1 U11299 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9463) );
  OR2_X1 U11300 ( .A1(n10120), .A2(n9463), .ZN(n9464) );
  NAND4_X1 U11301 ( .A1(n9467), .A2(n9466), .A3(n9465), .A4(n9464), .ZN(n14406) );
  XNOR2_X1 U11302 ( .A(n11979), .B(n14406), .ZN(n10193) );
  OR2_X1 U11303 ( .A1(n11979), .A2(n14406), .ZN(n9468) );
  XNOR2_X1 U11304 ( .A(n9470), .B(n9469), .ZN(n10884) );
  NAND2_X1 U11305 ( .A1(n10884), .A2(n10135), .ZN(n9477) );
  NOR2_X1 U11306 ( .A1(n9473), .A2(n9560), .ZN(n9471) );
  MUX2_X1 U11307 ( .A(n9560), .B(n9471), .S(P2_IR_REG_7__SCAN_IN), .Z(n9475)
         );
  INV_X1 U11308 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11309 ( .A1(n9473), .A2(n9472), .ZN(n9505) );
  INV_X1 U11310 ( .A(n9505), .ZN(n9474) );
  INV_X1 U11311 ( .A(n16118), .ZN(n11116) );
  AOI22_X1 U11312 ( .A1(n9754), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9678), .B2(
        n11116), .ZN(n9476) );
  NAND2_X1 U11313 ( .A1(n9477), .A2(n9476), .ZN(n12021) );
  NAND2_X1 U11314 ( .A1(n9906), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9486) );
  INV_X1 U11315 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9478) );
  OR2_X1 U11316 ( .A1(n10117), .A2(n9478), .ZN(n9485) );
  INV_X1 U11317 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U11318 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  NAND2_X1 U11319 ( .A1(n9494), .A2(n9481), .ZN(n13166) );
  OR2_X1 U11320 ( .A1(n9802), .A2(n13166), .ZN(n9484) );
  INV_X1 U11321 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9482) );
  OR2_X1 U11322 ( .A1(n10118), .A2(n9482), .ZN(n9483) );
  NAND4_X1 U11323 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n14405) );
  XNOR2_X1 U11324 ( .A(n12021), .B(n14405), .ZN(n10194) );
  NAND2_X1 U11325 ( .A1(n12021), .A2(n14405), .ZN(n9487) );
  NAND2_X1 U11326 ( .A1(n12011), .A2(n9487), .ZN(n11879) );
  XNOR2_X1 U11327 ( .A(n9489), .B(n9488), .ZN(n10888) );
  NAND2_X1 U11328 ( .A1(n10888), .A2(n10135), .ZN(n9492) );
  NAND2_X1 U11329 ( .A1(n9505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9490) );
  XNOR2_X1 U11330 ( .A(n9490), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U11331 ( .A1(n9754), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9678), .B2(
        n11119), .ZN(n9491) );
  NAND2_X1 U11332 ( .A1(n9492), .A2(n9491), .ZN(n12050) );
  NAND2_X1 U11333 ( .A1(n9906), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9499) );
  INV_X1 U11334 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11118) );
  OR2_X1 U11335 ( .A1(n10117), .A2(n11118), .ZN(n9498) );
  NAND2_X1 U11336 ( .A1(n9494), .A2(n9493), .ZN(n9495) );
  NAND2_X1 U11337 ( .A1(n9510), .A2(n9495), .ZN(n12059) );
  OR2_X1 U11338 ( .A1(n9802), .A2(n12059), .ZN(n9497) );
  INV_X1 U11339 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11880) );
  OR2_X1 U11340 ( .A1(n10118), .A2(n11880), .ZN(n9496) );
  NAND4_X1 U11341 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n14404) );
  XNOR2_X1 U11342 ( .A(n12050), .B(n14404), .ZN(n11878) );
  INV_X1 U11343 ( .A(n11878), .ZN(n9500) );
  NAND2_X1 U11344 ( .A1(n11879), .A2(n9500), .ZN(n9502) );
  NAND2_X1 U11345 ( .A1(n12050), .A2(n14404), .ZN(n9501) );
  NAND2_X1 U11346 ( .A1(n9502), .A2(n9501), .ZN(n12103) );
  NAND2_X1 U11347 ( .A1(n10941), .A2(n10135), .ZN(n9507) );
  NAND2_X1 U11348 ( .A1(n9558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U11349 ( .A(n9521), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U11350 ( .A1(n9754), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9678), .B2(
        n11231), .ZN(n9506) );
  NAND2_X1 U11351 ( .A1(n9906), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9516) );
  INV_X1 U11352 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9508) );
  OR2_X1 U11353 ( .A1(n10117), .A2(n9508), .ZN(n9515) );
  INV_X1 U11354 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U11355 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  NAND2_X1 U11356 ( .A1(n9528), .A2(n9511), .ZN(n12109) );
  OR2_X1 U11357 ( .A1(n9802), .A2(n12109), .ZN(n9514) );
  INV_X1 U11358 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9512) );
  OR2_X1 U11359 ( .A1(n10118), .A2(n9512), .ZN(n9513) );
  NAND4_X1 U11360 ( .A1(n9516), .A2(n9515), .A3(n9514), .A4(n9513), .ZN(n14403) );
  XNOR2_X1 U11361 ( .A(n12259), .B(n12408), .ZN(n12102) );
  NAND2_X1 U11362 ( .A1(n12103), .A2(n12102), .ZN(n9518) );
  NAND2_X1 U11363 ( .A1(n12259), .A2(n14403), .ZN(n9517) );
  XNOR2_X1 U11364 ( .A(n9520), .B(n9519), .ZN(n10946) );
  NAND2_X1 U11365 ( .A1(n10946), .A2(n10135), .ZN(n9526) );
  NAND2_X1 U11366 ( .A1(n9521), .A2(n9555), .ZN(n9522) );
  NAND2_X1 U11367 ( .A1(n9522), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U11368 ( .A1(n9523), .A2(n9556), .ZN(n9540) );
  OR2_X1 U11369 ( .A1(n9523), .A2(n9556), .ZN(n9524) );
  AOI22_X1 U11370 ( .A1(n9754), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n16187), 
        .B2(n9678), .ZN(n9525) );
  NAND2_X1 U11371 ( .A1(n9906), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9533) );
  INV_X1 U11372 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11234) );
  OR2_X1 U11373 ( .A1(n10117), .A2(n11234), .ZN(n9532) );
  NAND2_X1 U11374 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  NAND2_X1 U11375 ( .A1(n9546), .A2(n9529), .ZN(n12352) );
  OR2_X1 U11376 ( .A1(n9802), .A2(n12352), .ZN(n9531) );
  INV_X1 U11377 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11229) );
  OR2_X1 U11378 ( .A1(n10118), .A2(n11229), .ZN(n9530) );
  NAND4_X1 U11379 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n14402) );
  AND2_X1 U11380 ( .A1(n12400), .A2(n14402), .ZN(n9534) );
  OR2_X1 U11381 ( .A1(n12400), .A2(n14402), .ZN(n9535) );
  NAND2_X1 U11382 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND2_X1 U11383 ( .A1(n9539), .A2(n9538), .ZN(n10986) );
  NAND2_X1 U11384 ( .A1(n10986), .A2(n10135), .ZN(n9543) );
  NAND2_X1 U11385 ( .A1(n9540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9541) );
  XNOR2_X1 U11386 ( .A(n9541), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U11387 ( .A1(n11236), .A2(n9678), .B1(n9754), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U11388 ( .A1(n9388), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9551) );
  INV_X1 U11389 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9544) );
  OR2_X1 U11390 ( .A1(n10120), .A2(n9544), .ZN(n9550) );
  INV_X1 U11391 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U11392 ( .A1(n9546), .A2(n9545), .ZN(n9547) );
  NAND2_X1 U11393 ( .A1(n9569), .A2(n9547), .ZN(n12491) );
  OR2_X1 U11394 ( .A1(n9802), .A2(n12491), .ZN(n9549) );
  INV_X1 U11395 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12322) );
  OR2_X1 U11396 ( .A1(n10118), .A2(n12322), .ZN(n9548) );
  NAND4_X1 U11397 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n14401) );
  XNOR2_X1 U11398 ( .A(n12487), .B(n12691), .ZN(n12320) );
  NAND2_X1 U11399 ( .A1(n12487), .A2(n14401), .ZN(n9552) );
  XNOR2_X1 U11400 ( .A(n9553), .B(n8502), .ZN(n11085) );
  NAND2_X1 U11401 ( .A1(n11085), .A2(n10135), .ZN(n9567) );
  INV_X1 U11402 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9554) );
  NAND3_X1 U11403 ( .A1(n9556), .A2(n9555), .A3(n9554), .ZN(n9557) );
  NOR2_X1 U11404 ( .A1(n9562), .A2(n9560), .ZN(n9559) );
  MUX2_X1 U11405 ( .A(n9560), .B(n9559), .S(P2_IR_REG_12__SCAN_IN), .Z(n9564)
         );
  INV_X1 U11406 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9561) );
  NAND2_X1 U11407 ( .A1(n9562), .A2(n9561), .ZN(n9592) );
  INV_X1 U11408 ( .A(n9592), .ZN(n9563) );
  OAI22_X1 U11409 ( .A1(n11318), .A2(n8042), .B1(n10137), .B2(n11128), .ZN(
        n9565) );
  INV_X1 U11410 ( .A(n9565), .ZN(n9566) );
  NAND2_X1 U11411 ( .A1(n9906), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9574) );
  INV_X1 U11412 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11314) );
  OR2_X1 U11413 ( .A1(n10117), .A2(n11314), .ZN(n9573) );
  NAND2_X1 U11414 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  NAND2_X1 U11415 ( .A1(n9582), .A2(n9570), .ZN(n16456) );
  OR2_X1 U11416 ( .A1(n9802), .A2(n16456), .ZN(n9572) );
  INV_X1 U11417 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n16457) );
  OR2_X1 U11418 ( .A1(n10118), .A2(n16457), .ZN(n9571) );
  NAND4_X1 U11419 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(n14400) );
  XNOR2_X1 U11420 ( .A(n16462), .B(n14400), .ZN(n10197) );
  NAND2_X1 U11421 ( .A1(n16462), .A2(n14400), .ZN(n9575) );
  NAND2_X1 U11422 ( .A1(n11182), .A2(n10135), .ZN(n9580) );
  NAND2_X1 U11423 ( .A1(n9592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U11424 ( .A(n9578), .B(P2_IR_REG_13__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U11425 ( .A1(n12067), .A2(n9678), .B1(n9754), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U11426 ( .A1(n9582), .A2(n9581), .ZN(n9583) );
  NAND2_X1 U11427 ( .A1(n9597), .A2(n9583), .ZN(n12777) );
  OR2_X1 U11428 ( .A1(n9802), .A2(n12777), .ZN(n9588) );
  NAND2_X1 U11429 ( .A1(n9685), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9587) );
  INV_X1 U11430 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12071) );
  OR2_X1 U11431 ( .A1(n10118), .A2(n12071), .ZN(n9586) );
  INV_X1 U11432 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9584) );
  OR2_X1 U11433 ( .A1(n10120), .A2(n9584), .ZN(n9585) );
  NAND4_X1 U11434 ( .A1(n9588), .A2(n9587), .A3(n9586), .A4(n9585), .ZN(n14399) );
  OR2_X1 U11435 ( .A1(n12990), .A2(n14399), .ZN(n9589) );
  XNOR2_X1 U11436 ( .A(n9591), .B(n9590), .ZN(n11378) );
  NAND2_X1 U11437 ( .A1(n11378), .A2(n10135), .ZN(n9595) );
  NAND2_X1 U11438 ( .A1(n9610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9593) );
  XNOR2_X1 U11439 ( .A(n9593), .B(P2_IR_REG_14__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U11440 ( .A1(n16158), .A2(n9678), .B1(n9754), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9594) );
  INV_X1 U11441 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11442 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  NAND2_X1 U11443 ( .A1(n9617), .A2(n9598), .ZN(n12881) );
  NAND2_X1 U11444 ( .A1(n9905), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9599) );
  OAI21_X1 U11445 ( .B1(n12881), .B2(n9802), .A(n9599), .ZN(n9603) );
  INV_X1 U11446 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9600) );
  NOR2_X1 U11447 ( .A1(n10120), .A2(n9600), .ZN(n9602) );
  INV_X1 U11448 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12068) );
  NOR2_X1 U11449 ( .A1(n10117), .A2(n12068), .ZN(n9601) );
  INV_X1 U11450 ( .A(n14398), .ZN(n13064) );
  XNOR2_X1 U11451 ( .A(n14732), .B(n13064), .ZN(n12883) );
  NAND2_X1 U11452 ( .A1(n12884), .A2(n12883), .ZN(n9605) );
  NAND2_X1 U11453 ( .A1(n14732), .A2(n14398), .ZN(n9604) );
  NAND2_X1 U11454 ( .A1(n9605), .A2(n9604), .ZN(n13072) );
  INV_X1 U11455 ( .A(n13072), .ZN(n9627) );
  OR2_X1 U11456 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  NAND2_X1 U11457 ( .A1(n9609), .A2(n9608), .ZN(n11561) );
  NAND2_X1 U11458 ( .A1(n11561), .A2(n10135), .ZN(n9615) );
  OAI21_X1 U11459 ( .B1(n9610), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9612) );
  INV_X1 U11460 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9611) );
  XNOR2_X1 U11461 ( .A(n9612), .B(n9611), .ZN(n12273) );
  OAI22_X1 U11462 ( .A1(n12273), .A2(n8042), .B1(n10137), .B2(n11562), .ZN(
        n9613) );
  INV_X1 U11463 ( .A(n9613), .ZN(n9614) );
  INV_X1 U11464 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9625) );
  INV_X1 U11465 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U11466 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  NAND2_X1 U11467 ( .A1(n9636), .A2(n9618), .ZN(n13063) );
  OR2_X1 U11468 ( .A1(n13063), .A2(n9802), .ZN(n9624) );
  INV_X1 U11469 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9619) );
  OR2_X1 U11470 ( .A1(n10117), .A2(n9619), .ZN(n9622) );
  INV_X1 U11471 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9620) );
  OR2_X1 U11472 ( .A1(n10118), .A2(n9620), .ZN(n9621) );
  AND2_X1 U11473 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  OAI211_X1 U11474 ( .C1(n10120), .C2(n9625), .A(n9624), .B(n9623), .ZN(n14397) );
  XNOR2_X1 U11475 ( .A(n14728), .B(n14397), .ZN(n13073) );
  OR2_X1 U11476 ( .A1(n14728), .A2(n14397), .ZN(n9628) );
  XNOR2_X1 U11477 ( .A(n9630), .B(n9629), .ZN(n11718) );
  NAND2_X1 U11478 ( .A1(n11718), .A2(n10135), .ZN(n9634) );
  NAND2_X1 U11479 ( .A1(n9631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9632) );
  XNOR2_X1 U11480 ( .A(n9632), .B(P2_IR_REG_16__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U11481 ( .A1(n9754), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9678), 
        .B2(n12518), .ZN(n9633) );
  NAND2_X1 U11482 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NAND2_X1 U11483 ( .A1(n9648), .A2(n9637), .ZN(n13155) );
  AOI22_X1 U11484 ( .A1(n9685), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9906), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U11485 ( .A1(n9905), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9638) );
  OAI211_X1 U11486 ( .C1(n13155), .C2(n9802), .A(n9639), .B(n9638), .ZN(n14396) );
  XNOR2_X1 U11487 ( .A(n14719), .B(n14396), .ZN(n13086) );
  INV_X1 U11488 ( .A(n13086), .ZN(n13089) );
  NAND2_X1 U11489 ( .A1(n14719), .A2(n14396), .ZN(n9640) );
  NAND2_X1 U11490 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U11491 ( .A1(n9644), .A2(n9643), .ZN(n11822) );
  NAND2_X1 U11492 ( .A1(n11822), .A2(n10135), .ZN(n9646) );
  NAND2_X1 U11493 ( .A1(n9819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U11494 ( .A(n9657), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U11495 ( .A1(n9754), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9678), 
        .B2(n12832), .ZN(n9645) );
  INV_X1 U11496 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14633) );
  INV_X1 U11497 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U11498 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  NAND2_X1 U11499 ( .A1(n9683), .A2(n9649), .ZN(n14632) );
  OR2_X1 U11500 ( .A1(n14632), .A2(n9802), .ZN(n9651) );
  AOI22_X1 U11501 ( .A1(n9685), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9906), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n9650) );
  OAI211_X1 U11502 ( .C1(n10118), .C2(n14633), .A(n9651), .B(n9650), .ZN(
        n14601) );
  INV_X1 U11503 ( .A(n14601), .ZN(n13156) );
  XNOR2_X1 U11504 ( .A(n14714), .B(n13156), .ZN(n14636) );
  INV_X1 U11505 ( .A(n14636), .ZN(n9652) );
  OR2_X1 U11506 ( .A1(n14714), .A2(n14601), .ZN(n9653) );
  NAND2_X1 U11507 ( .A1(n9654), .A2(n9653), .ZN(n14608) );
  NAND2_X1 U11508 ( .A1(n12164), .A2(n10135), .ZN(n9661) );
  INV_X1 U11509 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U11510 ( .A1(n9657), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U11511 ( .A1(n9658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9659) );
  XNOR2_X1 U11512 ( .A(n9659), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U11513 ( .A1(n9754), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9678), 
        .B2(n12827), .ZN(n9660) );
  XNOR2_X1 U11514 ( .A(n9683), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U11515 ( .A1(n14612), .A2(n9789), .ZN(n9667) );
  INV_X1 U11516 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U11517 ( .A1(n9906), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U11518 ( .A1(n9685), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9662) );
  OAI211_X1 U11519 ( .C1(n9664), .C2(n9391), .A(n9663), .B(n9662), .ZN(n9665)
         );
  INV_X1 U11520 ( .A(n9665), .ZN(n9666) );
  NAND2_X1 U11521 ( .A1(n9667), .A2(n9666), .ZN(n14582) );
  XNOR2_X1 U11522 ( .A(n14709), .B(n14582), .ZN(n10200) );
  OR2_X1 U11523 ( .A1(n14709), .A2(n14582), .ZN(n9668) );
  NAND2_X1 U11524 ( .A1(n9670), .A2(n9669), .ZN(n9672) );
  XNOR2_X1 U11525 ( .A(n9672), .B(n9671), .ZN(n12381) );
  NAND2_X1 U11526 ( .A1(n12381), .A2(n10135), .ZN(n9680) );
  INV_X1 U11527 ( .A(n9673), .ZN(n9674) );
  OAI21_X2 U11528 ( .B1(n9819), .B2(n9674), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9676) );
  NAND2_X1 U11529 ( .A1(n9676), .A2(n9675), .ZN(n9834) );
  AOI22_X1 U11530 ( .A1(n9754), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n14444), 
        .B2(n9678), .ZN(n9679) );
  INV_X1 U11531 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9682) );
  INV_X1 U11532 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9681) );
  OAI21_X1 U11533 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  AND2_X1 U11534 ( .A1(n9684), .A2(n9697), .ZN(n14591) );
  NAND2_X1 U11535 ( .A1(n14591), .A2(n9789), .ZN(n9691) );
  INV_X1 U11536 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U11537 ( .A1(n9906), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9687) );
  NAND2_X1 U11538 ( .A1(n9685), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9686) );
  OAI211_X1 U11539 ( .C1(n9688), .C2(n10118), .A(n9687), .B(n9686), .ZN(n9689)
         );
  INV_X1 U11540 ( .A(n9689), .ZN(n9690) );
  NAND2_X1 U11541 ( .A1(n9691), .A2(n9690), .ZN(n14605) );
  XNOR2_X1 U11542 ( .A(n14704), .B(n14605), .ZN(n10202) );
  NAND2_X1 U11543 ( .A1(n14704), .A2(n14605), .ZN(n9692) );
  XNOR2_X1 U11544 ( .A(n9694), .B(n9693), .ZN(n12596) );
  NAND2_X1 U11545 ( .A1(n12596), .A2(n10135), .ZN(n9696) );
  OR2_X1 U11546 ( .A1(n10137), .A2(n13174), .ZN(n9695) );
  NAND2_X2 U11547 ( .A1(n9696), .A2(n9695), .ZN(n14700) );
  INV_X1 U11548 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14354) );
  NAND2_X1 U11549 ( .A1(n9697), .A2(n14354), .ZN(n9698) );
  NAND2_X1 U11550 ( .A1(n9710), .A2(n9698), .ZN(n14572) );
  OR2_X1 U11551 ( .A1(n14572), .A2(n9802), .ZN(n9704) );
  INV_X1 U11552 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U11553 ( .A1(n9906), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U11554 ( .A1(n9905), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9699) );
  OAI211_X1 U11555 ( .C1(n10117), .C2(n9701), .A(n9700), .B(n9699), .ZN(n9702)
         );
  INV_X1 U11556 ( .A(n9702), .ZN(n9703) );
  NAND2_X1 U11557 ( .A1(n9704), .A2(n9703), .ZN(n14584) );
  AND2_X1 U11558 ( .A1(n14700), .A2(n14584), .ZN(n9705) );
  XNOR2_X1 U11559 ( .A(n9707), .B(n9706), .ZN(n12728) );
  NAND2_X1 U11560 ( .A1(n12728), .A2(n10135), .ZN(n9709) );
  OR2_X1 U11561 ( .A1(n10137), .A2(n12733), .ZN(n9708) );
  NAND2_X1 U11562 ( .A1(n9710), .A2(n14319), .ZN(n9711) );
  AND2_X1 U11563 ( .A1(n9727), .A2(n9711), .ZN(n14318) );
  NAND2_X1 U11564 ( .A1(n14318), .A2(n9789), .ZN(n9717) );
  INV_X1 U11565 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9714) );
  NAND2_X1 U11566 ( .A1(n9905), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U11567 ( .A1(n9906), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9712) );
  OAI211_X1 U11568 ( .C1(n10117), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9715)
         );
  INV_X1 U11569 ( .A(n9715), .ZN(n9716) );
  NAND2_X1 U11570 ( .A1(n9717), .A2(n9716), .ZN(n14538) );
  NOR2_X1 U11571 ( .A1(n14690), .A2(n14538), .ZN(n9718) );
  NAND2_X1 U11572 ( .A1(n14690), .A2(n14538), .ZN(n9719) );
  NAND2_X1 U11573 ( .A1(n10599), .A2(n9722), .ZN(n9738) );
  INV_X1 U11574 ( .A(n10599), .ZN(n9724) );
  OR2_X1 U11575 ( .A1(n10137), .A2(n12843), .ZN(n9725) );
  NAND2_X2 U11576 ( .A1(n9726), .A2(n9725), .ZN(n14686) );
  INV_X1 U11577 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14361) );
  NAND2_X1 U11578 ( .A1(n9727), .A2(n14361), .ZN(n9728) );
  NAND2_X1 U11579 ( .A1(n9744), .A2(n9728), .ZN(n14542) );
  OR2_X1 U11580 ( .A1(n14542), .A2(n9802), .ZN(n9734) );
  INV_X1 U11581 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U11582 ( .A1(n9906), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U11583 ( .A1(n9905), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9729) );
  OAI211_X1 U11584 ( .C1(n10117), .C2(n9731), .A(n9730), .B(n9729), .ZN(n9732)
         );
  INV_X1 U11585 ( .A(n9732), .ZN(n9733) );
  NAND2_X1 U11586 ( .A1(n9734), .A2(n9733), .ZN(n14552) );
  INV_X1 U11587 ( .A(n14552), .ZN(n14321) );
  NAND2_X1 U11588 ( .A1(n14686), .A2(n14552), .ZN(n9735) );
  NAND2_X1 U11589 ( .A1(n9736), .A2(SI_22_), .ZN(n9737) );
  XNOR2_X1 U11590 ( .A(n9739), .B(SI_23_), .ZN(n9740) );
  NAND2_X1 U11591 ( .A1(n13028), .A2(n10135), .ZN(n9743) );
  NAND2_X1 U11592 ( .A1(n9754), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U11593 ( .A1(n9744), .A2(n14286), .ZN(n9745) );
  AND2_X1 U11594 ( .A1(n9758), .A2(n9745), .ZN(n14529) );
  NAND2_X1 U11595 ( .A1(n14529), .A2(n9789), .ZN(n9751) );
  INV_X1 U11596 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U11597 ( .A1(n9906), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U11598 ( .A1(n9905), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9746) );
  OAI211_X1 U11599 ( .C1(n10117), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9749)
         );
  INV_X1 U11600 ( .A(n9749), .ZN(n9750) );
  NAND2_X1 U11601 ( .A1(n9751), .A2(n9750), .ZN(n14537) );
  OR2_X1 U11602 ( .A1(n14530), .A2(n14537), .ZN(n10205) );
  NAND2_X1 U11603 ( .A1(n14530), .A2(n14537), .ZN(n10204) );
  XNOR2_X1 U11604 ( .A(n9753), .B(n9752), .ZN(n13032) );
  NAND2_X1 U11605 ( .A1(n13032), .A2(n10135), .ZN(n9756) );
  NAND2_X1 U11606 ( .A1(n9754), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9755) );
  INV_X1 U11607 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U11608 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  NAND2_X1 U11609 ( .A1(n9786), .A2(n9759), .ZN(n14345) );
  OR2_X1 U11610 ( .A1(n14345), .A2(n9802), .ZN(n9765) );
  INV_X1 U11611 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9762) );
  NAND2_X1 U11612 ( .A1(n9906), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11613 ( .A1(n9905), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9760) );
  OAI211_X1 U11614 ( .C1(n10117), .C2(n9762), .A(n9761), .B(n9760), .ZN(n9763)
         );
  INV_X1 U11615 ( .A(n9763), .ZN(n9764) );
  XNOR2_X1 U11616 ( .A(n14675), .B(n14523), .ZN(n14502) );
  INV_X1 U11617 ( .A(n14502), .ZN(n14510) );
  NAND2_X1 U11618 ( .A1(n14511), .A2(n14510), .ZN(n14509) );
  NAND2_X1 U11619 ( .A1(n14675), .A2(n14523), .ZN(n9766) );
  NAND2_X1 U11620 ( .A1(n14509), .A2(n9766), .ZN(n14486) );
  XNOR2_X1 U11621 ( .A(n9768), .B(n9767), .ZN(n13102) );
  NAND2_X1 U11622 ( .A1(n13102), .A2(n10135), .ZN(n9770) );
  OR2_X1 U11623 ( .A1(n10137), .A2(n13107), .ZN(n9769) );
  XNOR2_X1 U11624 ( .A(n9786), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U11625 ( .A1(n14493), .A2(n9789), .ZN(n9776) );
  INV_X1 U11626 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U11627 ( .A1(n9906), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U11628 ( .A1(n9905), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9771) );
  OAI211_X1 U11629 ( .C1(n10117), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9774)
         );
  INV_X1 U11630 ( .A(n9774), .ZN(n9775) );
  OR2_X1 U11631 ( .A1(n14671), .A2(n14474), .ZN(n9777) );
  NAND2_X1 U11632 ( .A1(n14486), .A2(n9777), .ZN(n9779) );
  NAND2_X1 U11633 ( .A1(n14671), .A2(n14474), .ZN(n9778) );
  XNOR2_X1 U11634 ( .A(n9781), .B(n9780), .ZN(n14779) );
  NAND2_X1 U11635 ( .A1(n14779), .A2(n10135), .ZN(n9783) );
  OR2_X1 U11636 ( .A1(n10137), .A2(n14782), .ZN(n9782) );
  OAI21_X1 U11637 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9788) );
  AND2_X1 U11638 ( .A1(n9788), .A2(n9787), .ZN(n14478) );
  NAND2_X1 U11639 ( .A1(n14478), .A2(n9789), .ZN(n9795) );
  INV_X1 U11640 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U11641 ( .A1(n9906), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U11642 ( .A1(n9905), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9790) );
  OAI211_X1 U11643 ( .C1(n10117), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9793)
         );
  INV_X1 U11644 ( .A(n9793), .ZN(n9794) );
  NAND2_X1 U11645 ( .A1(n9795), .A2(n9794), .ZN(n14395) );
  XNOR2_X1 U11646 ( .A(n14658), .B(n14388), .ZN(n14467) );
  NAND2_X1 U11647 ( .A1(n14439), .A2(n14438), .ZN(n14437) );
  MUX2_X1 U11648 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n7434), .Z(n10104) );
  XNOR2_X1 U11649 ( .A(n10104), .B(n15633), .ZN(n10105) );
  NAND2_X1 U11650 ( .A1(n14768), .A2(n10135), .ZN(n9801) );
  INV_X1 U11651 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14769) );
  OR2_X1 U11652 ( .A1(n10137), .A2(n14769), .ZN(n9800) );
  OR2_X1 U11653 ( .A1(n9920), .A2(n9802), .ZN(n9808) );
  INV_X1 U11654 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U11655 ( .A1(n9906), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U11656 ( .A1(n9905), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9803) );
  OAI211_X1 U11657 ( .C1(n10117), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9806)
         );
  INV_X1 U11658 ( .A(n9806), .ZN(n9807) );
  NAND2_X1 U11659 ( .A1(n9808), .A2(n9807), .ZN(n14449) );
  XNOR2_X1 U11660 ( .A(n14649), .B(n14449), .ZN(n10209) );
  NOR4_X1 U11661 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9817) );
  NOR4_X1 U11662 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9812) );
  NOR4_X1 U11663 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9811) );
  NOR4_X1 U11664 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9810) );
  NOR4_X1 U11665 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9809) );
  NAND4_X1 U11666 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(n9813)
         );
  NOR4_X1 U11667 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        n9814), .A4(n9813), .ZN(n9816) );
  NOR4_X1 U11668 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9815) );
  NAND3_X1 U11669 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9833) );
  NAND2_X1 U11670 ( .A1(n9827), .A2(n9826), .ZN(n9822) );
  XNOR2_X1 U11671 ( .A(n13035), .B(P2_B_REG_SCAN_IN), .ZN(n9828) );
  INV_X1 U11672 ( .A(n9852), .ZN(n16035) );
  AND2_X1 U11673 ( .A1(n9833), .A2(n16035), .ZN(n11159) );
  INV_X1 U11674 ( .A(n9835), .ZN(n9843) );
  NAND2_X1 U11675 ( .A1(n9839), .A2(n9836), .ZN(n9837) );
  NAND2_X1 U11676 ( .A1(n13175), .A2(n14508), .ZN(n11161) );
  XNOR2_X1 U11677 ( .A(n9839), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9856) );
  AND2_X1 U11678 ( .A1(n11161), .A2(n10182), .ZN(n10124) );
  AND2_X1 U11679 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n9842) );
  NAND2_X1 U11680 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n9840) );
  AOI22_X1 U11681 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(n9560), .B1(n9840), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U11682 ( .A1(n10124), .A2(n10217), .ZN(n11172) );
  INV_X1 U11683 ( .A(n11172), .ZN(n9845) );
  NOR2_X1 U11684 ( .A1(n11159), .A2(n9845), .ZN(n11193) );
  NAND2_X1 U11685 ( .A1(n14781), .A2(n13105), .ZN(n9846) );
  OAI21_X1 U11686 ( .B1(n9852), .B2(P2_D_REG_1__SCAN_IN), .A(n9846), .ZN(
        n11190) );
  INV_X1 U11687 ( .A(n11190), .ZN(n9853) );
  NAND2_X1 U11688 ( .A1(n9847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9849) );
  INV_X1 U11689 ( .A(n10827), .ZN(n11170) );
  NAND2_X1 U11690 ( .A1(n14781), .A2(n13035), .ZN(n9851) );
  AND3_X1 U11691 ( .A1(n9853), .A2(n16041), .A3(n16040), .ZN(n9854) );
  NAND2_X1 U11692 ( .A1(n11193), .A2(n9854), .ZN(n11749) );
  AND2_X1 U11693 ( .A1(n11148), .A2(n14444), .ZN(n9857) );
  NAND2_X1 U11694 ( .A1(n16458), .A2(n9857), .ZN(n14593) );
  NAND2_X2 U11695 ( .A1(n9858), .A2(n14508), .ZN(n14586) );
  INV_X1 U11696 ( .A(n14586), .ZN(n14522) );
  NAND2_X1 U11697 ( .A1(n16458), .A2(n14522), .ZN(n9859) );
  OR2_X1 U11698 ( .A1(n14411), .A2(n11211), .ZN(n9860) );
  NAND2_X1 U11699 ( .A1(n9861), .A2(n9860), .ZN(n11281) );
  NAND2_X1 U11700 ( .A1(n11281), .A2(n11280), .ZN(n9863) );
  INV_X1 U11701 ( .A(n11279), .ZN(n11539) );
  OR2_X1 U11702 ( .A1(n9929), .A2(n11539), .ZN(n9862) );
  OR2_X1 U11703 ( .A1(n14409), .A2(n11995), .ZN(n9864) );
  NAND2_X1 U11704 ( .A1(n11397), .A2(n9866), .ZN(n9868) );
  NAND2_X1 U11705 ( .A1(n7437), .A2(n11404), .ZN(n9867) );
  AND2_X1 U11706 ( .A1(n11517), .A2(n11841), .ZN(n9870) );
  INV_X1 U11707 ( .A(n14406), .ZN(n11868) );
  NAND2_X1 U11708 ( .A1(n11979), .A2(n11868), .ZN(n9871) );
  INV_X1 U11709 ( .A(n14405), .ZN(n12060) );
  NAND2_X1 U11710 ( .A1(n12014), .A2(n12021), .ZN(n9872) );
  INV_X1 U11711 ( .A(n12102), .ZN(n9874) );
  NAND2_X1 U11712 ( .A1(n12101), .A2(n9874), .ZN(n9876) );
  OR2_X1 U11713 ( .A1(n12259), .A2(n12408), .ZN(n9875) );
  INV_X1 U11714 ( .A(n14402), .ZN(n12316) );
  NOR2_X1 U11715 ( .A1(n12400), .A2(n12316), .ZN(n9877) );
  NAND2_X1 U11716 ( .A1(n12400), .A2(n12316), .ZN(n9878) );
  INV_X1 U11717 ( .A(n14400), .ZN(n12783) );
  OR2_X1 U11718 ( .A1(n16462), .A2(n12783), .ZN(n9879) );
  INV_X1 U11719 ( .A(n14399), .ZN(n12949) );
  NAND2_X1 U11720 ( .A1(n12990), .A2(n12949), .ZN(n9880) );
  NAND2_X1 U11721 ( .A1(n12785), .A2(n9880), .ZN(n9882) );
  OR2_X1 U11722 ( .A1(n12990), .A2(n12949), .ZN(n9881) );
  NAND2_X1 U11723 ( .A1(n9882), .A2(n9881), .ZN(n12878) );
  NOR2_X1 U11724 ( .A1(n14732), .A2(n13064), .ZN(n9883) );
  INV_X1 U11725 ( .A(n14732), .ZN(n12955) );
  INV_X1 U11726 ( .A(n14397), .ZN(n13157) );
  OR2_X1 U11727 ( .A1(n14728), .A2(n13157), .ZN(n9884) );
  INV_X1 U11728 ( .A(n14396), .ZN(n14622) );
  NOR2_X1 U11729 ( .A1(n14719), .A2(n14622), .ZN(n9885) );
  INV_X1 U11730 ( .A(n14719), .ZN(n13163) );
  INV_X1 U11731 ( .A(n14582), .ZN(n14624) );
  NAND2_X1 U11732 ( .A1(n14709), .A2(n14624), .ZN(n9886) );
  NAND2_X1 U11733 ( .A1(n14599), .A2(n9886), .ZN(n9888) );
  OR2_X1 U11734 ( .A1(n14709), .A2(n14624), .ZN(n9887) );
  NAND2_X1 U11735 ( .A1(n9888), .A2(n9887), .ZN(n14579) );
  INV_X1 U11736 ( .A(n14605), .ZN(n14568) );
  OR2_X1 U11737 ( .A1(n14704), .A2(n14568), .ZN(n9889) );
  INV_X1 U11738 ( .A(n14584), .ZN(n14320) );
  NAND2_X1 U11739 ( .A1(n14700), .A2(n14320), .ZN(n9891) );
  OR2_X1 U11740 ( .A1(n14700), .A2(n14320), .ZN(n9890) );
  NAND2_X1 U11741 ( .A1(n9891), .A2(n9890), .ZN(n14566) );
  OR2_X1 U11742 ( .A1(n14690), .A2(n14569), .ZN(n10188) );
  NAND2_X1 U11743 ( .A1(n14550), .A2(n10188), .ZN(n9892) );
  NAND2_X1 U11744 ( .A1(n14690), .A2(n14569), .ZN(n10187) );
  NAND2_X1 U11745 ( .A1(n9892), .A2(n10187), .ZN(n14536) );
  AND2_X1 U11746 ( .A1(n14686), .A2(n14321), .ZN(n9894) );
  OR2_X1 U11747 ( .A1(n14686), .A2(n14321), .ZN(n9893) );
  INV_X1 U11748 ( .A(n14537), .ZN(n14363) );
  NOR2_X1 U11749 ( .A1(n14530), .A2(n14363), .ZN(n9895) );
  INV_X1 U11750 ( .A(n14530), .ZN(n14679) );
  NAND2_X1 U11751 ( .A1(n14503), .A2(n14502), .ZN(n9897) );
  INV_X1 U11752 ( .A(n14523), .ZN(n14288) );
  NAND2_X1 U11753 ( .A1(n14675), .A2(n14288), .ZN(n9896) );
  XNOR2_X1 U11754 ( .A(n14671), .B(n14474), .ZN(n14487) );
  INV_X1 U11755 ( .A(n14474), .ZN(n9898) );
  NAND2_X1 U11756 ( .A1(n14671), .A2(n9898), .ZN(n9899) );
  INV_X1 U11757 ( .A(n14395), .ZN(n14459) );
  XNOR2_X1 U11758 ( .A(n14664), .B(n14459), .ZN(n14481) );
  INV_X1 U11759 ( .A(n14481), .ZN(n14472) );
  INV_X1 U11760 ( .A(n14467), .ZN(n14455) );
  INV_X1 U11761 ( .A(n14438), .ZN(n14447) );
  NAND2_X1 U11762 ( .A1(n14448), .A2(n14447), .ZN(n14446) );
  NAND2_X1 U11763 ( .A1(n14446), .A2(n9900), .ZN(n9902) );
  INV_X1 U11764 ( .A(n13175), .ZN(n10190) );
  NAND2_X1 U11765 ( .A1(n10190), .A2(n10182), .ZN(n9903) );
  NAND2_X1 U11766 ( .A1(n10217), .A2(n14444), .ZN(n10125) );
  INV_X1 U11767 ( .A(n11076), .ZN(n11071) );
  NAND2_X1 U11768 ( .A1(n14457), .A2(n14600), .ZN(n9914) );
  INV_X1 U11769 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U11770 ( .A1(n9905), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U11771 ( .A1(n9906), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U11772 ( .C1(n10117), .C2(n9909), .A(n9908), .B(n9907), .ZN(n14394) );
  INV_X1 U11773 ( .A(P2_B_REG_SCAN_IN), .ZN(n9911) );
  OR2_X1 U11774 ( .A1(n14778), .A2(n9911), .ZN(n9912) );
  AND2_X1 U11775 ( .A1(n14583), .A2(n9912), .ZN(n14424) );
  INV_X2 U11776 ( .A(n16458), .ZN(n14598) );
  INV_X1 U11777 ( .A(n14728), .ZN(n13082) );
  INV_X1 U11778 ( .A(n16462), .ZN(n12697) );
  NAND2_X1 U11779 ( .A1(n11211), .A2(n16298), .ZN(n11278) );
  INV_X1 U11780 ( .A(n12021), .ZN(n13167) );
  INV_X1 U11781 ( .A(n12050), .ZN(n16370) );
  NAND2_X1 U11782 ( .A1(n12020), .A2(n16370), .ZN(n12108) );
  INV_X1 U11783 ( .A(n12487), .ZN(n12324) );
  NAND2_X1 U11784 ( .A1(n13082), .A2(n13077), .ZN(n13096) );
  INV_X1 U11785 ( .A(n14675), .ZN(n14514) );
  OR2_X2 U11786 ( .A1(n14499), .A2(n14671), .ZN(n14491) );
  INV_X1 U11787 ( .A(n14658), .ZN(n14465) );
  INV_X1 U11788 ( .A(n11749), .ZN(n9917) );
  INV_X1 U11789 ( .A(n14649), .ZN(n9923) );
  INV_X1 U11790 ( .A(n10182), .ZN(n12731) );
  NAND2_X1 U11791 ( .A1(n10190), .A2(n12731), .ZN(n10179) );
  INV_X1 U11792 ( .A(n10179), .ZN(n9918) );
  NAND2_X1 U11793 ( .A1(n9918), .A2(n7660), .ZN(n11175) );
  INV_X1 U11794 ( .A(n11175), .ZN(n9919) );
  INV_X1 U11795 ( .A(n9920), .ZN(n9921) );
  INV_X1 U11796 ( .A(n16455), .ZN(n14611) );
  AOI22_X1 U11797 ( .A1(n9921), .A2(n14611), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14598), .ZN(n9922) );
  OAI21_X1 U11798 ( .B1(n9923), .B2(n14631), .A(n9922), .ZN(n9924) );
  AND2_X1 U11799 ( .A1(n11279), .A2(n9959), .ZN(n9928) );
  NAND2_X1 U11800 ( .A1(n9929), .A2(n10148), .ZN(n9932) );
  NAND2_X1 U11801 ( .A1(n11279), .A2(n9956), .ZN(n9931) );
  NAND2_X1 U11802 ( .A1(n9932), .A2(n9931), .ZN(n9950) );
  NAND2_X1 U11803 ( .A1(n9933), .A2(n10148), .ZN(n9935) );
  NAND2_X1 U11804 ( .A1(n9935), .A2(n9934), .ZN(n9946) );
  AOI22_X1 U11805 ( .A1(n9951), .A2(n9950), .B1(n9947), .B2(n9946), .ZN(n9949)
         );
  NAND2_X1 U11806 ( .A1(n9937), .A2(n9930), .ZN(n9942) );
  INV_X1 U11807 ( .A(n9938), .ZN(n9939) );
  NAND2_X1 U11808 ( .A1(n11148), .A2(n9939), .ZN(n9940) );
  NAND2_X1 U11809 ( .A1(n9941), .A2(n9940), .ZN(n9945) );
  OAI211_X1 U11810 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9948)
         );
  NAND2_X1 U11811 ( .A1(n9949), .A2(n9948), .ZN(n9955) );
  INV_X1 U11812 ( .A(n9950), .ZN(n9953) );
  INV_X1 U11813 ( .A(n9951), .ZN(n9952) );
  NAND2_X1 U11814 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  NAND2_X1 U11815 ( .A1(n9955), .A2(n9954), .ZN(n9963) );
  NAND2_X1 U11816 ( .A1(n14409), .A2(n9956), .ZN(n9958) );
  NAND2_X1 U11817 ( .A1(n11249), .A2(n10148), .ZN(n9957) );
  NAND2_X1 U11818 ( .A1(n9958), .A2(n9957), .ZN(n9964) );
  NAND2_X1 U11819 ( .A1(n9963), .A2(n9964), .ZN(n9962) );
  NAND2_X1 U11820 ( .A1(n14409), .A2(n10148), .ZN(n9960) );
  OAI21_X1 U11821 ( .B1(n10153), .B2(n11995), .A(n9960), .ZN(n9961) );
  NAND2_X1 U11822 ( .A1(n9962), .A2(n9961), .ZN(n9968) );
  INV_X1 U11823 ( .A(n9963), .ZN(n9966) );
  INV_X1 U11824 ( .A(n9964), .ZN(n9965) );
  NAND2_X1 U11825 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  NAND2_X1 U11826 ( .A1(n11404), .A2(n9956), .ZN(n9970) );
  NAND2_X1 U11827 ( .A1(n14408), .A2(n10148), .ZN(n9969) );
  NAND2_X1 U11828 ( .A1(n9970), .A2(n9969), .ZN(n9972) );
  AOI22_X1 U11829 ( .A1(n10153), .A2(n11404), .B1(n14408), .B2(n9956), .ZN(
        n9971) );
  NAND2_X1 U11830 ( .A1(n11517), .A2(n10153), .ZN(n9975) );
  NAND2_X1 U11831 ( .A1(n14407), .A2(n9956), .ZN(n9974) );
  NAND2_X1 U11832 ( .A1(n9975), .A2(n9974), .ZN(n9977) );
  AOI22_X1 U11833 ( .A1(n11517), .A2(n9930), .B1(n10153), .B2(n14407), .ZN(
        n9976) );
  NAND2_X1 U11834 ( .A1(n11979), .A2(n10176), .ZN(n9980) );
  NAND2_X1 U11835 ( .A1(n14406), .A2(n10153), .ZN(n9979) );
  NAND2_X1 U11836 ( .A1(n9980), .A2(n9979), .ZN(n9982) );
  AOI22_X1 U11837 ( .A1(n11979), .A2(n10148), .B1(n10176), .B2(n14406), .ZN(
        n9981) );
  NAND2_X1 U11838 ( .A1(n12021), .A2(n10153), .ZN(n9985) );
  NAND2_X1 U11839 ( .A1(n14405), .A2(n10176), .ZN(n9984) );
  NAND2_X1 U11840 ( .A1(n9985), .A2(n9984), .ZN(n9987) );
  AOI22_X1 U11841 ( .A1(n12021), .A2(n10176), .B1(n10153), .B2(n14405), .ZN(
        n9986) );
  NAND2_X1 U11842 ( .A1(n12050), .A2(n10176), .ZN(n9990) );
  NAND2_X1 U11843 ( .A1(n14404), .A2(n10153), .ZN(n9989) );
  NAND2_X1 U11844 ( .A1(n9990), .A2(n9989), .ZN(n9992) );
  AOI22_X1 U11845 ( .A1(n12050), .A2(n10148), .B1(n10176), .B2(n14404), .ZN(
        n9991) );
  NAND2_X1 U11846 ( .A1(n12259), .A2(n10153), .ZN(n9995) );
  NAND2_X1 U11847 ( .A1(n14403), .A2(n10176), .ZN(n9994) );
  NAND2_X1 U11848 ( .A1(n9995), .A2(n9994), .ZN(n9999) );
  NAND2_X1 U11849 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  NAND2_X1 U11850 ( .A1(n12259), .A2(n10176), .ZN(n9996) );
  OAI21_X1 U11851 ( .B1(n12408), .B2(n10176), .A(n9996), .ZN(n9997) );
  NAND2_X1 U11852 ( .A1(n12400), .A2(n10176), .ZN(n10002) );
  NAND2_X1 U11853 ( .A1(n14402), .A2(n10153), .ZN(n10001) );
  NAND2_X1 U11854 ( .A1(n10002), .A2(n10001), .ZN(n10004) );
  AOI22_X1 U11855 ( .A1(n12400), .A2(n10153), .B1(n10176), .B2(n14402), .ZN(
        n10003) );
  NAND2_X1 U11856 ( .A1(n12487), .A2(n10153), .ZN(n10006) );
  NAND2_X1 U11857 ( .A1(n14401), .A2(n10176), .ZN(n10005) );
  NAND2_X1 U11858 ( .A1(n10006), .A2(n10005), .ZN(n10010) );
  NAND2_X1 U11859 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  AOI22_X1 U11860 ( .A1(n12487), .A2(n10176), .B1(n10153), .B2(n14401), .ZN(
        n10007) );
  INV_X1 U11861 ( .A(n10007), .ZN(n10008) );
  NAND2_X1 U11862 ( .A1(n10009), .A2(n10008), .ZN(n10013) );
  NAND2_X1 U11863 ( .A1(n16462), .A2(n10176), .ZN(n10015) );
  NAND2_X1 U11864 ( .A1(n14400), .A2(n10148), .ZN(n10014) );
  NAND2_X1 U11865 ( .A1(n10015), .A2(n10014), .ZN(n10020) );
  NAND2_X1 U11866 ( .A1(n10019), .A2(n10020), .ZN(n10018) );
  NAND2_X1 U11867 ( .A1(n16462), .A2(n10148), .ZN(n10016) );
  OAI21_X1 U11868 ( .B1(n10153), .B2(n12783), .A(n10016), .ZN(n10017) );
  NAND2_X1 U11869 ( .A1(n10018), .A2(n10017), .ZN(n10024) );
  NAND2_X1 U11870 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  NAND2_X1 U11871 ( .A1(n12990), .A2(n10153), .ZN(n10026) );
  NAND2_X1 U11872 ( .A1(n14399), .A2(n10176), .ZN(n10025) );
  NAND2_X1 U11873 ( .A1(n10026), .A2(n10025), .ZN(n10028) );
  AOI22_X1 U11874 ( .A1(n12990), .A2(n10176), .B1(n10153), .B2(n14399), .ZN(
        n10027) );
  NAND2_X1 U11875 ( .A1(n14732), .A2(n10176), .ZN(n10030) );
  NAND2_X1 U11876 ( .A1(n14398), .A2(n10148), .ZN(n10029) );
  NAND2_X1 U11877 ( .A1(n10030), .A2(n10029), .ZN(n10035) );
  NAND2_X1 U11878 ( .A1(n14732), .A2(n10153), .ZN(n10032) );
  NAND2_X1 U11879 ( .A1(n14398), .A2(n10176), .ZN(n10031) );
  NAND2_X1 U11880 ( .A1(n10032), .A2(n10031), .ZN(n10033) );
  NAND2_X1 U11881 ( .A1(n10034), .A2(n10033), .ZN(n10037) );
  NAND2_X1 U11882 ( .A1(n14728), .A2(n10153), .ZN(n10039) );
  NAND2_X1 U11883 ( .A1(n14397), .A2(n10176), .ZN(n10038) );
  NAND2_X1 U11884 ( .A1(n10039), .A2(n10038), .ZN(n10041) );
  AOI22_X1 U11885 ( .A1(n14728), .A2(n10176), .B1(n10153), .B2(n14397), .ZN(
        n10040) );
  NAND2_X1 U11886 ( .A1(n14719), .A2(n10176), .ZN(n10043) );
  NAND2_X1 U11887 ( .A1(n14396), .A2(n10153), .ZN(n10042) );
  NAND2_X1 U11888 ( .A1(n10043), .A2(n10042), .ZN(n10045) );
  AOI22_X1 U11889 ( .A1(n14719), .A2(n10153), .B1(n10176), .B2(n14396), .ZN(
        n10044) );
  NAND2_X1 U11890 ( .A1(n14714), .A2(n10153), .ZN(n10048) );
  NAND2_X1 U11891 ( .A1(n14601), .A2(n10176), .ZN(n10047) );
  NAND2_X1 U11892 ( .A1(n10048), .A2(n10047), .ZN(n10052) );
  NAND2_X1 U11893 ( .A1(n14714), .A2(n10176), .ZN(n10049) );
  OAI21_X1 U11894 ( .B1(n13156), .B2(n10176), .A(n10049), .ZN(n10050) );
  NAND2_X1 U11895 ( .A1(n14709), .A2(n10176), .ZN(n10054) );
  NAND2_X1 U11896 ( .A1(n14582), .A2(n10153), .ZN(n10053) );
  AOI22_X1 U11897 ( .A1(n14709), .A2(n10153), .B1(n10176), .B2(n14582), .ZN(
        n10055) );
  INV_X1 U11898 ( .A(n10055), .ZN(n10056) );
  NAND2_X1 U11899 ( .A1(n14704), .A2(n10153), .ZN(n10058) );
  NAND2_X1 U11900 ( .A1(n14605), .A2(n10176), .ZN(n10057) );
  NAND2_X1 U11901 ( .A1(n10058), .A2(n10057), .ZN(n10064) );
  NAND2_X1 U11902 ( .A1(n10063), .A2(n10064), .ZN(n10062) );
  NAND2_X1 U11903 ( .A1(n14704), .A2(n10176), .ZN(n10060) );
  NAND2_X1 U11904 ( .A1(n14605), .A2(n10153), .ZN(n10059) );
  NAND2_X1 U11905 ( .A1(n10060), .A2(n10059), .ZN(n10061) );
  NAND2_X1 U11906 ( .A1(n10062), .A2(n10061), .ZN(n10068) );
  INV_X1 U11907 ( .A(n10063), .ZN(n10066) );
  INV_X1 U11908 ( .A(n10064), .ZN(n10065) );
  NAND2_X1 U11909 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND2_X1 U11910 ( .A1(n14700), .A2(n10176), .ZN(n10070) );
  NAND2_X1 U11911 ( .A1(n14584), .A2(n10153), .ZN(n10069) );
  NAND2_X1 U11912 ( .A1(n10070), .A2(n10069), .ZN(n10073) );
  AOI22_X1 U11913 ( .A1(n14700), .A2(n10153), .B1(n10176), .B2(n14584), .ZN(
        n10071) );
  AOI21_X1 U11914 ( .B1(n10074), .B2(n10073), .A(n10071), .ZN(n10072) );
  NAND2_X1 U11915 ( .A1(n14690), .A2(n10153), .ZN(n10076) );
  NAND2_X1 U11916 ( .A1(n14538), .A2(n10176), .ZN(n10075) );
  NAND2_X1 U11917 ( .A1(n14690), .A2(n10176), .ZN(n10077) );
  OAI21_X1 U11918 ( .B1(n14569), .B2(n10176), .A(n10077), .ZN(n10078) );
  NAND2_X1 U11919 ( .A1(n14686), .A2(n10176), .ZN(n10080) );
  NAND2_X1 U11920 ( .A1(n14552), .A2(n10153), .ZN(n10079) );
  NAND2_X1 U11921 ( .A1(n10080), .A2(n10079), .ZN(n10082) );
  AOI22_X1 U11922 ( .A1(n14686), .A2(n10153), .B1(n10176), .B2(n14552), .ZN(
        n10081) );
  NAND2_X1 U11923 ( .A1(n14530), .A2(n10148), .ZN(n10085) );
  NAND2_X1 U11924 ( .A1(n14537), .A2(n10176), .ZN(n10084) );
  NAND2_X1 U11925 ( .A1(n10085), .A2(n10084), .ZN(n10090) );
  NAND2_X1 U11926 ( .A1(n10089), .A2(n10090), .ZN(n10088) );
  NAND2_X1 U11927 ( .A1(n14530), .A2(n10176), .ZN(n10086) );
  OAI21_X1 U11928 ( .B1(n14363), .B2(n10176), .A(n10086), .ZN(n10087) );
  INV_X1 U11929 ( .A(n10089), .ZN(n10092) );
  INV_X1 U11930 ( .A(n10090), .ZN(n10091) );
  NAND2_X1 U11931 ( .A1(n14675), .A2(n10176), .ZN(n10094) );
  NAND2_X1 U11932 ( .A1(n14523), .A2(n10153), .ZN(n10093) );
  AOI22_X1 U11933 ( .A1(n14675), .A2(n10153), .B1(n10176), .B2(n14523), .ZN(
        n10095) );
  NAND2_X1 U11934 ( .A1(n14671), .A2(n10153), .ZN(n10097) );
  NAND2_X1 U11935 ( .A1(n14474), .A2(n10176), .ZN(n10096) );
  NAND2_X1 U11936 ( .A1(n10097), .A2(n10096), .ZN(n10102) );
  AND2_X1 U11937 ( .A1(n14395), .A2(n10153), .ZN(n10098) );
  AOI21_X1 U11938 ( .B1(n14664), .B2(n10176), .A(n10098), .ZN(n10172) );
  NAND2_X1 U11939 ( .A1(n14664), .A2(n10148), .ZN(n10100) );
  NAND2_X1 U11940 ( .A1(n14395), .A2(n10176), .ZN(n10099) );
  NAND2_X1 U11941 ( .A1(n10100), .A2(n10099), .ZN(n10171) );
  AOI22_X1 U11942 ( .A1(n14671), .A2(n10176), .B1(n10153), .B2(n14474), .ZN(
        n10101) );
  MUX2_X1 U11943 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7434), .Z(n10107) );
  NAND2_X1 U11944 ( .A1(n10107), .A2(SI_30_), .ZN(n10130) );
  OAI21_X1 U11945 ( .B1(SI_30_), .B2(n10107), .A(n10130), .ZN(n10110) );
  INV_X1 U11946 ( .A(n10110), .ZN(n10108) );
  NAND2_X1 U11947 ( .A1(n10109), .A2(n10108), .ZN(n10131) );
  INV_X1 U11948 ( .A(n10109), .ZN(n10111) );
  NAND2_X1 U11949 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  NAND2_X1 U11950 ( .A1(n10131), .A2(n10112), .ZN(n15618) );
  OR2_X1 U11951 ( .A1(n15618), .A2(n10113), .ZN(n10115) );
  INV_X1 U11952 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13456) );
  OR2_X1 U11953 ( .A1(n10137), .A2(n13456), .ZN(n10114) );
  INV_X1 U11954 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10116) );
  OR2_X1 U11955 ( .A1(n10117), .A2(n10116), .ZN(n10123) );
  INV_X1 U11956 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14427) );
  OR2_X1 U11957 ( .A1(n10118), .A2(n14427), .ZN(n10122) );
  INV_X1 U11958 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10119) );
  OR2_X1 U11959 ( .A1(n10120), .A2(n10119), .ZN(n10121) );
  AND3_X1 U11960 ( .A1(n10123), .A2(n10122), .A3(n10121), .ZN(n14426) );
  INV_X1 U11961 ( .A(n14426), .ZN(n10939) );
  NAND2_X1 U11962 ( .A1(n10939), .A2(n10176), .ZN(n10177) );
  OAI211_X1 U11963 ( .C1(n10190), .C2(n10125), .A(n10177), .B(n10124), .ZN(
        n10126) );
  AND2_X1 U11964 ( .A1(n10126), .A2(n14394), .ZN(n10127) );
  AOI21_X1 U11965 ( .B1(n14645), .B2(n10153), .A(n10127), .ZN(n10158) );
  NAND2_X1 U11966 ( .A1(n14645), .A2(n10176), .ZN(n10129) );
  NAND2_X1 U11967 ( .A1(n14394), .A2(n10148), .ZN(n10128) );
  NAND2_X1 U11968 ( .A1(n10129), .A2(n10128), .ZN(n10157) );
  AND2_X1 U11969 ( .A1(n10158), .A2(n10157), .ZN(n10173) );
  NAND2_X1 U11970 ( .A1(n10131), .A2(n10130), .ZN(n10134) );
  MUX2_X1 U11971 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7434), .Z(n10132) );
  XNOR2_X1 U11972 ( .A(n10132), .B(SI_31_), .ZN(n10133) );
  NAND2_X1 U11973 ( .A1(n10701), .A2(n10135), .ZN(n10139) );
  INV_X1 U11974 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10136) );
  OR2_X1 U11975 ( .A1(n10137), .A2(n10136), .ZN(n10138) );
  XNOR2_X1 U11976 ( .A(n10152), .B(n14426), .ZN(n10186) );
  AND2_X1 U11977 ( .A1(n14457), .A2(n10153), .ZN(n10140) );
  AOI21_X1 U11978 ( .B1(n14655), .B2(n10176), .A(n10140), .ZN(n10161) );
  NAND2_X1 U11979 ( .A1(n14655), .A2(n10148), .ZN(n10142) );
  NAND2_X1 U11980 ( .A1(n14457), .A2(n10176), .ZN(n10141) );
  NAND2_X1 U11981 ( .A1(n10142), .A2(n10141), .ZN(n10160) );
  AND2_X1 U11982 ( .A1(n14449), .A2(n10176), .ZN(n10143) );
  AOI21_X1 U11983 ( .B1(n14649), .B2(n10153), .A(n10143), .ZN(n10156) );
  NAND2_X1 U11984 ( .A1(n14649), .A2(n10176), .ZN(n10145) );
  NAND2_X1 U11985 ( .A1(n14449), .A2(n10148), .ZN(n10144) );
  NAND2_X1 U11986 ( .A1(n10145), .A2(n10144), .ZN(n10155) );
  NAND2_X1 U11987 ( .A1(n10156), .A2(n10155), .ZN(n10159) );
  OAI21_X1 U11988 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10146) );
  AND2_X1 U11989 ( .A1(n14475), .A2(n10176), .ZN(n10147) );
  AOI21_X1 U11990 ( .B1(n14658), .B2(n10153), .A(n10147), .ZN(n10166) );
  NAND2_X1 U11991 ( .A1(n14658), .A2(n10176), .ZN(n10150) );
  NAND2_X1 U11992 ( .A1(n14475), .A2(n10148), .ZN(n10149) );
  NAND2_X1 U11993 ( .A1(n10150), .A2(n10149), .ZN(n10165) );
  AND2_X1 U11994 ( .A1(n10166), .A2(n10165), .ZN(n10151) );
  INV_X1 U11995 ( .A(n10152), .ZN(n10175) );
  MUX2_X1 U11996 ( .A(n10153), .B(n10939), .S(n10175), .Z(n10154) );
  OAI21_X1 U11997 ( .B1(n14426), .B2(n10176), .A(n10154), .ZN(n10169) );
  OAI22_X1 U11998 ( .A1(n10158), .A2(n10157), .B1(n10156), .B2(n10155), .ZN(
        n10168) );
  INV_X1 U11999 ( .A(n10159), .ZN(n10164) );
  INV_X1 U12000 ( .A(n10160), .ZN(n10163) );
  INV_X1 U12001 ( .A(n10161), .ZN(n10162) );
  NOR4_X1 U12002 ( .A1(n10186), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10167) );
  MUX2_X1 U12003 ( .A(n10176), .B(n10939), .S(n10175), .Z(n10178) );
  AOI22_X1 U12004 ( .A1(n11148), .A2(n7660), .B1(n14508), .B2(n10179), .ZN(
        n10180) );
  INV_X1 U12005 ( .A(n10180), .ZN(n10181) );
  NOR2_X1 U12006 ( .A1(n10213), .A2(n10181), .ZN(n10221) );
  MUX2_X1 U12007 ( .A(n10217), .B(n10182), .S(n10190), .Z(n10183) );
  NAND2_X1 U12008 ( .A1(n10183), .A2(n14444), .ZN(n10184) );
  INV_X1 U12009 ( .A(n13024), .ZN(n10216) );
  NAND2_X1 U12010 ( .A1(n10185), .A2(n13024), .ZN(n10220) );
  NAND2_X1 U12011 ( .A1(n10188), .A2(n10187), .ZN(n14553) );
  XOR2_X1 U12012 ( .A(n14402), .B(n12400), .Z(n12345) );
  INV_X1 U12013 ( .A(n10189), .ZN(n11221) );
  NOR2_X1 U12014 ( .A1(n11223), .A2(n11221), .ZN(n16300) );
  NAND4_X1 U12015 ( .A1(n16300), .A2(n10190), .A3(n11280), .A4(n11198), .ZN(
        n10192) );
  XNOR2_X1 U12016 ( .A(n11517), .B(n11841), .ZN(n11473) );
  NOR4_X1 U12017 ( .A1(n10192), .A2(n11473), .A3(n11396), .A4(n10191), .ZN(
        n10195) );
  NAND4_X1 U12018 ( .A1(n11878), .A2(n10195), .A3(n10194), .A4(n10193), .ZN(
        n10196) );
  NOR4_X1 U12019 ( .A1(n12345), .A2(n12320), .A3(n12102), .A4(n10196), .ZN(
        n10198) );
  XNOR2_X1 U12020 ( .A(n12990), .B(n14399), .ZN(n12784) );
  NAND4_X1 U12021 ( .A1(n13073), .A2(n10198), .A3(n12784), .A4(n10197), .ZN(
        n10199) );
  NOR3_X1 U12022 ( .A1(n14636), .A2(n12883), .A3(n10199), .ZN(n10201) );
  NAND4_X1 U12023 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n13086), .ZN(
        n10203) );
  NOR4_X1 U12024 ( .A1(n14545), .A2(n14553), .A3(n14566), .A4(n10203), .ZN(
        n10206) );
  NAND2_X1 U12025 ( .A1(n10205), .A2(n10204), .ZN(n14520) );
  NAND4_X1 U12026 ( .A1(n14487), .A2(n10206), .A3(n14502), .A4(n14520), .ZN(
        n10207) );
  NOR4_X1 U12027 ( .A1(n14438), .A2(n14467), .A3(n14481), .A4(n10207), .ZN(
        n10210) );
  XNOR2_X1 U12028 ( .A(n14645), .B(n14394), .ZN(n10208) );
  NAND4_X1 U12029 ( .A1(n8003), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10211) );
  XOR2_X1 U12030 ( .A(n14508), .B(n10211), .Z(n10212) );
  INV_X1 U12031 ( .A(n11161), .ZN(n11165) );
  INV_X1 U12032 ( .A(n14778), .ZN(n10214) );
  NAND4_X1 U12033 ( .A1(n14600), .A2(n11165), .A3(n10214), .A4(n16041), .ZN(
        n10215) );
  OAI211_X1 U12034 ( .C1(n10217), .C2(n10216), .A(n10215), .B(P2_B_REG_SCAN_IN), .ZN(n10218) );
  OAI211_X1 U12035 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        P2_U3328) );
  NOR2_X1 U12036 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n10225) );
  NOR2_X1 U12037 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n10226) );
  NAND3_X1 U12038 ( .A1(n10226), .A2(n16023), .A3(n16024), .ZN(n10227) );
  NOR2_X2 U12039 ( .A1(n10261), .A2(n10227), .ZN(n10269) );
  NAND2_X1 U12040 ( .A1(n10232), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U12041 ( .A1(n10687), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10238) );
  AND2_X4 U12042 ( .A1(n15616), .A2(n15621), .ZN(n10710) );
  XNOR2_X2 U12043 ( .A(n10245), .B(P1_IR_REG_30__SCAN_IN), .ZN(n10234) );
  INV_X1 U12044 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n15457) );
  NAND2_X1 U12045 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10242) );
  MUX2_X1 U12046 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10242), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n10244) );
  INV_X1 U12047 ( .A(n10293), .ZN(n10243) );
  NAND2_X1 U12048 ( .A1(n11291), .A2(n16330), .ZN(n11296) );
  AOI22_X1 U12049 ( .A1(n10252), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(P1_REG0_REG_0__SCAN_IN), .ZN(n10250) );
  INV_X1 U12050 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U12051 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n10246) );
  OAI21_X1 U12052 ( .B1(n10247), .B2(P1_IR_REG_30__SCAN_IN), .A(n10246), .ZN(
        n10248) );
  NAND2_X1 U12053 ( .A1(n10245), .A2(n10248), .ZN(n10249) );
  OAI21_X1 U12054 ( .B1(n10245), .B2(n10250), .A(n10249), .ZN(n10251) );
  NAND2_X1 U12055 ( .A1(n10251), .A2(n15621), .ZN(n10260) );
  AOI22_X1 U12056 ( .A1(n10252), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n10256) );
  INV_X1 U12057 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U12058 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .ZN(n10253) );
  OAI21_X1 U12059 ( .B1(n11011), .B2(P1_IR_REG_30__SCAN_IN), .A(n10253), .ZN(
        n10254) );
  NAND2_X1 U12060 ( .A1(n10245), .A2(n10254), .ZN(n10255) );
  OAI21_X1 U12061 ( .B1(n10245), .B2(n10256), .A(n10255), .ZN(n10258) );
  NAND2_X1 U12062 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  NAND2_X1 U12063 ( .A1(n10260), .A2(n10259), .ZN(n15061) );
  NAND2_X1 U12064 ( .A1(n10272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10264) );
  INV_X1 U12065 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n16195) );
  INV_X1 U12066 ( .A(SI_0_), .ZN(n10266) );
  OAI21_X1 U12067 ( .B1(n10831), .B2(n10266), .A(n10265), .ZN(n10267) );
  NAND2_X1 U12068 ( .A1(n10268), .A2(n10267), .ZN(n15631) );
  MUX2_X1 U12069 ( .A(n16195), .B(n15631), .S(n10892), .Z(n11303) );
  NAND2_X1 U12070 ( .A1(n10229), .A2(n10269), .ZN(n10777) );
  AND2_X1 U12071 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n10271) );
  NAND2_X1 U12072 ( .A1(n10272), .A2(n10271), .ZN(n10277) );
  INV_X1 U12073 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10273) );
  NAND3_X1 U12074 ( .A1(n16024), .A2(n10273), .A3(P1_IR_REG_22__SCAN_IN), .ZN(
        n10275) );
  XNOR2_X1 U12075 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .ZN(
        n10274) );
  NAND2_X1 U12076 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NAND2_X1 U12077 ( .A1(n10278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U12078 ( .A1(n15629), .A2(n15414), .ZN(n11055) );
  NAND2_X1 U12079 ( .A1(n11055), .A2(n10280), .ZN(n10281) );
  NAND2_X1 U12080 ( .A1(n11033), .A2(n10727), .ZN(n11056) );
  NAND2_X1 U12081 ( .A1(n10709), .A2(n11056), .ZN(n10720) );
  OAI211_X1 U12082 ( .C1(n15061), .C2(n11053), .A(n11303), .B(n10358), .ZN(
        n10285) );
  NAND3_X1 U12083 ( .A1(n15061), .A2(n11053), .A3(n10358), .ZN(n10284) );
  INV_X1 U12084 ( .A(n15061), .ZN(n15452) );
  INV_X1 U12085 ( .A(n11303), .ZN(n15462) );
  NAND3_X1 U12086 ( .A1(n15452), .A2(n15462), .A3(n7436), .ZN(n10283) );
  NAND3_X1 U12087 ( .A1(n10285), .A2(n10284), .A3(n10283), .ZN(n10297) );
  NOR2_X1 U12088 ( .A1(n11296), .A2(n10297), .ZN(n10300) );
  MUX2_X1 U12089 ( .A(n15060), .B(n7438), .S(n10358), .Z(n10299) );
  INV_X1 U12090 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11461) );
  OR2_X1 U12091 ( .A1(n10690), .A2(n11461), .ZN(n10289) );
  INV_X1 U12092 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10894) );
  OR2_X1 U12093 ( .A1(n10303), .A2(n10894), .ZN(n10288) );
  NAND2_X1 U12094 ( .A1(n10710), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10287) );
  INV_X1 U12095 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11459) );
  OR2_X1 U12096 ( .A1(n10691), .A2(n11459), .ZN(n10286) );
  INV_X1 U12097 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10836) );
  OR2_X1 U12098 ( .A1(n10322), .A2(n10836), .ZN(n10296) );
  INV_X1 U12099 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10291) );
  NOR2_X1 U12100 ( .A1(n10293), .A2(n10291), .ZN(n10290) );
  MUX2_X1 U12101 ( .A(n10291), .B(n10290), .S(P1_IR_REG_2__SCAN_IN), .Z(n10292) );
  INV_X1 U12102 ( .A(n10292), .ZN(n10294) );
  NAND2_X1 U12103 ( .A1(n10294), .A2(n10409), .ZN(n15086) );
  OR2_X1 U12104 ( .A1(n10892), .A2(n15086), .ZN(n10295) );
  NAND3_X1 U12105 ( .A1(n10297), .A2(n7438), .A3(n15060), .ZN(n10298) );
  OAI211_X1 U12106 ( .C1(n10300), .C2(n10299), .A(n11297), .B(n10298), .ZN(
        n10313) );
  INV_X1 U12107 ( .A(n15449), .ZN(n11302) );
  INV_X1 U12108 ( .A(n11372), .ZN(n11462) );
  AOI21_X1 U12109 ( .B1(n11302), .B2(n10358), .A(n11462), .ZN(n10302) );
  AOI21_X1 U12110 ( .B1(n15449), .B2(n7436), .A(n11372), .ZN(n10301) );
  NAND2_X1 U12111 ( .A1(n10710), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U12112 ( .A1(n10331), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10306) );
  OR2_X1 U12113 ( .A1(n10690), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10305) );
  INV_X1 U12114 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10895) );
  OR2_X1 U12115 ( .A1(n10303), .A2(n10895), .ZN(n10304) );
  NAND2_X1 U12116 ( .A1(n10409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10308) );
  INV_X4 U12117 ( .A(n10309), .ZN(n10702) );
  NAND2_X1 U12118 ( .A1(n10842), .A2(n10702), .ZN(n10311) );
  INV_X1 U12119 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10853) );
  OR2_X1 U12120 ( .A1(n10322), .A2(n10853), .ZN(n10310) );
  XNOR2_X1 U12121 ( .A(n15058), .B(n10314), .ZN(n11289) );
  OAI21_X1 U12122 ( .B1(n15058), .B2(n10358), .A(n10314), .ZN(n10317) );
  NAND2_X1 U12123 ( .A1(n15058), .A2(n10358), .ZN(n10315) );
  NAND2_X1 U12124 ( .A1(n10315), .A2(n11436), .ZN(n10316) );
  NAND2_X1 U12125 ( .A1(n10317), .A2(n10316), .ZN(n10326) );
  NAND2_X1 U12126 ( .A1(n10710), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12127 ( .A1(n7431), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12128 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10332) );
  OAI21_X1 U12129 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n10332), .ZN(n11711) );
  OR2_X1 U12130 ( .A1(n10690), .A2(n11711), .ZN(n10319) );
  INV_X1 U12131 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11529) );
  OR2_X1 U12132 ( .A1(n10691), .A2(n11529), .ZN(n10318) );
  INV_X2 U12134 ( .A(n7723), .ZN(n10559) );
  NAND2_X1 U12135 ( .A1(n10339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10323) );
  XNOR2_X1 U12136 ( .A(n10323), .B(P1_IR_REG_4__SCAN_IN), .ZN(n15117) );
  AOI22_X1 U12137 ( .A1(n10560), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n10559), 
        .B2(n15117), .ZN(n10324) );
  XNOR2_X1 U12138 ( .A(n15057), .B(n11715), .ZN(n11544) );
  OAI21_X1 U12139 ( .B1(n15057), .B2(n7436), .A(n11715), .ZN(n10329) );
  NAND2_X1 U12140 ( .A1(n15057), .A2(n7436), .ZN(n10327) );
  NAND2_X1 U12141 ( .A1(n10327), .A2(n11696), .ZN(n10328) );
  NAND2_X1 U12142 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  NAND2_X1 U12143 ( .A1(n10710), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10338) );
  NAND2_X1 U12144 ( .A1(n7433), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10337) );
  AND2_X1 U12145 ( .A1(n10332), .A2(n11736), .ZN(n10333) );
  NOR2_X1 U12146 ( .A1(n10332), .A2(n11736), .ZN(n10350) );
  OR2_X1 U12147 ( .A1(n10333), .A2(n10350), .ZN(n11737) );
  OR2_X1 U12148 ( .A1(n10690), .A2(n11737), .ZN(n10336) );
  INV_X1 U12149 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10334) );
  OR2_X1 U12150 ( .A1(n10714), .A2(n10334), .ZN(n10335) );
  NAND4_X1 U12151 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n15056) );
  NAND2_X1 U12152 ( .A1(n10854), .A2(n10702), .ZN(n10344) );
  INV_X1 U12153 ( .A(n10339), .ZN(n10341) );
  INV_X1 U12154 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U12155 ( .A1(n10341), .A2(n10340), .ZN(n10346) );
  NAND2_X1 U12156 ( .A1(n10346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10342) );
  XNOR2_X1 U12157 ( .A(n10342), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U12158 ( .A1(n10560), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10559), 
        .B2(n10927), .ZN(n10343) );
  NAND2_X1 U12159 ( .A1(n10344), .A2(n10343), .ZN(n11890) );
  MUX2_X1 U12160 ( .A(n15056), .B(n11890), .S(n10358), .Z(n10356) );
  MUX2_X1 U12161 ( .A(n15056), .B(n11890), .S(n7436), .Z(n10345) );
  NAND2_X1 U12162 ( .A1(n10878), .A2(n10702), .ZN(n10349) );
  NAND2_X1 U12163 ( .A1(n10370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10347) );
  XNOR2_X1 U12164 ( .A(n10347), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U12165 ( .A1(n10560), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10559), 
        .B2(n10954), .ZN(n10348) );
  NAND2_X1 U12166 ( .A1(n7431), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U12167 ( .A1(n10710), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U12168 ( .A1(n10350), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10363) );
  OR2_X1 U12169 ( .A1(n10350), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12170 ( .A1(n10363), .A2(n10351), .ZN(n11940) );
  OR2_X1 U12171 ( .A1(n10690), .A2(n11940), .ZN(n10353) );
  INV_X1 U12172 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11939) );
  OR2_X1 U12173 ( .A1(n10691), .A2(n11939), .ZN(n10352) );
  NAND4_X1 U12174 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n15055) );
  XNOR2_X1 U12175 ( .A(n12029), .B(n15055), .ZN(n11888) );
  AND2_X1 U12176 ( .A1(n15055), .A2(n7436), .ZN(n10360) );
  OAI21_X1 U12177 ( .B1(n7436), .B2(n15055), .A(n12029), .ZN(n10359) );
  OAI21_X1 U12178 ( .B1(n10360), .B2(n12029), .A(n10359), .ZN(n10361) );
  NAND2_X1 U12179 ( .A1(n10710), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10369) );
  NAND2_X1 U12180 ( .A1(n7433), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U12181 ( .A1(n10363), .A2(n10362), .ZN(n10364) );
  NAND2_X1 U12182 ( .A1(n10380), .A2(n10364), .ZN(n12042) );
  OR2_X1 U12183 ( .A1(n10690), .A2(n12042), .ZN(n10367) );
  INV_X1 U12184 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10365) );
  OR2_X1 U12185 ( .A1(n10714), .A2(n10365), .ZN(n10366) );
  NAND4_X1 U12186 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n15054) );
  NAND2_X1 U12187 ( .A1(n10884), .A2(n10702), .ZN(n10374) );
  INV_X1 U12188 ( .A(n10370), .ZN(n10371) );
  INV_X1 U12189 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n15995) );
  NAND2_X1 U12190 ( .A1(n10371), .A2(n15995), .ZN(n10386) );
  NAND2_X1 U12191 ( .A1(n10386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10372) );
  XNOR2_X1 U12192 ( .A(n10372), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U12193 ( .A1(n10560), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10559), 
        .B2(n10955), .ZN(n10373) );
  NAND2_X1 U12194 ( .A1(n10374), .A2(n10373), .ZN(n16350) );
  MUX2_X1 U12195 ( .A(n15054), .B(n16350), .S(n10358), .Z(n10377) );
  MUX2_X1 U12196 ( .A(n15054), .B(n16350), .S(n7436), .Z(n10375) );
  NAND2_X1 U12197 ( .A1(n7431), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U12198 ( .A1(n10710), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U12199 ( .A1(n10380), .A2(n10379), .ZN(n10381) );
  NAND2_X1 U12200 ( .A1(n10399), .A2(n10381), .ZN(n12193) );
  OR2_X1 U12201 ( .A1(n10690), .A2(n12193), .ZN(n10383) );
  INV_X1 U12202 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n12095) );
  OR2_X1 U12203 ( .A1(n10691), .A2(n12095), .ZN(n10382) );
  NAND4_X1 U12204 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n15053) );
  NAND2_X1 U12205 ( .A1(n10888), .A2(n10702), .ZN(n10389) );
  OAI21_X1 U12206 ( .B1(n10386), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10387) );
  XNOR2_X1 U12207 ( .A(n10387), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U12208 ( .A1(n10560), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10559), 
        .B2(n10996), .ZN(n10388) );
  NAND2_X1 U12209 ( .A1(n10389), .A2(n10388), .ZN(n16359) );
  MUX2_X1 U12210 ( .A(n15053), .B(n16359), .S(n7436), .Z(n10393) );
  NAND2_X1 U12211 ( .A1(n10392), .A2(n10393), .ZN(n10391) );
  MUX2_X1 U12212 ( .A(n15053), .B(n16359), .S(n10650), .Z(n10390) );
  NAND2_X1 U12213 ( .A1(n10391), .A2(n10390), .ZN(n10397) );
  INV_X1 U12214 ( .A(n10393), .ZN(n10394) );
  NAND2_X1 U12215 ( .A1(n10395), .A2(n10394), .ZN(n10396) );
  NAND2_X1 U12216 ( .A1(n10710), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10406) );
  NAND2_X1 U12217 ( .A1(n7433), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10405) );
  INV_X1 U12218 ( .A(n10417), .ZN(n10401) );
  NAND2_X1 U12219 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  NAND2_X1 U12220 ( .A1(n10401), .A2(n10400), .ZN(n12507) );
  OR2_X1 U12221 ( .A1(n10690), .A2(n12507), .ZN(n10404) );
  INV_X1 U12222 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10402) );
  OR2_X1 U12223 ( .A1(n10714), .A2(n10402), .ZN(n10403) );
  NAND4_X1 U12224 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n15052) );
  NAND2_X1 U12225 ( .A1(n10941), .A2(n10702), .ZN(n10413) );
  NAND2_X1 U12226 ( .A1(n10407), .A2(n10408), .ZN(n10410) );
  OR2_X1 U12227 ( .A1(n10410), .A2(n10409), .ZN(n10424) );
  NAND2_X1 U12228 ( .A1(n10424), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10411) );
  XNOR2_X1 U12229 ( .A(n10411), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U12230 ( .A1(n10560), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10559), 
        .B2(n11335), .ZN(n10412) );
  MUX2_X1 U12231 ( .A(n15052), .B(n12496), .S(n7436), .Z(n10414) );
  NAND2_X1 U12232 ( .A1(n10710), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U12233 ( .A1(n7433), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10422) );
  NAND2_X1 U12234 ( .A1(n10417), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10431) );
  OR2_X1 U12235 ( .A1(n10417), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U12236 ( .A1(n10431), .A2(n10418), .ZN(n12563) );
  OR2_X1 U12237 ( .A1(n10690), .A2(n12563), .ZN(n10421) );
  INV_X1 U12238 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10419) );
  OR2_X1 U12239 ( .A1(n10714), .A2(n10419), .ZN(n10420) );
  NAND4_X1 U12240 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n15051) );
  NAND2_X1 U12241 ( .A1(n10946), .A2(n10702), .ZN(n10427) );
  OAI21_X1 U12242 ( .B1(n10424), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10425) );
  XNOR2_X1 U12243 ( .A(n10425), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U12244 ( .A1(n10560), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10559), 
        .B2(n11347), .ZN(n10426) );
  MUX2_X1 U12245 ( .A(n15051), .B(n12567), .S(n7436), .Z(n10429) );
  MUX2_X1 U12246 ( .A(n15051), .B(n12567), .S(n10650), .Z(n10428) );
  NAND2_X1 U12247 ( .A1(n7431), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U12248 ( .A1(n10710), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U12249 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  NAND2_X1 U12250 ( .A1(n10446), .A2(n10432), .ZN(n12708) );
  OR2_X1 U12251 ( .A1(n10690), .A2(n12708), .ZN(n10435) );
  INV_X1 U12252 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10433) );
  OR2_X1 U12253 ( .A1(n10691), .A2(n10433), .ZN(n10434) );
  NAND4_X1 U12254 ( .A1(n10437), .A2(n10436), .A3(n10435), .A4(n10434), .ZN(
        n15050) );
  NAND2_X1 U12255 ( .A1(n10986), .A2(n10702), .ZN(n10441) );
  NAND2_X1 U12256 ( .A1(n10453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10439) );
  XNOR2_X1 U12257 ( .A(n10439), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U12258 ( .A1(n10560), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10559), 
        .B2(n11604), .ZN(n10440) );
  MUX2_X1 U12259 ( .A(n15050), .B(n12712), .S(n10650), .Z(n10444) );
  MUX2_X1 U12260 ( .A(n15050), .B(n12712), .S(n7436), .Z(n10442) );
  NAND2_X1 U12261 ( .A1(n7431), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12262 ( .A1(n10710), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10451) );
  INV_X1 U12263 ( .A(n10461), .ZN(n10448) );
  NAND2_X1 U12264 ( .A1(n10446), .A2(n10445), .ZN(n10447) );
  NAND2_X1 U12265 ( .A1(n10448), .A2(n10447), .ZN(n12855) );
  OR2_X1 U12266 ( .A1(n10690), .A2(n12855), .ZN(n10450) );
  INV_X1 U12267 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12614) );
  OR2_X1 U12268 ( .A1(n10691), .A2(n12614), .ZN(n10449) );
  NAND4_X1 U12269 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n15049) );
  NAND2_X1 U12270 ( .A1(n11085), .A2(n10702), .ZN(n10455) );
  NOR2_X1 U12271 ( .A1(n10453), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10499) );
  OR2_X1 U12272 ( .A1(n10499), .A2(n10291), .ZN(n10467) );
  XNOR2_X1 U12273 ( .A(n10467), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U12274 ( .A1(n10560), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10559), 
        .B2(n11815), .ZN(n10454) );
  MUX2_X1 U12275 ( .A(n15049), .B(n12851), .S(n7436), .Z(n10458) );
  MUX2_X1 U12276 ( .A(n15049), .B(n12851), .S(n10650), .Z(n10456) );
  NAND2_X1 U12277 ( .A1(n10457), .A2(n10456), .ZN(n10460) );
  NAND2_X1 U12278 ( .A1(n7431), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U12279 ( .A1(n10710), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U12280 ( .A1(n7433), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U12281 ( .A1(n10461), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10476) );
  OR2_X1 U12282 ( .A1(n10461), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12283 ( .A1(n10476), .A2(n10462), .ZN(n12965) );
  OR2_X1 U12284 ( .A1(n10690), .A2(n12965), .ZN(n10463) );
  NAND4_X1 U12285 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n15048) );
  NAND2_X1 U12286 ( .A1(n11182), .A2(n10702), .ZN(n10472) );
  AOI21_X1 U12287 ( .B1(n10467), .B2(n16006), .A(n10291), .ZN(n10468) );
  NAND2_X1 U12288 ( .A1(n10468), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n10470) );
  INV_X1 U12289 ( .A(n10468), .ZN(n10469) );
  NAND2_X1 U12290 ( .A1(n10469), .A2(n16007), .ZN(n10483) );
  AOI22_X1 U12291 ( .A1(n10560), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n10559), 
        .B2(n12393), .ZN(n10471) );
  MUX2_X1 U12292 ( .A(n15048), .B(n12967), .S(n10650), .Z(n10474) );
  MUX2_X1 U12293 ( .A(n15048), .B(n12967), .S(n7436), .Z(n10473) );
  INV_X1 U12294 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U12295 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U12296 ( .A1(n10490), .A2(n10477), .ZN(n12764) );
  OR2_X1 U12297 ( .A1(n12764), .A2(n10690), .ZN(n10482) );
  NAND2_X1 U12298 ( .A1(n7431), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10481) );
  INV_X1 U12299 ( .A(n10710), .ZN(n10689) );
  INV_X1 U12300 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10478) );
  OR2_X1 U12301 ( .A1(n10689), .A2(n10478), .ZN(n10480) );
  INV_X1 U12302 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12620) );
  OR2_X1 U12303 ( .A1(n10691), .A2(n12620), .ZN(n10479) );
  NAND4_X1 U12304 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n15047) );
  NAND2_X1 U12305 ( .A1(n11378), .A2(n10702), .ZN(n10486) );
  NAND2_X1 U12306 ( .A1(n10483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10484) );
  XNOR2_X1 U12307 ( .A(n10484), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U12308 ( .A1(n10560), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n10559), 
        .B2(n12394), .ZN(n10485) );
  MUX2_X1 U12309 ( .A(n15047), .B(n15579), .S(n7436), .Z(n10488) );
  MUX2_X1 U12310 ( .A(n15047), .B(n15579), .S(n10650), .Z(n10487) );
  INV_X1 U12311 ( .A(n10488), .ZN(n10489) );
  AND2_X1 U12312 ( .A1(n10490), .A2(n15034), .ZN(n10491) );
  OR2_X1 U12313 ( .A1(n10491), .A2(n10507), .ZN(n15035) );
  INV_X1 U12314 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10492) );
  OR2_X1 U12315 ( .A1(n10689), .A2(n10492), .ZN(n10495) );
  INV_X1 U12316 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10493) );
  OR2_X1 U12317 ( .A1(n10714), .A2(n10493), .ZN(n10494) );
  AND2_X1 U12318 ( .A1(n10495), .A2(n10494), .ZN(n10497) );
  INV_X1 U12319 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12983) );
  OR2_X1 U12320 ( .A1(n10691), .A2(n12983), .ZN(n10496) );
  OAI211_X1 U12321 ( .C1(n15035), .C2(n10690), .A(n10497), .B(n10496), .ZN(
        n15175) );
  NAND2_X1 U12322 ( .A1(n11561), .A2(n10702), .ZN(n10502) );
  INV_X1 U12323 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n16013) );
  AND3_X1 U12324 ( .A1(n16006), .A2(n16007), .A3(n16013), .ZN(n10498) );
  AND2_X1 U12325 ( .A1(n10499), .A2(n10498), .ZN(n10511) );
  OR2_X1 U12326 ( .A1(n10511), .A2(n10291), .ZN(n10500) );
  XNOR2_X1 U12327 ( .A(n10500), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U12328 ( .A1(n10560), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10559), 
        .B2(n12805), .ZN(n10501) );
  MUX2_X1 U12329 ( .A(n15175), .B(n15571), .S(n10650), .Z(n10505) );
  MUX2_X1 U12330 ( .A(n15571), .B(n15175), .S(n10650), .Z(n10503) );
  INV_X1 U12331 ( .A(n10505), .ZN(n10506) );
  NOR2_X1 U12332 ( .A1(n10507), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10508) );
  OR2_X1 U12333 ( .A1(n10521), .A2(n10508), .ZN(n15429) );
  AOI22_X1 U12334 ( .A1(n7431), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n10710), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n10510) );
  OR2_X1 U12335 ( .A1(n10691), .A2(n12801), .ZN(n10509) );
  OAI211_X1 U12336 ( .C1(n15429), .C2(n10690), .A(n10510), .B(n10509), .ZN(
        n15177) );
  NAND2_X1 U12337 ( .A1(n11718), .A2(n10702), .ZN(n10517) );
  INV_X1 U12338 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n16012) );
  AND2_X1 U12339 ( .A1(n10511), .A2(n16012), .ZN(n10514) );
  NOR2_X1 U12340 ( .A1(n10514), .A2(n10291), .ZN(n10512) );
  MUX2_X1 U12341 ( .A(n10291), .B(n10512), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n10513) );
  INV_X1 U12342 ( .A(n10513), .ZN(n10515) );
  INV_X1 U12343 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U12344 ( .A1(n10514), .A2(n16017), .ZN(n10542) );
  AOI22_X1 U12345 ( .A1(n10560), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12808), 
        .B2(n10559), .ZN(n10516) );
  MUX2_X1 U12346 ( .A(n15177), .B(n15562), .S(n7436), .Z(n10520) );
  MUX2_X1 U12347 ( .A(n15177), .B(n15562), .S(n10650), .Z(n10518) );
  OR2_X1 U12348 ( .A1(n10521), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U12349 ( .A1(n10534), .A2(n10522), .ZN(n14975) );
  AOI22_X1 U12350 ( .A1(n10710), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n7433), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n10524) );
  INV_X1 U12351 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15131) );
  OR2_X1 U12352 ( .A1(n10714), .A2(n15131), .ZN(n10523) );
  OAI211_X1 U12353 ( .C1(n14975), .C2(n10690), .A(n10524), .B(n10523), .ZN(
        n15385) );
  NAND2_X1 U12354 ( .A1(n11822), .A2(n10702), .ZN(n10528) );
  NAND2_X1 U12355 ( .A1(n10542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10525) );
  INV_X1 U12356 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n16018) );
  XNOR2_X1 U12357 ( .A(n10525), .B(n16018), .ZN(n15130) );
  INV_X1 U12358 ( .A(n15130), .ZN(n10526) );
  AOI22_X1 U12359 ( .A1(n10560), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n10526), 
        .B2(n10559), .ZN(n10527) );
  MUX2_X1 U12360 ( .A(n15385), .B(n15555), .S(n10650), .Z(n10531) );
  MUX2_X1 U12361 ( .A(n15555), .B(n15385), .S(n10650), .Z(n10529) );
  NAND2_X1 U12362 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND2_X1 U12363 ( .A1(n10553), .A2(n10535), .ZN(n15394) );
  OR2_X1 U12364 ( .A1(n15394), .A2(n10690), .ZN(n10541) );
  INV_X1 U12365 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U12366 ( .A1(n10710), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n10537) );
  INV_X1 U12367 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15393) );
  OR2_X1 U12368 ( .A1(n10691), .A2(n15393), .ZN(n10536) );
  OAI211_X1 U12369 ( .C1(n10538), .C2(n10714), .A(n10537), .B(n10536), .ZN(
        n10539) );
  INV_X1 U12370 ( .A(n10539), .ZN(n10540) );
  NAND2_X1 U12371 ( .A1(n10541), .A2(n10540), .ZN(n15370) );
  NAND2_X1 U12372 ( .A1(n12164), .A2(n10702), .ZN(n10545) );
  OAI21_X1 U12373 ( .B1(n10542), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10543) );
  XNOR2_X1 U12374 ( .A(n10543), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U12375 ( .A1(n10560), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n15145), 
        .B2(n10559), .ZN(n10544) );
  MUX2_X1 U12376 ( .A(n15370), .B(n15396), .S(n7436), .Z(n10548) );
  MUX2_X1 U12377 ( .A(n15370), .B(n15396), .S(n10650), .Z(n10546) );
  NAND2_X1 U12378 ( .A1(n10547), .A2(n10546), .ZN(n10551) );
  INV_X1 U12379 ( .A(n10548), .ZN(n10549) );
  NAND2_X1 U12380 ( .A1(n7495), .A2(n10549), .ZN(n10550) );
  NAND2_X1 U12381 ( .A1(n10551), .A2(n10550), .ZN(n10564) );
  INV_X1 U12382 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U12383 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  NAND2_X1 U12384 ( .A1(n10567), .A2(n10554), .ZN(n15375) );
  INV_X1 U12385 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U12386 ( .A1(n7433), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n10556) );
  NAND2_X1 U12387 ( .A1(n10710), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n10555) );
  OAI211_X1 U12388 ( .C1(n10714), .C2(n15142), .A(n10556), .B(n10555), .ZN(
        n10557) );
  INV_X1 U12389 ( .A(n10557), .ZN(n10558) );
  OAI21_X1 U12390 ( .B1(n15375), .B2(n10690), .A(n10558), .ZN(n15387) );
  NAND2_X1 U12391 ( .A1(n12381), .A2(n10702), .ZN(n10562) );
  AOI22_X1 U12392 ( .A1(n10560), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15414), 
        .B2(n10559), .ZN(n10561) );
  MUX2_X1 U12393 ( .A(n15387), .B(n15538), .S(n10650), .Z(n10565) );
  MUX2_X1 U12394 ( .A(n15387), .B(n15538), .S(n7436), .Z(n10563) );
  INV_X1 U12395 ( .A(n10565), .ZN(n10566) );
  INV_X1 U12396 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14995) );
  NOR2_X1 U12397 ( .A1(n10580), .A2(n8499), .ZN(n15357) );
  NAND2_X1 U12398 ( .A1(n15357), .A2(n10568), .ZN(n10574) );
  INV_X1 U12399 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U12400 ( .A1(n7433), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U12401 ( .A1(n10710), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n10569) );
  OAI211_X1 U12402 ( .C1(n10714), .C2(n10571), .A(n10570), .B(n10569), .ZN(
        n10572) );
  INV_X1 U12403 ( .A(n10572), .ZN(n10573) );
  NAND2_X1 U12404 ( .A1(n10574), .A2(n10573), .ZN(n15369) );
  NAND2_X1 U12405 ( .A1(n12596), .A2(n10702), .ZN(n10576) );
  OR2_X1 U12406 ( .A1(n10322), .A2(n12598), .ZN(n10575) );
  MUX2_X1 U12407 ( .A(n15369), .B(n15533), .S(n7436), .Z(n10579) );
  MUX2_X1 U12408 ( .A(n15369), .B(n15533), .S(n10650), .Z(n10577) );
  NOR2_X1 U12409 ( .A1(n10580), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n10581) );
  OR2_X1 U12410 ( .A1(n10592), .A2(n10581), .ZN(n14948) );
  INV_X1 U12411 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U12412 ( .A1(n10710), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U12413 ( .A1(n7433), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n10582) );
  OAI211_X1 U12414 ( .C1(n10714), .C2(n10584), .A(n10583), .B(n10582), .ZN(
        n10585) );
  INV_X1 U12415 ( .A(n10585), .ZN(n10586) );
  NAND2_X1 U12416 ( .A1(n12728), .A2(n10702), .ZN(n10588) );
  OR2_X1 U12417 ( .A1(n10322), .A2(n12730), .ZN(n10587) );
  MUX2_X1 U12418 ( .A(n15319), .B(n15528), .S(n7436), .Z(n10589) );
  NOR2_X1 U12419 ( .A1(n10592), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n10593) );
  OR2_X1 U12420 ( .A1(n10605), .A2(n10593), .ZN(n15003) );
  INV_X1 U12421 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U12422 ( .A1(n10710), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U12423 ( .A1(n7433), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n10594) );
  OAI211_X1 U12424 ( .C1(n10714), .C2(n10596), .A(n10595), .B(n10594), .ZN(
        n10597) );
  INV_X1 U12425 ( .A(n10597), .ZN(n10598) );
  MUX2_X1 U12426 ( .A(n15333), .B(n15522), .S(n7436), .Z(n10602) );
  MUX2_X1 U12427 ( .A(n15333), .B(n15522), .S(n10650), .Z(n10600) );
  NAND2_X1 U12428 ( .A1(n10601), .A2(n10600), .ZN(n10604) );
  INV_X1 U12429 ( .A(n10602), .ZN(n10603) );
  OR2_X1 U12430 ( .A1(n10605), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U12431 ( .A1(n10605), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U12432 ( .A1(n10606), .A2(n10616), .ZN(n15309) );
  INV_X1 U12433 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U12434 ( .A1(n7433), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U12435 ( .A1(n10710), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n10607) );
  OAI211_X1 U12436 ( .C1(n10714), .C2(n10609), .A(n10608), .B(n10607), .ZN(
        n10610) );
  INV_X1 U12437 ( .A(n10610), .ZN(n10611) );
  OR2_X1 U12438 ( .A1(n10322), .A2(n13031), .ZN(n10612) );
  MUX2_X1 U12439 ( .A(n15320), .B(n15517), .S(n7436), .Z(n10613) );
  INV_X1 U12440 ( .A(n10614), .ZN(n10615) );
  NAND2_X1 U12441 ( .A1(n7431), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U12442 ( .A1(n10710), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n10620) );
  OAI21_X1 U12443 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n10617), .A(n10629), 
        .ZN(n15296) );
  OR2_X1 U12444 ( .A1(n10690), .A2(n15296), .ZN(n10619) );
  INV_X1 U12445 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15297) );
  OR2_X1 U12446 ( .A1(n10691), .A2(n15297), .ZN(n10618) );
  NAND4_X1 U12447 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n15183) );
  NAND2_X1 U12448 ( .A1(n13032), .A2(n10702), .ZN(n10623) );
  INV_X1 U12449 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13034) );
  OR2_X1 U12450 ( .A1(n10322), .A2(n13034), .ZN(n10622) );
  MUX2_X1 U12451 ( .A(n15183), .B(n15509), .S(n7436), .Z(n10626) );
  MUX2_X1 U12452 ( .A(n15183), .B(n15509), .S(n10650), .Z(n10624) );
  NAND2_X1 U12453 ( .A1(n10625), .A2(n10624), .ZN(n10628) );
  NAND2_X1 U12454 ( .A1(n10628), .A2(n10627), .ZN(n10639) );
  NAND2_X1 U12455 ( .A1(n10710), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U12456 ( .A1(n7433), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n10634) );
  NAND2_X1 U12457 ( .A1(n10630), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n10642) );
  OAI21_X1 U12458 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n10630), .A(n10642), 
        .ZN(n15279) );
  OR2_X1 U12459 ( .A1(n10690), .A2(n15279), .ZN(n10633) );
  INV_X1 U12460 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10631) );
  OR2_X1 U12461 ( .A1(n10714), .A2(n10631), .ZN(n10632) );
  NAND4_X1 U12462 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n15290) );
  NAND2_X1 U12463 ( .A1(n13102), .A2(n10702), .ZN(n10637) );
  OR2_X1 U12464 ( .A1(n10322), .A2(n7719), .ZN(n10636) );
  MUX2_X1 U12465 ( .A(n15290), .B(n15501), .S(n10650), .Z(n10640) );
  MUX2_X1 U12466 ( .A(n15290), .B(n15501), .S(n7436), .Z(n10638) );
  INV_X1 U12467 ( .A(n10640), .ZN(n10641) );
  NAND2_X1 U12468 ( .A1(n10710), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U12469 ( .A1(n7431), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U12470 ( .A1(n10643), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n10659) );
  OAI21_X1 U12471 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n10643), .A(n10659), 
        .ZN(n15262) );
  OR2_X1 U12472 ( .A1(n10690), .A2(n15262), .ZN(n10645) );
  INV_X1 U12473 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15263) );
  OR2_X1 U12474 ( .A1(n10691), .A2(n15263), .ZN(n10644) );
  NAND4_X1 U12475 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n15046) );
  NAND2_X1 U12476 ( .A1(n14779), .A2(n10702), .ZN(n10649) );
  OR2_X1 U12477 ( .A1(n10322), .A2(n7735), .ZN(n10648) );
  MUX2_X1 U12478 ( .A(n15046), .B(n15495), .S(n7436), .Z(n10654) );
  MUX2_X1 U12479 ( .A(n15046), .B(n15495), .S(n10650), .Z(n10651) );
  NAND2_X1 U12480 ( .A1(n10652), .A2(n10651), .ZN(n10658) );
  INV_X1 U12481 ( .A(n10653), .ZN(n10656) );
  INV_X1 U12482 ( .A(n10654), .ZN(n10655) );
  NAND2_X1 U12483 ( .A1(n10656), .A2(n10655), .ZN(n10657) );
  NAND2_X1 U12484 ( .A1(n10658), .A2(n10657), .ZN(n10668) );
  NAND2_X1 U12485 ( .A1(n7431), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n10664) );
  NAND2_X1 U12486 ( .A1(n10710), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n10663) );
  INV_X1 U12487 ( .A(n10659), .ZN(n10660) );
  NAND2_X1 U12488 ( .A1(n10660), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n10671) );
  OAI21_X1 U12489 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n10660), .A(n10671), 
        .ZN(n15250) );
  OR2_X1 U12490 ( .A1(n10690), .A2(n15250), .ZN(n10662) );
  INV_X1 U12491 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n15251) );
  OR2_X1 U12492 ( .A1(n10691), .A2(n15251), .ZN(n10661) );
  NAND2_X1 U12493 ( .A1(n14776), .A2(n10702), .ZN(n10666) );
  OR2_X1 U12494 ( .A1(n10322), .A2(n15624), .ZN(n10665) );
  NAND2_X2 U12495 ( .A1(n10666), .A2(n10665), .ZN(n15489) );
  MUX2_X1 U12496 ( .A(n15217), .B(n15489), .S(n10358), .Z(n10669) );
  MUX2_X1 U12497 ( .A(n15217), .B(n15489), .S(n7436), .Z(n10667) );
  INV_X1 U12498 ( .A(n10669), .ZN(n10670) );
  NAND2_X1 U12499 ( .A1(n7431), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U12500 ( .A1(n10710), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n10675) );
  INV_X1 U12501 ( .A(n10671), .ZN(n10672) );
  NAND2_X1 U12502 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n10672), .ZN(n15206) );
  OAI21_X1 U12503 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n10672), .A(n15206), 
        .ZN(n15228) );
  OR2_X1 U12504 ( .A1(n10690), .A2(n15228), .ZN(n10674) );
  INV_X1 U12505 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15229) );
  OR2_X1 U12506 ( .A1(n10691), .A2(n15229), .ZN(n10673) );
  NAND4_X1 U12507 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n15201) );
  NAND2_X1 U12508 ( .A1(n14772), .A2(n10702), .ZN(n10678) );
  OR2_X1 U12509 ( .A1(n10322), .A2(n7738), .ZN(n10677) );
  MUX2_X1 U12510 ( .A(n15201), .B(n15483), .S(n7436), .Z(n10682) );
  MUX2_X1 U12511 ( .A(n15201), .B(n15483), .S(n10358), .Z(n10679) );
  NAND2_X1 U12512 ( .A1(n10680), .A2(n10679), .ZN(n10686) );
  INV_X1 U12513 ( .A(n10681), .ZN(n10684) );
  INV_X1 U12514 ( .A(n10682), .ZN(n10683) );
  NAND2_X1 U12515 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  NAND2_X1 U12516 ( .A1(n10686), .A2(n10685), .ZN(n10700) );
  NAND2_X1 U12517 ( .A1(n7431), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n10695) );
  INV_X1 U12518 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10688) );
  OR2_X1 U12519 ( .A1(n10689), .A2(n10688), .ZN(n10694) );
  OR2_X1 U12520 ( .A1(n10690), .A2(n15206), .ZN(n10693) );
  INV_X1 U12521 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15207) );
  OR2_X1 U12522 ( .A1(n10691), .A2(n15207), .ZN(n10692) );
  NAND2_X1 U12523 ( .A1(n14768), .A2(n10702), .ZN(n10697) );
  INV_X1 U12524 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15619) );
  OR2_X1 U12525 ( .A1(n10322), .A2(n15619), .ZN(n10696) );
  MUX2_X1 U12526 ( .A(n15216), .B(n15477), .S(n10358), .Z(n10699) );
  MUX2_X1 U12527 ( .A(n15211), .B(n14941), .S(n10358), .Z(n10698) );
  INV_X1 U12528 ( .A(n10771), .ZN(n10726) );
  NAND2_X1 U12529 ( .A1(n10701), .A2(n10702), .ZN(n10705) );
  INV_X1 U12530 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10703) );
  OR2_X1 U12531 ( .A1(n10322), .A2(n10703), .ZN(n10704) );
  INV_X1 U12532 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10708) );
  NAND2_X1 U12533 ( .A1(n7433), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10707) );
  NAND2_X1 U12534 ( .A1(n10710), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10706) );
  OAI211_X1 U12535 ( .C1(n10714), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n15164) );
  XNOR2_X1 U12536 ( .A(n15165), .B(n15164), .ZN(n10728) );
  INV_X1 U12537 ( .A(n10709), .ZN(n10715) );
  INV_X1 U12538 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U12539 ( .A1(n7433), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U12540 ( .A1(n10710), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n10711) );
  OAI211_X1 U12541 ( .C1(n10714), .C2(n10713), .A(n10712), .B(n10711), .ZN(
        n15475) );
  OAI21_X1 U12542 ( .B1(n15164), .B2(n10715), .A(n15475), .ZN(n10716) );
  INV_X1 U12543 ( .A(n10716), .ZN(n10719) );
  OR2_X1 U12544 ( .A1(n15618), .A2(n10309), .ZN(n10718) );
  INV_X1 U12545 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15617) );
  OR2_X1 U12546 ( .A1(n10322), .A2(n15617), .ZN(n10717) );
  MUX2_X1 U12547 ( .A(n10719), .B(n15171), .S(n10358), .Z(n10763) );
  INV_X1 U12548 ( .A(n10763), .ZN(n10724) );
  INV_X1 U12549 ( .A(n10720), .ZN(n10721) );
  OAI21_X1 U12550 ( .B1(n15164), .B2(n10721), .A(n15475), .ZN(n10722) );
  INV_X1 U12551 ( .A(n10722), .ZN(n10723) );
  MUX2_X1 U12552 ( .A(n15171), .B(n10723), .S(n10358), .Z(n10762) );
  NAND2_X1 U12553 ( .A1(n10724), .A2(n10762), .ZN(n10754) );
  OR2_X1 U12554 ( .A1(n11053), .A2(n15157), .ZN(n11565) );
  NAND2_X1 U12555 ( .A1(n11033), .A2(n15629), .ZN(n11048) );
  INV_X1 U12556 ( .A(n15629), .ZN(n11052) );
  NAND2_X1 U12557 ( .A1(n12597), .A2(n11052), .ZN(n11058) );
  NAND2_X1 U12558 ( .A1(n11048), .A2(n11058), .ZN(n10725) );
  AND2_X1 U12559 ( .A1(n11565), .A2(n10725), .ZN(n10752) );
  NAND3_X1 U12560 ( .A1(n10728), .A2(n10754), .A3(n10752), .ZN(n10769) );
  INV_X1 U12561 ( .A(n11033), .ZN(n12729) );
  NAND2_X1 U12562 ( .A1(n12729), .A2(n10727), .ZN(n11043) );
  INV_X1 U12563 ( .A(n11043), .ZN(n10760) );
  XOR2_X1 U12564 ( .A(n15475), .B(n15171), .Z(n10743) );
  XNOR2_X1 U12565 ( .A(n15483), .B(n15201), .ZN(n15185) );
  OR2_X1 U12566 ( .A1(n15495), .A2(n15243), .ZN(n10729) );
  NAND2_X1 U12567 ( .A1(n15238), .A2(n10729), .ZN(n15184) );
  XNOR2_X1 U12568 ( .A(n15509), .B(n15183), .ZN(n15288) );
  XNOR2_X1 U12569 ( .A(n15329), .B(n15197), .ZN(n15317) );
  NAND2_X1 U12570 ( .A1(n15533), .A2(n15182), .ZN(n10730) );
  NAND2_X1 U12571 ( .A1(n15196), .A2(n10730), .ZN(n15352) );
  XNOR2_X1 U12572 ( .A(n15396), .B(n15411), .ZN(n15382) );
  INV_X1 U12573 ( .A(n15387), .ZN(n15193) );
  XNOR2_X1 U12574 ( .A(n15538), .B(n15193), .ZN(n15365) );
  XNOR2_X1 U12575 ( .A(n15555), .B(n15385), .ZN(n15405) );
  INV_X1 U12576 ( .A(n15175), .ZN(n15186) );
  XNOR2_X1 U12577 ( .A(n15571), .B(n15186), .ZN(n15187) );
  XNOR2_X1 U12578 ( .A(n12967), .B(n14896), .ZN(n12758) );
  XNOR2_X1 U12579 ( .A(n12851), .B(n12722), .ZN(n12601) );
  XNOR2_X1 U12580 ( .A(n12712), .B(n15050), .ZN(n12460) );
  XNOR2_X1 U12581 ( .A(n16359), .B(n12508), .ZN(n12087) );
  INV_X1 U12582 ( .A(n15054), .ZN(n12195) );
  OR2_X1 U12583 ( .A1(n16350), .A2(n12195), .ZN(n12090) );
  NAND2_X1 U12584 ( .A1(n16350), .A2(n12195), .ZN(n10731) );
  NAND2_X1 U12585 ( .A1(n15462), .A2(n15452), .ZN(n11290) );
  NAND2_X1 U12586 ( .A1(n11303), .A2(n15061), .ZN(n10732) );
  AND2_X1 U12587 ( .A1(n11290), .A2(n10732), .ZN(n11745) );
  NAND4_X1 U12588 ( .A1(n11294), .A2(n11297), .A3(n11289), .A4(n11745), .ZN(
        n10733) );
  INV_X1 U12589 ( .A(n11544), .ZN(n11433) );
  NOR2_X1 U12590 ( .A1(n10733), .A2(n11433), .ZN(n10734) );
  XNOR2_X1 U12591 ( .A(n11890), .B(n15056), .ZN(n11547) );
  NAND4_X1 U12592 ( .A1(n12031), .A2(n10734), .A3(n11888), .A4(n11547), .ZN(
        n10735) );
  NOR2_X1 U12593 ( .A1(n12087), .A2(n10735), .ZN(n10736) );
  XNOR2_X1 U12594 ( .A(n12567), .B(n15051), .ZN(n12294) );
  XNOR2_X1 U12595 ( .A(n12496), .B(n15052), .ZN(n12123) );
  NAND4_X1 U12596 ( .A1(n12460), .A2(n10736), .A3(n12294), .A4(n12123), .ZN(
        n10737) );
  NOR4_X1 U12597 ( .A1(n15187), .A2(n12758), .A3(n12601), .A4(n10737), .ZN(
        n10738) );
  XNOR2_X1 U12598 ( .A(n15562), .B(n15177), .ZN(n15421) );
  XNOR2_X1 U12599 ( .A(n15579), .B(n15047), .ZN(n12761) );
  NAND4_X1 U12600 ( .A1(n15405), .A2(n10738), .A3(n15421), .A4(n12761), .ZN(
        n10739) );
  NOR4_X1 U12601 ( .A1(n15352), .A2(n15382), .A3(n15365), .A4(n10739), .ZN(
        n10740) );
  XNOR2_X1 U12602 ( .A(n15528), .B(n15319), .ZN(n15340) );
  NAND4_X1 U12603 ( .A1(n15288), .A2(n15317), .A3(n10740), .A4(n15340), .ZN(
        n10741) );
  NOR3_X1 U12604 ( .A1(n15184), .A2(n15302), .A3(n10741), .ZN(n10742) );
  XNOR2_X1 U12605 ( .A(n15501), .B(n15290), .ZN(n15274) );
  XNOR2_X1 U12606 ( .A(n7444), .B(n15414), .ZN(n10759) );
  NOR2_X1 U12607 ( .A1(n15164), .A2(n10752), .ZN(n10744) );
  OR2_X1 U12608 ( .A1(n15164), .A2(n10358), .ZN(n10748) );
  MUX2_X1 U12609 ( .A(n10752), .B(n10744), .S(n10748), .Z(n10757) );
  INV_X1 U12610 ( .A(n10752), .ZN(n10765) );
  NAND2_X1 U12611 ( .A1(n15164), .A2(n10765), .ZN(n10745) );
  NAND2_X1 U12612 ( .A1(n15164), .A2(n10358), .ZN(n10747) );
  MUX2_X1 U12613 ( .A(n10765), .B(n10745), .S(n10747), .Z(n10746) );
  OAI21_X1 U12614 ( .B1(n15165), .B2(n10746), .A(n11043), .ZN(n10756) );
  OR2_X1 U12615 ( .A1(n15165), .A2(n10747), .ZN(n10751) );
  INV_X1 U12616 ( .A(n10748), .ZN(n10749) );
  NAND2_X1 U12617 ( .A1(n15165), .A2(n10749), .ZN(n10750) );
  AND2_X1 U12618 ( .A1(n10751), .A2(n10750), .ZN(n10766) );
  INV_X1 U12619 ( .A(n10766), .ZN(n10753) );
  NOR3_X1 U12620 ( .A1(n10754), .A2(n10753), .A3(n10752), .ZN(n10755) );
  AOI211_X1 U12621 ( .C1(n15165), .C2(n10757), .A(n10756), .B(n10755), .ZN(
        n10758) );
  AOI21_X1 U12622 ( .B1(n10760), .B2(n10759), .A(n10758), .ZN(n10774) );
  INV_X1 U12623 ( .A(n10761), .ZN(n10767) );
  INV_X1 U12624 ( .A(n10762), .ZN(n10764) );
  NAND2_X1 U12625 ( .A1(n10764), .A2(n10763), .ZN(n10768) );
  NAND4_X1 U12626 ( .A1(n10766), .A2(n10768), .A3(n11043), .A4(n10765), .ZN(
        n10770) );
  OAI22_X1 U12627 ( .A1(n10771), .A2(n10770), .B1(n10769), .B2(n10768), .ZN(
        n10772) );
  NOR4_X2 U12628 ( .A1(n10775), .A2(n10774), .A3(n10773), .A4(n10772), .ZN(
        n10790) );
  NAND2_X1 U12629 ( .A1(n10777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10776) );
  XNOR2_X1 U12630 ( .A(n10776), .B(n7625), .ZN(n11039) );
  INV_X1 U12631 ( .A(n11039), .ZN(n10891) );
  NAND2_X1 U12632 ( .A1(n10891), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13029) );
  NAND2_X1 U12633 ( .A1(n10781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10782) );
  NOR2_X1 U12634 ( .A1(n13033), .A2(n15628), .ZN(n10785) );
  OR2_X1 U12635 ( .A1(n11048), .A2(n11034), .ZN(n11046) );
  NAND2_X1 U12636 ( .A1(n15609), .A2(n11046), .ZN(n11062) );
  NOR3_X1 U12637 ( .A1(n11062), .A2(n15622), .A3(n15451), .ZN(n10788) );
  OAI21_X1 U12638 ( .B1(n13029), .B2(n15629), .A(P1_B_REG_SCAN_IN), .ZN(n10787) );
  OAI21_X1 U12639 ( .B1(n10790), .B2(n13029), .A(n10789), .ZN(P1_U3242) );
  AOI22_X1 U12640 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n14775), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n7738), .ZN(n10800) );
  INV_X1 U12641 ( .A(n10800), .ZN(n10794) );
  XNOR2_X1 U12642 ( .A(n10799), .B(n10794), .ZN(n13181) );
  NAND2_X1 U12643 ( .A1(n13181), .A2(n13458), .ZN(n10796) );
  XNOR2_X1 U12644 ( .A(n13866), .B(n13607), .ZN(n13859) );
  NAND2_X1 U12645 ( .A1(n13280), .A2(n13316), .ZN(n13856) );
  NAND2_X1 U12646 ( .A1(n13866), .A2(n13656), .ZN(n10798) );
  NAND2_X1 U12647 ( .A1(n13858), .A2(n10798), .ZN(n10809) );
  OAI22_X1 U12648 ( .A1(n15619), .A2(n14769), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13192) );
  INV_X1 U12649 ( .A(n13192), .ZN(n10801) );
  XNOR2_X1 U12650 ( .A(n13191), .B(n10801), .ZN(n14236) );
  NOR2_X1 U12651 ( .A1(n8954), .A2(n15633), .ZN(n10802) );
  NAND2_X1 U12652 ( .A1(n13849), .A2(n10803), .ZN(n11927) );
  INV_X1 U12653 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10806) );
  NAND2_X1 U12654 ( .A1(n8960), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U12655 ( .A1(n10810), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U12656 ( .C1(n8800), .C2(n10806), .A(n10805), .B(n10804), .ZN(
        n10807) );
  INV_X1 U12657 ( .A(n10807), .ZN(n10808) );
  NAND2_X1 U12658 ( .A1(n11927), .A2(n10808), .ZN(n13860) );
  NOR2_X1 U12659 ( .A1(n13188), .A2(n13860), .ZN(n13466) );
  XNOR2_X1 U12660 ( .A(n10809), .B(n13617), .ZN(n10818) );
  INV_X1 U12661 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n10813) );
  NAND2_X1 U12662 ( .A1(n8960), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U12663 ( .A1(n10810), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10811) );
  OAI211_X1 U12664 ( .C1(n8800), .C2(n10813), .A(n10812), .B(n10811), .ZN(
        n10814) );
  INV_X1 U12665 ( .A(n10814), .ZN(n10815) );
  AND2_X1 U12666 ( .A1(n11927), .A2(n10815), .ZN(n13465) );
  INV_X1 U12667 ( .A(P3_B_REG_SCAN_IN), .ZN(n10816) );
  OAI21_X1 U12668 ( .B1(n13183), .B2(n10816), .A(n16313), .ZN(n13850) );
  OAI22_X1 U12669 ( .A1(n13607), .A2(n14092), .B1(n13465), .B2(n13850), .ZN(
        n10817) );
  NAND2_X1 U12670 ( .A1(n10819), .A2(n13595), .ZN(n13865) );
  INV_X1 U12671 ( .A(n13859), .ZN(n13864) );
  NAND2_X1 U12672 ( .A1(n13866), .A2(n13607), .ZN(n13609) );
  NAND2_X1 U12673 ( .A1(n13863), .A2(n13609), .ZN(n13469) );
  NAND2_X1 U12674 ( .A1(n13185), .A2(n10821), .ZN(n10824) );
  NAND2_X1 U12675 ( .A1(n10824), .A2(n16473), .ZN(n10823) );
  INV_X1 U12676 ( .A(n16473), .ZN(n10822) );
  NAND2_X1 U12677 ( .A1(n10826), .A2(n8494), .ZN(P3_U3456) );
  AND2_X1 U12678 ( .A1(n11171), .A2(n10827), .ZN(n11066) );
  INV_X1 U12679 ( .A(n10828), .ZN(n10829) );
  INV_X2 U12680 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U12681 ( .A1(n7434), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14229) );
  INV_X2 U12682 ( .A(n14229), .ZN(n13194) );
  OAI222_X1 U12683 ( .A1(n12245), .A2(P3_U3151), .B1(n13194), .B2(n10832), 
        .C1(n7764), .C2(n14237), .ZN(P3_U3289) );
  INV_X1 U12684 ( .A(n10833), .ZN(n10835) );
  INV_X1 U12685 ( .A(SI_9_), .ZN(n10834) );
  OAI222_X1 U12686 ( .A1(n13194), .A2(n10835), .B1(n14237), .B2(n10834), .C1(
        n16279), .C2(P3_U3151), .ZN(P3_U3286) );
  NOR2_X1 U12687 ( .A1(n7434), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15612) );
  OAI222_X1 U12688 ( .A1(n7555), .A2(n10836), .B1(n15627), .B2(n10840), .C1(
        P1_U3086), .C2(n15086), .ZN(P1_U3353) );
  INV_X1 U12689 ( .A(n10837), .ZN(n10845) );
  AND2_X1 U12690 ( .A1(n7434), .A2(P2_U3088), .ZN(n14771) );
  INV_X2 U12691 ( .A(n14771), .ZN(n14780) );
  AND2_X1 U12692 ( .A1(n10838), .A2(P2_U3088), .ZN(n13025) );
  AOI22_X1 U12693 ( .A1(n16078), .A2(P2_STATE_REG_SCAN_IN), .B1(n13025), .B2(
        P1_DATAO_REG_4__SCAN_IN), .ZN(n10839) );
  OAI21_X1 U12694 ( .B1(n10845), .B2(n14780), .A(n10839), .ZN(P2_U3323) );
  INV_X2 U12695 ( .A(n13025), .ZN(n14783) );
  INV_X1 U12696 ( .A(n11106), .ZN(n16042) );
  OAI222_X1 U12697 ( .A1(n14783), .A2(n10841), .B1(n14780), .B2(n10840), .C1(
        P2_U3088), .C2(n16042), .ZN(P2_U3325) );
  INV_X1 U12698 ( .A(n10842), .ZN(n10852) );
  OAI222_X1 U12699 ( .A1(n14783), .A2(n10843), .B1(n14780), .B2(n10852), .C1(
        P2_U3088), .C2(n16067), .ZN(P2_U3324) );
  INV_X1 U12700 ( .A(n15117), .ZN(n10844) );
  OAI222_X1 U12701 ( .A1(n7555), .A2(n8010), .B1(n15627), .B2(n10845), .C1(
        P1_U3086), .C2(n10844), .ZN(P1_U3351) );
  INV_X1 U12702 ( .A(n14419), .ZN(n10846) );
  OAI222_X1 U12703 ( .A1(n14783), .A2(n10847), .B1(n14780), .B2(n10851), .C1(
        P2_U3088), .C2(n10846), .ZN(P2_U3326) );
  INV_X1 U12704 ( .A(n10848), .ZN(n10850) );
  INV_X1 U12705 ( .A(SI_10_), .ZN(n10849) );
  OAI222_X1 U12706 ( .A1(n13194), .A2(n10850), .B1(n14237), .B2(n10849), .C1(
        n12900), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U12707 ( .A1(n8360), .A2(n7555), .B1(n15627), .B2(n10851), .C1(
        P1_U3086), .C2(n15067), .ZN(P1_U3354) );
  OAI222_X1 U12708 ( .A1(n7555), .A2(n10853), .B1(n15627), .B2(n10852), .C1(
        P1_U3086), .C2(n15098), .ZN(P1_U3352) );
  INV_X1 U12709 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10855) );
  INV_X1 U12710 ( .A(n10854), .ZN(n10856) );
  INV_X1 U12711 ( .A(n10927), .ZN(n10920) );
  OAI222_X1 U12712 ( .A1(n7555), .A2(n10855), .B1(n15627), .B2(n10856), .C1(
        P1_U3086), .C2(n10920), .ZN(P1_U3350) );
  INV_X1 U12713 ( .A(n11112), .ZN(n16094) );
  OAI222_X1 U12714 ( .A1(n14783), .A2(n10857), .B1(n14780), .B2(n10856), .C1(
        P2_U3088), .C2(n16094), .ZN(P2_U3322) );
  INV_X1 U12715 ( .A(n10858), .ZN(n10859) );
  INV_X1 U12716 ( .A(n13111), .ZN(n12909) );
  OAI222_X1 U12717 ( .A1(n13194), .A2(n10859), .B1(n14237), .B2(n15857), .C1(
        n12909), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12718 ( .A(n10860), .ZN(n10862) );
  INV_X1 U12719 ( .A(SI_7_), .ZN(n10861) );
  INV_X1 U12720 ( .A(n12246), .ZN(n12363) );
  OAI222_X1 U12721 ( .A1(n13194), .A2(n10862), .B1(n14237), .B2(n10861), .C1(
        n12363), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12722 ( .A1(P3_U3151), .A2(n12672), .B1(n14237), .B2(n10864), 
        .C1(n13194), .C2(n10863), .ZN(P3_U3287) );
  OAI222_X1 U12723 ( .A1(n13194), .A2(n10866), .B1(n14237), .B2(n10865), .C1(
        n11509), .C2(P3_U3151), .ZN(P3_U3294) );
  INV_X1 U12724 ( .A(n11664), .ZN(n11636) );
  INV_X1 U12725 ( .A(n10867), .ZN(n10868) );
  OAI222_X1 U12726 ( .A1(n11636), .A2(P3_U3151), .B1(n13194), .B2(n10868), 
        .C1(n15873), .C2(n14237), .ZN(P3_U3293) );
  INV_X1 U12727 ( .A(n10869), .ZN(n10871) );
  INV_X1 U12728 ( .A(SI_4_), .ZN(n10870) );
  OAI222_X1 U12729 ( .A1(n11780), .A2(P3_U3151), .B1(n13194), .B2(n10871), 
        .C1(n10870), .C2(n14237), .ZN(P3_U3291) );
  INV_X1 U12730 ( .A(n11677), .ZN(n11667) );
  INV_X1 U12731 ( .A(n10872), .ZN(n10874) );
  INV_X1 U12732 ( .A(SI_3_), .ZN(n10873) );
  OAI222_X1 U12733 ( .A1(n11667), .A2(P3_U3151), .B1(n13194), .B2(n10874), 
        .C1(n10873), .C2(n14237), .ZN(P3_U3292) );
  INV_X1 U12734 ( .A(n10875), .ZN(n10877) );
  INV_X1 U12735 ( .A(SI_5_), .ZN(n10876) );
  OAI222_X1 U12736 ( .A1(n8149), .A2(P3_U3151), .B1(n13194), .B2(n10877), .C1(
        n10876), .C2(n14237), .ZN(P3_U3290) );
  INV_X1 U12737 ( .A(n10878), .ZN(n10880) );
  OAI222_X1 U12738 ( .A1(n14783), .A2(n10879), .B1(n14780), .B2(n10880), .C1(
        P2_U3088), .C2(n16106), .ZN(P2_U3321) );
  INV_X1 U12739 ( .A(n10954), .ZN(n10935) );
  OAI222_X1 U12740 ( .A1(n7555), .A2(n10881), .B1(n15627), .B2(n10880), .C1(
        P1_U3086), .C2(n10935), .ZN(P1_U3349) );
  INV_X1 U12741 ( .A(n10882), .ZN(n10883) );
  INV_X1 U12742 ( .A(n13694), .ZN(n13701) );
  OAI222_X1 U12743 ( .A1(n13194), .A2(n10883), .B1(n14237), .B2(n15856), .C1(
        n13701), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12744 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10885) );
  INV_X1 U12745 ( .A(n10884), .ZN(n10886) );
  OAI222_X1 U12746 ( .A1(n14783), .A2(n10885), .B1(n14780), .B2(n10886), .C1(
        P2_U3088), .C2(n16118), .ZN(P2_U3320) );
  INV_X1 U12747 ( .A(n10955), .ZN(n10980) );
  OAI222_X1 U12748 ( .A1(n7555), .A2(n10887), .B1(n15627), .B2(n10886), .C1(
        P1_U3086), .C2(n10980), .ZN(P1_U3348) );
  INV_X1 U12749 ( .A(n10888), .ZN(n10936) );
  AOI22_X1 U12750 ( .A1(n10996), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n15625), .ZN(n10889) );
  OAI21_X1 U12751 ( .B1(n10936), .B2(n15627), .A(n10889), .ZN(P1_U3347) );
  INV_X1 U12752 ( .A(n15609), .ZN(n10890) );
  NAND2_X1 U12753 ( .A1(n10890), .A2(n13029), .ZN(n10912) );
  OR2_X1 U12754 ( .A1(n11048), .A2(n10891), .ZN(n10893) );
  AND2_X1 U12755 ( .A1(n10893), .A2(n7723), .ZN(n10910) );
  NAND2_X1 U12756 ( .A1(n10912), .A2(n10910), .ZN(n16199) );
  INV_X1 U12757 ( .A(n15622), .ZN(n16194) );
  MUX2_X1 U12758 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10334), .S(n10927), .Z(
        n10899) );
  MUX2_X1 U12759 ( .A(n10894), .B(P1_REG1_REG_2__SCAN_IN), .S(n15086), .Z(
        n15083) );
  INV_X1 U12760 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n16335) );
  MUX2_X1 U12761 ( .A(n16335), .B(P1_REG1_REG_1__SCAN_IN), .S(n15067), .Z(
        n15065) );
  AND2_X1 U12762 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15066) );
  NAND2_X1 U12763 ( .A1(n15065), .A2(n15066), .ZN(n15064) );
  OAI21_X1 U12764 ( .B1(n16335), .B2(n15067), .A(n15064), .ZN(n15082) );
  NAND2_X1 U12765 ( .A1(n15083), .A2(n15082), .ZN(n15101) );
  OR2_X1 U12766 ( .A1(n15086), .A2(n10894), .ZN(n15100) );
  NAND2_X1 U12767 ( .A1(n15101), .A2(n15100), .ZN(n10897) );
  MUX2_X1 U12768 ( .A(n10895), .B(P1_REG1_REG_3__SCAN_IN), .S(n15098), .Z(
        n10896) );
  NAND2_X1 U12769 ( .A1(n10897), .A2(n10896), .ZN(n15114) );
  OR2_X1 U12770 ( .A1(n15098), .A2(n10895), .ZN(n15113) );
  INV_X1 U12771 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11470) );
  MUX2_X1 U12772 ( .A(n11470), .B(P1_REG1_REG_4__SCAN_IN), .S(n15117), .Z(
        n15112) );
  NAND2_X1 U12773 ( .A1(n10898), .A2(n10899), .ZN(n10926) );
  OAI21_X1 U12774 ( .B1(n10899), .B2(n10898), .A(n10926), .ZN(n10917) );
  INV_X1 U12775 ( .A(n15073), .ZN(n15077) );
  OR2_X1 U12776 ( .A1(n16199), .A2(n15077), .ZN(n15149) );
  OR2_X1 U12777 ( .A1(n15073), .A2(n15622), .ZN(n10900) );
  MUX2_X1 U12778 ( .A(n11459), .B(P1_REG2_REG_2__SCAN_IN), .S(n15086), .Z(
        n15081) );
  MUX2_X1 U12779 ( .A(n15457), .B(P1_REG2_REG_1__SCAN_IN), .S(n15067), .Z(
        n15063) );
  AND2_X1 U12780 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15075) );
  NAND2_X1 U12781 ( .A1(n15063), .A2(n15075), .ZN(n15062) );
  OAI21_X1 U12782 ( .B1(n15457), .B2(n15067), .A(n15062), .ZN(n15080) );
  NAND2_X1 U12783 ( .A1(n15081), .A2(n15080), .ZN(n15096) );
  OR2_X1 U12784 ( .A1(n15086), .A2(n11459), .ZN(n15095) );
  NAND2_X1 U12785 ( .A1(n15096), .A2(n15095), .ZN(n10903) );
  INV_X1 U12786 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10901) );
  MUX2_X1 U12787 ( .A(n10901), .B(P1_REG2_REG_3__SCAN_IN), .S(n15098), .Z(
        n10902) );
  NAND2_X1 U12788 ( .A1(n10903), .A2(n10902), .ZN(n15108) );
  OR2_X1 U12789 ( .A1(n15098), .A2(n10901), .ZN(n15107) );
  NAND2_X1 U12790 ( .A1(n15108), .A2(n15107), .ZN(n10905) );
  MUX2_X1 U12791 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11529), .S(n15117), .Z(
        n10904) );
  NAND2_X1 U12792 ( .A1(n10905), .A2(n10904), .ZN(n15110) );
  NAND2_X1 U12793 ( .A1(n15117), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10907) );
  INV_X1 U12794 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10919) );
  MUX2_X1 U12795 ( .A(n10919), .B(P1_REG2_REG_5__SCAN_IN), .S(n10927), .Z(
        n10906) );
  AOI21_X1 U12796 ( .B1(n15110), .B2(n10907), .A(n10906), .ZN(n10923) );
  INV_X1 U12797 ( .A(n10923), .ZN(n10909) );
  NAND3_X1 U12798 ( .A1(n15110), .A2(n10907), .A3(n10906), .ZN(n10908) );
  NAND3_X1 U12799 ( .A1(n15154), .A2(n10909), .A3(n10908), .ZN(n10915) );
  INV_X1 U12800 ( .A(n10910), .ZN(n10911) );
  AND2_X1 U12801 ( .A1(n10912), .A2(n10911), .ZN(n16197) );
  AND2_X1 U12802 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10913) );
  AOI21_X1 U12803 ( .B1(n16197), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10913), .ZN(
        n10914) );
  OAI211_X1 U12804 ( .C1(n15149), .C2(n10920), .A(n10915), .B(n10914), .ZN(
        n10916) );
  AOI21_X1 U12805 ( .B1(n15155), .B2(n10917), .A(n10916), .ZN(n10918) );
  INV_X1 U12806 ( .A(n10918), .ZN(P1_U3248) );
  NOR2_X1 U12807 ( .A1(n10920), .A2(n10919), .ZN(n10922) );
  MUX2_X1 U12808 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11939), .S(n10954), .Z(
        n10921) );
  OAI21_X1 U12809 ( .B1(n10923), .B2(n10922), .A(n10921), .ZN(n10975) );
  OR3_X1 U12810 ( .A1(n10923), .A2(n10922), .A3(n10921), .ZN(n10924) );
  NAND3_X1 U12811 ( .A1(n15154), .A2(n10975), .A3(n10924), .ZN(n10934) );
  NAND2_X1 U12812 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11835) );
  INV_X1 U12813 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10925) );
  MUX2_X1 U12814 ( .A(n10925), .B(P1_REG1_REG_6__SCAN_IN), .S(n10954), .Z(
        n10929) );
  OAI21_X1 U12815 ( .B1(n10927), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10926), .ZN(
        n10928) );
  AOI211_X1 U12816 ( .C1(n10929), .C2(n10928), .A(n10949), .B(n12627), .ZN(
        n10930) );
  INV_X1 U12817 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U12818 ( .A1(n11835), .A2(n10931), .ZN(n10932) );
  AOI21_X1 U12819 ( .B1(n16197), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10932), .ZN(
        n10933) );
  OAI211_X1 U12820 ( .C1(n15149), .C2(n10935), .A(n10934), .B(n10933), .ZN(
        P1_U3249) );
  INV_X1 U12821 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10937) );
  INV_X1 U12822 ( .A(n11119), .ZN(n16131) );
  OAI222_X1 U12823 ( .A1(n14783), .A2(n10937), .B1(n14780), .B2(n10936), .C1(
        P2_U3088), .C2(n16131), .ZN(P2_U3319) );
  NOR2_X1 U12824 ( .A1(n16197), .A2(n15059), .ZN(P1_U3085) );
  OAI222_X1 U12825 ( .A1(n13697), .A2(P3_U3151), .B1(n13194), .B2(n10938), 
        .C1(n15855), .C2(n14237), .ZN(P3_U3282) );
  NAND2_X1 U12826 ( .A1(n10939), .A2(P2_U3947), .ZN(n10940) );
  OAI21_X1 U12827 ( .B1(n10703), .B2(P2_U3947), .A(n10940), .ZN(P2_U3562) );
  INV_X1 U12828 ( .A(n10941), .ZN(n10944) );
  INV_X1 U12829 ( .A(n11335), .ZN(n11328) );
  OAI222_X1 U12830 ( .A1(n7555), .A2(n10942), .B1(n15627), .B2(n10944), .C1(
        P1_U3086), .C2(n11328), .ZN(P1_U3346) );
  INV_X1 U12831 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10945) );
  INV_X1 U12832 ( .A(n11231), .ZN(n10943) );
  OAI222_X1 U12833 ( .A1(n14783), .A2(n10945), .B1(n14780), .B2(n10944), .C1(
        P2_U3088), .C2(n10943), .ZN(P2_U3318) );
  INV_X1 U12834 ( .A(n10946), .ZN(n10982) );
  AOI22_X1 U12835 ( .A1(n11347), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15625), .ZN(n10947) );
  OAI21_X1 U12836 ( .B1(n10982), .B2(n15627), .A(n10947), .ZN(P1_U3345) );
  OAI222_X1 U12837 ( .A1(n13194), .A2(n10948), .B1(n14237), .B2(n15851), .C1(
        n13734), .C2(P3_U3151), .ZN(P3_U3281) );
  AOI21_X1 U12838 ( .B1(n10954), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10949), .ZN(
        n10967) );
  MUX2_X1 U12839 ( .A(n10365), .B(P1_REG1_REG_7__SCAN_IN), .S(n10955), .Z(
        n10966) );
  AOI21_X1 U12840 ( .B1(n10955), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10965), .ZN(
        n10951) );
  INV_X1 U12841 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n16366) );
  MUX2_X1 U12842 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n16366), .S(n10996), .Z(
        n10950) );
  NOR2_X1 U12843 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  OAI21_X1 U12844 ( .B1(n10952), .B2(n10999), .A(n15155), .ZN(n10964) );
  INV_X1 U12845 ( .A(n15149), .ZN(n15118) );
  INV_X1 U12846 ( .A(n16197), .ZN(n15162) );
  INV_X1 U12847 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U12848 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n12194) );
  OAI21_X1 U12849 ( .B1(n15162), .B2(n10953), .A(n12194), .ZN(n10962) );
  NAND2_X1 U12850 ( .A1(n10954), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10974) );
  INV_X1 U12851 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10956) );
  MUX2_X1 U12852 ( .A(n10956), .B(P1_REG2_REG_7__SCAN_IN), .S(n10955), .Z(
        n10973) );
  AOI21_X1 U12853 ( .B1(n10975), .B2(n10974), .A(n10973), .ZN(n10972) );
  NOR2_X1 U12854 ( .A1(n10980), .A2(n10956), .ZN(n10958) );
  MUX2_X1 U12855 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n12095), .S(n10996), .Z(
        n10957) );
  OAI21_X1 U12856 ( .B1(n10972), .B2(n10958), .A(n10957), .ZN(n10994) );
  INV_X1 U12857 ( .A(n10994), .ZN(n10960) );
  NOR3_X1 U12858 ( .A1(n10972), .A2(n10958), .A3(n10957), .ZN(n10959) );
  NOR3_X1 U12859 ( .A1(n10960), .A2(n10959), .A3(n15150), .ZN(n10961) );
  AOI211_X1 U12860 ( .C1(n15118), .C2(n10996), .A(n10962), .B(n10961), .ZN(
        n10963) );
  NAND2_X1 U12861 ( .A1(n10964), .A2(n10963), .ZN(P1_U3251) );
  AND2_X1 U12862 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11974) );
  INV_X1 U12863 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10970) );
  AOI211_X1 U12864 ( .C1(n10967), .C2(n10966), .A(n12627), .B(n10965), .ZN(
        n10968) );
  INV_X1 U12865 ( .A(n10968), .ZN(n10969) );
  OAI21_X1 U12866 ( .B1(n10970), .B2(n15162), .A(n10969), .ZN(n10971) );
  NOR2_X1 U12867 ( .A1(n11974), .A2(n10971), .ZN(n10979) );
  INV_X1 U12868 ( .A(n10972), .ZN(n10977) );
  NAND3_X1 U12869 ( .A1(n10975), .A2(n10974), .A3(n10973), .ZN(n10976) );
  NAND3_X1 U12870 ( .A1(n10977), .A2(n15154), .A3(n10976), .ZN(n10978) );
  OAI211_X1 U12871 ( .C1(n15149), .C2(n10980), .A(n10979), .B(n10978), .ZN(
        P1_U3250) );
  INV_X1 U12872 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10983) );
  INV_X1 U12873 ( .A(n16187), .ZN(n10981) );
  OAI222_X1 U12874 ( .A1(n14783), .A2(n10983), .B1(n14780), .B2(n10982), .C1(
        P2_U3088), .C2(n10981), .ZN(P2_U3317) );
  AND2_X1 U12875 ( .A1(n10985), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12876 ( .A1(n10985), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12877 ( .A1(n10985), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12878 ( .A1(n10985), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12879 ( .A1(n10985), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12880 ( .A1(n10985), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12881 ( .A1(n10985), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12882 ( .A1(n10985), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12883 ( .A1(n10985), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12884 ( .A1(n10985), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12885 ( .A1(n10985), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12886 ( .A1(n10985), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12887 ( .A1(n10985), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12888 ( .A1(n10985), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12889 ( .A1(n10985), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12890 ( .A1(n10985), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12891 ( .A1(n10985), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12892 ( .A1(n10985), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12893 ( .A1(n10985), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12894 ( .A1(n10985), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12895 ( .A1(n10985), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12896 ( .A1(n10985), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12897 ( .A1(n10985), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12898 ( .A1(n10985), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12899 ( .A1(n10985), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12900 ( .A1(n10985), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12901 ( .A1(n10985), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12902 ( .A1(n10985), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12903 ( .A1(n10985), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12904 ( .A1(n10985), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  INV_X1 U12905 ( .A(n10986), .ZN(n10989) );
  AOI22_X1 U12906 ( .A1(n11604), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n15625), .ZN(n10987) );
  OAI21_X1 U12907 ( .B1(n10989), .B2(n15627), .A(n10987), .ZN(P1_U3344) );
  NAND2_X1 U12908 ( .A1(n15164), .A2(n15059), .ZN(n10988) );
  OAI21_X1 U12909 ( .B1(n10136), .B2(n15059), .A(n10988), .ZN(P1_U3591) );
  INV_X1 U12910 ( .A(n11236), .ZN(n16145) );
  OAI222_X1 U12911 ( .A1(n14783), .A2(n10990), .B1(n14780), .B2(n10989), .C1(
        P2_U3088), .C2(n16145), .ZN(P2_U3316) );
  OAI222_X1 U12912 ( .A1(n13194), .A2(n10991), .B1(n14237), .B2(n15850), .C1(
        n13773), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U12913 ( .A1(n10996), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10993) );
  INV_X1 U12914 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12131) );
  MUX2_X1 U12915 ( .A(n12131), .B(P1_REG2_REG_9__SCAN_IN), .S(n11335), .Z(
        n10992) );
  AOI21_X1 U12916 ( .B1(n10994), .B2(n10993), .A(n10992), .ZN(n11352) );
  NAND3_X1 U12917 ( .A1(n10994), .A2(n10993), .A3(n10992), .ZN(n10995) );
  NAND2_X1 U12918 ( .A1(n10995), .A2(n15154), .ZN(n11005) );
  NOR2_X1 U12919 ( .A1(n10996), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10997) );
  MUX2_X1 U12920 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10402), .S(n11335), .Z(
        n10998) );
  INV_X1 U12921 ( .A(n11334), .ZN(n11001) );
  NOR3_X1 U12922 ( .A1(n10999), .A2(n10998), .A3(n10997), .ZN(n11000) );
  OAI21_X1 U12923 ( .B1(n11001), .B2(n11000), .A(n15155), .ZN(n11004) );
  AND2_X1 U12924 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12510) );
  NOR2_X1 U12925 ( .A1(n15149), .A2(n11328), .ZN(n11002) );
  AOI211_X1 U12926 ( .C1(n16197), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n12510), .B(
        n11002), .ZN(n11003) );
  OAI211_X1 U12927 ( .C1(n11352), .C2(n11005), .A(n11004), .B(n11003), .ZN(
        P1_U3252) );
  INV_X1 U12928 ( .A(n11053), .ZN(n11006) );
  AND2_X2 U12929 ( .A1(n11006), .A2(n11040), .ZN(n11694) );
  INV_X1 U12930 ( .A(n11040), .ZN(n11007) );
  NAND2_X1 U12931 ( .A1(n11007), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n11010) );
  INV_X1 U12932 ( .A(n16428), .ZN(n11008) );
  NAND2_X1 U12933 ( .A1(n11008), .A2(n15157), .ZN(n11525) );
  AND2_X2 U12934 ( .A1(n11525), .A2(n11013), .ZN(n12699) );
  NAND2_X1 U12935 ( .A1(n12699), .A2(n15061), .ZN(n11009) );
  OAI211_X1 U12936 ( .C1(n11303), .C2(n11968), .A(n11010), .B(n11009), .ZN(
        n11132) );
  NOR2_X1 U12937 ( .A1(n11040), .A2(n11011), .ZN(n11012) );
  AOI21_X1 U12938 ( .B1(n15061), .B2(n11694), .A(n11012), .ZN(n11015) );
  OR2_X1 U12939 ( .A1(n11303), .A2(n11695), .ZN(n11014) );
  NAND2_X1 U12940 ( .A1(n11015), .A2(n11014), .ZN(n11131) );
  XNOR2_X1 U12941 ( .A(n11132), .B(n11131), .ZN(n15076) );
  NAND2_X1 U12942 ( .A1(n13033), .A2(P1_B_REG_SCAN_IN), .ZN(n11018) );
  INV_X1 U12943 ( .A(n15628), .ZN(n11029) );
  OAI21_X1 U12944 ( .B1(n13033), .B2(P1_B_REG_SCAN_IN), .A(n11029), .ZN(n11016) );
  INV_X1 U12945 ( .A(n11016), .ZN(n11017) );
  NOR4_X1 U12946 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n11027) );
  NOR4_X1 U12947 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n11026) );
  OR4_X1 U12948 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n11024) );
  NOR4_X1 U12949 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n11022) );
  NOR4_X1 U12950 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n11021) );
  NOR4_X1 U12951 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n11020) );
  NOR4_X1 U12952 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n11019) );
  NAND4_X1 U12953 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(
        n11023) );
  NOR4_X1 U12954 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n11024), .A4(n11023), .ZN(n11025) );
  AND3_X1 U12955 ( .A1(n11027), .A2(n11026), .A3(n11025), .ZN(n11028) );
  NOR2_X1 U12956 ( .A1(n15608), .A2(n11028), .ZN(n11061) );
  OR2_X1 U12957 ( .A1(n15608), .A2(P1_D_REG_1__SCAN_IN), .ZN(n11030) );
  OR2_X1 U12958 ( .A1(n13103), .A2(n11029), .ZN(n15610) );
  NAND2_X1 U12959 ( .A1(n11030), .A2(n15610), .ZN(n11450) );
  NOR2_X1 U12960 ( .A1(n11061), .A2(n11450), .ZN(n11032) );
  NAND2_X1 U12961 ( .A1(n13033), .A2(n15628), .ZN(n15611) );
  AND2_X1 U12962 ( .A1(n11032), .A2(n11184), .ZN(n11037) );
  AND2_X1 U12963 ( .A1(n11037), .A2(n15609), .ZN(n11047) );
  OR2_X1 U12964 ( .A1(n11033), .A2(n15629), .ZN(n11059) );
  INV_X1 U12965 ( .A(n11048), .ZN(n11035) );
  NOR2_X1 U12966 ( .A1(n16358), .A2(n11035), .ZN(n11036) );
  INV_X1 U12967 ( .A(n11037), .ZN(n11038) );
  NAND2_X1 U12968 ( .A1(n16326), .A2(n15414), .ZN(n11063) );
  NAND2_X1 U12969 ( .A1(n11038), .A2(n11063), .ZN(n11042) );
  AND3_X1 U12970 ( .A1(n11046), .A2(n11040), .A3(n11039), .ZN(n11041) );
  NAND2_X1 U12971 ( .A1(n11042), .A2(n11041), .ZN(n11710) );
  NOR2_X1 U12972 ( .A1(n11710), .A2(P1_U3086), .ZN(n11267) );
  INV_X1 U12973 ( .A(n11267), .ZN(n11143) );
  NOR2_X1 U12974 ( .A1(n11043), .A2(n15629), .ZN(n11460) );
  NAND2_X1 U12975 ( .A1(n11047), .A2(n11460), .ZN(n11045) );
  INV_X1 U12976 ( .A(n11063), .ZN(n11044) );
  AOI22_X1 U12977 ( .A1(n11143), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n15462), 
        .B2(n15042), .ZN(n11050) );
  NAND2_X1 U12978 ( .A1(n15029), .A2(n15448), .ZN(n15037) );
  INV_X1 U12979 ( .A(n15037), .ZN(n15006) );
  NAND2_X1 U12980 ( .A1(n15006), .A2(n15060), .ZN(n11049) );
  OAI211_X1 U12981 ( .C1(n15076), .C2(n15044), .A(n11050), .B(n11049), .ZN(
        P1_U3232) );
  NAND2_X1 U12982 ( .A1(n15629), .A2(n15157), .ZN(n11051) );
  OR2_X1 U12983 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  NAND2_X1 U12984 ( .A1(n11130), .A2(n11054), .ZN(n11456) );
  OR2_X1 U12985 ( .A1(n11456), .A2(n15414), .ZN(n11301) );
  NOR2_X1 U12986 ( .A1(n15445), .A2(n15584), .ZN(n11057) );
  OAI22_X1 U12987 ( .A1(n11291), .A2(n15410), .B1(n11745), .B2(n11057), .ZN(
        n11747) );
  OAI22_X1 U12988 ( .A1(n11745), .A2(n16353), .B1(n11303), .B2(n11059), .ZN(
        n11060) );
  NOR2_X1 U12989 ( .A1(n11747), .A2(n11060), .ZN(n11187) );
  OR2_X1 U12990 ( .A1(n11062), .A2(n11061), .ZN(n11453) );
  NAND2_X1 U12991 ( .A1(n11450), .A2(n11063), .ZN(n11064) );
  NOR2_X1 U12992 ( .A1(n11453), .A2(n11064), .ZN(n11185) );
  AND2_X2 U12993 ( .A1(n11185), .A2(n11451), .ZN(n16338) );
  OR2_X1 U12994 ( .A1(n16338), .A2(n10247), .ZN(n11065) );
  OAI21_X1 U12995 ( .B1(n11187), .B2(n16447), .A(n11065), .ZN(P1_U3459) );
  INV_X1 U12996 ( .A(n11066), .ZN(n11070) );
  NAND2_X1 U12997 ( .A1(n11162), .A2(n11171), .ZN(n11068) );
  NAND2_X1 U12998 ( .A1(n11068), .A2(n8042), .ZN(n11069) );
  AND2_X1 U12999 ( .A1(n11070), .A2(n11069), .ZN(n11082) );
  NAND2_X1 U13000 ( .A1(n11071), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14773) );
  INV_X1 U13001 ( .A(n14773), .ZN(n11072) );
  INV_X1 U13002 ( .A(n11074), .ZN(n11073) );
  OR2_X1 U13003 ( .A1(n11073), .A2(n14778), .ZN(n16182) );
  AND2_X1 U13004 ( .A1(n11074), .A2(n14778), .ZN(n16163) );
  NAND2_X1 U13005 ( .A1(n16163), .A2(n11075), .ZN(n11078) );
  NAND2_X1 U13006 ( .A1(n11077), .A2(n11076), .ZN(n16043) );
  OAI211_X1 U13007 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n16182), .A(n11078), .B(
        n16168), .ZN(n11081) );
  INV_X1 U13008 ( .A(n16163), .ZN(n16177) );
  OAI22_X1 U13009 ( .A1(n16177), .A2(n11075), .B1(n9379), .B2(n16182), .ZN(
        n11080) );
  MUX2_X1 U13010 ( .A(n11081), .B(n11080), .S(n11079), .Z(n11084) );
  AND2_X1 U13011 ( .A1(n11082), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16055) );
  OAI22_X1 U13012 ( .A1(n16191), .A2(n16201), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11931), .ZN(n11083) );
  OR2_X1 U13013 ( .A1(n11084), .A2(n11083), .ZN(P2_U3214) );
  INV_X1 U13014 ( .A(n11085), .ZN(n11129) );
  AOI22_X1 U13015 ( .A1(n11815), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15625), .ZN(n11086) );
  OAI21_X1 U13016 ( .B1(n11129), .B2(n15627), .A(n11086), .ZN(P1_U3343) );
  INV_X1 U13017 ( .A(n11087), .ZN(n11089) );
  INV_X1 U13018 ( .A(SI_16_), .ZN(n11088) );
  OAI222_X1 U13019 ( .A1(n13194), .A2(n11089), .B1(n14237), .B2(n11088), .C1(
        n13794), .C2(P3_U3151), .ZN(P3_U3279) );
  MUX2_X1 U13020 ( .A(n9512), .B(P2_REG2_REG_9__SCAN_IN), .S(n11231), .Z(
        n11102) );
  XNOR2_X1 U13021 ( .A(n11106), .B(n11535), .ZN(n16047) );
  XNOR2_X1 U13022 ( .A(n14419), .B(n11090), .ZN(n14418) );
  AND2_X1 U13023 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14417) );
  NAND2_X1 U13024 ( .A1(n14418), .A2(n14417), .ZN(n14416) );
  NAND2_X1 U13025 ( .A1(n14419), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U13026 ( .A1(n14416), .A2(n11091), .ZN(n16046) );
  NAND2_X1 U13027 ( .A1(n16047), .A2(n16046), .ZN(n16045) );
  NAND2_X1 U13028 ( .A1(n11106), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U13029 ( .A1(n16045), .A2(n11092), .ZN(n16062) );
  XNOR2_X1 U13030 ( .A(n16067), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n16063) );
  NAND2_X1 U13031 ( .A1(n16062), .A2(n16063), .ZN(n16061) );
  OR2_X1 U13032 ( .A1(n16067), .A2(n11093), .ZN(n11094) );
  NAND2_X1 U13033 ( .A1(n16061), .A2(n11094), .ZN(n16073) );
  XNOR2_X1 U13034 ( .A(n16078), .B(n11751), .ZN(n16074) );
  NAND2_X1 U13035 ( .A1(n16073), .A2(n16074), .ZN(n16072) );
  NAND2_X1 U13036 ( .A1(n16078), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13037 ( .A1(n16072), .A2(n11095), .ZN(n16087) );
  MUX2_X1 U13038 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11516), .S(n11112), .Z(
        n16088) );
  NAND2_X1 U13039 ( .A1(n16087), .A2(n16088), .ZN(n16086) );
  NAND2_X1 U13040 ( .A1(n11112), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U13041 ( .A1(n16086), .A2(n11096), .ZN(n16099) );
  XNOR2_X1 U13042 ( .A(n16106), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n16100) );
  NAND2_X1 U13043 ( .A1(n16099), .A2(n16100), .ZN(n16098) );
  NAND2_X1 U13044 ( .A1(n11114), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13045 ( .A1(n16098), .A2(n11097), .ZN(n16111) );
  MUX2_X1 U13046 ( .A(n9482), .B(P2_REG2_REG_7__SCAN_IN), .S(n16118), .Z(
        n16112) );
  NAND2_X1 U13047 ( .A1(n16111), .A2(n16112), .ZN(n16110) );
  NAND2_X1 U13048 ( .A1(n11116), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11098) );
  NAND2_X1 U13049 ( .A1(n16110), .A2(n11098), .ZN(n16125) );
  XNOR2_X1 U13050 ( .A(n11119), .B(n11880), .ZN(n16124) );
  NAND2_X1 U13051 ( .A1(n16125), .A2(n16124), .ZN(n16123) );
  NAND2_X1 U13052 ( .A1(n11119), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n11099) );
  NAND2_X1 U13053 ( .A1(n16123), .A2(n11099), .ZN(n11101) );
  OR2_X1 U13054 ( .A1(n11101), .A2(n11102), .ZN(n11228) );
  INV_X1 U13055 ( .A(n11228), .ZN(n11100) );
  AOI21_X1 U13056 ( .B1(n11102), .B2(n11101), .A(n11100), .ZN(n11127) );
  INV_X1 U13057 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n11103) );
  NAND2_X1 U13058 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n12224) );
  OAI21_X1 U13059 ( .B1(n16191), .B2(n11103), .A(n12224), .ZN(n11125) );
  INV_X1 U13060 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11104) );
  XNOR2_X1 U13061 ( .A(n11106), .B(n11104), .ZN(n16051) );
  XNOR2_X1 U13062 ( .A(n14419), .B(n7574), .ZN(n14415) );
  AND2_X1 U13063 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14414) );
  NAND2_X1 U13064 ( .A1(n14415), .A2(n14414), .ZN(n14413) );
  NAND2_X1 U13065 ( .A1(n14419), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U13066 ( .A1(n14413), .A2(n11105), .ZN(n16050) );
  NAND2_X1 U13067 ( .A1(n16051), .A2(n16050), .ZN(n16049) );
  NAND2_X1 U13068 ( .A1(n11106), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U13069 ( .A1(n16049), .A2(n11107), .ZN(n16059) );
  XNOR2_X1 U13070 ( .A(n16067), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n16060) );
  NAND2_X1 U13071 ( .A1(n16059), .A2(n16060), .ZN(n16058) );
  INV_X1 U13072 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11108) );
  OR2_X1 U13073 ( .A1(n16067), .A2(n11108), .ZN(n11109) );
  NAND2_X1 U13074 ( .A1(n16058), .A2(n11109), .ZN(n16076) );
  INV_X1 U13075 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11110) );
  XNOR2_X1 U13076 ( .A(n16078), .B(n11110), .ZN(n16077) );
  NAND2_X1 U13077 ( .A1(n16076), .A2(n16077), .ZN(n16075) );
  NAND2_X1 U13078 ( .A1(n16078), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U13079 ( .A1(n16075), .A2(n11111), .ZN(n16090) );
  MUX2_X1 U13080 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9439), .S(n11112), .Z(
        n16091) );
  NAND2_X1 U13081 ( .A1(n16090), .A2(n16091), .ZN(n16089) );
  NAND2_X1 U13082 ( .A1(n11112), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U13083 ( .A1(n16089), .A2(n11113), .ZN(n16102) );
  XNOR2_X1 U13084 ( .A(n16106), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n16103) );
  NAND2_X1 U13085 ( .A1(n16102), .A2(n16103), .ZN(n16101) );
  NAND2_X1 U13086 ( .A1(n11114), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11115) );
  NAND2_X1 U13087 ( .A1(n16101), .A2(n11115), .ZN(n16114) );
  MUX2_X1 U13088 ( .A(n9478), .B(P2_REG1_REG_7__SCAN_IN), .S(n16118), .Z(
        n16115) );
  NAND2_X1 U13089 ( .A1(n16114), .A2(n16115), .ZN(n16113) );
  NAND2_X1 U13090 ( .A1(n11116), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11117) );
  NAND2_X1 U13091 ( .A1(n16113), .A2(n11117), .ZN(n16128) );
  XNOR2_X1 U13092 ( .A(n11119), .B(n11118), .ZN(n16127) );
  NAND2_X1 U13093 ( .A1(n16128), .A2(n16127), .ZN(n16126) );
  NAND2_X1 U13094 ( .A1(n11119), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U13095 ( .A1(n16126), .A2(n11120), .ZN(n11122) );
  MUX2_X1 U13096 ( .A(n9508), .B(P2_REG1_REG_9__SCAN_IN), .S(n11231), .Z(
        n11121) );
  OR2_X1 U13097 ( .A1(n11122), .A2(n11121), .ZN(n11233) );
  NAND2_X1 U13098 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  AOI21_X1 U13099 ( .B1(n11233), .B2(n11123), .A(n16177), .ZN(n11124) );
  AOI211_X1 U13100 ( .C1(n16188), .C2(n11231), .A(n11125), .B(n11124), .ZN(
        n11126) );
  OAI21_X1 U13101 ( .B1(n11127), .B2(n16182), .A(n11126), .ZN(P2_U3223) );
  OAI222_X1 U13102 ( .A1(n14780), .A2(n11129), .B1(n11318), .B2(P2_U3088), 
        .C1(n11128), .C2(n14783), .ZN(P2_U3315) );
  AND2_X1 U13103 ( .A1(n7438), .A2(n11694), .ZN(n11133) );
  AOI21_X1 U13104 ( .B1(n15060), .B2(n12699), .A(n11133), .ZN(n11137) );
  NAND2_X1 U13105 ( .A1(n7438), .A2(n11013), .ZN(n11135) );
  NAND2_X1 U13106 ( .A1(n11136), .A2(n11137), .ZN(n11262) );
  INV_X1 U13107 ( .A(n11263), .ZN(n11140) );
  AOI21_X1 U13108 ( .B1(n11142), .B2(n11141), .A(n11140), .ZN(n11147) );
  AOI22_X1 U13109 ( .A1(n11143), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7438), .B2(
        n15042), .ZN(n11146) );
  NAND2_X1 U13110 ( .A1(n15029), .A2(n15386), .ZN(n15038) );
  INV_X1 U13111 ( .A(n15038), .ZN(n11144) );
  AOI22_X1 U13112 ( .A1(n11144), .A2(n15061), .B1(n15006), .B2(n15449), .ZN(
        n11145) );
  OAI211_X1 U13113 ( .C1(n11147), .C2(n15044), .A(n11146), .B(n11145), .ZN(
        P1_U3222) );
  INV_X1 U13114 ( .A(n11148), .ZN(n11149) );
  XNOR2_X1 U13115 ( .A(n14242), .B(n12000), .ZN(n11150) );
  INV_X1 U13116 ( .A(n14242), .ZN(n14254) );
  AOI22_X1 U13117 ( .A1(n11197), .A2(n14305), .B1(n14254), .B2(n16298), .ZN(
        n11207) );
  INV_X1 U13118 ( .A(n11152), .ZN(n11153) );
  AND2_X1 U13119 ( .A1(n9929), .A2(n14265), .ZN(n11155) );
  AOI21_X1 U13120 ( .B1(n11155), .B2(n11154), .A(n11156), .ZN(n11217) );
  INV_X1 U13121 ( .A(n11156), .ZN(n11157) );
  XNOR2_X1 U13122 ( .A(n11995), .B(n14242), .ZN(n11384) );
  NAND2_X1 U13123 ( .A1(n14409), .A2(n14305), .ZN(n11383) );
  XNOR2_X1 U13124 ( .A(n11384), .B(n11383), .ZN(n11385) );
  XNOR2_X1 U13125 ( .A(n11386), .B(n11385), .ZN(n11180) );
  OR2_X1 U13126 ( .A1(n16040), .A2(n11190), .ZN(n11158) );
  NOR2_X1 U13127 ( .A1(n11159), .A2(n11158), .ZN(n11168) );
  INV_X1 U13128 ( .A(n11166), .ZN(n11176) );
  NAND2_X1 U13129 ( .A1(n11161), .A2(n11160), .ZN(n16407) );
  INV_X1 U13130 ( .A(n11162), .ZN(n11163) );
  NAND2_X1 U13131 ( .A1(n16407), .A2(n11163), .ZN(n11164) );
  INV_X1 U13132 ( .A(n9929), .ZN(n11167) );
  INV_X1 U13133 ( .A(n14600), .ZN(n14621) );
  INV_X1 U13134 ( .A(n14583), .ZN(n14623) );
  OAI22_X1 U13135 ( .A1(n11167), .A2(n14621), .B1(n7437), .B2(n14623), .ZN(
        n11252) );
  AOI22_X1 U13136 ( .A1(n14328), .A2(n11252), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11179) );
  INV_X1 U13137 ( .A(n11168), .ZN(n11169) );
  NAND2_X1 U13138 ( .A1(n11169), .A2(n11191), .ZN(n11174) );
  AND3_X1 U13139 ( .A1(n11172), .A2(n11171), .A3(n11170), .ZN(n11173) );
  NAND2_X1 U13140 ( .A1(n11174), .A2(n11173), .ZN(n11203) );
  INV_X1 U13141 ( .A(n14373), .ZN(n14385) );
  INV_X1 U13142 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11991) );
  OR2_X1 U13143 ( .A1(n11176), .A2(n11175), .ZN(n11177) );
  AOI22_X1 U13144 ( .A1(n14385), .A2(n11991), .B1(n14375), .B2(n11249), .ZN(
        n11178) );
  OAI211_X1 U13145 ( .C1(n11180), .C2(n14377), .A(n11179), .B(n11178), .ZN(
        P2_U3190) );
  OAI222_X1 U13146 ( .A1(n13194), .A2(n11181), .B1(n14237), .B2(n15657), .C1(
        n13803), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13147 ( .A(n11182), .ZN(n11188) );
  INV_X1 U13148 ( .A(n12067), .ZN(n12072) );
  INV_X1 U13149 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n11183) );
  OAI222_X1 U13150 ( .A1(n14780), .A2(n11188), .B1(n12072), .B2(P2_U3088), 
        .C1(n11183), .C2(n14783), .ZN(P2_U3314) );
  INV_X1 U13151 ( .A(n16446), .ZN(n16444) );
  NAND2_X1 U13152 ( .A1(n16444), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11186) );
  OAI21_X1 U13153 ( .B1(n11187), .B2(n16444), .A(n11186), .ZN(P1_U3528) );
  INV_X1 U13154 ( .A(n12393), .ZN(n12385) );
  OAI222_X1 U13155 ( .A1(n7555), .A2(n11189), .B1(n15627), .B2(n11188), .C1(
        n12385), .C2(P1_U3086), .ZN(P1_U3342) );
  AND2_X1 U13156 ( .A1(n11190), .A2(n16041), .ZN(n16033) );
  INV_X2 U13157 ( .A(n16414), .ZN(n14760) );
  XNOR2_X1 U13158 ( .A(n11198), .B(n11223), .ZN(n11196) );
  NAND2_X1 U13159 ( .A1(n14412), .A2(n14600), .ZN(n11195) );
  NAND2_X1 U13160 ( .A1(n9929), .A2(n14604), .ZN(n11194) );
  NAND2_X1 U13161 ( .A1(n11195), .A2(n11194), .ZN(n11204) );
  AOI21_X1 U13162 ( .B1(n11196), .B2(n14603), .A(n11204), .ZN(n12007) );
  XNOR2_X1 U13163 ( .A(n11198), .B(n11197), .ZN(n12005) );
  INV_X1 U13164 ( .A(n14739), .ZN(n16374) );
  OAI211_X1 U13165 ( .C1(n11211), .C2(n16298), .A(n14734), .B(n11278), .ZN(
        n12003) );
  OAI21_X1 U13166 ( .B1(n11211), .B2(n16407), .A(n12003), .ZN(n11200) );
  AOI21_X1 U13167 ( .B1(n12005), .B2(n16374), .A(n11200), .ZN(n11201) );
  NAND2_X1 U13168 ( .A1(n12007), .A2(n11201), .ZN(n11256) );
  NAND2_X1 U13169 ( .A1(n14760), .A2(n11256), .ZN(n11202) );
  OAI21_X1 U13170 ( .B1(n14760), .B2(n9368), .A(n11202), .ZN(P2_U3433) );
  INV_X1 U13171 ( .A(n14375), .ZN(n14393) );
  NOR2_X1 U13172 ( .A1(n11203), .A2(P2_U3088), .ZN(n11226) );
  INV_X1 U13173 ( .A(n11226), .ZN(n11214) );
  AOI22_X1 U13174 ( .A1(n11214), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n14328), 
        .B2(n11204), .ZN(n11210) );
  OAI21_X1 U13175 ( .B1(n11207), .B2(n11206), .A(n11205), .ZN(n11208) );
  NAND2_X1 U13176 ( .A1(n14382), .A2(n11208), .ZN(n11209) );
  OAI211_X1 U13177 ( .C1(n11211), .C2(n14393), .A(n11210), .B(n11209), .ZN(
        P2_U3194) );
  NAND2_X1 U13178 ( .A1(n14411), .A2(n14600), .ZN(n11213) );
  NAND2_X1 U13179 ( .A1(n14409), .A2(n14604), .ZN(n11212) );
  NAND2_X1 U13180 ( .A1(n11213), .A2(n11212), .ZN(n11282) );
  AOI22_X1 U13181 ( .A1(n11214), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n14328), 
        .B2(n11282), .ZN(n11220) );
  OAI21_X1 U13182 ( .B1(n11217), .B2(n11216), .A(n11215), .ZN(n11218) );
  NAND2_X1 U13183 ( .A1(n11218), .A2(n14382), .ZN(n11219) );
  OAI211_X1 U13184 ( .C1(n11539), .C2(n14393), .A(n11220), .B(n11219), .ZN(
        P2_U3209) );
  INV_X1 U13185 ( .A(n14387), .ZN(n14370) );
  AOI22_X1 U13186 ( .A1(n14370), .A2(n14411), .B1(n7635), .B2(n14375), .ZN(
        n11225) );
  MUX2_X1 U13187 ( .A(n7635), .B(n11221), .S(n14305), .Z(n11222) );
  OAI21_X1 U13188 ( .B1(n11223), .B2(n11222), .A(n14382), .ZN(n11224) );
  OAI211_X1 U13189 ( .C1(n11226), .C2(n11931), .A(n11225), .B(n11224), .ZN(
        P2_U3204) );
  OR2_X1 U13190 ( .A1(n11231), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U13191 ( .A1(n11228), .A2(n11227), .ZN(n16183) );
  MUX2_X1 U13192 ( .A(n11229), .B(P2_REG2_REG_10__SCAN_IN), .S(n16187), .Z(
        n16184) );
  OR2_X1 U13193 ( .A1(n16183), .A2(n16184), .ZN(n16180) );
  NAND2_X1 U13194 ( .A1(n16187), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11230) );
  AND2_X1 U13195 ( .A1(n16180), .A2(n11230), .ZN(n16137) );
  XNOR2_X1 U13196 ( .A(n11236), .B(n12322), .ZN(n16138) );
  NAND2_X1 U13197 ( .A1(n16137), .A2(n16138), .ZN(n16136) );
  OAI21_X1 U13198 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n11236), .A(n16136), 
        .ZN(n11317) );
  XOR2_X1 U13199 ( .A(n11318), .B(n11317), .Z(n11319) );
  XOR2_X1 U13200 ( .A(n16457), .B(n11319), .Z(n11245) );
  INV_X1 U13201 ( .A(n11318), .ZN(n11243) );
  NAND2_X1 U13202 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12690)
         );
  OAI21_X1 U13203 ( .B1(n16191), .B2(n16230), .A(n12690), .ZN(n11242) );
  MUX2_X1 U13204 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11314), .S(n11318), .Z(
        n11239) );
  INV_X1 U13205 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11237) );
  OR2_X1 U13206 ( .A1(n11231), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11232) );
  NAND2_X1 U13207 ( .A1(n11233), .A2(n11232), .ZN(n16178) );
  MUX2_X1 U13208 ( .A(n11234), .B(P2_REG1_REG_10__SCAN_IN), .S(n16187), .Z(
        n16179) );
  OR2_X1 U13209 ( .A1(n16178), .A2(n16179), .ZN(n16175) );
  NAND2_X1 U13210 ( .A1(n16187), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U13211 ( .A1(n16175), .A2(n11235), .ZN(n16142) );
  MUX2_X1 U13212 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11237), .S(n11236), .Z(
        n16141) );
  NAND2_X1 U13213 ( .A1(n16142), .A2(n16141), .ZN(n16140) );
  OAI21_X1 U13214 ( .B1(n16145), .B2(n11237), .A(n16140), .ZN(n11238) );
  NOR2_X1 U13215 ( .A1(n11238), .A2(n11239), .ZN(n11313) );
  AOI21_X1 U13216 ( .B1(n11239), .B2(n11238), .A(n11313), .ZN(n11240) );
  NOR2_X1 U13217 ( .A1(n11240), .A2(n16177), .ZN(n11241) );
  AOI211_X1 U13218 ( .C1(n16188), .C2(n11243), .A(n11242), .B(n11241), .ZN(
        n11244) );
  OAI21_X1 U13219 ( .B1(n11245), .B2(n16182), .A(n11244), .ZN(P2_U3226) );
  INV_X1 U13220 ( .A(n16040), .ZN(n11246) );
  XNOR2_X1 U13221 ( .A(n11248), .B(n11250), .ZN(n11990) );
  INV_X2 U13222 ( .A(n16407), .ZN(n14733) );
  AOI211_X1 U13223 ( .C1(n11249), .C2(n11276), .A(n14692), .B(n11401), .ZN(
        n11992) );
  AOI21_X1 U13224 ( .B1(n14733), .B2(n11249), .A(n11992), .ZN(n11254) );
  XNOR2_X1 U13225 ( .A(n11251), .B(n11250), .ZN(n11253) );
  AOI21_X1 U13226 ( .B1(n11253), .B2(n14603), .A(n11252), .ZN(n11999) );
  OAI211_X1 U13227 ( .C1(n14739), .C2(n11990), .A(n11254), .B(n11999), .ZN(
        n11272) );
  NAND2_X1 U13228 ( .A1(n11272), .A2(n16413), .ZN(n11255) );
  OAI21_X1 U13229 ( .B1(n16413), .B2(n11108), .A(n11255), .ZN(P2_U3502) );
  NAND2_X1 U13230 ( .A1(n16413), .A2(n11256), .ZN(n11257) );
  OAI21_X1 U13231 ( .B1(n16413), .B2(n7574), .A(n11257), .ZN(P2_U3500) );
  NAND2_X1 U13232 ( .A1(n15449), .A2(n11694), .ZN(n11259) );
  NAND2_X1 U13233 ( .A1(n11372), .A2(n14856), .ZN(n11258) );
  NAND2_X1 U13234 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  XNOR2_X1 U13235 ( .A(n11260), .B(n11130), .ZN(n11680) );
  AND2_X1 U13236 ( .A1(n11372), .A2(n11694), .ZN(n11261) );
  AOI21_X1 U13237 ( .B1(n15449), .B2(n12699), .A(n11261), .ZN(n11681) );
  XNOR2_X1 U13238 ( .A(n11680), .B(n11681), .ZN(n11266) );
  NAND2_X1 U13239 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  OAI21_X1 U13240 ( .B1(n11266), .B2(n11265), .A(n11684), .ZN(n11270) );
  OAI22_X1 U13241 ( .A1(n15026), .A2(n11462), .B1(n11267), .B2(n11461), .ZN(
        n11269) );
  INV_X1 U13242 ( .A(n15058), .ZN(n11712) );
  OAI22_X1 U13243 ( .A1(n11291), .A2(n15038), .B1(n15037), .B2(n11712), .ZN(
        n11268) );
  AOI211_X1 U13244 ( .C1(n11270), .C2(n15012), .A(n11269), .B(n11268), .ZN(
        n11271) );
  INV_X1 U13245 ( .A(n11271), .ZN(P1_U3237) );
  NAND2_X1 U13246 ( .A1(n11272), .A2(n14760), .ZN(n11273) );
  OAI21_X1 U13247 ( .B1(n14760), .B2(n9406), .A(n11273), .ZN(P2_U3439) );
  XNOR2_X1 U13248 ( .A(n11275), .B(n11274), .ZN(n11541) );
  INV_X1 U13249 ( .A(n11541), .ZN(n11285) );
  INV_X1 U13250 ( .A(n11276), .ZN(n11277) );
  AOI211_X1 U13251 ( .C1(n11279), .C2(n11278), .A(n14692), .B(n11277), .ZN(
        n11537) );
  AOI21_X1 U13252 ( .B1(n14733), .B2(n11279), .A(n11537), .ZN(n11284) );
  XNOR2_X1 U13253 ( .A(n11281), .B(n11280), .ZN(n11283) );
  AOI21_X1 U13254 ( .B1(n11283), .B2(n14603), .A(n11282), .ZN(n11543) );
  OAI211_X1 U13255 ( .C1(n14739), .C2(n11285), .A(n11284), .B(n11543), .ZN(
        n14741) );
  NAND2_X1 U13256 ( .A1(n14741), .A2(n14760), .ZN(n11286) );
  OAI21_X1 U13257 ( .B1(n14760), .B2(n9389), .A(n11286), .ZN(P2_U3436) );
  INV_X1 U13258 ( .A(n11287), .ZN(n11288) );
  INV_X1 U13259 ( .A(n13827), .ZN(n13816) );
  OAI222_X1 U13260 ( .A1(n13194), .A2(n11288), .B1(n14237), .B2(n15843), .C1(
        n13816), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13261 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n11308) );
  INV_X1 U13262 ( .A(n11289), .ZN(n11299) );
  INV_X1 U13263 ( .A(n11290), .ZN(n15447) );
  NAND2_X1 U13264 ( .A1(n11291), .A2(n7438), .ZN(n11366) );
  NAND2_X1 U13265 ( .A1(n15446), .A2(n11366), .ZN(n11292) );
  NAND2_X1 U13266 ( .A1(n11292), .A2(n11297), .ZN(n11369) );
  NAND2_X1 U13267 ( .A1(n11302), .A2(n11372), .ZN(n11293) );
  XNOR2_X1 U13268 ( .A(n11299), .B(n11438), .ZN(n11727) );
  INV_X1 U13269 ( .A(n11294), .ZN(n11295) );
  OR2_X1 U13270 ( .A1(n11303), .A2(n15452), .ZN(n15441) );
  NAND2_X1 U13271 ( .A1(n11295), .A2(n15441), .ZN(n15444) );
  NAND2_X1 U13272 ( .A1(n15444), .A2(n11296), .ZN(n11364) );
  INV_X1 U13273 ( .A(n11297), .ZN(n11367) );
  NAND2_X1 U13274 ( .A1(n11364), .A2(n11367), .ZN(n11363) );
  NAND2_X1 U13275 ( .A1(n11302), .A2(n11462), .ZN(n11298) );
  NAND2_X1 U13276 ( .A1(n11363), .A2(n11298), .ZN(n11300) );
  NAND2_X1 U13277 ( .A1(n11300), .A2(n11299), .ZN(n11432) );
  OAI21_X1 U13278 ( .B1(n11300), .B2(n11299), .A(n11432), .ZN(n11725) );
  INV_X1 U13279 ( .A(n15057), .ZN(n11697) );
  OAI22_X1 U13280 ( .A1(n11697), .A2(n15410), .B1(n11302), .B2(n15451), .ZN(
        n14915) );
  INV_X1 U13281 ( .A(n14915), .ZN(n11304) );
  NAND2_X1 U13282 ( .A1(n16330), .A2(n11303), .ZN(n16328) );
  OAI211_X1 U13283 ( .C1(n11371), .C2(n11436), .A(n16326), .B(n11445), .ZN(
        n11723) );
  OAI211_X1 U13284 ( .C1(n11436), .C2(n16437), .A(n11304), .B(n11723), .ZN(
        n11305) );
  AOI21_X1 U13285 ( .B1(n11725), .B2(n15568), .A(n11305), .ZN(n11306) );
  OAI21_X1 U13286 ( .B1(n15567), .B2(n11727), .A(n11306), .ZN(n11427) );
  NAND2_X1 U13287 ( .A1(n11427), .A2(n16338), .ZN(n11307) );
  OAI21_X1 U13288 ( .B1(n16338), .B2(n11308), .A(n11307), .ZN(P1_U3468) );
  INV_X1 U13289 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U13290 ( .A1(n13484), .A2(P3_U3897), .ZN(n11309) );
  OAI21_X1 U13291 ( .B1(P3_U3897), .B2(n11310), .A(n11309), .ZN(P3_U3492) );
  INV_X1 U13292 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n11312) );
  NAND2_X1 U13293 ( .A1(n14046), .A2(P3_U3897), .ZN(n11311) );
  OAI21_X1 U13294 ( .B1(P3_U3897), .B2(n11312), .A(n11311), .ZN(P3_U3506) );
  AOI21_X1 U13295 ( .B1(n11318), .B2(n11314), .A(n11313), .ZN(n11316) );
  INV_X1 U13296 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12996) );
  MUX2_X1 U13297 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n12996), .S(n12067), .Z(
        n11315) );
  AND2_X1 U13298 ( .A1(n11316), .A2(n11315), .ZN(n12066) );
  OAI21_X1 U13299 ( .B1(n11316), .B2(n11315), .A(n16163), .ZN(n11325) );
  AOI22_X1 U13300 ( .A1(n11319), .A2(n16457), .B1(n11318), .B2(n11317), .ZN(
        n11321) );
  XOR2_X1 U13301 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n12067), .Z(n11320) );
  NAND2_X1 U13302 ( .A1(n11321), .A2(n11320), .ZN(n12070) );
  INV_X1 U13303 ( .A(n16182), .ZN(n16171) );
  OAI211_X1 U13304 ( .C1(n11321), .C2(n11320), .A(n12070), .B(n16171), .ZN(
        n11324) );
  AND2_X1 U13305 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12779) );
  NOR2_X1 U13306 ( .A1(n16168), .A2(n12072), .ZN(n11322) );
  AOI211_X1 U13307 ( .C1(n16055), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n12779), 
        .B(n11322), .ZN(n11323) );
  OAI211_X1 U13308 ( .C1(n12066), .C2(n11325), .A(n11324), .B(n11323), .ZN(
        P2_U3227) );
  INV_X1 U13309 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n11327) );
  NAND2_X1 U13310 ( .A1(n13134), .A2(P3_U3897), .ZN(n11326) );
  OAI21_X1 U13311 ( .B1(P3_U3897), .B2(n11327), .A(n11326), .ZN(P3_U3501) );
  NOR2_X1 U13312 ( .A1(n11328), .A2(n12131), .ZN(n11346) );
  INV_X1 U13313 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11329) );
  MUX2_X1 U13314 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11329), .S(n11347), .Z(
        n11330) );
  OAI21_X1 U13315 ( .B1(n11352), .B2(n11346), .A(n11330), .ZN(n11350) );
  NAND2_X1 U13316 ( .A1(n11347), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11332) );
  MUX2_X1 U13317 ( .A(n10433), .B(P1_REG2_REG_11__SCAN_IN), .S(n11604), .Z(
        n11331) );
  AOI21_X1 U13318 ( .B1(n11350), .B2(n11332), .A(n11331), .ZN(n11599) );
  NAND3_X1 U13319 ( .A1(n11350), .A2(n11332), .A3(n11331), .ZN(n11333) );
  NAND2_X1 U13320 ( .A1(n11333), .A2(n15154), .ZN(n11343) );
  OAI21_X1 U13321 ( .B1(n11335), .B2(P1_REG1_REG_9__SCAN_IN), .A(n11334), .ZN(
        n11354) );
  MUX2_X1 U13322 ( .A(n10419), .B(P1_REG1_REG_10__SCAN_IN), .S(n11347), .Z(
        n11355) );
  INV_X1 U13323 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n16433) );
  MUX2_X1 U13324 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n16433), .S(n11604), .Z(
        n11336) );
  NOR2_X1 U13325 ( .A1(n11337), .A2(n11336), .ZN(n11338) );
  OAI21_X1 U13326 ( .B1(n11338), .B2(n11607), .A(n15155), .ZN(n11342) );
  NAND2_X1 U13327 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n12707)
         );
  OAI21_X1 U13328 ( .B1(n15162), .B2(n11339), .A(n12707), .ZN(n11340) );
  AOI21_X1 U13329 ( .B1(n11604), .B2(n15118), .A(n11340), .ZN(n11341) );
  OAI211_X1 U13330 ( .C1(n11599), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        P1_U3254) );
  INV_X1 U13331 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n11345) );
  NAND2_X1 U13332 ( .A1(n13981), .A2(P3_U3897), .ZN(n11344) );
  OAI21_X1 U13333 ( .B1(P3_U3897), .B2(n11345), .A(n11344), .ZN(P3_U3509) );
  INV_X1 U13334 ( .A(n11347), .ZN(n11361) );
  INV_X1 U13335 ( .A(n11346), .ZN(n11349) );
  MUX2_X1 U13336 ( .A(n11329), .B(P1_REG2_REG_10__SCAN_IN), .S(n11347), .Z(
        n11348) );
  NAND2_X1 U13337 ( .A1(n11349), .A2(n11348), .ZN(n11351) );
  OAI211_X1 U13338 ( .C1(n11352), .C2(n11351), .A(n11350), .B(n15154), .ZN(
        n11360) );
  NAND2_X1 U13339 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n12562)
         );
  AOI211_X1 U13340 ( .C1(n11355), .C2(n11354), .A(n11353), .B(n12627), .ZN(
        n11356) );
  INV_X1 U13341 ( .A(n11356), .ZN(n11357) );
  NAND2_X1 U13342 ( .A1(n12562), .A2(n11357), .ZN(n11358) );
  AOI21_X1 U13343 ( .B1(n16197), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11358), 
        .ZN(n11359) );
  OAI211_X1 U13344 ( .C1(n15149), .C2(n11361), .A(n11360), .B(n11359), .ZN(
        P1_U3253) );
  NAND2_X1 U13345 ( .A1(n14537), .A2(P2_U3947), .ZN(n11362) );
  OAI21_X1 U13346 ( .B1(n13031), .B2(P2_U3947), .A(n11362), .ZN(P2_U3554) );
  INV_X1 U13347 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11375) );
  OAI21_X1 U13348 ( .B1(n11364), .B2(n11367), .A(n11363), .ZN(n11365) );
  INV_X1 U13349 ( .A(n11365), .ZN(n11467) );
  NAND3_X1 U13350 ( .A1(n15446), .A2(n11367), .A3(n11366), .ZN(n11368) );
  NAND2_X1 U13351 ( .A1(n11369), .A2(n11368), .ZN(n11370) );
  AOI222_X1 U13352 ( .A1(n15584), .A2(n11370), .B1(n15058), .B2(n15448), .C1(
        n15060), .C2(n15386), .ZN(n11458) );
  AOI211_X1 U13353 ( .C1(n11372), .C2(n16328), .A(n16428), .B(n11371), .ZN(
        n11464) );
  AOI21_X1 U13354 ( .B1(n15563), .B2(n11372), .A(n11464), .ZN(n11373) );
  OAI211_X1 U13355 ( .C1(n16425), .C2(n11467), .A(n11458), .B(n11373), .ZN(
        n11376) );
  NAND2_X1 U13356 ( .A1(n11376), .A2(n16338), .ZN(n11374) );
  OAI21_X1 U13357 ( .B1(n16338), .B2(n11375), .A(n11374), .ZN(P1_U3465) );
  NAND2_X1 U13358 ( .A1(n11376), .A2(n16446), .ZN(n11377) );
  OAI21_X1 U13359 ( .B1(n16446), .B2(n10894), .A(n11377), .ZN(P1_U3530) );
  INV_X1 U13360 ( .A(n11378), .ZN(n11381) );
  INV_X1 U13361 ( .A(n16158), .ZN(n11379) );
  OAI222_X1 U13362 ( .A1(n14783), .A2(n11380), .B1(n14780), .B2(n11381), .C1(
        P2_U3088), .C2(n11379), .ZN(P2_U3313) );
  INV_X1 U13363 ( .A(n12394), .ZN(n12622) );
  OAI222_X1 U13364 ( .A1(n7555), .A2(n11382), .B1(n15627), .B2(n11381), .C1(
        P1_U3086), .C2(n12622), .ZN(P1_U3341) );
  XNOR2_X1 U13365 ( .A(n11404), .B(n14254), .ZN(n11388) );
  NAND2_X1 U13366 ( .A1(n11388), .A2(n11387), .ZN(n11413) );
  OAI21_X1 U13367 ( .B1(n11388), .B2(n11387), .A(n11413), .ZN(n11389) );
  AOI21_X1 U13368 ( .B1(n11390), .B2(n11389), .A(n11415), .ZN(n11394) );
  NAND2_X1 U13369 ( .A1(n14328), .A2(n14600), .ZN(n14362) );
  INV_X1 U13370 ( .A(n14362), .ZN(n14390) );
  NAND2_X1 U13371 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n16083) );
  OAI21_X1 U13372 ( .B1(n14373), .B2(n11750), .A(n16083), .ZN(n11392) );
  OAI22_X1 U13373 ( .A1(n11841), .A2(n14387), .B1(n14393), .B2(n11752), .ZN(
        n11391) );
  AOI211_X1 U13374 ( .C1(n14390), .C2(n14409), .A(n11392), .B(n11391), .ZN(
        n11393) );
  OAI21_X1 U13375 ( .B1(n11394), .B2(n14377), .A(n11393), .ZN(P2_U3202) );
  XNOR2_X1 U13376 ( .A(n11395), .B(n11396), .ZN(n11756) );
  INV_X1 U13377 ( .A(n11756), .ZN(n11406) );
  XNOR2_X1 U13378 ( .A(n11397), .B(n11396), .ZN(n11399) );
  AOI22_X1 U13379 ( .A1(n14600), .A2(n14409), .B1(n14407), .B2(n14604), .ZN(
        n11398) );
  OAI21_X1 U13380 ( .B1(n11399), .B2(n14619), .A(n11398), .ZN(n11400) );
  AOI21_X1 U13381 ( .B1(n14522), .B2(n11756), .A(n11400), .ZN(n11759) );
  INV_X1 U13382 ( .A(n11401), .ZN(n11403) );
  INV_X1 U13383 ( .A(n11477), .ZN(n11402) );
  AOI21_X1 U13384 ( .B1(n11404), .B2(n11403), .A(n11402), .ZN(n11755) );
  AOI22_X1 U13385 ( .A1(n11755), .A2(n14734), .B1(n14733), .B2(n11404), .ZN(
        n11405) );
  OAI211_X1 U13386 ( .C1(n16299), .C2(n11406), .A(n11759), .B(n11405), .ZN(
        n11408) );
  NAND2_X1 U13387 ( .A1(n11408), .A2(n16413), .ZN(n11407) );
  OAI21_X1 U13388 ( .B1(n16413), .B2(n11110), .A(n11407), .ZN(P2_U3503) );
  INV_X1 U13389 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11410) );
  NAND2_X1 U13390 ( .A1(n11408), .A2(n14760), .ZN(n11409) );
  OAI21_X1 U13391 ( .B1(n14760), .B2(n11410), .A(n11409), .ZN(P2_U3442) );
  INV_X1 U13392 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U13393 ( .A1(n13389), .A2(P3_U3897), .ZN(n11411) );
  OAI21_X1 U13394 ( .B1(P3_U3897), .B2(n11412), .A(n11411), .ZN(P3_U3514) );
  INV_X1 U13395 ( .A(n11413), .ZN(n11414) );
  XNOR2_X1 U13396 ( .A(n11517), .B(n14254), .ZN(n11417) );
  NAND2_X1 U13397 ( .A1(n14407), .A2(n14305), .ZN(n11416) );
  NAND2_X1 U13398 ( .A1(n11417), .A2(n11416), .ZN(n11613) );
  OAI21_X1 U13399 ( .B1(n11417), .B2(n11416), .A(n11613), .ZN(n11418) );
  AOI21_X1 U13400 ( .B1(n11419), .B2(n11418), .A(n11615), .ZN(n11426) );
  NAND2_X1 U13401 ( .A1(n14408), .A2(n14600), .ZN(n11421) );
  NAND2_X1 U13402 ( .A1(n14406), .A2(n14604), .ZN(n11420) );
  NAND2_X1 U13403 ( .A1(n11421), .A2(n11420), .ZN(n11474) );
  NAND2_X1 U13404 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n16096) );
  INV_X1 U13405 ( .A(n16096), .ZN(n11422) );
  AOI21_X1 U13406 ( .B1(n14328), .B2(n11474), .A(n11422), .ZN(n11423) );
  OAI21_X1 U13407 ( .B1(n11518), .B2(n14373), .A(n11423), .ZN(n11424) );
  AOI21_X1 U13408 ( .B1(n11517), .B2(n14375), .A(n11424), .ZN(n11425) );
  OAI21_X1 U13409 ( .B1(n11426), .B2(n14377), .A(n11425), .ZN(P2_U3199) );
  NAND2_X1 U13410 ( .A1(n11427), .A2(n16446), .ZN(n11428) );
  OAI21_X1 U13411 ( .B1(n16446), .B2(n10895), .A(n11428), .ZN(P1_U3531) );
  INV_X1 U13412 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n11430) );
  NAND2_X1 U13413 ( .A1(n8598), .A2(P3_U3897), .ZN(n11429) );
  OAI21_X1 U13414 ( .B1(P3_U3897), .B2(n11430), .A(n11429), .ZN(P3_U3493) );
  INV_X1 U13415 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U13416 ( .A1(n11712), .A2(n11436), .ZN(n11431) );
  NAND2_X1 U13417 ( .A1(n11432), .A2(n11431), .ZN(n11434) );
  NAND2_X1 U13418 ( .A1(n11434), .A2(n11433), .ZN(n11549) );
  OAI21_X1 U13419 ( .B1(n11434), .B2(n11433), .A(n11549), .ZN(n11435) );
  INV_X1 U13420 ( .A(n11435), .ZN(n11533) );
  NAND2_X1 U13421 ( .A1(n15058), .A2(n11436), .ZN(n11437) );
  NAND2_X1 U13422 ( .A1(n11438), .A2(n11437), .ZN(n11440) );
  NAND2_X1 U13423 ( .A1(n11712), .A2(n10314), .ZN(n11439) );
  XNOR2_X1 U13424 ( .A(n11545), .B(n11544), .ZN(n11441) );
  NAND2_X1 U13425 ( .A1(n11441), .A2(n15584), .ZN(n11443) );
  AOI22_X1 U13426 ( .A1(n15386), .A2(n15058), .B1(n15056), .B2(n15448), .ZN(
        n11442) );
  NAND2_X1 U13427 ( .A1(n11443), .A2(n11442), .ZN(n11526) );
  INV_X1 U13428 ( .A(n11526), .ZN(n11447) );
  INV_X1 U13429 ( .A(n11552), .ZN(n11444) );
  AOI21_X1 U13430 ( .B1(n11715), .B2(n11445), .A(n11444), .ZN(n11527) );
  AOI22_X1 U13431 ( .A1(n11527), .A2(n16326), .B1(n15563), .B2(n11715), .ZN(
        n11446) );
  OAI211_X1 U13432 ( .C1(n11533), .C2(n16425), .A(n11447), .B(n11446), .ZN(
        n11468) );
  NAND2_X1 U13433 ( .A1(n11468), .A2(n16338), .ZN(n11448) );
  OAI21_X1 U13434 ( .B1(n16338), .B2(n11449), .A(n11448), .ZN(P1_U3471) );
  INV_X1 U13435 ( .A(n11450), .ZN(n11452) );
  NAND2_X1 U13436 ( .A1(n11452), .A2(n11451), .ZN(n11454) );
  INV_X1 U13437 ( .A(n15205), .ZN(n11455) );
  INV_X2 U13438 ( .A(n15432), .ZN(n15356) );
  INV_X1 U13439 ( .A(n11456), .ZN(n11457) );
  NAND2_X1 U13440 ( .A1(n15430), .A2(n11457), .ZN(n15342) );
  MUX2_X1 U13441 ( .A(n11459), .B(n11458), .S(n15430), .Z(n11466) );
  AND2_X1 U13442 ( .A1(n15205), .A2(n15157), .ZN(n15437) );
  OAI22_X1 U13443 ( .A1(n15434), .A2(n11462), .B1(n15428), .B2(n11461), .ZN(
        n11463) );
  AOI21_X1 U13444 ( .B1(n11464), .B2(n15437), .A(n11463), .ZN(n11465) );
  OAI211_X1 U13445 ( .C1(n11467), .C2(n15342), .A(n11466), .B(n11465), .ZN(
        P1_U3291) );
  NAND2_X1 U13446 ( .A1(n11468), .A2(n16446), .ZN(n11469) );
  OAI21_X1 U13447 ( .B1(n16446), .B2(n11470), .A(n11469), .ZN(P1_U3532) );
  XOR2_X1 U13448 ( .A(n11473), .B(n11471), .Z(n11524) );
  XOR2_X1 U13449 ( .A(n11473), .B(n11472), .Z(n11475) );
  AOI21_X1 U13450 ( .B1(n11475), .B2(n14603), .A(n11474), .ZN(n11515) );
  INV_X1 U13451 ( .A(n11847), .ZN(n11476) );
  AOI211_X1 U13452 ( .C1(n11517), .C2(n11477), .A(n14692), .B(n11476), .ZN(
        n11521) );
  AOI21_X1 U13453 ( .B1(n14733), .B2(n11517), .A(n11521), .ZN(n11478) );
  OAI211_X1 U13454 ( .C1(n11524), .C2(n14739), .A(n11515), .B(n11478), .ZN(
        n11480) );
  NAND2_X1 U13455 ( .A1(n11480), .A2(n16413), .ZN(n11479) );
  OAI21_X1 U13456 ( .B1(n16413), .B2(n9439), .A(n11479), .ZN(P2_U3504) );
  INV_X1 U13457 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U13458 ( .A1(n11480), .A2(n14760), .ZN(n11481) );
  OAI21_X1 U13459 ( .B1(n14760), .B2(n11482), .A(n11481), .ZN(P2_U3445) );
  NOR2_X1 U13460 ( .A1(n11483), .A2(P3_U3151), .ZN(n12256) );
  OR2_X1 U13461 ( .A1(n11595), .A2(n12256), .ZN(n11502) );
  NAND2_X1 U13462 ( .A1(n13605), .A2(n11483), .ZN(n11484) );
  NAND2_X1 U13463 ( .A1(n7432), .A2(n11484), .ZN(n11501) );
  INV_X1 U13464 ( .A(n11501), .ZN(n11486) );
  NAND2_X1 U13465 ( .A1(n11502), .A2(n11486), .ZN(n11495) );
  INV_X2 U13466 ( .A(P3_U3897), .ZN(n13666) );
  MUX2_X1 U13467 ( .A(n11495), .B(n13666), .S(n13648), .Z(n16278) );
  MUX2_X1 U13468 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13775), .Z(n16257) );
  INV_X1 U13469 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n16264) );
  NOR2_X1 U13470 ( .A1(n16257), .A2(n16264), .ZN(n16262) );
  OAI21_X1 U13471 ( .B1(n11487), .B2(n16262), .A(n11641), .ZN(n11507) );
  NAND2_X1 U13472 ( .A1(P3_U3897), .A2(n13183), .ZN(n16259) );
  NOR2_X2 U13473 ( .A1(n11495), .A2(n11488), .ZN(n13840) );
  NOR2_X1 U13474 ( .A1(n11915), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11489) );
  NAND2_X1 U13475 ( .A1(n8592), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11620) );
  INV_X1 U13476 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11490) );
  OR2_X1 U13477 ( .A1(n11491), .A2(n11490), .ZN(n11621) );
  NAND2_X1 U13478 ( .A1(n11491), .A2(n11490), .ZN(n11492) );
  NAND2_X1 U13479 ( .A1(n11621), .A2(n11492), .ZN(n11493) );
  NAND2_X1 U13480 ( .A1(n13840), .A2(n11493), .ZN(n11505) );
  NOR2_X1 U13481 ( .A1(n11496), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11497) );
  NAND2_X1 U13482 ( .A1(n8592), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n11625) );
  OAI21_X1 U13483 ( .B1(n11509), .B2(n11497), .A(n11625), .ZN(n11498) );
  NAND2_X1 U13484 ( .A1(n11498), .A2(n8568), .ZN(n11499) );
  NAND2_X1 U13485 ( .A1(n11626), .A2(n11499), .ZN(n11500) );
  NAND2_X1 U13486 ( .A1(n13847), .A2(n11500), .ZN(n11504) );
  AND2_X1 U13487 ( .A1(n11502), .A2(n11501), .ZN(n16037) );
  AOI22_X1 U13488 ( .A1(n16037), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11503) );
  NAND3_X1 U13489 ( .A1(n11505), .A2(n11504), .A3(n11503), .ZN(n11506) );
  AOI21_X1 U13490 ( .B1(n11507), .B2(n16272), .A(n11506), .ZN(n11508) );
  OAI21_X1 U13491 ( .B1(n11509), .B2(n16278), .A(n11508), .ZN(P3_U3183) );
  NAND2_X1 U13492 ( .A1(n15320), .A2(n15059), .ZN(n11510) );
  OAI21_X1 U13493 ( .B1(n15059), .B2(n11511), .A(n11510), .ZN(P1_U3583) );
  INV_X1 U13494 ( .A(n11512), .ZN(n11513) );
  OAI222_X1 U13495 ( .A1(P3_U3151), .A2(n13837), .B1(n14237), .B2(n11514), 
        .C1(n13194), .C2(n11513), .ZN(P3_U3276) );
  MUX2_X1 U13496 ( .A(n11516), .B(n11515), .S(n16458), .Z(n11523) );
  INV_X1 U13497 ( .A(n11517), .ZN(n11519) );
  OAI22_X1 U13498 ( .A1(n14631), .A2(n11519), .B1(n11518), .B2(n16455), .ZN(
        n11520) );
  AOI21_X1 U13499 ( .B1(n11521), .B2(n14596), .A(n11520), .ZN(n11522) );
  OAI211_X1 U13500 ( .C1(n14638), .C2(n11524), .A(n11523), .B(n11522), .ZN(
        P2_U3260) );
  INV_X1 U13501 ( .A(n11525), .ZN(n11937) );
  AOI21_X1 U13502 ( .B1(n11937), .B2(n11527), .A(n11526), .ZN(n11528) );
  MUX2_X1 U13503 ( .A(n11529), .B(n11528), .S(n15430), .Z(n11532) );
  INV_X1 U13504 ( .A(n11711), .ZN(n11530) );
  INV_X1 U13505 ( .A(n15428), .ZN(n15458) );
  AOI22_X1 U13506 ( .A1(n15459), .A2(n11715), .B1(n11530), .B2(n15458), .ZN(
        n11531) );
  OAI211_X1 U13507 ( .C1(n11533), .C2(n15342), .A(n11532), .B(n11531), .ZN(
        P1_U3289) );
  OAI22_X1 U13508 ( .A1(n16458), .A2(n11535), .B1(n11534), .B2(n16455), .ZN(
        n11536) );
  AOI21_X1 U13509 ( .B1(n14596), .B2(n11537), .A(n11536), .ZN(n11538) );
  OAI21_X1 U13510 ( .B1(n11539), .B2(n14631), .A(n11538), .ZN(n11540) );
  AOI21_X1 U13511 ( .B1(n11541), .B2(n14617), .A(n11540), .ZN(n11542) );
  OAI21_X1 U13512 ( .B1(n14598), .B2(n11543), .A(n11542), .ZN(P2_U3263) );
  INV_X1 U13513 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U13514 ( .A1(n11697), .A2(n11715), .ZN(n11546) );
  XNOR2_X1 U13515 ( .A(n11894), .B(n11550), .ZN(n11576) );
  NAND2_X1 U13516 ( .A1(n11697), .A2(n11696), .ZN(n11548) );
  NAND2_X1 U13517 ( .A1(n11549), .A2(n11548), .ZN(n11551) );
  NAND2_X1 U13518 ( .A1(n11551), .A2(n11550), .ZN(n11887) );
  OAI21_X1 U13519 ( .B1(n11551), .B2(n11550), .A(n11887), .ZN(n11574) );
  AOI21_X1 U13520 ( .B1(n11552), .B2(n11890), .A(n16428), .ZN(n11553) );
  NAND2_X1 U13521 ( .A1(n11553), .A2(n11901), .ZN(n11568) );
  NAND2_X1 U13522 ( .A1(n15055), .A2(n15448), .ZN(n11555) );
  NAND2_X1 U13523 ( .A1(n15057), .A2(n15386), .ZN(n11554) );
  NAND2_X1 U13524 ( .A1(n11555), .A2(n11554), .ZN(n11740) );
  AOI21_X1 U13525 ( .B1(n16358), .B2(n11890), .A(n11740), .ZN(n11556) );
  NAND2_X1 U13526 ( .A1(n11568), .A2(n11556), .ZN(n11557) );
  AOI21_X1 U13527 ( .B1(n11574), .B2(n15568), .A(n11557), .ZN(n11558) );
  OAI21_X1 U13528 ( .B1(n15567), .B2(n11576), .A(n11558), .ZN(n15589) );
  NAND2_X1 U13529 ( .A1(n15589), .A2(n16338), .ZN(n11559) );
  OAI21_X1 U13530 ( .B1(n16338), .B2(n11560), .A(n11559), .ZN(P1_U3474) );
  INV_X1 U13531 ( .A(n11561), .ZN(n11563) );
  OAI222_X1 U13532 ( .A1(n14783), .A2(n11562), .B1(n14780), .B2(n11563), .C1(
        P2_U3088), .C2(n12273), .ZN(P2_U3312) );
  INV_X1 U13533 ( .A(n12805), .ZN(n12629) );
  OAI222_X1 U13534 ( .A1(n7555), .A2(n11564), .B1(n15627), .B2(n11563), .C1(
        P1_U3086), .C2(n12629), .ZN(P1_U3340) );
  AND2_X1 U13535 ( .A1(n15430), .A2(n15584), .ZN(n15269) );
  INV_X1 U13536 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U13537 ( .A1(n15430), .A2(n11566), .ZN(n12127) );
  NAND2_X1 U13538 ( .A1(n15430), .A2(n15445), .ZN(n11567) );
  NAND2_X1 U13539 ( .A1(n12127), .A2(n11567), .ZN(n15224) );
  INV_X1 U13540 ( .A(n15437), .ZN(n15168) );
  NOR2_X1 U13541 ( .A1(n11568), .A2(n15168), .ZN(n11573) );
  INV_X1 U13542 ( .A(n11890), .ZN(n11891) );
  INV_X1 U13543 ( .A(n11740), .ZN(n11569) );
  MUX2_X1 U13544 ( .A(n11569), .B(n10919), .S(n15356), .Z(n11571) );
  OR2_X1 U13545 ( .A1(n15428), .A2(n11737), .ZN(n11570) );
  OAI211_X1 U13546 ( .C1(n11891), .C2(n15434), .A(n11571), .B(n11570), .ZN(
        n11572) );
  AOI211_X1 U13547 ( .C1(n11574), .C2(n15224), .A(n11573), .B(n11572), .ZN(
        n11575) );
  OAI21_X1 U13548 ( .B1(n11576), .B2(n15440), .A(n11575), .ZN(P1_U3288) );
  NAND2_X1 U13549 ( .A1(n11594), .A2(n11587), .ZN(n11582) );
  INV_X1 U13550 ( .A(n11577), .ZN(n11581) );
  NAND2_X1 U13551 ( .A1(n11592), .A2(n11578), .ZN(n11580) );
  NAND4_X1 U13552 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  NAND2_X1 U13553 ( .A1(n11583), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11585) );
  NAND2_X1 U13554 ( .A1(n11595), .A2(n11762), .ZN(n11803) );
  INV_X1 U13555 ( .A(n11803), .ZN(n13649) );
  AOI21_X1 U13556 ( .B1(n11592), .B2(n13649), .A(n12256), .ZN(n11584) );
  NAND2_X1 U13557 ( .A1(n13447), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11808) );
  INV_X1 U13558 ( .A(n11808), .ZN(n13205) );
  NAND2_X1 U13559 ( .A1(n16312), .A2(n11855), .ZN(n13486) );
  INV_X1 U13560 ( .A(n13486), .ZN(n11586) );
  OR2_X1 U13561 ( .A1(n11586), .A2(n16306), .ZN(n13619) );
  NAND2_X1 U13562 ( .A1(n11587), .A2(n16467), .ZN(n11589) );
  OAI22_X1 U13563 ( .A1(n11594), .A2(n11589), .B1(n11592), .B2(n11588), .ZN(
        n11590) );
  INV_X1 U13564 ( .A(n11802), .ZN(n11591) );
  NOR2_X1 U13565 ( .A1(n11803), .A2(n11591), .ZN(n11593) );
  INV_X1 U13566 ( .A(n11592), .ZN(n11804) );
  NAND2_X1 U13567 ( .A1(n11594), .A2(n13645), .ZN(n11596) );
  AND2_X1 U13568 ( .A1(n11595), .A2(n16418), .ZN(n11914) );
  OAI22_X1 U13569 ( .A1(n12154), .A2(n13446), .B1(n11855), .B2(n13453), .ZN(
        n11597) );
  AOI21_X1 U13570 ( .B1(n13619), .B2(n13442), .A(n11597), .ZN(n11598) );
  OAI21_X1 U13571 ( .B1(n13205), .B2(n16263), .A(n11598), .ZN(P3_U3172) );
  MUX2_X1 U13572 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12614), .S(n11815), .Z(
        n11601) );
  AOI21_X1 U13573 ( .B1(n11604), .B2(P1_REG2_REG_11__SCAN_IN), .A(n11599), 
        .ZN(n11600) );
  NAND2_X1 U13574 ( .A1(n11600), .A2(n11601), .ZN(n11814) );
  OAI21_X1 U13575 ( .B1(n11601), .B2(n11600), .A(n11814), .ZN(n11611) );
  NAND2_X1 U13576 ( .A1(n15118), .A2(n11815), .ZN(n11602) );
  NAND2_X1 U13577 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12856)
         );
  OAI211_X1 U13578 ( .C1(n11603), .C2(n15162), .A(n11602), .B(n12856), .ZN(
        n11610) );
  NOR2_X1 U13579 ( .A1(n11604), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11605) );
  INV_X1 U13580 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n16445) );
  MUX2_X1 U13581 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n16445), .S(n11815), .Z(
        n11606) );
  OAI21_X1 U13582 ( .B1(n11607), .B2(n11605), .A(n11606), .ZN(n11811) );
  OR3_X1 U13583 ( .A1(n11607), .A2(n11606), .A3(n11605), .ZN(n11608) );
  AOI21_X1 U13584 ( .B1(n11811), .B2(n11608), .A(n12627), .ZN(n11609) );
  AOI211_X1 U13585 ( .C1(n15154), .C2(n11611), .A(n11610), .B(n11609), .ZN(
        n11612) );
  INV_X1 U13586 ( .A(n11612), .ZN(P1_U3255) );
  INV_X1 U13587 ( .A(n11613), .ZN(n11614) );
  XNOR2_X1 U13588 ( .A(n11979), .B(n14306), .ZN(n11859) );
  NAND2_X1 U13589 ( .A1(n14406), .A2(n14305), .ZN(n11858) );
  XNOR2_X1 U13590 ( .A(n11859), .B(n11858), .ZN(n11861) );
  XNOR2_X1 U13591 ( .A(n11862), .B(n11861), .ZN(n11619) );
  AOI22_X1 U13592 ( .A1(n14370), .A2(n14405), .B1(n14390), .B2(n14407), .ZN(
        n11616) );
  NAND2_X1 U13593 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n16108) );
  OAI211_X1 U13594 ( .C1(n11980), .C2(n14373), .A(n11616), .B(n16108), .ZN(
        n11617) );
  AOI21_X1 U13595 ( .B1(n11979), .B2(n14375), .A(n11617), .ZN(n11618) );
  OAI21_X1 U13596 ( .B1(n11619), .B2(n14377), .A(n11618), .ZN(P2_U3211) );
  NAND2_X1 U13597 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  OAI21_X1 U13598 ( .B1(n11623), .B2(n11622), .A(n11659), .ZN(n11624) );
  NAND2_X1 U13599 ( .A1(n13840), .A2(n11624), .ZN(n11633) );
  XNOR2_X1 U13600 ( .A(n11664), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U13601 ( .A1(n11628), .A2(n11627), .ZN(n11666) );
  OAI21_X1 U13602 ( .B1(n11628), .B2(n11627), .A(n11666), .ZN(n11629) );
  NAND2_X1 U13603 ( .A1(n13847), .A2(n11629), .ZN(n11632) );
  NOR2_X1 U13604 ( .A1(n16340), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11630) );
  AOI21_X1 U13605 ( .B1(n16037), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n11630), .ZN(
        n11631) );
  NAND3_X1 U13606 ( .A1(n11633), .A2(n11632), .A3(n11631), .ZN(n11645) );
  INV_X1 U13607 ( .A(n11634), .ZN(n11640) );
  INV_X1 U13608 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11663) );
  MUX2_X1 U13609 ( .A(n11657), .B(n11663), .S(n13775), .Z(n11635) );
  NAND2_X1 U13610 ( .A1(n11635), .A2(n11664), .ZN(n11647) );
  INV_X1 U13611 ( .A(n11635), .ZN(n11637) );
  NAND2_X1 U13612 ( .A1(n11637), .A2(n11636), .ZN(n11638) );
  NAND2_X1 U13613 ( .A1(n11647), .A2(n11638), .ZN(n11639) );
  AOI21_X1 U13614 ( .B1(n11641), .B2(n11640), .A(n11639), .ZN(n11654) );
  INV_X1 U13615 ( .A(n11654), .ZN(n11643) );
  NAND3_X1 U13616 ( .A1(n11641), .A2(n11640), .A3(n11639), .ZN(n11642) );
  AOI21_X1 U13617 ( .B1(n11643), .B2(n11642), .A(n16259), .ZN(n11644) );
  AOI211_X1 U13618 ( .C1(n13813), .C2(n11664), .A(n11645), .B(n11644), .ZN(
        n11646) );
  INV_X1 U13619 ( .A(n11646), .ZN(P3_U3184) );
  INV_X1 U13620 ( .A(n11647), .ZN(n11653) );
  INV_X1 U13621 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11648) );
  MUX2_X1 U13622 ( .A(n8147), .B(n11648), .S(n13775), .Z(n11649) );
  NAND2_X1 U13623 ( .A1(n11649), .A2(n11677), .ZN(n13667) );
  INV_X1 U13624 ( .A(n11649), .ZN(n11650) );
  NAND2_X1 U13625 ( .A1(n11650), .A2(n11667), .ZN(n11651) );
  AND2_X1 U13626 ( .A1(n13667), .A2(n11651), .ZN(n11652) );
  INV_X1 U13627 ( .A(n13669), .ZN(n11656) );
  NOR3_X1 U13628 ( .A1(n11654), .A2(n11653), .A3(n11652), .ZN(n11655) );
  OAI21_X1 U13629 ( .B1(n11656), .B2(n11655), .A(n16272), .ZN(n11679) );
  OR2_X1 U13630 ( .A1(n11664), .A2(n11657), .ZN(n11658) );
  NAND2_X1 U13631 ( .A1(n11659), .A2(n11658), .ZN(n11660) );
  OAI21_X1 U13632 ( .B1(n11661), .B2(P3_REG2_REG_3__SCAN_IN), .A(n13683), .ZN(
        n11662) );
  NAND2_X1 U13633 ( .A1(n13840), .A2(n11662), .ZN(n11675) );
  OR2_X1 U13634 ( .A1(n11664), .A2(n11663), .ZN(n11665) );
  NAND2_X1 U13635 ( .A1(n11666), .A2(n11665), .ZN(n11668) );
  NAND2_X1 U13636 ( .A1(n11668), .A2(n11667), .ZN(n13673) );
  OR2_X1 U13637 ( .A1(n11668), .A2(n11667), .ZN(n11669) );
  OAI21_X1 U13638 ( .B1(n11670), .B2(P3_REG1_REG_3__SCAN_IN), .A(n13675), .ZN(
        n11671) );
  NAND2_X1 U13639 ( .A1(n13847), .A2(n11671), .ZN(n11674) );
  INV_X1 U13640 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11672) );
  NOR2_X1 U13641 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11672), .ZN(n12147) );
  AOI21_X1 U13642 ( .B1(n16037), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n12147), .ZN(
        n11673) );
  NAND3_X1 U13643 ( .A1(n11675), .A2(n11674), .A3(n11673), .ZN(n11676) );
  AOI21_X1 U13644 ( .B1(n11677), .B2(n13813), .A(n11676), .ZN(n11678) );
  NAND2_X1 U13645 ( .A1(n11679), .A2(n11678), .ZN(P3_U3185) );
  INV_X1 U13646 ( .A(n11680), .ZN(n11682) );
  NAND2_X1 U13647 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  NAND2_X1 U13648 ( .A1(n15058), .A2(n11694), .ZN(n11686) );
  NAND2_X1 U13649 ( .A1(n10314), .A2(n14856), .ZN(n11685) );
  NAND2_X1 U13650 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  XNOR2_X1 U13651 ( .A(n11687), .B(n11130), .ZN(n11690) );
  AOI22_X1 U13652 ( .A1(n15058), .A2(n14817), .B1(n11694), .B2(n10314), .ZN(
        n11688) );
  XNOR2_X1 U13653 ( .A(n11690), .B(n11688), .ZN(n14914) );
  INV_X1 U13654 ( .A(n11688), .ZN(n11689) );
  NAND2_X1 U13655 ( .A1(n11690), .A2(n11689), .ZN(n11699) );
  NAND2_X1 U13656 ( .A1(n15057), .A2(n14817), .ZN(n11692) );
  NAND2_X1 U13657 ( .A1(n11715), .A2(n11694), .ZN(n11691) );
  AND2_X1 U13658 ( .A1(n11692), .A2(n11691), .ZN(n11700) );
  AND2_X1 U13659 ( .A1(n11699), .A2(n11700), .ZN(n11693) );
  INV_X1 U13660 ( .A(n14856), .ZN(n14932) );
  OAI22_X1 U13661 ( .A1(n11697), .A2(n14935), .B1(n11696), .B2(n14932), .ZN(
        n11698) );
  XNOR2_X1 U13662 ( .A(n11698), .B(n11130), .ZN(n11706) );
  NAND2_X1 U13663 ( .A1(n11708), .A2(n11706), .ZN(n11703) );
  NAND2_X1 U13664 ( .A1(n14912), .A2(n11699), .ZN(n11702) );
  INV_X1 U13665 ( .A(n11700), .ZN(n11701) );
  NAND2_X1 U13666 ( .A1(n11702), .A2(n11701), .ZN(n11704) );
  INV_X1 U13667 ( .A(n11735), .ZN(n11709) );
  INV_X1 U13668 ( .A(n11703), .ZN(n11705) );
  NAND2_X1 U13669 ( .A1(n11705), .A2(n11704), .ZN(n11707) );
  AOI22_X1 U13670 ( .A1(n11709), .A2(n11708), .B1(n11707), .B2(n11706), .ZN(
        n11717) );
  NAND2_X1 U13671 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15119) );
  OAI21_X1 U13672 ( .B1(n15036), .B2(n11711), .A(n15119), .ZN(n11714) );
  INV_X1 U13673 ( .A(n15056), .ZN(n11889) );
  OAI22_X1 U13674 ( .A1(n11712), .A2(n15038), .B1(n15037), .B2(n11889), .ZN(
        n11713) );
  AOI211_X1 U13675 ( .C1(n11715), .C2(n15042), .A(n11714), .B(n11713), .ZN(
        n11716) );
  OAI21_X1 U13676 ( .B1(n11717), .B2(n15044), .A(n11716), .ZN(P1_U3230) );
  INV_X1 U13677 ( .A(n11718), .ZN(n11760) );
  INV_X1 U13678 ( .A(n12518), .ZN(n12280) );
  OAI222_X1 U13679 ( .A1(n14780), .A2(n11760), .B1(n12280), .B2(P2_U3088), 
        .C1(n11719), .C2(n14783), .ZN(P2_U3311) );
  INV_X1 U13680 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15090) );
  AOI21_X1 U13681 ( .B1(n15458), .B2(n15090), .A(n14915), .ZN(n11720) );
  MUX2_X1 U13682 ( .A(n10901), .B(n11720), .S(n15430), .Z(n11722) );
  NAND2_X1 U13683 ( .A1(n15459), .A2(n10314), .ZN(n11721) );
  OAI211_X1 U13684 ( .C1(n11723), .C2(n15168), .A(n11722), .B(n11721), .ZN(
        n11724) );
  AOI21_X1 U13685 ( .B1(n11725), .B2(n15425), .A(n11724), .ZN(n11726) );
  OAI21_X1 U13686 ( .B1(n11727), .B2(n15440), .A(n11726), .ZN(P1_U3290) );
  NAND2_X1 U13687 ( .A1(n11890), .A2(n14856), .ZN(n11729) );
  NAND2_X1 U13688 ( .A1(n15056), .A2(n11694), .ZN(n11728) );
  NAND2_X1 U13689 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  XNOR2_X1 U13690 ( .A(n11730), .B(n12183), .ZN(n11732) );
  AOI22_X1 U13691 ( .A1(n11890), .A2(n14831), .B1(n14817), .B2(n15056), .ZN(
        n11731) );
  NOR2_X1 U13692 ( .A1(n11732), .A2(n11731), .ZN(n11829) );
  NAND2_X1 U13693 ( .A1(n11732), .A2(n11731), .ZN(n11828) );
  INV_X1 U13694 ( .A(n11828), .ZN(n11733) );
  NOR2_X1 U13695 ( .A1(n11829), .A2(n11733), .ZN(n11734) );
  XNOR2_X1 U13696 ( .A(n11735), .B(n11734), .ZN(n11742) );
  OAI22_X1 U13697 ( .A1(n15036), .A2(n11737), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11736), .ZN(n11739) );
  NOR2_X1 U13698 ( .A1(n15026), .A2(n11891), .ZN(n11738) );
  AOI211_X1 U13699 ( .C1(n15029), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        n11741) );
  OAI21_X1 U13700 ( .B1(n11742), .B2(n15044), .A(n11741), .ZN(P1_U3227) );
  NAND2_X1 U13701 ( .A1(n15205), .A2(n11937), .ZN(n15398) );
  INV_X1 U13702 ( .A(n15398), .ZN(n15463) );
  OAI21_X1 U13703 ( .B1(n15459), .B2(n15463), .A(n15462), .ZN(n11744) );
  AOI22_X1 U13704 ( .A1(n15356), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15458), .ZN(n11743) );
  OAI211_X1 U13705 ( .C1(n11745), .C2(n12127), .A(n11744), .B(n11743), .ZN(
        n11746) );
  AOI21_X1 U13706 ( .B1(n15430), .B2(n11747), .A(n11746), .ZN(n11748) );
  INV_X1 U13707 ( .A(n11748), .ZN(P1_U3293) );
  OR2_X1 U13708 ( .A1(n11749), .A2(n14305), .ZN(n14561) );
  OAI22_X1 U13709 ( .A1(n16458), .A2(n11751), .B1(n11750), .B2(n16455), .ZN(
        n11754) );
  NOR2_X1 U13710 ( .A1(n14631), .A2(n11752), .ZN(n11753) );
  AOI211_X1 U13711 ( .C1(n11755), .C2(n16452), .A(n11754), .B(n11753), .ZN(
        n11758) );
  INV_X1 U13712 ( .A(n14593), .ZN(n16453) );
  NAND2_X1 U13713 ( .A1(n16453), .A2(n11756), .ZN(n11757) );
  OAI211_X1 U13714 ( .C1(n14598), .C2(n11759), .A(n11758), .B(n11757), .ZN(
        P2_U3261) );
  INV_X1 U13715 ( .A(n12808), .ZN(n13016) );
  OAI222_X1 U13716 ( .A1(n7555), .A2(n11761), .B1(n15627), .B2(n11760), .C1(
        n13016), .C2(P1_U3086), .ZN(P1_U3339) );
  NOR2_X1 U13717 ( .A1(n11762), .A2(n16418), .ZN(n11764) );
  AND2_X1 U13718 ( .A1(n13484), .A2(n16313), .ZN(n11763) );
  AOI21_X1 U13719 ( .B1(n13619), .B2(n11764), .A(n11763), .ZN(n11916) );
  OAI22_X1 U13720 ( .A1(n14164), .A2(n11855), .B1(n16473), .B2(n11496), .ZN(
        n11765) );
  INV_X1 U13721 ( .A(n11765), .ZN(n11766) );
  OAI21_X1 U13722 ( .B1(n11916), .B2(n10822), .A(n11766), .ZN(P3_U3459) );
  MUX2_X1 U13723 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13775), .Z(n11767) );
  INV_X1 U13724 ( .A(n11767), .ZN(n11768) );
  XNOR2_X1 U13725 ( .A(n11767), .B(n11780), .ZN(n13668) );
  INV_X1 U13726 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11770) );
  MUX2_X1 U13727 ( .A(n11770), .B(n11769), .S(n13775), .Z(n11771) );
  NOR2_X1 U13728 ( .A1(n11771), .A2(n11776), .ZN(n11773) );
  AND2_X1 U13729 ( .A1(n11771), .A2(n11776), .ZN(n11945) );
  OAI21_X1 U13730 ( .B1(n11773), .B2(n11945), .A(n11772), .ZN(n11774) );
  OAI21_X1 U13731 ( .B1(n7850), .B2(n11945), .A(n11774), .ZN(n11775) );
  NAND2_X1 U13732 ( .A1(n11775), .A2(n16272), .ZN(n11791) );
  XNOR2_X1 U13733 ( .A(n11780), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n13682) );
  OAI21_X1 U13734 ( .B1(n11778), .B2(P3_REG2_REG_5__SCAN_IN), .A(n11957), .ZN(
        n11789) );
  INV_X1 U13735 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11779) );
  XNOR2_X1 U13736 ( .A(n11780), .B(n11779), .ZN(n13672) );
  NAND2_X1 U13737 ( .A1(n11780), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U13738 ( .A1(n13677), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U13739 ( .A1(n11782), .A2(n8149), .ZN(n11951) );
  OAI21_X1 U13740 ( .B1(n11783), .B2(P3_REG1_REG_5__SCAN_IN), .A(n11953), .ZN(
        n11784) );
  NAND2_X1 U13741 ( .A1(n13847), .A2(n11784), .ZN(n11786) );
  NOR2_X1 U13742 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15902), .ZN(n12337) );
  INV_X1 U13743 ( .A(n12337), .ZN(n11785) );
  OAI211_X1 U13744 ( .C1(n16292), .C2(n11787), .A(n11786), .B(n11785), .ZN(
        n11788) );
  AOI21_X1 U13745 ( .B1(n13840), .B2(n11789), .A(n11788), .ZN(n11790) );
  OAI211_X1 U13746 ( .C1(n16278), .C2(n8149), .A(n11791), .B(n11790), .ZN(
        P3_U3187) );
  NAND2_X1 U13747 ( .A1(n11792), .A2(n11793), .ZN(n11797) );
  XNOR2_X1 U13748 ( .A(n11799), .B(n13484), .ZN(n13196) );
  NAND2_X1 U13749 ( .A1(n13265), .A2(n11855), .ZN(n11798) );
  NAND2_X1 U13750 ( .A1(n11799), .A2(n12154), .ZN(n11800) );
  NAND2_X1 U13751 ( .A1(n13195), .A2(n11800), .ZN(n12137) );
  XNOR2_X1 U13752 ( .A(n13265), .B(n11801), .ZN(n12138) );
  XNOR2_X1 U13753 ( .A(n12138), .B(n8598), .ZN(n12136) );
  XOR2_X1 U13754 ( .A(n12137), .B(n12136), .Z(n11810) );
  INV_X1 U13755 ( .A(n13442), .ZN(n13421) );
  NOR2_X1 U13756 ( .A1(n11803), .A2(n11802), .ZN(n11805) );
  AOI22_X1 U13757 ( .A1(n13450), .A2(n13484), .B1(n13665), .B2(n13439), .ZN(
        n11806) );
  OAI21_X1 U13758 ( .B1(n16342), .B2(n13453), .A(n11806), .ZN(n11807) );
  AOI21_X1 U13759 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n11808), .A(n11807), .ZN(
        n11809) );
  OAI21_X1 U13760 ( .B1(n11810), .B2(n13421), .A(n11809), .ZN(P3_U3177) );
  OAI21_X1 U13761 ( .B1(n11815), .B2(P1_REG1_REG_12__SCAN_IN), .A(n11811), 
        .ZN(n11813) );
  INV_X1 U13762 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n12825) );
  MUX2_X1 U13763 ( .A(n12825), .B(P1_REG1_REG_13__SCAN_IN), .S(n12393), .Z(
        n11812) );
  AOI211_X1 U13764 ( .C1(n11813), .C2(n11812), .A(n12627), .B(n12392), .ZN(
        n11821) );
  OAI21_X1 U13765 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n11815), .A(n11814), 
        .ZN(n11817) );
  INV_X1 U13766 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n12384) );
  MUX2_X1 U13767 ( .A(n12384), .B(P1_REG2_REG_13__SCAN_IN), .S(n12393), .Z(
        n11816) );
  NOR2_X1 U13768 ( .A1(n11817), .A2(n11816), .ZN(n12391) );
  AOI211_X1 U13769 ( .C1(n11817), .C2(n11816), .A(n15150), .B(n12391), .ZN(
        n11820) );
  NAND2_X1 U13770 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12963)
         );
  NAND2_X1 U13771 ( .A1(n16197), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11818) );
  OAI211_X1 U13772 ( .C1(n15149), .C2(n12385), .A(n12963), .B(n11818), .ZN(
        n11819) );
  OR3_X1 U13773 ( .A1(n11821), .A2(n11820), .A3(n11819), .ZN(P1_U3256) );
  INV_X1 U13774 ( .A(n11822), .ZN(n11824) );
  OAI222_X1 U13775 ( .A1(n7555), .A2(n11823), .B1(n15627), .B2(n11824), .C1(
        P1_U3086), .C2(n15130), .ZN(P1_U3338) );
  INV_X1 U13776 ( .A(n12832), .ZN(n12522) );
  OAI222_X1 U13777 ( .A1(n14783), .A2(n11825), .B1(n14780), .B2(n11824), .C1(
        P2_U3088), .C2(n12522), .ZN(P2_U3310) );
  INV_X1 U13778 ( .A(n11826), .ZN(n11827) );
  OAI222_X1 U13779 ( .A1(n11794), .A2(P3_U3151), .B1(n13194), .B2(n11827), 
        .C1(n15839), .C2(n14237), .ZN(P3_U3275) );
  OAI21_X2 U13780 ( .B1(n11830), .B2(n11829), .A(n11828), .ZN(n11967) );
  NAND2_X1 U13781 ( .A1(n12029), .A2(n11013), .ZN(n11832) );
  NAND2_X1 U13782 ( .A1(n15055), .A2(n11694), .ZN(n11831) );
  NAND2_X1 U13783 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  XNOR2_X1 U13784 ( .A(n11833), .B(n12183), .ZN(n11964) );
  AND2_X1 U13785 ( .A1(n15055), .A2(n12699), .ZN(n11834) );
  AOI21_X1 U13786 ( .B1(n12029), .B2(n11694), .A(n11834), .ZN(n11965) );
  XNOR2_X1 U13787 ( .A(n11964), .B(n11965), .ZN(n11966) );
  XNOR2_X1 U13788 ( .A(n11967), .B(n11966), .ZN(n11839) );
  OAI21_X1 U13789 ( .B1(n15036), .B2(n11940), .A(n11835), .ZN(n11837) );
  OAI22_X1 U13790 ( .A1(n11889), .A2(n15038), .B1(n15037), .B2(n12195), .ZN(
        n11836) );
  AOI211_X1 U13791 ( .C1(n12029), .C2(n15042), .A(n11837), .B(n11836), .ZN(
        n11838) );
  OAI21_X1 U13792 ( .B1(n11839), .B2(n15044), .A(n11838), .ZN(P1_U3239) );
  INV_X1 U13793 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11851) );
  OAI21_X1 U13794 ( .B1(n7548), .B2(n11842), .A(n11840), .ZN(n11987) );
  INV_X1 U13795 ( .A(n11987), .ZN(n11849) );
  OAI22_X1 U13796 ( .A1(n12060), .A2(n14623), .B1(n11841), .B2(n14621), .ZN(
        n11846) );
  AOI21_X1 U13797 ( .B1(n11844), .B2(n11843), .A(n14619), .ZN(n11845) );
  AOI211_X1 U13798 ( .C1(n14522), .C2(n11987), .A(n11846), .B(n11845), .ZN(
        n11989) );
  AOI21_X1 U13799 ( .B1(n11979), .B2(n11847), .A(n12018), .ZN(n11982) );
  AOI22_X1 U13800 ( .A1(n11982), .A2(n14734), .B1(n14733), .B2(n11979), .ZN(
        n11848) );
  OAI211_X1 U13801 ( .C1(n11849), .C2(n16299), .A(n11989), .B(n11848), .ZN(
        n11852) );
  NAND2_X1 U13802 ( .A1(n11852), .A2(n16413), .ZN(n11850) );
  OAI21_X1 U13803 ( .B1(n16413), .B2(n11851), .A(n11850), .ZN(P2_U3505) );
  NAND2_X1 U13804 ( .A1(n11852), .A2(n14760), .ZN(n11853) );
  OAI21_X1 U13805 ( .B1(n14760), .B2(n9463), .A(n11853), .ZN(P2_U3448) );
  INV_X1 U13806 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11854) );
  OAI22_X1 U13807 ( .A1(n14221), .A2(n11855), .B1(n16476), .B2(n11854), .ZN(
        n11856) );
  INV_X1 U13808 ( .A(n11856), .ZN(n11857) );
  OAI21_X1 U13809 ( .B1(n11916), .B2(n16483), .A(n11857), .ZN(P3_U3390) );
  INV_X1 U13810 ( .A(n11858), .ZN(n11860) );
  AND2_X1 U13811 ( .A1(n14405), .A2(n14305), .ZN(n11864) );
  XNOR2_X1 U13812 ( .A(n12021), .B(n14306), .ZN(n11863) );
  NOR2_X1 U13813 ( .A1(n11863), .A2(n11864), .ZN(n12053) );
  AOI21_X1 U13814 ( .B1(n11864), .B2(n11863), .A(n12053), .ZN(n11865) );
  NAND2_X1 U13815 ( .A1(n11866), .A2(n11865), .ZN(n12055) );
  OAI21_X1 U13816 ( .B1(n11866), .B2(n11865), .A(n12055), .ZN(n11867) );
  NAND2_X1 U13817 ( .A1(n11867), .A2(n14382), .ZN(n11873) );
  INV_X1 U13818 ( .A(n13166), .ZN(n11871) );
  NAND2_X1 U13819 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n16120) );
  INV_X1 U13820 ( .A(n16120), .ZN(n11870) );
  INV_X1 U13821 ( .A(n14404), .ZN(n12225) );
  OAI22_X1 U13822 ( .A1(n12225), .A2(n14387), .B1(n14362), .B2(n11868), .ZN(
        n11869) );
  AOI211_X1 U13823 ( .C1(n11871), .C2(n14385), .A(n11870), .B(n11869), .ZN(
        n11872) );
  OAI211_X1 U13824 ( .C1(n13167), .C2(n14393), .A(n11873), .B(n11872), .ZN(
        P2_U3185) );
  XNOR2_X1 U13825 ( .A(n11874), .B(n11878), .ZN(n11875) );
  NAND2_X1 U13826 ( .A1(n11875), .A2(n14603), .ZN(n11877) );
  AOI22_X1 U13827 ( .A1(n14600), .A2(n14405), .B1(n14403), .B2(n14604), .ZN(
        n11876) );
  NAND2_X1 U13828 ( .A1(n11877), .A2(n11876), .ZN(n16371) );
  INV_X1 U13829 ( .A(n16371), .ZN(n11885) );
  XNOR2_X1 U13830 ( .A(n11879), .B(n11878), .ZN(n16373) );
  INV_X1 U13831 ( .A(n14596), .ZN(n12355) );
  OAI211_X1 U13832 ( .C1(n12020), .C2(n16370), .A(n14734), .B(n12108), .ZN(
        n16369) );
  OAI22_X1 U13833 ( .A1(n16458), .A2(n11880), .B1(n12059), .B2(n16455), .ZN(
        n11881) );
  AOI21_X1 U13834 ( .B1(n16463), .B2(n12050), .A(n11881), .ZN(n11882) );
  OAI21_X1 U13835 ( .B1(n12355), .B2(n16369), .A(n11882), .ZN(n11883) );
  AOI21_X1 U13836 ( .B1(n16373), .B2(n14617), .A(n11883), .ZN(n11884) );
  OAI21_X1 U13837 ( .B1(n11885), .B2(n14598), .A(n11884), .ZN(P2_U3257) );
  INV_X1 U13838 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11906) );
  OR2_X1 U13839 ( .A1(n15056), .A2(n11890), .ZN(n11886) );
  XNOR2_X1 U13840 ( .A(n12027), .B(n7867), .ZN(n11897) );
  INV_X1 U13841 ( .A(n11897), .ZN(n11944) );
  AND2_X1 U13842 ( .A1(n11890), .A2(n11889), .ZN(n11893) );
  NAND2_X1 U13843 ( .A1(n11891), .A2(n15056), .ZN(n11892) );
  INV_X1 U13844 ( .A(n12033), .ZN(n11895) );
  AOI21_X1 U13845 ( .B1(n7867), .B2(n11896), .A(n11895), .ZN(n11900) );
  AOI22_X1 U13846 ( .A1(n15386), .A2(n15056), .B1(n15054), .B2(n15448), .ZN(
        n11899) );
  NAND2_X1 U13847 ( .A1(n11897), .A2(n15445), .ZN(n11898) );
  OAI211_X1 U13848 ( .C1(n11900), .C2(n15567), .A(n11899), .B(n11898), .ZN(
        n11935) );
  INV_X1 U13849 ( .A(n11935), .ZN(n11904) );
  AND2_X1 U13850 ( .A1(n11901), .A2(n12029), .ZN(n11902) );
  NOR2_X1 U13851 ( .A1(n12039), .A2(n11902), .ZN(n11936) );
  AOI22_X1 U13852 ( .A1(n11936), .A2(n16326), .B1(n15563), .B2(n12029), .ZN(
        n11903) );
  OAI211_X1 U13853 ( .C1(n16353), .C2(n11944), .A(n11904), .B(n11903), .ZN(
        n15588) );
  NAND2_X1 U13854 ( .A1(n15588), .A2(n16338), .ZN(n11905) );
  OAI21_X1 U13855 ( .B1(n16338), .B2(n11906), .A(n11905), .ZN(P1_U3477) );
  AND2_X1 U13856 ( .A1(n11907), .A2(n11912), .ZN(n11908) );
  NOR2_X1 U13857 ( .A1(n11909), .A2(n11908), .ZN(n11911) );
  MUX2_X1 U13858 ( .A(n11916), .B(n11915), .S(n16348), .Z(n11921) );
  INV_X1 U13859 ( .A(n11917), .ZN(n11918) );
  NOR2_X1 U13860 ( .A1(n16467), .A2(n12431), .ZN(n16319) );
  AOI22_X1 U13861 ( .A1(n16384), .A2(n11919), .B1(n16382), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U13862 ( .A1(n11921), .A2(n11920), .ZN(P3_U3233) );
  INV_X1 U13863 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11929) );
  INV_X1 U13864 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U13865 ( .A1(n10810), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U13866 ( .A1(n8611), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11922) );
  OAI211_X1 U13867 ( .C1(n8800), .C2(n11924), .A(n11923), .B(n11922), .ZN(
        n11925) );
  INV_X1 U13868 ( .A(n11925), .ZN(n11926) );
  NAND2_X1 U13869 ( .A1(n11927), .A2(n11926), .ZN(n13612) );
  NAND2_X1 U13870 ( .A1(n13612), .A2(P3_U3897), .ZN(n11928) );
  OAI21_X1 U13871 ( .B1(P3_U3897), .B2(n11929), .A(n11928), .ZN(P3_U3522) );
  AOI21_X1 U13872 ( .B1(n14619), .B2(n14586), .A(n16300), .ZN(n11930) );
  AOI21_X1 U13873 ( .B1(n14583), .B2(n14411), .A(n11930), .ZN(n16296) );
  OAI22_X1 U13874 ( .A1(n16296), .A2(n14598), .B1(n11931), .B2(n16455), .ZN(
        n11932) );
  AOI21_X1 U13875 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14598), .A(n11932), .ZN(
        n11934) );
  OAI21_X1 U13876 ( .B1(n16463), .B2(n16452), .A(n7635), .ZN(n11933) );
  OAI211_X1 U13877 ( .C1(n16300), .C2(n14593), .A(n11934), .B(n11933), .ZN(
        P2_U3265) );
  AOI21_X1 U13878 ( .B1(n11937), .B2(n11936), .A(n11935), .ZN(n11938) );
  MUX2_X1 U13879 ( .A(n11939), .B(n11938), .S(n15430), .Z(n11943) );
  INV_X1 U13880 ( .A(n11940), .ZN(n11941) );
  AOI22_X1 U13881 ( .A1(n15459), .A2(n12029), .B1(n11941), .B2(n15458), .ZN(
        n11942) );
  OAI211_X1 U13882 ( .C1(n11944), .C2(n12127), .A(n11943), .B(n11942), .ZN(
        P1_U3287) );
  MUX2_X1 U13883 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13775), .Z(n12231) );
  XNOR2_X1 U13884 ( .A(n12231), .B(n12245), .ZN(n11946) );
  AOI21_X1 U13885 ( .B1(n11947), .B2(n11946), .A(n12232), .ZN(n11963) );
  INV_X1 U13886 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11948) );
  NOR2_X1 U13887 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11948), .ZN(n12640) );
  XNOR2_X1 U13888 ( .A(n12245), .B(n12445), .ZN(n11950) );
  NAND2_X1 U13889 ( .A1(n11949), .A2(n11950), .ZN(n12236) );
  INV_X1 U13890 ( .A(n11950), .ZN(n11952) );
  NAND3_X1 U13891 ( .A1(n11953), .A2(n11952), .A3(n11951), .ZN(n11954) );
  AOI21_X1 U13892 ( .B1(n12236), .B2(n11954), .A(n16285), .ZN(n11955) );
  AOI211_X1 U13893 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n16037), .A(n12640), .B(
        n11955), .ZN(n11960) );
  XNOR2_X1 U13894 ( .A(n12245), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11956) );
  AND3_X1 U13895 ( .A1(n11957), .A2(n11956), .A3(n7456), .ZN(n11958) );
  OAI21_X1 U13896 ( .B1(n12244), .B2(n11958), .A(n13840), .ZN(n11959) );
  OAI211_X1 U13897 ( .C1(n16278), .C2(n12245), .A(n11960), .B(n11959), .ZN(
        n11961) );
  INV_X1 U13898 ( .A(n11961), .ZN(n11962) );
  OAI21_X1 U13899 ( .B1(n11963), .B2(n16259), .A(n11962), .ZN(P3_U3188) );
  NAND2_X1 U13900 ( .A1(n16350), .A2(n14856), .ZN(n11970) );
  NAND2_X1 U13901 ( .A1(n15054), .A2(n14831), .ZN(n11969) );
  NAND2_X1 U13902 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  XNOR2_X1 U13903 ( .A(n11971), .B(n11130), .ZN(n12186) );
  AND2_X1 U13904 ( .A1(n15054), .A2(n14817), .ZN(n11972) );
  AOI21_X1 U13905 ( .B1(n16350), .B2(n14831), .A(n11972), .ZN(n12185) );
  XNOR2_X1 U13906 ( .A(n12186), .B(n12185), .ZN(n12188) );
  XNOR2_X1 U13907 ( .A(n12189), .B(n12188), .ZN(n11978) );
  INV_X1 U13908 ( .A(n12042), .ZN(n11975) );
  INV_X1 U13909 ( .A(n15055), .ZN(n12028) );
  OAI22_X1 U13910 ( .A1(n12028), .A2(n15038), .B1(n15037), .B2(n12508), .ZN(
        n11973) );
  AOI211_X1 U13911 ( .C1(n15017), .C2(n11975), .A(n11974), .B(n11973), .ZN(
        n11977) );
  NAND2_X1 U13912 ( .A1(n16350), .A2(n15042), .ZN(n11976) );
  OAI211_X1 U13913 ( .C1(n11978), .C2(n15044), .A(n11977), .B(n11976), .ZN(
        P1_U3213) );
  INV_X1 U13914 ( .A(n11979), .ZN(n11985) );
  INV_X1 U13915 ( .A(n11980), .ZN(n11981) );
  AOI22_X1 U13916 ( .A1(n14598), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n11981), 
        .B2(n14611), .ZN(n11984) );
  NAND2_X1 U13917 ( .A1(n11982), .A2(n16452), .ZN(n11983) );
  OAI211_X1 U13918 ( .C1(n11985), .C2(n14631), .A(n11984), .B(n11983), .ZN(
        n11986) );
  AOI21_X1 U13919 ( .B1(n11987), .B2(n16453), .A(n11986), .ZN(n11988) );
  OAI21_X1 U13920 ( .B1(n11989), .B2(n14598), .A(n11988), .ZN(P2_U3259) );
  INV_X1 U13921 ( .A(n11990), .ZN(n11997) );
  AOI22_X1 U13922 ( .A1(n14598), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n14611), 
        .B2(n11991), .ZN(n11994) );
  NAND2_X1 U13923 ( .A1(n14596), .A2(n11992), .ZN(n11993) );
  OAI211_X1 U13924 ( .C1(n11995), .C2(n14631), .A(n11994), .B(n11993), .ZN(
        n11996) );
  AOI21_X1 U13925 ( .B1(n11997), .B2(n14617), .A(n11996), .ZN(n11998) );
  OAI21_X1 U13926 ( .B1(n14598), .B2(n11999), .A(n11998), .ZN(P2_U3262) );
  AOI22_X1 U13927 ( .A1(n14598), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14611), .ZN(n12002) );
  NAND2_X1 U13928 ( .A1(n16463), .A2(n12000), .ZN(n12001) );
  OAI211_X1 U13929 ( .C1(n12355), .C2(n12003), .A(n12002), .B(n12001), .ZN(
        n12004) );
  AOI21_X1 U13930 ( .B1(n12005), .B2(n14617), .A(n12004), .ZN(n12006) );
  OAI21_X1 U13931 ( .B1(n14598), .B2(n12007), .A(n12006), .ZN(P2_U3264) );
  INV_X1 U13932 ( .A(n12008), .ZN(n12009) );
  OAI222_X1 U13933 ( .A1(P3_U3151), .A2(n13487), .B1(n14237), .B2(n12010), 
        .C1(n13194), .C2(n12009), .ZN(P3_U3274) );
  OAI21_X1 U13934 ( .B1(n12012), .B2(n12013), .A(n12011), .ZN(n13171) );
  XNOR2_X1 U13935 ( .A(n12014), .B(n12013), .ZN(n12017) );
  OR2_X1 U13936 ( .A1(n13171), .A2(n14586), .ZN(n12016) );
  AOI22_X1 U13937 ( .A1(n14604), .A2(n14404), .B1(n14406), .B2(n14600), .ZN(
        n12015) );
  OAI211_X1 U13938 ( .C1(n14619), .C2(n12017), .A(n12016), .B(n12015), .ZN(
        n13164) );
  INV_X1 U13939 ( .A(n13164), .ZN(n12024) );
  NOR2_X1 U13940 ( .A1(n12018), .A2(n13167), .ZN(n12019) );
  OR2_X1 U13941 ( .A1(n12020), .A2(n12019), .ZN(n13165) );
  INV_X1 U13942 ( .A(n13165), .ZN(n12022) );
  AOI22_X1 U13943 ( .A1(n12022), .A2(n14734), .B1(n14733), .B2(n12021), .ZN(
        n12023) );
  OAI211_X1 U13944 ( .C1(n16299), .C2(n13171), .A(n12024), .B(n12023), .ZN(
        n12047) );
  NAND2_X1 U13945 ( .A1(n12047), .A2(n16413), .ZN(n12025) );
  OAI21_X1 U13946 ( .B1(n16413), .B2(n9478), .A(n12025), .ZN(P2_U3506) );
  INV_X1 U13947 ( .A(n12029), .ZN(n12026) );
  XNOR2_X1 U13948 ( .A(n12085), .B(n12084), .ZN(n12038) );
  INV_X1 U13949 ( .A(n12038), .ZN(n16354) );
  OAI22_X1 U13950 ( .A1(n12028), .A2(n15451), .B1(n12508), .B2(n15410), .ZN(
        n12037) );
  NAND2_X1 U13951 ( .A1(n12029), .A2(n12028), .ZN(n12032) );
  AND2_X1 U13952 ( .A1(n12031), .A2(n12032), .ZN(n12030) );
  INV_X1 U13953 ( .A(n12091), .ZN(n12035) );
  AOI21_X1 U13954 ( .B1(n12033), .B2(n12032), .A(n12031), .ZN(n12034) );
  NOR3_X1 U13955 ( .A1(n12035), .A2(n12034), .A3(n15567), .ZN(n12036) );
  AOI211_X1 U13956 ( .C1(n15445), .C2(n12038), .A(n12037), .B(n12036), .ZN(
        n16352) );
  MUX2_X1 U13957 ( .A(n10956), .B(n16352), .S(n15430), .Z(n12046) );
  INV_X1 U13958 ( .A(n12039), .ZN(n12041) );
  INV_X1 U13959 ( .A(n16350), .ZN(n12043) );
  NAND2_X1 U13960 ( .A1(n12039), .A2(n12043), .ZN(n12128) );
  INV_X1 U13961 ( .A(n12128), .ZN(n12040) );
  AOI211_X1 U13962 ( .C1(n16350), .C2(n12041), .A(n16428), .B(n12040), .ZN(
        n16349) );
  OAI22_X1 U13963 ( .A1(n12043), .A2(n15434), .B1(n15428), .B2(n12042), .ZN(
        n12044) );
  AOI21_X1 U13964 ( .B1(n16349), .B2(n15437), .A(n12044), .ZN(n12045) );
  OAI211_X1 U13965 ( .C1(n16354), .C2(n12127), .A(n12046), .B(n12045), .ZN(
        P1_U3286) );
  INV_X1 U13966 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U13967 ( .A1(n12047), .A2(n14760), .ZN(n12048) );
  OAI21_X1 U13968 ( .B1(n14760), .B2(n12049), .A(n12048), .ZN(P2_U3451) );
  AND2_X1 U13969 ( .A1(n14404), .A2(n14305), .ZN(n12052) );
  XNOR2_X1 U13970 ( .A(n12050), .B(n14306), .ZN(n12051) );
  NOR2_X1 U13971 ( .A1(n12051), .A2(n12052), .ZN(n12218) );
  AOI21_X1 U13972 ( .B1(n12052), .B2(n12051), .A(n12218), .ZN(n12057) );
  INV_X1 U13973 ( .A(n12053), .ZN(n12054) );
  OAI21_X1 U13974 ( .B1(n12057), .B2(n12056), .A(n12220), .ZN(n12058) );
  NAND2_X1 U13975 ( .A1(n12058), .A2(n14382), .ZN(n12065) );
  INV_X1 U13976 ( .A(n12059), .ZN(n12063) );
  NAND2_X1 U13977 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n16133) );
  INV_X1 U13978 ( .A(n16133), .ZN(n12062) );
  OAI22_X1 U13979 ( .A1(n12060), .A2(n14362), .B1(n14387), .B2(n12408), .ZN(
        n12061) );
  AOI211_X1 U13980 ( .C1(n12063), .C2(n14385), .A(n12062), .B(n12061), .ZN(
        n12064) );
  OAI211_X1 U13981 ( .C1(n16370), .C2(n14393), .A(n12065), .B(n12064), .ZN(
        P2_U3193) );
  AOI21_X1 U13982 ( .B1(n12067), .B2(P2_REG1_REG_13__SCAN_IN), .A(n12066), 
        .ZN(n16155) );
  MUX2_X1 U13983 ( .A(n12068), .B(P2_REG1_REG_14__SCAN_IN), .S(n16158), .Z(
        n16154) );
  NOR2_X1 U13984 ( .A1(n16155), .A2(n16154), .ZN(n16153) );
  AOI21_X1 U13985 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n16158), .A(n16153), 
        .ZN(n12274) );
  XNOR2_X1 U13986 ( .A(n12274), .B(n12273), .ZN(n12069) );
  NOR2_X1 U13987 ( .A1(n9619), .A2(n12069), .ZN(n12275) );
  AOI211_X1 U13988 ( .C1(n12069), .C2(n9619), .A(n12275), .B(n16177), .ZN(
        n12078) );
  OAI21_X1 U13989 ( .B1(n12072), .B2(n12071), .A(n12070), .ZN(n16150) );
  INV_X1 U13990 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12073) );
  MUX2_X1 U13991 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n12073), .S(n16158), .Z(
        n16149) );
  AOI21_X1 U13992 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n16158), .A(n16151), 
        .ZN(n12268) );
  XNOR2_X1 U13993 ( .A(n12268), .B(n12273), .ZN(n12074) );
  NOR2_X1 U13994 ( .A1(n9620), .A2(n12074), .ZN(n12269) );
  AOI211_X1 U13995 ( .C1(n12074), .C2(n9620), .A(n12269), .B(n16182), .ZN(
        n12077) );
  AND2_X1 U13996 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13066) );
  AOI21_X1 U13997 ( .B1(n16055), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n13066), 
        .ZN(n12075) );
  OAI21_X1 U13998 ( .B1(n12273), .B2(n16168), .A(n12075), .ZN(n12076) );
  OR3_X1 U13999 ( .A1(n12078), .A2(n12077), .A3(n12076), .ZN(P2_U3229) );
  NOR2_X1 U14000 ( .A1(n14237), .A2(SI_22_), .ZN(n12079) );
  AOI21_X1 U14001 ( .B1(n12080), .B2(P3_STATE_REG_SCAN_IN), .A(n12079), .ZN(
        n12081) );
  OAI21_X1 U14002 ( .B1(n12082), .B2(n13194), .A(n12081), .ZN(n12083) );
  INV_X1 U14003 ( .A(n12083), .ZN(P3_U3273) );
  OR2_X1 U14004 ( .A1(n16350), .A2(n15054), .ZN(n12086) );
  NAND2_X1 U14005 ( .A1(n12088), .A2(n12119), .ZN(n12089) );
  INV_X1 U14006 ( .A(n16363), .ZN(n12100) );
  NAND2_X1 U14007 ( .A1(n12091), .A2(n12090), .ZN(n12120) );
  XNOR2_X1 U14008 ( .A(n12120), .B(n12119), .ZN(n12093) );
  AOI22_X1 U14009 ( .A1(n15386), .A2(n15054), .B1(n15052), .B2(n15448), .ZN(
        n12092) );
  OAI21_X1 U14010 ( .B1(n12093), .B2(n15567), .A(n12092), .ZN(n12094) );
  AOI21_X1 U14011 ( .B1(n16363), .B2(n15445), .A(n12094), .ZN(n16365) );
  MUX2_X1 U14012 ( .A(n12095), .B(n16365), .S(n15430), .Z(n12099) );
  INV_X1 U14013 ( .A(n16359), .ZN(n12201) );
  XNOR2_X1 U14014 ( .A(n12128), .B(n12201), .ZN(n12096) );
  AND2_X1 U14015 ( .A1(n12096), .A2(n16326), .ZN(n16361) );
  OAI22_X1 U14016 ( .A1(n12201), .A2(n15434), .B1(n12193), .B2(n15428), .ZN(
        n12097) );
  AOI21_X1 U14017 ( .B1(n16361), .B2(n15437), .A(n12097), .ZN(n12098) );
  OAI211_X1 U14018 ( .C1(n12100), .C2(n12127), .A(n12099), .B(n12098), .ZN(
        P1_U3285) );
  XNOR2_X1 U14019 ( .A(n12101), .B(n12102), .ZN(n12106) );
  XNOR2_X1 U14020 ( .A(n12103), .B(n12102), .ZN(n12263) );
  AOI22_X1 U14021 ( .A1(n14600), .A2(n14404), .B1(n14402), .B2(n14604), .ZN(
        n12104) );
  OAI21_X1 U14022 ( .B1(n12263), .B2(n14586), .A(n12104), .ZN(n12105) );
  AOI21_X1 U14023 ( .B1(n12106), .B2(n14603), .A(n12105), .ZN(n12262) );
  INV_X1 U14024 ( .A(n12107), .ZN(n12351) );
  AOI21_X1 U14025 ( .B1(n12259), .B2(n12108), .A(n12351), .ZN(n12260) );
  INV_X1 U14026 ( .A(n12109), .ZN(n12228) );
  AOI22_X1 U14027 ( .A1(n14598), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n12228), 
        .B2(n14611), .ZN(n12110) );
  OAI21_X1 U14028 ( .B1(n7598), .B2(n14631), .A(n12110), .ZN(n12112) );
  NOR2_X1 U14029 ( .A1(n12263), .A2(n14593), .ZN(n12111) );
  AOI211_X1 U14030 ( .C1(n12260), .C2(n16452), .A(n12112), .B(n12111), .ZN(
        n12113) );
  OAI21_X1 U14031 ( .B1(n14598), .B2(n12262), .A(n12113), .ZN(P2_U3256) );
  NAND2_X1 U14032 ( .A1(n16359), .A2(n15053), .ZN(n12114) );
  NAND2_X1 U14033 ( .A1(n12117), .A2(n12123), .ZN(n12118) );
  NAND2_X1 U14034 ( .A1(n12285), .A2(n12118), .ZN(n16394) );
  NAND2_X1 U14035 ( .A1(n12120), .A2(n12119), .ZN(n12122) );
  OR2_X1 U14036 ( .A1(n16359), .A2(n12508), .ZN(n12121) );
  NAND2_X1 U14037 ( .A1(n12122), .A2(n12121), .ZN(n12291) );
  XNOR2_X1 U14038 ( .A(n12291), .B(n12123), .ZN(n12125) );
  AOI22_X1 U14039 ( .A1(n15386), .A2(n15053), .B1(n15051), .B2(n15448), .ZN(
        n12124) );
  OAI21_X1 U14040 ( .B1(n12125), .B2(n15567), .A(n12124), .ZN(n12126) );
  AOI21_X1 U14041 ( .B1(n16394), .B2(n15445), .A(n12126), .ZN(n16396) );
  OR2_X1 U14042 ( .A1(n12128), .A2(n16359), .ZN(n12129) );
  AND2_X1 U14043 ( .A1(n12129), .A2(n12496), .ZN(n12130) );
  OR2_X1 U14044 ( .A1(n12130), .A2(n12286), .ZN(n16392) );
  OAI22_X1 U14045 ( .A1(n15430), .A2(n12131), .B1(n12507), .B2(n15428), .ZN(
        n12132) );
  AOI21_X1 U14046 ( .B1(n12496), .B2(n15459), .A(n12132), .ZN(n12133) );
  OAI21_X1 U14047 ( .B1(n16392), .B2(n15398), .A(n12133), .ZN(n12134) );
  AOI21_X1 U14048 ( .B1(n16394), .B2(n15460), .A(n12134), .ZN(n12135) );
  OAI21_X1 U14049 ( .B1(n16396), .B2(n15356), .A(n12135), .ZN(P1_U3284) );
  XNOR2_X1 U14050 ( .A(n7663), .B(n12432), .ZN(n12202) );
  XNOR2_X1 U14051 ( .A(n12202), .B(n13665), .ZN(n12145) );
  NAND2_X1 U14052 ( .A1(n12137), .A2(n12136), .ZN(n12140) );
  NAND2_X1 U14053 ( .A1(n12138), .A2(n13200), .ZN(n12139) );
  INV_X1 U14054 ( .A(n12144), .ZN(n12142) );
  INV_X1 U14055 ( .A(n12204), .ZN(n12143) );
  AOI211_X1 U14056 ( .C1(n12145), .C2(n12144), .A(n13421), .B(n12143), .ZN(
        n12151) );
  AOI22_X1 U14057 ( .A1(n13418), .A2(n12146), .B1(n8598), .B2(n13450), .ZN(
        n12149) );
  AOI21_X1 U14058 ( .B1(n13664), .B2(n13439), .A(n12147), .ZN(n12148) );
  OAI211_X1 U14059 ( .C1(n13447), .C2(P3_REG3_REG_3__SCAN_IN), .A(n12149), .B(
        n12148), .ZN(n12150) );
  OR2_X1 U14060 ( .A1(n12151), .A2(n12150), .ZN(P3_U3158) );
  XNOR2_X1 U14061 ( .A(n12152), .B(n13489), .ZN(n12157) );
  OAI21_X1 U14062 ( .B1(n12153), .B2(n13489), .A(n13494), .ZN(n16345) );
  OAI22_X1 U14063 ( .A1(n12154), .A2(n14092), .B1(n12210), .B2(n14090), .ZN(
        n12155) );
  AOI21_X1 U14064 ( .B1(n16345), .B2(n12302), .A(n12155), .ZN(n12156) );
  OAI21_X1 U14065 ( .B1(n14005), .B2(n12157), .A(n12156), .ZN(n16343) );
  INV_X1 U14066 ( .A(n16343), .ZN(n12163) );
  INV_X1 U14067 ( .A(n14223), .ZN(n12937) );
  INV_X1 U14068 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n12158) );
  OAI22_X1 U14069 ( .A1(n14221), .A2(n16342), .B1(n16476), .B2(n12158), .ZN(
        n12159) );
  AOI21_X1 U14070 ( .B1(n16345), .B2(n12937), .A(n12159), .ZN(n12160) );
  OAI21_X1 U14071 ( .B1(n12163), .B2(n16483), .A(n12160), .ZN(P3_U3396) );
  INV_X1 U14072 ( .A(n14165), .ZN(n12933) );
  OAI22_X1 U14073 ( .A1(n14164), .A2(n16342), .B1(n16473), .B2(n11663), .ZN(
        n12161) );
  AOI21_X1 U14074 ( .B1(n16345), .B2(n12933), .A(n12161), .ZN(n12162) );
  OAI21_X1 U14075 ( .B1(n12163), .B2(n10822), .A(n12162), .ZN(P3_U3461) );
  INV_X1 U14076 ( .A(n12164), .ZN(n12182) );
  AOI22_X1 U14077 ( .A1(n15145), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15625), .ZN(n12165) );
  OAI21_X1 U14078 ( .B1(n12182), .B2(n15627), .A(n12165), .ZN(P1_U3337) );
  OR2_X1 U14079 ( .A1(n12166), .A2(n13628), .ZN(n12167) );
  NAND2_X1 U14080 ( .A1(n12168), .A2(n12167), .ZN(n12436) );
  NAND2_X1 U14081 ( .A1(n12436), .A2(n12302), .ZN(n12174) );
  OR2_X1 U14082 ( .A1(n12169), .A2(n13628), .ZN(n12304) );
  NAND2_X1 U14083 ( .A1(n12169), .A2(n13628), .ZN(n12170) );
  NAND3_X1 U14084 ( .A1(n12304), .A2(n16309), .A3(n12170), .ZN(n12172) );
  AOI22_X1 U14085 ( .A1(n16311), .A2(n8598), .B1(n13664), .B2(n16313), .ZN(
        n12171) );
  AND2_X1 U14086 ( .A1(n12172), .A2(n12171), .ZN(n12173) );
  NAND2_X1 U14087 ( .A1(n12174), .A2(n12173), .ZN(n12433) );
  INV_X1 U14088 ( .A(n12433), .ZN(n12180) );
  INV_X1 U14089 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n12175) );
  OAI22_X1 U14090 ( .A1(n14221), .A2(n12432), .B1(n16476), .B2(n12175), .ZN(
        n12176) );
  AOI21_X1 U14091 ( .B1(n12436), .B2(n12937), .A(n12176), .ZN(n12177) );
  OAI21_X1 U14092 ( .B1(n12180), .B2(n16483), .A(n12177), .ZN(P3_U3399) );
  OAI22_X1 U14093 ( .A1(n14164), .A2(n12432), .B1(n16473), .B2(n11648), .ZN(
        n12178) );
  AOI21_X1 U14094 ( .B1(n12436), .B2(n12933), .A(n12178), .ZN(n12179) );
  OAI21_X1 U14095 ( .B1(n12180), .B2(n10822), .A(n12179), .ZN(P3_U3462) );
  INV_X1 U14096 ( .A(n12827), .ZN(n16167) );
  OAI222_X1 U14097 ( .A1(n14780), .A2(n12182), .B1(n16167), .B2(P2_U3088), 
        .C1(n12181), .C2(n14783), .ZN(P2_U3309) );
  AOI22_X1 U14098 ( .A1(n16359), .A2(n14831), .B1(n14817), .B2(n15053), .ZN(
        n12501) );
  AOI22_X1 U14099 ( .A1(n16359), .A2(n14856), .B1(n11694), .B2(n15053), .ZN(
        n12184) );
  XNOR2_X1 U14100 ( .A(n12184), .B(n11130), .ZN(n12500) );
  XOR2_X1 U14101 ( .A(n12501), .B(n12500), .Z(n12191) );
  INV_X1 U14102 ( .A(n12185), .ZN(n12187) );
  OAI21_X1 U14103 ( .B1(n12191), .B2(n12190), .A(n12503), .ZN(n12192) );
  NAND2_X1 U14104 ( .A1(n12192), .A2(n15012), .ZN(n12200) );
  INV_X1 U14105 ( .A(n12193), .ZN(n12198) );
  INV_X1 U14106 ( .A(n12194), .ZN(n12197) );
  INV_X1 U14107 ( .A(n15052), .ZN(n12564) );
  OAI22_X1 U14108 ( .A1(n12195), .A2(n15038), .B1(n15037), .B2(n12564), .ZN(
        n12196) );
  AOI211_X1 U14109 ( .C1(n12198), .C2(n15017), .A(n12197), .B(n12196), .ZN(
        n12199) );
  OAI211_X1 U14110 ( .C1(n12201), .C2(n15026), .A(n12200), .B(n12199), .ZN(
        P1_U3221) );
  XNOR2_X1 U14111 ( .A(n13265), .B(n12427), .ZN(n12330) );
  XNOR2_X1 U14112 ( .A(n12330), .B(n13664), .ZN(n12208) );
  NAND2_X1 U14113 ( .A1(n12202), .A2(n13665), .ZN(n12203) );
  INV_X1 U14114 ( .A(n12334), .ZN(n12206) );
  AOI21_X1 U14115 ( .B1(n12208), .B2(n12207), .A(n12206), .ZN(n12215) );
  INV_X1 U14116 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n12209) );
  NOR2_X1 U14117 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12209), .ZN(n13679) );
  INV_X1 U14118 ( .A(n13450), .ZN(n13406) );
  OAI22_X1 U14119 ( .A1(n12210), .A2(n13406), .B1(n12427), .B2(n13453), .ZN(
        n12211) );
  AOI211_X1 U14120 ( .C1(n13439), .C2(n13663), .A(n13679), .B(n12211), .ZN(
        n12214) );
  INV_X1 U14121 ( .A(n13447), .ZN(n13414) );
  INV_X1 U14122 ( .A(n12212), .ZN(n12475) );
  NAND2_X1 U14123 ( .A1(n13414), .A2(n12475), .ZN(n12213) );
  OAI211_X1 U14124 ( .C1(n12215), .C2(n13421), .A(n12214), .B(n12213), .ZN(
        P3_U3170) );
  AND2_X1 U14125 ( .A1(n14403), .A2(n14305), .ZN(n12217) );
  XNOR2_X1 U14126 ( .A(n12259), .B(n14306), .ZN(n12216) );
  NOR2_X1 U14127 ( .A1(n12216), .A2(n12217), .ZN(n12403) );
  AOI21_X1 U14128 ( .B1(n12217), .B2(n12216), .A(n12403), .ZN(n12222) );
  INV_X1 U14129 ( .A(n12218), .ZN(n12219) );
  OAI21_X1 U14130 ( .B1(n12222), .B2(n12221), .A(n12404), .ZN(n12223) );
  NAND2_X1 U14131 ( .A1(n12223), .A2(n14382), .ZN(n12230) );
  INV_X1 U14132 ( .A(n12224), .ZN(n12227) );
  OAI22_X1 U14133 ( .A1(n12225), .A2(n14362), .B1(n14387), .B2(n12316), .ZN(
        n12226) );
  AOI211_X1 U14134 ( .C1(n12228), .C2(n14385), .A(n12227), .B(n12226), .ZN(
        n12229) );
  OAI211_X1 U14135 ( .C1(n7598), .C2(n14393), .A(n12230), .B(n12229), .ZN(
        P2_U3203) );
  MUX2_X1 U14136 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13775), .Z(n12364) );
  XOR2_X1 U14137 ( .A(n12246), .B(n12364), .Z(n12365) );
  INV_X1 U14138 ( .A(n12245), .ZN(n12234) );
  INV_X1 U14139 ( .A(n12231), .ZN(n12233) );
  XOR2_X1 U14140 ( .A(n12365), .B(n12366), .Z(n12254) );
  NAND2_X1 U14141 ( .A1(n12245), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n12235) );
  NOR2_X1 U14142 ( .A1(n12237), .A2(n12363), .ZN(n12238) );
  NAND2_X1 U14143 ( .A1(n12239), .A2(n8672), .ZN(n12241) );
  INV_X1 U14144 ( .A(n12370), .ZN(n12240) );
  NAND2_X1 U14145 ( .A1(n12241), .A2(n12240), .ZN(n12252) );
  INV_X1 U14146 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12242) );
  NOR2_X1 U14147 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12242), .ZN(n12592) );
  AOI21_X1 U14148 ( .B1(n16037), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12592), .ZN(
        n12243) );
  OAI21_X1 U14149 ( .B1(n16278), .B2(n12363), .A(n12243), .ZN(n12251) );
  AOI21_X1 U14150 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n12245), .A(n12244), .ZN(
        n12247) );
  INV_X1 U14151 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n12551) );
  AOI21_X1 U14152 ( .B1(n12248), .B2(n12551), .A(n12359), .ZN(n12249) );
  NOR2_X1 U14153 ( .A1(n12249), .A2(n16280), .ZN(n12250) );
  AOI211_X1 U14154 ( .C1(n13847), .C2(n12252), .A(n12251), .B(n12250), .ZN(
        n12253) );
  OAI21_X1 U14155 ( .B1(n12254), .B2(n16259), .A(n12253), .ZN(P3_U3189) );
  NAND2_X1 U14156 ( .A1(n12255), .A2(n14229), .ZN(n12257) );
  INV_X1 U14157 ( .A(n12256), .ZN(n13653) );
  OAI211_X1 U14158 ( .C1(n12258), .C2(n14237), .A(n12257), .B(n13653), .ZN(
        P3_U3272) );
  AOI22_X1 U14159 ( .A1(n12260), .A2(n14734), .B1(n14733), .B2(n12259), .ZN(
        n12261) );
  OAI211_X1 U14160 ( .C1(n12263), .C2(n16299), .A(n12262), .B(n12261), .ZN(
        n12265) );
  NAND2_X1 U14161 ( .A1(n12265), .A2(n16413), .ZN(n12264) );
  OAI21_X1 U14162 ( .B1(n16413), .B2(n9508), .A(n12264), .ZN(P2_U3508) );
  INV_X1 U14163 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U14164 ( .A1(n12265), .A2(n14760), .ZN(n12266) );
  OAI21_X1 U14165 ( .B1(n14760), .B2(n12267), .A(n12266), .ZN(P2_U3457) );
  NOR2_X1 U14166 ( .A1(n12268), .A2(n12273), .ZN(n12270) );
  NOR2_X1 U14167 ( .A1(n12270), .A2(n12269), .ZN(n12272) );
  XNOR2_X1 U14168 ( .A(n12518), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n12271) );
  NOR2_X1 U14169 ( .A1(n12272), .A2(n12271), .ZN(n12514) );
  AOI211_X1 U14170 ( .C1(n12272), .C2(n12271), .A(n16182), .B(n12514), .ZN(
        n12283) );
  NOR2_X1 U14171 ( .A1(n12274), .A2(n12273), .ZN(n12276) );
  NOR2_X1 U14172 ( .A1(n12276), .A2(n12275), .ZN(n12278) );
  XNOR2_X1 U14173 ( .A(n12518), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n12277) );
  NOR2_X1 U14174 ( .A1(n12278), .A2(n12277), .ZN(n12517) );
  AOI211_X1 U14175 ( .C1(n12278), .C2(n12277), .A(n16177), .B(n12517), .ZN(
        n12282) );
  AND2_X1 U14176 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13159) );
  AOI21_X1 U14177 ( .B1(n16055), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13159), 
        .ZN(n12279) );
  OAI21_X1 U14178 ( .B1(n12280), .B2(n16168), .A(n12279), .ZN(n12281) );
  OR3_X1 U14179 ( .A1(n12283), .A2(n12282), .A3(n12281), .ZN(P2_U3230) );
  OR2_X1 U14180 ( .A1(n12496), .A2(n15052), .ZN(n12284) );
  NAND2_X1 U14181 ( .A1(n12285), .A2(n12284), .ZN(n12457) );
  INV_X1 U14182 ( .A(n12294), .ZN(n12456) );
  XNOR2_X1 U14183 ( .A(n12457), .B(n12456), .ZN(n12414) );
  INV_X1 U14184 ( .A(n12567), .ZN(n12560) );
  OAI21_X1 U14185 ( .B1(n12286), .B2(n12560), .A(n16326), .ZN(n12287) );
  OR2_X1 U14186 ( .A1(n12287), .A2(n12611), .ZN(n12289) );
  NAND2_X1 U14187 ( .A1(n15050), .A2(n15448), .ZN(n12288) );
  AND2_X1 U14188 ( .A1(n12289), .A2(n12288), .ZN(n12419) );
  NOR2_X1 U14189 ( .A1(n12496), .A2(n12564), .ZN(n12290) );
  NAND2_X1 U14190 ( .A1(n12496), .A2(n12564), .ZN(n12292) );
  NAND2_X1 U14191 ( .A1(n7545), .A2(n12456), .ZN(n12416) );
  NAND3_X1 U14192 ( .A1(n12416), .A2(n15269), .A3(n12452), .ZN(n12298) );
  AND2_X1 U14193 ( .A1(n15052), .A2(n15386), .ZN(n12415) );
  OAI22_X1 U14194 ( .A1(n15430), .A2(n11329), .B1(n12563), .B2(n15428), .ZN(
        n12296) );
  NOR2_X1 U14195 ( .A1(n12560), .A2(n15434), .ZN(n12295) );
  AOI211_X1 U14196 ( .C1(n12415), .C2(n15432), .A(n12296), .B(n12295), .ZN(
        n12297) );
  OAI211_X1 U14197 ( .C1(n12419), .C2(n15168), .A(n12298), .B(n12297), .ZN(
        n12299) );
  AOI21_X1 U14198 ( .B1(n12414), .B2(n15224), .A(n12299), .ZN(n12300) );
  INV_X1 U14199 ( .A(n12300), .ZN(P1_U3283) );
  XNOR2_X1 U14200 ( .A(n12301), .B(n13503), .ZN(n12426) );
  NAND2_X1 U14201 ( .A1(n12426), .A2(n12302), .ZN(n12310) );
  NAND2_X1 U14202 ( .A1(n12304), .A2(n12303), .ZN(n12306) );
  NAND2_X1 U14203 ( .A1(n12306), .A2(n13624), .ZN(n12305) );
  OAI211_X1 U14204 ( .C1(n12306), .C2(n13624), .A(n12305), .B(n16309), .ZN(
        n12308) );
  AOI22_X1 U14205 ( .A1(n16313), .A2(n13663), .B1(n13665), .B2(n16311), .ZN(
        n12307) );
  AND2_X1 U14206 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  NAND2_X1 U14207 ( .A1(n12310), .A2(n12309), .ZN(n12425) );
  INV_X1 U14208 ( .A(n12425), .ZN(n12474) );
  INV_X1 U14209 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n12311) );
  OAI22_X1 U14210 ( .A1(n14221), .A2(n12427), .B1(n16476), .B2(n12311), .ZN(
        n12312) );
  AOI21_X1 U14211 ( .B1(n12426), .B2(n12937), .A(n12312), .ZN(n12313) );
  OAI21_X1 U14212 ( .B1(n12474), .B2(n16483), .A(n12313), .ZN(P3_U3402) );
  XNOR2_X1 U14213 ( .A(n12315), .B(n12314), .ZN(n12317) );
  OAI22_X1 U14214 ( .A1(n12316), .A2(n14621), .B1(n12783), .B2(n14623), .ZN(
        n12488) );
  AOI21_X1 U14215 ( .B1(n12317), .B2(n14603), .A(n12488), .ZN(n12468) );
  INV_X1 U14216 ( .A(n12318), .ZN(n12321) );
  OAI21_X1 U14217 ( .B1(n12321), .B2(n12320), .A(n12319), .ZN(n12469) );
  OAI22_X1 U14218 ( .A1(n16458), .A2(n12322), .B1(n12491), .B2(n16455), .ZN(
        n12323) );
  AOI21_X1 U14219 ( .B1(n12487), .B2(n16463), .A(n12323), .ZN(n12327) );
  OAI21_X1 U14220 ( .B1(n12349), .B2(n12324), .A(n14734), .ZN(n12325) );
  NOR2_X1 U14221 ( .A1(n12325), .A2(n12742), .ZN(n12466) );
  NAND2_X1 U14222 ( .A1(n12466), .A2(n14596), .ZN(n12326) );
  OAI211_X1 U14223 ( .C1(n12469), .C2(n14638), .A(n12327), .B(n12326), .ZN(
        n12328) );
  INV_X1 U14224 ( .A(n12328), .ZN(n12329) );
  OAI21_X1 U14225 ( .B1(n14598), .B2(n12468), .A(n12329), .ZN(P2_U3254) );
  INV_X1 U14226 ( .A(n12330), .ZN(n12332) );
  NAND2_X1 U14227 ( .A1(n12332), .A2(n12331), .ZN(n12333) );
  NAND2_X1 U14228 ( .A1(n12334), .A2(n12333), .ZN(n12579) );
  XNOR2_X1 U14229 ( .A(n13265), .B(n12336), .ZN(n12581) );
  XNOR2_X1 U14230 ( .A(n12581), .B(n13663), .ZN(n12578) );
  XNOR2_X1 U14231 ( .A(n12335), .B(n12578), .ZN(n12341) );
  AOI22_X1 U14232 ( .A1(n13418), .A2(n12336), .B1(n13664), .B2(n13450), .ZN(
        n12339) );
  AOI21_X1 U14233 ( .B1(n13662), .B2(n13439), .A(n12337), .ZN(n12338) );
  OAI211_X1 U14234 ( .C1(n13447), .C2(n12531), .A(n12339), .B(n12338), .ZN(
        n12340) );
  AOI21_X1 U14235 ( .B1(n12341), .B2(n13442), .A(n12340), .ZN(n12342) );
  INV_X1 U14236 ( .A(n12342), .ZN(P3_U3167) );
  XOR2_X1 U14237 ( .A(n12343), .B(n12345), .Z(n12348) );
  XOR2_X1 U14238 ( .A(n12345), .B(n12344), .Z(n16411) );
  OAI22_X1 U14239 ( .A1(n12691), .A2(n14623), .B1(n12408), .B2(n14621), .ZN(
        n12346) );
  AOI21_X1 U14240 ( .B1(n16411), .B2(n14522), .A(n12346), .ZN(n12347) );
  OAI21_X1 U14241 ( .B1(n14619), .B2(n12348), .A(n12347), .ZN(n16409) );
  INV_X1 U14242 ( .A(n16409), .ZN(n12358) );
  INV_X1 U14243 ( .A(n12400), .ZN(n16408) );
  INV_X1 U14244 ( .A(n12349), .ZN(n12350) );
  OAI211_X1 U14245 ( .C1(n16408), .C2(n12351), .A(n12350), .B(n14734), .ZN(
        n16406) );
  INV_X1 U14246 ( .A(n12352), .ZN(n12411) );
  AOI22_X1 U14247 ( .A1(n14598), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12411), 
        .B2(n14611), .ZN(n12354) );
  NAND2_X1 U14248 ( .A1(n16463), .A2(n12400), .ZN(n12353) );
  OAI211_X1 U14249 ( .C1(n16406), .C2(n12355), .A(n12354), .B(n12353), .ZN(
        n12356) );
  AOI21_X1 U14250 ( .B1(n16411), .B2(n16453), .A(n12356), .ZN(n12357) );
  OAI21_X1 U14251 ( .B1(n12358), .B2(n14598), .A(n12357), .ZN(P2_U3255) );
  NAND2_X1 U14252 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n12672), .ZN(n12360) );
  OAI21_X1 U14253 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n12672), .A(n12360), .ZN(
        n12361) );
  AOI21_X1 U14254 ( .B1(n12362), .B2(n12361), .A(n12663), .ZN(n12380) );
  MUX2_X1 U14255 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13775), .Z(n12652) );
  XOR2_X1 U14256 ( .A(n12672), .B(n12652), .Z(n12655) );
  XNOR2_X1 U14257 ( .A(n12656), .B(n12655), .ZN(n12367) );
  NAND2_X1 U14258 ( .A1(n12367), .A2(n16272), .ZN(n12379) );
  INV_X1 U14259 ( .A(n12672), .ZN(n12654) );
  NOR2_X1 U14260 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15892), .ZN(n13328) );
  INV_X1 U14261 ( .A(n13328), .ZN(n12368) );
  OAI21_X1 U14262 ( .B1(n16292), .B2(n12369), .A(n12368), .ZN(n12377) );
  NAND2_X1 U14263 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n12672), .ZN(n12372) );
  OAI21_X1 U14264 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n12672), .A(n12372), .ZN(
        n12373) );
  AOI21_X1 U14265 ( .B1(n12374), .B2(n12373), .A(n12674), .ZN(n12375) );
  NOR2_X1 U14266 ( .A1(n12375), .A2(n16285), .ZN(n12376) );
  AOI211_X1 U14267 ( .C1(n13813), .C2(n12654), .A(n12377), .B(n12376), .ZN(
        n12378) );
  OAI211_X1 U14268 ( .C1(n12380), .C2(n16280), .A(n12379), .B(n12378), .ZN(
        P3_U3190) );
  INV_X1 U14269 ( .A(n12381), .ZN(n12383) );
  OAI222_X1 U14270 ( .A1(n14783), .A2(n12382), .B1(n14780), .B2(n12383), .C1(
        P2_U3088), .C2(n14508), .ZN(P2_U3308) );
  OAI222_X1 U14271 ( .A1(n7555), .A2(n8186), .B1(n15627), .B2(n12383), .C1(
        P1_U3086), .C2(n15157), .ZN(P1_U3336) );
  MUX2_X1 U14272 ( .A(n12620), .B(P1_REG2_REG_14__SCAN_IN), .S(n12394), .Z(
        n12387) );
  NOR2_X1 U14273 ( .A1(n12385), .A2(n12384), .ZN(n12389) );
  INV_X1 U14274 ( .A(n12389), .ZN(n12386) );
  NAND2_X1 U14275 ( .A1(n12387), .A2(n12386), .ZN(n12390) );
  MUX2_X1 U14276 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n12620), .S(n12394), .Z(
        n12388) );
  OAI21_X1 U14277 ( .B1(n12391), .B2(n12389), .A(n12388), .ZN(n12619) );
  OAI211_X1 U14278 ( .C1(n12391), .C2(n12390), .A(n12619), .B(n15154), .ZN(
        n12399) );
  NAND2_X1 U14279 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14895)
         );
  AOI21_X1 U14280 ( .B1(n12393), .B2(P1_REG1_REG_13__SCAN_IN), .A(n12392), 
        .ZN(n12623) );
  XOR2_X1 U14281 ( .A(n12394), .B(n12623), .Z(n12625) );
  XNOR2_X1 U14282 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n12625), .ZN(n12395) );
  NAND2_X1 U14283 ( .A1(n15155), .A2(n12395), .ZN(n12396) );
  NAND2_X1 U14284 ( .A1(n14895), .A2(n12396), .ZN(n12397) );
  AOI21_X1 U14285 ( .B1(n16197), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n12397), 
        .ZN(n12398) );
  OAI211_X1 U14286 ( .C1(n15149), .C2(n12622), .A(n12399), .B(n12398), .ZN(
        P1_U3257) );
  AND2_X1 U14287 ( .A1(n14402), .A2(n14305), .ZN(n12402) );
  XNOR2_X1 U14288 ( .A(n12400), .B(n14306), .ZN(n12401) );
  NOR2_X1 U14289 ( .A1(n12401), .A2(n12402), .ZN(n12482) );
  AOI21_X1 U14290 ( .B1(n12402), .B2(n12401), .A(n12482), .ZN(n12406) );
  OAI21_X1 U14291 ( .B1(n12406), .B2(n12405), .A(n12484), .ZN(n12407) );
  NAND2_X1 U14292 ( .A1(n12407), .A2(n14382), .ZN(n12413) );
  NAND2_X1 U14293 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n16189)
         );
  INV_X1 U14294 ( .A(n16189), .ZN(n12410) );
  OAI22_X1 U14295 ( .A1(n12691), .A2(n14387), .B1(n14362), .B2(n12408), .ZN(
        n12409) );
  AOI211_X1 U14296 ( .C1(n12411), .C2(n14385), .A(n12410), .B(n12409), .ZN(
        n12412) );
  OAI211_X1 U14297 ( .C1(n16408), .C2(n14393), .A(n12413), .B(n12412), .ZN(
        P2_U3189) );
  INV_X1 U14298 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n12422) );
  NAND2_X1 U14299 ( .A1(n12414), .A2(n15568), .ZN(n12420) );
  AOI21_X1 U14300 ( .B1(n12567), .B2(n16358), .A(n12415), .ZN(n12418) );
  NAND3_X1 U14301 ( .A1(n12416), .A2(n15584), .A3(n12452), .ZN(n12417) );
  NAND4_X1 U14302 ( .A1(n12420), .A2(n12419), .A3(n12418), .A4(n12417), .ZN(
        n12423) );
  NAND2_X1 U14303 ( .A1(n12423), .A2(n16338), .ZN(n12421) );
  OAI21_X1 U14304 ( .B1(n16338), .B2(n12422), .A(n12421), .ZN(P1_U3489) );
  NAND2_X1 U14305 ( .A1(n12423), .A2(n16446), .ZN(n12424) );
  OAI21_X1 U14306 ( .B1(n16446), .B2(n10419), .A(n12424), .ZN(P1_U3538) );
  MUX2_X1 U14307 ( .A(n12425), .B(P3_REG1_REG_4__SCAN_IN), .S(n10822), .Z(
        n12429) );
  INV_X1 U14308 ( .A(n12426), .ZN(n12479) );
  OAI22_X1 U14309 ( .A1(n12479), .A2(n14165), .B1(n12427), .B2(n14164), .ZN(
        n12428) );
  OR2_X1 U14310 ( .A1(n12429), .A2(n12428), .ZN(P3_U3463) );
  NAND2_X1 U14311 ( .A1(n12431), .A2(n12430), .ZN(n12526) );
  INV_X1 U14312 ( .A(n12526), .ZN(n16346) );
  NAND2_X1 U14313 ( .A1(n16386), .A2(n16346), .ZN(n14104) );
  INV_X1 U14314 ( .A(n14104), .ZN(n14084) );
  OAI22_X1 U14315 ( .A1(n14075), .A2(n12432), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n16339), .ZN(n12435) );
  MUX2_X1 U14316 ( .A(n12433), .B(P3_REG2_REG_3__SCAN_IN), .S(n16348), .Z(
        n12434) );
  AOI211_X1 U14317 ( .C1(n14084), .C2(n12436), .A(n12435), .B(n12434), .ZN(
        n12437) );
  INV_X1 U14318 ( .A(n12437), .ZN(P3_U3230) );
  OAI21_X1 U14319 ( .B1(n12439), .B2(n13621), .A(n12438), .ZN(n12650) );
  NAND2_X1 U14320 ( .A1(n12440), .A2(n13621), .ZN(n12441) );
  NAND3_X1 U14321 ( .A1(n12442), .A2(n16309), .A3(n12441), .ZN(n12444) );
  AOI22_X1 U14322 ( .A1(n16313), .A2(n13661), .B1(n13663), .B2(n16311), .ZN(
        n12443) );
  NAND2_X1 U14323 ( .A1(n12444), .A2(n12443), .ZN(n12647) );
  AOI21_X1 U14324 ( .B1(n10820), .B2(n12650), .A(n12647), .ZN(n12450) );
  INV_X1 U14325 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n12445) );
  OAI22_X1 U14326 ( .A1(n14164), .A2(n12646), .B1(n16473), .B2(n12445), .ZN(
        n12446) );
  INV_X1 U14327 ( .A(n12446), .ZN(n12447) );
  OAI21_X1 U14328 ( .B1(n12450), .B2(n10822), .A(n12447), .ZN(P3_U3465) );
  OAI22_X1 U14329 ( .A1(n14221), .A2(n12646), .B1(n16476), .B2(n8650), .ZN(
        n12448) );
  INV_X1 U14330 ( .A(n12448), .ZN(n12449) );
  OAI21_X1 U14331 ( .B1(n12450), .B2(n16483), .A(n12449), .ZN(P3_U3408) );
  INV_X1 U14332 ( .A(n15051), .ZN(n12709) );
  OR2_X1 U14333 ( .A1(n12567), .A2(n12709), .ZN(n12451) );
  XNOR2_X1 U14334 ( .A(n12605), .B(n12460), .ZN(n12453) );
  OAI222_X1 U14335 ( .A1(n15410), .A2(n12722), .B1(n15451), .B2(n12709), .C1(
        n12453), .C2(n15567), .ZN(n16430) );
  INV_X1 U14336 ( .A(n16430), .ZN(n12465) );
  OAI22_X1 U14337 ( .A1(n15430), .A2(n10433), .B1(n12708), .B2(n15428), .ZN(
        n12455) );
  XNOR2_X1 U14338 ( .A(n12611), .B(n16427), .ZN(n16429) );
  NOR2_X1 U14339 ( .A1(n16429), .A2(n15398), .ZN(n12454) );
  AOI211_X1 U14340 ( .C1(n15459), .C2(n12712), .A(n12455), .B(n12454), .ZN(
        n12464) );
  OR2_X1 U14341 ( .A1(n12567), .A2(n15051), .ZN(n12458) );
  AND2_X1 U14342 ( .A1(n12459), .A2(n12460), .ZN(n16426) );
  INV_X1 U14343 ( .A(n16426), .ZN(n12462) );
  NAND3_X1 U14344 ( .A1(n12462), .A2(n15425), .A3(n12600), .ZN(n12463) );
  OAI211_X1 U14345 ( .C1(n12465), .C2(n15356), .A(n12464), .B(n12463), .ZN(
        P1_U3282) );
  INV_X2 U14346 ( .A(n16412), .ZN(n16413) );
  AOI21_X1 U14347 ( .B1(n14733), .B2(n12487), .A(n12466), .ZN(n12467) );
  OAI211_X1 U14348 ( .C1(n12469), .C2(n14739), .A(n12468), .B(n12467), .ZN(
        n12471) );
  NAND2_X1 U14349 ( .A1(n12471), .A2(n16413), .ZN(n12470) );
  OAI21_X1 U14350 ( .B1(n16413), .B2(n11237), .A(n12470), .ZN(P2_U3510) );
  NAND2_X1 U14351 ( .A1(n12471), .A2(n14760), .ZN(n12472) );
  OAI21_X1 U14352 ( .B1(n14760), .B2(n9544), .A(n12472), .ZN(P2_U3463) );
  INV_X1 U14353 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n12473) );
  MUX2_X1 U14354 ( .A(n12474), .B(n12473), .S(n16348), .Z(n12478) );
  AOI22_X1 U14355 ( .A1(n16384), .A2(n12476), .B1(n16382), .B2(n12475), .ZN(
        n12477) );
  OAI211_X1 U14356 ( .C1(n12479), .C2(n14104), .A(n12478), .B(n12477), .ZN(
        P3_U3229) );
  AND2_X1 U14357 ( .A1(n14401), .A2(n14305), .ZN(n12481) );
  XNOR2_X1 U14358 ( .A(n12487), .B(n14306), .ZN(n12480) );
  NOR2_X1 U14359 ( .A1(n12480), .A2(n12481), .ZN(n12684) );
  AOI21_X1 U14360 ( .B1(n12481), .B2(n12480), .A(n12684), .ZN(n12486) );
  INV_X1 U14361 ( .A(n12482), .ZN(n12483) );
  OAI21_X1 U14362 ( .B1(n12486), .B2(n12485), .A(n12686), .ZN(n12493) );
  NAND2_X1 U14363 ( .A1(n12487), .A2(n14375), .ZN(n12490) );
  AOI22_X1 U14364 ( .A1(n14328), .A2(n12488), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12489) );
  OAI211_X1 U14365 ( .C1(n14373), .C2(n12491), .A(n12490), .B(n12489), .ZN(
        n12492) );
  AOI21_X1 U14366 ( .B1(n12493), .B2(n14382), .A(n12492), .ZN(n12494) );
  INV_X1 U14367 ( .A(n12494), .ZN(P2_U3208) );
  INV_X1 U14368 ( .A(n12496), .ZN(n16391) );
  AND2_X1 U14369 ( .A1(n15052), .A2(n14817), .ZN(n12495) );
  AOI21_X1 U14370 ( .B1(n12496), .B2(n14831), .A(n12495), .ZN(n12556) );
  NAND2_X1 U14371 ( .A1(n12496), .A2(n14856), .ZN(n12498) );
  NAND2_X1 U14372 ( .A1(n15052), .A2(n14831), .ZN(n12497) );
  NAND2_X1 U14373 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  XNOR2_X1 U14374 ( .A(n12499), .B(n11130), .ZN(n12557) );
  XOR2_X1 U14375 ( .A(n12556), .B(n12557), .Z(n12505) );
  AOI211_X1 U14376 ( .C1(n12505), .C2(n12504), .A(n15044), .B(n7543), .ZN(
        n12506) );
  INV_X1 U14377 ( .A(n12506), .ZN(n12513) );
  INV_X1 U14378 ( .A(n12507), .ZN(n12511) );
  OAI22_X1 U14379 ( .A1(n12508), .A2(n15038), .B1(n15037), .B2(n12709), .ZN(
        n12509) );
  AOI211_X1 U14380 ( .C1(n15017), .C2(n12511), .A(n12510), .B(n12509), .ZN(
        n12512) );
  OAI211_X1 U14381 ( .C1(n16391), .C2(n15026), .A(n12513), .B(n12512), .ZN(
        P1_U3231) );
  AOI21_X1 U14382 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n12518), .A(n12514), 
        .ZN(n12516) );
  XNOR2_X1 U14383 ( .A(n12832), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n12515) );
  NOR2_X1 U14384 ( .A1(n12516), .A2(n12515), .ZN(n12826) );
  AOI211_X1 U14385 ( .C1(n12516), .C2(n12515), .A(n16182), .B(n12826), .ZN(
        n12525) );
  AOI21_X1 U14386 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n12518), .A(n12517), 
        .ZN(n12520) );
  XNOR2_X1 U14387 ( .A(n12832), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n12519) );
  NOR2_X1 U14388 ( .A1(n12520), .A2(n12519), .ZN(n12831) );
  AOI211_X1 U14389 ( .C1(n12520), .C2(n12519), .A(n16177), .B(n12831), .ZN(
        n12524) );
  AND2_X1 U14390 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14338) );
  AOI21_X1 U14391 ( .B1(n16055), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n14338), 
        .ZN(n12521) );
  OAI21_X1 U14392 ( .B1(n12522), .B2(n16168), .A(n12521), .ZN(n12523) );
  OR3_X1 U14393 ( .A1(n12525), .A2(n12524), .A3(n12523), .ZN(P2_U3231) );
  NAND2_X1 U14394 ( .A1(n14097), .A2(n12526), .ZN(n16377) );
  XNOR2_X1 U14395 ( .A(n12527), .B(n13623), .ZN(n12537) );
  OAI21_X1 U14396 ( .B1(n12529), .B2(n13623), .A(n12528), .ZN(n12530) );
  AOI222_X1 U14397 ( .A1(n16309), .A2(n12530), .B1(n13662), .B2(n16313), .C1(
        n13664), .C2(n16311), .ZN(n12536) );
  INV_X1 U14398 ( .A(n12536), .ZN(n12534) );
  NOR2_X1 U14399 ( .A1(n16386), .A2(n11770), .ZN(n12533) );
  OAI22_X1 U14400 ( .A1(n14075), .A2(n12541), .B1(n12531), .B2(n16339), .ZN(
        n12532) );
  AOI211_X1 U14401 ( .C1(n12534), .C2(n16386), .A(n12533), .B(n12532), .ZN(
        n12535) );
  OAI21_X1 U14402 ( .B1(n14054), .B2(n12537), .A(n12535), .ZN(P3_U3228) );
  OAI21_X1 U14403 ( .B1(n14150), .B2(n12537), .A(n12536), .ZN(n12543) );
  OAI22_X1 U14404 ( .A1(n14164), .A2(n12541), .B1(n16473), .B2(n11769), .ZN(
        n12538) );
  AOI21_X1 U14405 ( .B1(n12543), .B2(n16473), .A(n12538), .ZN(n12539) );
  INV_X1 U14406 ( .A(n12539), .ZN(P3_U3464) );
  INV_X1 U14407 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n12540) );
  OAI22_X1 U14408 ( .A1(n14221), .A2(n12541), .B1(n16476), .B2(n12540), .ZN(
        n12542) );
  AOI21_X1 U14409 ( .B1(n12543), .B2(n16476), .A(n12542), .ZN(n12544) );
  INV_X1 U14410 ( .A(n12544), .ZN(P3_U3405) );
  OAI211_X1 U14411 ( .C1(n12546), .C2(n13622), .A(n12545), .B(n16309), .ZN(
        n12548) );
  AOI22_X1 U14412 ( .A1(n16311), .A2(n13662), .B1(n13660), .B2(n16313), .ZN(
        n12547) );
  NAND2_X1 U14413 ( .A1(n12548), .A2(n12547), .ZN(n12570) );
  INV_X1 U14414 ( .A(n12570), .ZN(n12555) );
  OAI21_X1 U14415 ( .B1(n12550), .B2(n13518), .A(n12549), .ZN(n12571) );
  NOR2_X1 U14416 ( .A1(n16386), .A2(n12551), .ZN(n12553) );
  OAI22_X1 U14417 ( .A1(n14075), .A2(n12589), .B1(n12595), .B2(n16339), .ZN(
        n12552) );
  AOI211_X1 U14418 ( .C1(n12571), .C2(n14039), .A(n12553), .B(n12552), .ZN(
        n12554) );
  OAI21_X1 U14419 ( .B1(n12555), .B2(n16348), .A(n12554), .ZN(P3_U3226) );
  INV_X1 U14420 ( .A(n12556), .ZN(n12558) );
  AND2_X1 U14421 ( .A1(n15051), .A2(n14817), .ZN(n12559) );
  AOI21_X1 U14422 ( .B1(n12567), .B2(n14831), .A(n12559), .ZN(n12702) );
  OAI22_X1 U14423 ( .A1(n12560), .A2(n14932), .B1(n12709), .B2(n14935), .ZN(
        n12561) );
  XNOR2_X1 U14424 ( .A(n12561), .B(n11130), .ZN(n12700) );
  XOR2_X1 U14425 ( .A(n12702), .B(n12700), .Z(n12703) );
  XNOR2_X1 U14426 ( .A(n12704), .B(n12703), .ZN(n12569) );
  OAI21_X1 U14427 ( .B1(n15036), .B2(n12563), .A(n12562), .ZN(n12566) );
  INV_X1 U14428 ( .A(n15050), .ZN(n12857) );
  OAI22_X1 U14429 ( .A1(n12564), .A2(n15038), .B1(n15037), .B2(n12857), .ZN(
        n12565) );
  AOI211_X1 U14430 ( .C1(n12567), .C2(n15042), .A(n12566), .B(n12565), .ZN(
        n12568) );
  OAI21_X1 U14431 ( .B1(n12569), .B2(n15044), .A(n12568), .ZN(P1_U3217) );
  AOI21_X1 U14432 ( .B1(n10820), .B2(n12571), .A(n12570), .ZN(n12577) );
  OAI22_X1 U14433 ( .A1(n14164), .A2(n12589), .B1(n16473), .B2(n8672), .ZN(
        n12572) );
  INV_X1 U14434 ( .A(n12572), .ZN(n12573) );
  OAI21_X1 U14435 ( .B1(n12577), .B2(n10822), .A(n12573), .ZN(P3_U3466) );
  INV_X1 U14436 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n12574) );
  OAI22_X1 U14437 ( .A1(n14221), .A2(n12589), .B1(n16476), .B2(n12574), .ZN(
        n12575) );
  INV_X1 U14438 ( .A(n12575), .ZN(n12576) );
  OAI21_X1 U14439 ( .B1(n12577), .B2(n16483), .A(n12576), .ZN(P3_U3411) );
  NAND2_X1 U14440 ( .A1(n12579), .A2(n12578), .ZN(n12583) );
  NAND2_X1 U14441 ( .A1(n12581), .A2(n12580), .ZN(n12582) );
  XNOR2_X1 U14442 ( .A(n7663), .B(n12646), .ZN(n12584) );
  XNOR2_X1 U14443 ( .A(n12584), .B(n13662), .ZN(n12638) );
  NAND2_X1 U14444 ( .A1(n12584), .A2(n13662), .ZN(n12585) );
  XNOR2_X1 U14445 ( .A(n7663), .B(n12586), .ZN(n12863) );
  XNOR2_X1 U14446 ( .A(n12863), .B(n13661), .ZN(n12587) );
  OAI211_X1 U14447 ( .C1(n12588), .C2(n12587), .A(n12866), .B(n13442), .ZN(
        n12594) );
  OAI22_X1 U14448 ( .A1(n12590), .A2(n13406), .B1(n13453), .B2(n12589), .ZN(
        n12591) );
  AOI211_X1 U14449 ( .C1(n13439), .C2(n13660), .A(n12592), .B(n12591), .ZN(
        n12593) );
  OAI211_X1 U14450 ( .C1(n12595), .C2(n13447), .A(n12594), .B(n12593), .ZN(
        P3_U3153) );
  INV_X1 U14451 ( .A(n12596), .ZN(n13176) );
  OAI222_X1 U14452 ( .A1(n7555), .A2(n12598), .B1(n15627), .B2(n13176), .C1(
        n12597), .C2(P1_U3086), .ZN(P1_U3335) );
  NAND2_X1 U14453 ( .A1(n12712), .A2(n15050), .ZN(n12599) );
  NAND2_X1 U14454 ( .A1(n12602), .A2(n12715), .ZN(n12603) );
  NAND2_X1 U14455 ( .A1(n12720), .A2(n12603), .ZN(n16441) );
  NAND2_X1 U14456 ( .A1(n12712), .A2(n12857), .ZN(n12604) );
  OR2_X1 U14457 ( .A1(n12712), .A2(n12857), .ZN(n12606) );
  NAND2_X1 U14458 ( .A1(n12607), .A2(n12606), .ZN(n12716) );
  XNOR2_X1 U14459 ( .A(n12716), .B(n12715), .ZN(n12609) );
  AOI22_X1 U14460 ( .A1(n15448), .A2(n15048), .B1(n15050), .B2(n15386), .ZN(
        n12608) );
  OAI21_X1 U14461 ( .B1(n12609), .B2(n15567), .A(n12608), .ZN(n12610) );
  AOI21_X1 U14462 ( .B1(n16441), .B2(n15445), .A(n12610), .ZN(n16443) );
  AOI21_X1 U14463 ( .B1(n12612), .B2(n12851), .A(n16428), .ZN(n12613) );
  NAND2_X1 U14464 ( .A1(n12613), .A2(n12721), .ZN(n16436) );
  OAI22_X1 U14465 ( .A1(n15430), .A2(n12614), .B1(n12855), .B2(n15428), .ZN(
        n12615) );
  AOI21_X1 U14466 ( .B1(n12851), .B2(n15459), .A(n12615), .ZN(n12616) );
  OAI21_X1 U14467 ( .B1(n16436), .B2(n15168), .A(n12616), .ZN(n12617) );
  AOI21_X1 U14468 ( .B1(n16441), .B2(n15460), .A(n12617), .ZN(n12618) );
  OAI21_X1 U14469 ( .B1(n16443), .B2(n15356), .A(n12618), .ZN(P1_U3281) );
  OAI21_X1 U14470 ( .B1(n12622), .B2(n12620), .A(n12619), .ZN(n12797) );
  XNOR2_X1 U14471 ( .A(n12797), .B(n12805), .ZN(n12621) );
  NOR2_X1 U14472 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n12621), .ZN(n12798) );
  AOI21_X1 U14473 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n12621), .A(n12798), 
        .ZN(n12634) );
  INV_X1 U14474 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n12624) );
  NOR2_X1 U14475 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n12626), .ZN(n12806) );
  AOI21_X1 U14476 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n12626), .A(n12806), 
        .ZN(n12628) );
  OR2_X1 U14477 ( .A1(n12628), .A2(n12627), .ZN(n12633) );
  NOR2_X1 U14478 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15034), .ZN(n12631) );
  NOR2_X1 U14479 ( .A1(n15149), .A2(n12629), .ZN(n12630) );
  AOI211_X1 U14480 ( .C1(n16197), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n12631), 
        .B(n12630), .ZN(n12632) );
  OAI211_X1 U14481 ( .C1(n12634), .C2(n15150), .A(n12633), .B(n12632), .ZN(
        P1_U3258) );
  INV_X1 U14482 ( .A(n12635), .ZN(n12636) );
  AOI211_X1 U14483 ( .C1(n12638), .C2(n12637), .A(n13421), .B(n12636), .ZN(
        n12644) );
  AOI22_X1 U14484 ( .A1(n13418), .A2(n12639), .B1(n13663), .B2(n13450), .ZN(
        n12642) );
  AOI21_X1 U14485 ( .B1(n13661), .B2(n13439), .A(n12640), .ZN(n12641) );
  OAI211_X1 U14486 ( .C1(n13447), .C2(n12645), .A(n12642), .B(n12641), .ZN(
        n12643) );
  OR2_X1 U14487 ( .A1(n12644), .A2(n12643), .ZN(P3_U3179) );
  OAI22_X1 U14488 ( .A1(n14075), .A2(n12646), .B1(n12645), .B2(n16339), .ZN(
        n12649) );
  MUX2_X1 U14489 ( .A(n12647), .B(P3_REG2_REG_6__SCAN_IN), .S(n16348), .Z(
        n12648) );
  AOI211_X1 U14490 ( .C1(n14039), .C2(n12650), .A(n12649), .B(n12648), .ZN(
        n12651) );
  INV_X1 U14491 ( .A(n12651), .ZN(P3_U3227) );
  MUX2_X1 U14492 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13775), .Z(n12888) );
  XNOR2_X1 U14493 ( .A(n12888), .B(n12900), .ZN(n12661) );
  MUX2_X1 U14494 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13775), .Z(n12657) );
  INV_X1 U14495 ( .A(n12657), .ZN(n12658) );
  INV_X1 U14496 ( .A(n12652), .ZN(n12653) );
  XNOR2_X1 U14497 ( .A(n12657), .B(n12659), .ZN(n16274) );
  NOR2_X1 U14498 ( .A1(n12660), .A2(n12661), .ZN(n12889) );
  AOI21_X1 U14499 ( .B1(n12661), .B2(n12660), .A(n12889), .ZN(n12681) );
  AOI22_X1 U14500 ( .A1(n12891), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n14099), 
        .B2(n12900), .ZN(n12668) );
  AND2_X1 U14501 ( .A1(n12672), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12662) );
  INV_X1 U14502 ( .A(n12664), .ZN(n12666) );
  INV_X1 U14503 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n16389) );
  OAI21_X1 U14504 ( .B1(n12665), .B2(n16279), .A(n12664), .ZN(n16277) );
  AOI21_X1 U14505 ( .B1(n12668), .B2(n12667), .A(n12901), .ZN(n12671) );
  NAND2_X1 U14506 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n13044)
         );
  INV_X1 U14507 ( .A(n13044), .ZN(n12669) );
  AOI21_X1 U14508 ( .B1(n16037), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12669), 
        .ZN(n12670) );
  OAI21_X1 U14509 ( .B1(n16280), .B2(n12671), .A(n12670), .ZN(n12679) );
  AND2_X1 U14510 ( .A1(n12672), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n12673) );
  INV_X1 U14511 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16270) );
  INV_X1 U14512 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n16403) );
  AOI22_X1 U14513 ( .A1(n12891), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n16403), 
        .B2(n12900), .ZN(n12675) );
  AOI21_X1 U14514 ( .B1(n12676), .B2(n12675), .A(n12895), .ZN(n12677) );
  NOR2_X1 U14515 ( .A1(n12677), .A2(n16285), .ZN(n12678) );
  AOI211_X1 U14516 ( .C1(n13813), .C2(n12891), .A(n12679), .B(n12678), .ZN(
        n12680) );
  OAI21_X1 U14517 ( .B1(n12681), .B2(n16259), .A(n12680), .ZN(P3_U3192) );
  AND2_X1 U14518 ( .A1(n14400), .A2(n14305), .ZN(n12683) );
  XNOR2_X1 U14519 ( .A(n16462), .B(n14306), .ZN(n12682) );
  NOR2_X1 U14520 ( .A1(n12682), .A2(n12683), .ZN(n12772) );
  AOI21_X1 U14521 ( .B1(n12683), .B2(n12682), .A(n12772), .ZN(n12688) );
  INV_X1 U14522 ( .A(n12684), .ZN(n12685) );
  OAI21_X1 U14523 ( .B1(n12688), .B2(n12687), .A(n12773), .ZN(n12689) );
  NAND2_X1 U14524 ( .A1(n12689), .A2(n14382), .ZN(n12696) );
  INV_X1 U14525 ( .A(n16456), .ZN(n12694) );
  INV_X1 U14526 ( .A(n12690), .ZN(n12693) );
  OAI22_X1 U14527 ( .A1(n12691), .A2(n14362), .B1(n14387), .B2(n12949), .ZN(
        n12692) );
  AOI211_X1 U14528 ( .C1(n12694), .C2(n14385), .A(n12693), .B(n12692), .ZN(
        n12695) );
  OAI211_X1 U14529 ( .C1(n12697), .C2(n14393), .A(n12696), .B(n12695), .ZN(
        P2_U3196) );
  OAI22_X1 U14530 ( .A1(n16427), .A2(n14932), .B1(n12857), .B2(n14935), .ZN(
        n12698) );
  XNOR2_X1 U14531 ( .A(n12698), .B(n11130), .ZN(n12846) );
  INV_X1 U14532 ( .A(n12699), .ZN(n14934) );
  OAI22_X1 U14533 ( .A1(n16427), .A2(n14935), .B1(n12857), .B2(n14934), .ZN(
        n12845) );
  XNOR2_X1 U14534 ( .A(n12846), .B(n12845), .ZN(n12706) );
  INV_X1 U14535 ( .A(n12700), .ZN(n12701) );
  AOI21_X1 U14536 ( .B1(n12706), .B2(n12705), .A(n12847), .ZN(n12714) );
  OAI21_X1 U14537 ( .B1(n15036), .B2(n12708), .A(n12707), .ZN(n12711) );
  OAI22_X1 U14538 ( .A1(n12709), .A2(n15038), .B1(n15037), .B2(n12722), .ZN(
        n12710) );
  AOI211_X1 U14539 ( .C1(n12712), .C2(n15042), .A(n12711), .B(n12710), .ZN(
        n12713) );
  OAI21_X1 U14540 ( .B1(n12714), .B2(n15044), .A(n12713), .ZN(P1_U3236) );
  NAND2_X1 U14541 ( .A1(n12716), .A2(n12715), .ZN(n12718) );
  OR2_X1 U14542 ( .A1(n12851), .A2(n12722), .ZN(n12717) );
  NAND2_X1 U14543 ( .A1(n12718), .A2(n12717), .ZN(n12759) );
  XOR2_X1 U14544 ( .A(n12758), .B(n12759), .Z(n12820) );
  OR2_X1 U14545 ( .A1(n12851), .A2(n15049), .ZN(n12719) );
  NAND2_X1 U14546 ( .A1(n12720), .A2(n12719), .ZN(n12753) );
  XNOR2_X1 U14547 ( .A(n12753), .B(n12758), .ZN(n12815) );
  NAND2_X1 U14548 ( .A1(n12815), .A2(n15425), .ZN(n12727) );
  AOI21_X1 U14549 ( .B1(n12967), .B2(n12721), .A(n7541), .ZN(n12817) );
  INV_X1 U14550 ( .A(n15047), .ZN(n15039) );
  OAI22_X1 U14551 ( .A1(n12722), .A2(n15451), .B1(n15039), .B2(n15410), .ZN(
        n12962) );
  OAI22_X1 U14552 ( .A1(n15430), .A2(n12384), .B1(n12965), .B2(n15428), .ZN(
        n12723) );
  AOI21_X1 U14553 ( .B1(n12962), .B2(n15432), .A(n12723), .ZN(n12724) );
  OAI21_X1 U14554 ( .B1(n8179), .B2(n15434), .A(n12724), .ZN(n12725) );
  AOI21_X1 U14555 ( .B1(n12817), .B2(n15463), .A(n12725), .ZN(n12726) );
  OAI211_X1 U14556 ( .C1(n12820), .C2(n15440), .A(n12727), .B(n12726), .ZN(
        P1_U3280) );
  INV_X1 U14557 ( .A(n12728), .ZN(n12732) );
  OAI222_X1 U14558 ( .A1(n7555), .A2(n12730), .B1(n15627), .B2(n12732), .C1(
        P1_U3086), .C2(n12729), .ZN(P1_U3334) );
  OAI222_X1 U14559 ( .A1(n14783), .A2(n12733), .B1(n14780), .B2(n12732), .C1(
        P2_U3088), .C2(n12731), .ZN(P2_U3306) );
  OAI21_X1 U14560 ( .B1(n12735), .B2(n12736), .A(n12734), .ZN(n16450) );
  AOI21_X1 U14561 ( .B1(n12737), .B2(n12736), .A(n14619), .ZN(n12741) );
  AOI22_X1 U14562 ( .A1(n14583), .A2(n14399), .B1(n14401), .B2(n14600), .ZN(
        n12738) );
  OAI21_X1 U14563 ( .B1(n16450), .B2(n14586), .A(n12738), .ZN(n12739) );
  AOI21_X1 U14564 ( .B1(n12741), .B2(n12740), .A(n12739), .ZN(n16459) );
  INV_X1 U14565 ( .A(n12742), .ZN(n12744) );
  INV_X1 U14566 ( .A(n12790), .ZN(n12743) );
  AOI21_X1 U14567 ( .B1(n16462), .B2(n12744), .A(n12743), .ZN(n16451) );
  AOI22_X1 U14568 ( .A1(n16451), .A2(n14734), .B1(n14733), .B2(n16462), .ZN(
        n12745) );
  OAI211_X1 U14569 ( .C1(n16299), .C2(n16450), .A(n16459), .B(n12745), .ZN(
        n12747) );
  NAND2_X1 U14570 ( .A1(n12747), .A2(n16413), .ZN(n12746) );
  OAI21_X1 U14571 ( .B1(n16413), .B2(n11314), .A(n12746), .ZN(P2_U3511) );
  INV_X1 U14572 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U14573 ( .A1(n12747), .A2(n14760), .ZN(n12748) );
  OAI21_X1 U14574 ( .B1(n14760), .B2(n12749), .A(n12748), .ZN(P2_U3466) );
  INV_X1 U14575 ( .A(n12750), .ZN(n12751) );
  OAI222_X1 U14576 ( .A1(n12752), .A2(P3_U3151), .B1(n14237), .B2(n15644), 
        .C1(n13194), .C2(n12751), .ZN(P3_U3270) );
  NAND2_X1 U14577 ( .A1(n12753), .A2(n12758), .ZN(n12755) );
  OR2_X1 U14578 ( .A1(n12967), .A2(n15048), .ZN(n12754) );
  NAND2_X1 U14579 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  NAND2_X1 U14580 ( .A1(n12756), .A2(n12761), .ZN(n12757) );
  NAND2_X1 U14581 ( .A1(n12971), .A2(n12757), .ZN(n15578) );
  NAND2_X1 U14582 ( .A1(n12967), .A2(n14896), .ZN(n12760) );
  OAI21_X1 U14583 ( .B1(n12762), .B2(n12761), .A(n12975), .ZN(n15585) );
  INV_X1 U14584 ( .A(n15579), .ZN(n14902) );
  OR2_X1 U14585 ( .A1(n14902), .A2(n7541), .ZN(n12763) );
  NAND2_X1 U14586 ( .A1(n12977), .A2(n12763), .ZN(n15582) );
  AOI22_X1 U14587 ( .A1(n15175), .A2(n15448), .B1(n15386), .B2(n15048), .ZN(
        n15581) );
  INV_X1 U14588 ( .A(n12764), .ZN(n14899) );
  AOI22_X1 U14589 ( .A1(n15356), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14899), 
        .B2(n15458), .ZN(n12765) );
  OAI21_X1 U14590 ( .B1(n15581), .B2(n15356), .A(n12765), .ZN(n12766) );
  AOI21_X1 U14591 ( .B1(n15579), .B2(n15459), .A(n12766), .ZN(n12767) );
  OAI21_X1 U14592 ( .B1(n15582), .B2(n15398), .A(n12767), .ZN(n12768) );
  AOI21_X1 U14593 ( .B1(n15585), .B2(n15269), .A(n12768), .ZN(n12769) );
  OAI21_X1 U14594 ( .B1(n15578), .B2(n15342), .A(n12769), .ZN(P1_U3279) );
  INV_X1 U14595 ( .A(n12990), .ZN(n12794) );
  AND2_X1 U14596 ( .A1(n14399), .A2(n14305), .ZN(n12771) );
  XNOR2_X1 U14597 ( .A(n12990), .B(n14306), .ZN(n12770) );
  NOR2_X1 U14598 ( .A1(n12770), .A2(n12771), .ZN(n12943) );
  AOI21_X1 U14599 ( .B1(n12771), .B2(n12770), .A(n12943), .ZN(n12775) );
  OAI21_X1 U14600 ( .B1(n12775), .B2(n12774), .A(n12945), .ZN(n12776) );
  NAND2_X1 U14601 ( .A1(n12776), .A2(n14382), .ZN(n12781) );
  INV_X1 U14602 ( .A(n12777), .ZN(n12791) );
  OAI22_X1 U14603 ( .A1(n12783), .A2(n14362), .B1(n14387), .B2(n13064), .ZN(
        n12778) );
  AOI211_X1 U14604 ( .C1(n12791), .C2(n14385), .A(n12779), .B(n12778), .ZN(
        n12780) );
  OAI211_X1 U14605 ( .C1(n12794), .C2(n14393), .A(n12781), .B(n12780), .ZN(
        P2_U3206) );
  XNOR2_X1 U14606 ( .A(n12782), .B(n12784), .ZN(n12989) );
  OAI22_X1 U14607 ( .A1(n13064), .A2(n14623), .B1(n12783), .B2(n14621), .ZN(
        n12788) );
  XNOR2_X1 U14608 ( .A(n12785), .B(n12784), .ZN(n12786) );
  NOR2_X1 U14609 ( .A1(n12786), .A2(n14619), .ZN(n12787) );
  AOI211_X1 U14610 ( .C1(n14522), .C2(n12989), .A(n12788), .B(n12787), .ZN(
        n12993) );
  INV_X1 U14611 ( .A(n12880), .ZN(n12789) );
  AOI21_X1 U14612 ( .B1(n12990), .B2(n12790), .A(n12789), .ZN(n12991) );
  NAND2_X1 U14613 ( .A1(n12991), .A2(n16452), .ZN(n12793) );
  AOI22_X1 U14614 ( .A1(n14598), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12791), 
        .B2(n14611), .ZN(n12792) );
  OAI211_X1 U14615 ( .C1(n12794), .C2(n14631), .A(n12793), .B(n12792), .ZN(
        n12795) );
  AOI21_X1 U14616 ( .B1(n12989), .B2(n16453), .A(n12795), .ZN(n12796) );
  OAI21_X1 U14617 ( .B1(n12993), .B2(n14598), .A(n12796), .ZN(P2_U3252) );
  NOR2_X1 U14618 ( .A1(n12805), .A2(n12797), .ZN(n12799) );
  NOR2_X1 U14619 ( .A1(n12799), .A2(n12798), .ZN(n12803) );
  INV_X1 U14620 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U14621 ( .A1(n12808), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13011) );
  INV_X1 U14622 ( .A(n13011), .ZN(n12800) );
  AOI21_X1 U14623 ( .B1(n12801), .B2(n13016), .A(n12800), .ZN(n12802) );
  NAND2_X1 U14624 ( .A1(n12802), .A2(n12803), .ZN(n13010) );
  OAI211_X1 U14625 ( .C1(n12803), .C2(n12802), .A(n15154), .B(n13010), .ZN(
        n12814) );
  NAND2_X1 U14626 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14965)
         );
  NOR2_X1 U14627 ( .A1(n12805), .A2(n12804), .ZN(n12807) );
  XOR2_X1 U14628 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12808), .Z(n12809) );
  NAND2_X1 U14629 ( .A1(n12809), .A2(n12810), .ZN(n13015) );
  OAI211_X1 U14630 ( .C1(n12810), .C2(n12809), .A(n15155), .B(n13015), .ZN(
        n12811) );
  NAND2_X1 U14631 ( .A1(n14965), .A2(n12811), .ZN(n12812) );
  AOI21_X1 U14632 ( .B1(n16197), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12812), 
        .ZN(n12813) );
  OAI211_X1 U14633 ( .C1(n15149), .C2(n13016), .A(n12814), .B(n12813), .ZN(
        P1_U3259) );
  INV_X1 U14634 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n12822) );
  NAND2_X1 U14635 ( .A1(n12815), .A2(n15568), .ZN(n12819) );
  NOR2_X1 U14636 ( .A1(n8179), .A2(n16437), .ZN(n12816) );
  AOI211_X1 U14637 ( .C1(n12817), .C2(n16326), .A(n12816), .B(n12962), .ZN(
        n12818) );
  OAI211_X1 U14638 ( .C1(n15567), .C2(n12820), .A(n12819), .B(n12818), .ZN(
        n12823) );
  NAND2_X1 U14639 ( .A1(n12823), .A2(n16338), .ZN(n12821) );
  OAI21_X1 U14640 ( .B1(n16338), .B2(n12822), .A(n12821), .ZN(P1_U3498) );
  NAND2_X1 U14641 ( .A1(n12823), .A2(n16446), .ZN(n12824) );
  OAI21_X1 U14642 ( .B1(n16446), .B2(n12825), .A(n12824), .ZN(P1_U3541) );
  MUX2_X1 U14643 ( .A(n9688), .B(P2_REG2_REG_19__SCAN_IN), .S(n14444), .Z(
        n12830) );
  AOI21_X1 U14644 ( .B1(n12832), .B2(P2_REG2_REG_17__SCAN_IN), .A(n12826), 
        .ZN(n12828) );
  XNOR2_X1 U14645 ( .A(n12828), .B(n12827), .ZN(n16162) );
  AOI22_X1 U14646 ( .A1(n16162), .A2(n9664), .B1(n12828), .B2(n16167), .ZN(
        n12829) );
  XOR2_X1 U14647 ( .A(n12830), .B(n12829), .Z(n12842) );
  AOI21_X1 U14648 ( .B1(n12832), .B2(P2_REG1_REG_17__SCAN_IN), .A(n12831), 
        .ZN(n12833) );
  NOR2_X1 U14649 ( .A1(n12833), .A2(n16167), .ZN(n12834) );
  AOI21_X1 U14650 ( .B1(n12833), .B2(n16167), .A(n12834), .ZN(n16165) );
  NAND2_X1 U14651 ( .A1(n16165), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n16164) );
  INV_X1 U14652 ( .A(n12834), .ZN(n12835) );
  NAND2_X1 U14653 ( .A1(n16164), .A2(n12835), .ZN(n12837) );
  XNOR2_X1 U14654 ( .A(n14444), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12836) );
  XNOR2_X1 U14655 ( .A(n12837), .B(n12836), .ZN(n12840) );
  AND2_X1 U14656 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14296) );
  AOI21_X1 U14657 ( .B1(n16055), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14296), 
        .ZN(n12838) );
  OAI21_X1 U14658 ( .B1(n14508), .B2(n16168), .A(n12838), .ZN(n12839) );
  AOI21_X1 U14659 ( .B1(n12840), .B2(n16163), .A(n12839), .ZN(n12841) );
  OAI21_X1 U14660 ( .B1(n12842), .B2(n16182), .A(n12841), .ZN(P2_U3233) );
  OAI222_X1 U14661 ( .A1(n14780), .A2(n12844), .B1(n7660), .B2(P2_U3088), .C1(
        n12843), .C2(n14783), .ZN(P2_U3305) );
  INV_X1 U14662 ( .A(n12851), .ZN(n16438) );
  INV_X1 U14663 ( .A(n12845), .ZN(n12849) );
  INV_X1 U14664 ( .A(n12846), .ZN(n12848) );
  AND2_X1 U14665 ( .A1(n15049), .A2(n14817), .ZN(n12850) );
  AOI21_X1 U14666 ( .B1(n12851), .B2(n11694), .A(n12850), .ZN(n12958) );
  AOI22_X1 U14667 ( .A1(n12851), .A2(n11013), .B1(n11694), .B2(n15049), .ZN(
        n12852) );
  XNOR2_X1 U14668 ( .A(n12852), .B(n11130), .ZN(n12957) );
  XOR2_X1 U14669 ( .A(n12958), .B(n12957), .Z(n12853) );
  OAI211_X1 U14670 ( .C1(n12854), .C2(n12853), .A(n12956), .B(n15012), .ZN(
        n12862) );
  INV_X1 U14671 ( .A(n12855), .ZN(n12860) );
  INV_X1 U14672 ( .A(n12856), .ZN(n12859) );
  OAI22_X1 U14673 ( .A1(n12857), .A2(n15038), .B1(n15037), .B2(n14896), .ZN(
        n12858) );
  AOI211_X1 U14674 ( .C1(n12860), .C2(n15017), .A(n12859), .B(n12858), .ZN(
        n12861) );
  OAI211_X1 U14675 ( .C1(n16438), .C2(n15026), .A(n12862), .B(n12861), .ZN(
        P1_U3224) );
  INV_X1 U14676 ( .A(n12863), .ZN(n12864) );
  NAND2_X1 U14677 ( .A1(n12864), .A2(n13661), .ZN(n12865) );
  XNOR2_X1 U14678 ( .A(n7663), .B(n13526), .ZN(n12867) );
  XNOR2_X1 U14679 ( .A(n12867), .B(n13660), .ZN(n13326) );
  INV_X1 U14680 ( .A(n12867), .ZN(n12868) );
  NAND2_X1 U14681 ( .A1(n12868), .A2(n13660), .ZN(n12869) );
  XNOR2_X1 U14682 ( .A(n7663), .B(n13006), .ZN(n13037) );
  XNOR2_X1 U14683 ( .A(n13037), .B(n13659), .ZN(n12871) );
  INV_X1 U14684 ( .A(n12871), .ZN(n12870) );
  NAND2_X1 U14685 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  AOI21_X1 U14686 ( .B1(n13040), .B2(n12873), .A(n13421), .ZN(n12877) );
  AOI22_X1 U14687 ( .A1(n13418), .A2(n16385), .B1(n13660), .B2(n13450), .ZN(
        n12875) );
  NOR2_X1 U14688 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15713), .ZN(n16288) );
  AOI21_X1 U14689 ( .B1(n13134), .B2(n13439), .A(n16288), .ZN(n12874) );
  OAI211_X1 U14690 ( .C1(n13447), .C2(n16381), .A(n12875), .B(n12874), .ZN(
        n12876) );
  OR2_X1 U14691 ( .A1(n12877), .A2(n12876), .ZN(P3_U3171) );
  XNOR2_X1 U14692 ( .A(n12878), .B(n12883), .ZN(n12879) );
  AOI222_X1 U14693 ( .A1(n14399), .A2(n14600), .B1(n14603), .B2(n12879), .C1(
        n14397), .C2(n14583), .ZN(n14737) );
  AOI21_X1 U14694 ( .B1(n14732), .B2(n12880), .A(n13077), .ZN(n14735) );
  INV_X1 U14695 ( .A(n12881), .ZN(n12952) );
  AOI22_X1 U14696 ( .A1(n14598), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12952), 
        .B2(n14611), .ZN(n12882) );
  OAI21_X1 U14697 ( .B1(n12955), .B2(n14631), .A(n12882), .ZN(n12886) );
  XNOR2_X1 U14698 ( .A(n12884), .B(n12883), .ZN(n14738) );
  NOR2_X1 U14699 ( .A1(n14738), .A2(n14638), .ZN(n12885) );
  AOI211_X1 U14700 ( .C1(n14735), .C2(n16452), .A(n12886), .B(n12885), .ZN(
        n12887) );
  OAI21_X1 U14701 ( .B1(n14737), .B2(n14598), .A(n12887), .ZN(P2_U3251) );
  INV_X1 U14702 ( .A(n12888), .ZN(n12890) );
  MUX2_X1 U14703 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13775), .Z(n13108) );
  XOR2_X1 U14704 ( .A(n13111), .B(n13108), .Z(n12892) );
  AOI21_X1 U14705 ( .B1(n12893), .B2(n12892), .A(n13109), .ZN(n12913) );
  AND2_X1 U14706 ( .A1(n12900), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U14707 ( .A1(n12896), .A2(n12909), .ZN(n13116) );
  INV_X1 U14708 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16422) );
  AOI21_X1 U14709 ( .B1(n12897), .B2(n16422), .A(n13117), .ZN(n12898) );
  NOR2_X1 U14710 ( .A1(n12898), .A2(n16285), .ZN(n12911) );
  INV_X1 U14711 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n12899) );
  NOR2_X1 U14712 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12899), .ZN(n13140) );
  AOI21_X1 U14713 ( .B1(n16037), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n13140), 
        .ZN(n12908) );
  NAND2_X1 U14714 ( .A1(n12900), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n12902) );
  NOR2_X1 U14715 ( .A1(n12903), .A2(n12909), .ZN(n12904) );
  AND2_X1 U14716 ( .A1(n12905), .A2(n13051), .ZN(n12906) );
  OAI21_X1 U14717 ( .B1(n13122), .B2(n12906), .A(n13840), .ZN(n12907) );
  OAI211_X1 U14718 ( .C1(n16278), .C2(n12909), .A(n12908), .B(n12907), .ZN(
        n12910) );
  NOR2_X1 U14719 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  OAI21_X1 U14720 ( .B1(n12913), .B2(n16259), .A(n12912), .ZN(P3_U3193) );
  INV_X1 U14721 ( .A(n12914), .ZN(n12915) );
  OAI222_X1 U14722 ( .A1(n12917), .A2(P3_U3151), .B1(n14237), .B2(n12916), 
        .C1(n13194), .C2(n12915), .ZN(P3_U3269) );
  OAI21_X1 U14723 ( .B1(n13630), .B2(n12919), .A(n12918), .ZN(n12926) );
  INV_X1 U14724 ( .A(n13659), .ZN(n14093) );
  OAI22_X1 U14725 ( .A1(n12920), .A2(n14092), .B1(n14093), .B2(n14090), .ZN(
        n12925) );
  OR2_X1 U14726 ( .A1(n12921), .A2(n13523), .ZN(n12922) );
  NOR2_X1 U14727 ( .A1(n12930), .A2(n14097), .ZN(n12924) );
  AOI211_X1 U14728 ( .C1(n16309), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        n12940) );
  OAI22_X1 U14729 ( .A1(n14075), .A2(n13527), .B1(n13329), .B2(n16339), .ZN(
        n12928) );
  NOR2_X1 U14730 ( .A1(n12930), .A2(n14104), .ZN(n12927) );
  AOI211_X1 U14731 ( .C1(n16348), .C2(P3_REG2_REG_8__SCAN_IN), .A(n12928), .B(
        n12927), .ZN(n12929) );
  OAI21_X1 U14732 ( .B1(n12940), .B2(n16348), .A(n12929), .ZN(P3_U3225) );
  INV_X1 U14733 ( .A(n12930), .ZN(n12938) );
  INV_X1 U14734 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12931) );
  OAI22_X1 U14735 ( .A1(n14164), .A2(n13527), .B1(n16473), .B2(n12931), .ZN(
        n12932) );
  AOI21_X1 U14736 ( .B1(n12938), .B2(n12933), .A(n12932), .ZN(n12934) );
  OAI21_X1 U14737 ( .B1(n12940), .B2(n10822), .A(n12934), .ZN(P3_U3467) );
  OAI22_X1 U14738 ( .A1(n14221), .A2(n13527), .B1(n16476), .B2(n12935), .ZN(
        n12936) );
  AOI21_X1 U14739 ( .B1(n12938), .B2(n12937), .A(n12936), .ZN(n12939) );
  OAI21_X1 U14740 ( .B1(n12940), .B2(n16483), .A(n12939), .ZN(P3_U3414) );
  AND2_X1 U14741 ( .A1(n14398), .A2(n14305), .ZN(n12942) );
  XNOR2_X1 U14742 ( .A(n14732), .B(n14306), .ZN(n12941) );
  NOR2_X1 U14743 ( .A1(n12941), .A2(n12942), .ZN(n13057) );
  AOI21_X1 U14744 ( .B1(n12942), .B2(n12941), .A(n13057), .ZN(n12947) );
  INV_X1 U14745 ( .A(n12943), .ZN(n12944) );
  OAI21_X1 U14746 ( .B1(n12947), .B2(n12946), .A(n13059), .ZN(n12948) );
  NAND2_X1 U14747 ( .A1(n12948), .A2(n14382), .ZN(n12954) );
  NAND2_X1 U14748 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n16159)
         );
  INV_X1 U14749 ( .A(n16159), .ZN(n12951) );
  OAI22_X1 U14750 ( .A1(n12949), .A2(n14362), .B1(n14387), .B2(n13157), .ZN(
        n12950) );
  AOI211_X1 U14751 ( .C1(n12952), .C2(n14385), .A(n12951), .B(n12950), .ZN(
        n12953) );
  OAI211_X1 U14752 ( .C1(n12955), .C2(n14393), .A(n12954), .B(n12953), .ZN(
        P2_U3187) );
  NAND2_X1 U14753 ( .A1(n12967), .A2(n11013), .ZN(n12960) );
  NAND2_X1 U14754 ( .A1(n15048), .A2(n14831), .ZN(n12959) );
  NAND2_X1 U14755 ( .A1(n12960), .A2(n12959), .ZN(n12961) );
  XNOR2_X1 U14756 ( .A(n12961), .B(n11130), .ZN(n14800) );
  AOI22_X1 U14757 ( .A1(n12967), .A2(n14831), .B1(n14817), .B2(n15048), .ZN(
        n14799) );
  XNOR2_X1 U14758 ( .A(n14800), .B(n14799), .ZN(n14802) );
  XNOR2_X1 U14759 ( .A(n14803), .B(n14802), .ZN(n12969) );
  NAND2_X1 U14760 ( .A1(n12962), .A2(n15029), .ZN(n12964) );
  OAI211_X1 U14761 ( .C1(n15036), .C2(n12965), .A(n12964), .B(n12963), .ZN(
        n12966) );
  AOI21_X1 U14762 ( .B1(n12967), .B2(n15042), .A(n12966), .ZN(n12968) );
  OAI21_X1 U14763 ( .B1(n12969), .B2(n15044), .A(n12968), .ZN(P1_U3234) );
  NAND2_X1 U14764 ( .A1(n15579), .A2(n15047), .ZN(n12970) );
  INV_X1 U14765 ( .A(n15187), .ZN(n12976) );
  NAND2_X1 U14766 ( .A1(n12972), .A2(n12976), .ZN(n12973) );
  NAND2_X1 U14767 ( .A1(n15176), .A2(n12973), .ZN(n15569) );
  INV_X1 U14768 ( .A(n15569), .ZN(n12988) );
  NAND2_X1 U14769 ( .A1(n15579), .A2(n15039), .ZN(n12974) );
  XNOR2_X1 U14770 ( .A(n15188), .B(n12976), .ZN(n15575) );
  AOI21_X1 U14771 ( .B1(n12977), .B2(n15571), .A(n16428), .ZN(n12978) );
  OR2_X2 U14772 ( .A1(n12977), .A2(n15571), .ZN(n15427) );
  NAND2_X1 U14773 ( .A1(n12978), .A2(n15427), .ZN(n15573) );
  NAND2_X1 U14774 ( .A1(n15177), .A2(n15448), .ZN(n12980) );
  NAND2_X1 U14775 ( .A1(n15047), .A2(n15386), .ZN(n12979) );
  NAND2_X1 U14776 ( .A1(n12980), .A2(n12979), .ZN(n15570) );
  NOR2_X1 U14777 ( .A1(n15035), .A2(n15428), .ZN(n12981) );
  OAI21_X1 U14778 ( .B1(n15570), .B2(n12981), .A(n15430), .ZN(n12982) );
  OAI21_X1 U14779 ( .B1(n15430), .B2(n12983), .A(n12982), .ZN(n12984) );
  AOI21_X1 U14780 ( .B1(n15571), .B2(n15459), .A(n12984), .ZN(n12985) );
  OAI21_X1 U14781 ( .B1(n15573), .B2(n15168), .A(n12985), .ZN(n12986) );
  AOI21_X1 U14782 ( .B1(n15575), .B2(n15269), .A(n12986), .ZN(n12987) );
  OAI21_X1 U14783 ( .B1(n12988), .B2(n15342), .A(n12987), .ZN(P1_U3278) );
  INV_X1 U14784 ( .A(n12989), .ZN(n12994) );
  AOI22_X1 U14785 ( .A1(n12991), .A2(n14734), .B1(n14733), .B2(n12990), .ZN(
        n12992) );
  OAI211_X1 U14786 ( .C1(n12994), .C2(n16299), .A(n12993), .B(n12992), .ZN(
        n12997) );
  NAND2_X1 U14787 ( .A1(n12997), .A2(n16413), .ZN(n12995) );
  OAI21_X1 U14788 ( .B1(n16413), .B2(n12996), .A(n12995), .ZN(P2_U3512) );
  NAND2_X1 U14789 ( .A1(n12997), .A2(n14760), .ZN(n12998) );
  OAI21_X1 U14790 ( .B1(n14760), .B2(n9584), .A(n12998), .ZN(P2_U3469) );
  OR2_X1 U14791 ( .A1(n7942), .A2(n13534), .ZN(n13525) );
  XNOR2_X1 U14792 ( .A(n13000), .B(n13525), .ZN(n16379) );
  XNOR2_X1 U14793 ( .A(n13001), .B(n13525), .ZN(n13002) );
  AOI222_X1 U14794 ( .A1(n16309), .A2(n13002), .B1(n13134), .B2(n16313), .C1(
        n13660), .C2(n16311), .ZN(n16378) );
  OAI21_X1 U14795 ( .B1(n14150), .B2(n16379), .A(n16378), .ZN(n13008) );
  OAI22_X1 U14796 ( .A1(n14164), .A2(n13006), .B1(n16473), .B2(n16270), .ZN(
        n13003) );
  AOI21_X1 U14797 ( .B1(n13008), .B2(n16473), .A(n13003), .ZN(n13004) );
  INV_X1 U14798 ( .A(n13004), .ZN(P3_U3468) );
  INV_X1 U14799 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n13005) );
  OAI22_X1 U14800 ( .A1(n14221), .A2(n13006), .B1(n16476), .B2(n13005), .ZN(
        n13007) );
  AOI21_X1 U14801 ( .B1(n13008), .B2(n16476), .A(n13007), .ZN(n13009) );
  INV_X1 U14802 ( .A(n13009), .ZN(P3_U3417) );
  NAND2_X1 U14803 ( .A1(n13011), .A2(n13010), .ZN(n13014) );
  INV_X1 U14804 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U14805 ( .A1(n15130), .A2(n15127), .ZN(n13012) );
  AOI21_X1 U14806 ( .B1(n15127), .B2(n15130), .A(n13012), .ZN(n13013) );
  NAND2_X1 U14807 ( .A1(n13013), .A2(n13014), .ZN(n15126) );
  OAI211_X1 U14808 ( .C1(n13014), .C2(n13013), .A(n15154), .B(n15126), .ZN(
        n13023) );
  NAND2_X1 U14809 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14976)
         );
  XNOR2_X1 U14810 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15130), .ZN(n13019) );
  INV_X1 U14811 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n13017) );
  OAI21_X1 U14812 ( .B1(n13017), .B2(n13016), .A(n13015), .ZN(n13018) );
  NAND2_X1 U14813 ( .A1(n13019), .A2(n13018), .ZN(n15129) );
  OAI211_X1 U14814 ( .C1(n13019), .C2(n13018), .A(n15155), .B(n15129), .ZN(
        n13020) );
  NAND2_X1 U14815 ( .A1(n14976), .A2(n13020), .ZN(n13021) );
  AOI21_X1 U14816 ( .B1(n16197), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n13021), 
        .ZN(n13022) );
  OAI211_X1 U14817 ( .C1(n15149), .C2(n15130), .A(n13023), .B(n13022), .ZN(
        P1_U3260) );
  INV_X1 U14818 ( .A(n13028), .ZN(n13027) );
  AOI21_X1 U14819 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13025), .A(n13024), 
        .ZN(n13026) );
  OAI21_X1 U14820 ( .B1(n13027), .B2(n14780), .A(n13026), .ZN(P2_U3304) );
  NAND2_X1 U14821 ( .A1(n13028), .A2(n15612), .ZN(n13030) );
  OAI211_X1 U14822 ( .C1(n13031), .C2(n7555), .A(n13030), .B(n13029), .ZN(
        P1_U3332) );
  INV_X1 U14823 ( .A(n13032), .ZN(n13036) );
  OAI222_X1 U14824 ( .A1(n7555), .A2(n13034), .B1(n15627), .B2(n13036), .C1(
        P1_U3086), .C2(n13033), .ZN(P1_U3331) );
  OAI222_X1 U14825 ( .A1(n14783), .A2(n7633), .B1(n14780), .B2(n13036), .C1(
        P2_U3088), .C2(n13035), .ZN(P2_U3303) );
  INV_X1 U14826 ( .A(n13037), .ZN(n13038) );
  NAND2_X1 U14827 ( .A1(n13038), .A2(n14093), .ZN(n13039) );
  XNOR2_X1 U14828 ( .A(n7663), .B(n14101), .ZN(n13133) );
  XNOR2_X1 U14829 ( .A(n13133), .B(n13134), .ZN(n13041) );
  NAND2_X1 U14830 ( .A1(n13042), .A2(n13041), .ZN(n13221) );
  OAI211_X1 U14831 ( .C1(n13042), .C2(n13041), .A(n13136), .B(n13442), .ZN(
        n13047) );
  NAND2_X1 U14832 ( .A1(n13659), .A2(n13450), .ZN(n13043) );
  OAI211_X1 U14833 ( .C1(n14091), .C2(n13446), .A(n13044), .B(n13043), .ZN(
        n13045) );
  AOI21_X1 U14834 ( .B1(n14101), .B2(n13418), .A(n13045), .ZN(n13046) );
  OAI211_X1 U14835 ( .C1(n14098), .C2(n13447), .A(n13047), .B(n13046), .ZN(
        P3_U3157) );
  XNOR2_X1 U14836 ( .A(n13048), .B(n13632), .ZN(n13049) );
  AOI222_X1 U14837 ( .A1(n16309), .A2(n13049), .B1(n13658), .B2(n16313), .C1(
        n13134), .C2(n16311), .ZN(n16421) );
  XNOR2_X1 U14838 ( .A(n13050), .B(n13632), .ZN(n16419) );
  NOR2_X1 U14839 ( .A1(n14075), .A2(n13147), .ZN(n13053) );
  OAI22_X1 U14840 ( .A1(n16386), .A2(n13051), .B1(n13139), .B2(n16339), .ZN(
        n13052) );
  AOI211_X1 U14841 ( .C1(n16419), .C2(n14039), .A(n13053), .B(n13052), .ZN(
        n13054) );
  OAI21_X1 U14842 ( .B1(n16421), .B2(n16348), .A(n13054), .ZN(P3_U3222) );
  AND2_X1 U14843 ( .A1(n14397), .A2(n14305), .ZN(n13056) );
  XNOR2_X1 U14844 ( .A(n14728), .B(n14306), .ZN(n13055) );
  NOR2_X1 U14845 ( .A1(n13055), .A2(n13056), .ZN(n13150) );
  AOI21_X1 U14846 ( .B1(n13056), .B2(n13055), .A(n13150), .ZN(n13061) );
  INV_X1 U14847 ( .A(n13057), .ZN(n13058) );
  OAI21_X1 U14848 ( .B1(n13061), .B2(n13060), .A(n13151), .ZN(n13062) );
  NAND2_X1 U14849 ( .A1(n13062), .A2(n14382), .ZN(n13068) );
  INV_X1 U14850 ( .A(n13063), .ZN(n13080) );
  OAI22_X1 U14851 ( .A1(n13064), .A2(n14362), .B1(n14387), .B2(n14622), .ZN(
        n13065) );
  AOI211_X1 U14852 ( .C1(n14385), .C2(n13080), .A(n13066), .B(n13065), .ZN(
        n13067) );
  OAI211_X1 U14853 ( .C1(n13082), .C2(n14393), .A(n13068), .B(n13067), .ZN(
        P2_U3213) );
  XNOR2_X1 U14854 ( .A(n7646), .B(n13073), .ZN(n13076) );
  INV_X1 U14855 ( .A(n13070), .ZN(n13071) );
  AOI21_X1 U14856 ( .B1(n13073), .B2(n13072), .A(n13071), .ZN(n14731) );
  AOI22_X1 U14857 ( .A1(n14396), .A2(n14583), .B1(n14600), .B2(n14398), .ZN(
        n13074) );
  OAI21_X1 U14858 ( .B1(n14731), .B2(n14586), .A(n13074), .ZN(n13075) );
  AOI21_X1 U14859 ( .B1(n14603), .B2(n13076), .A(n13075), .ZN(n14730) );
  INV_X1 U14860 ( .A(n13077), .ZN(n13079) );
  INV_X1 U14861 ( .A(n13096), .ZN(n13078) );
  AOI211_X1 U14862 ( .C1(n14728), .C2(n13079), .A(n14692), .B(n13078), .ZN(
        n14727) );
  AOI22_X1 U14863 ( .A1(n14598), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13080), 
        .B2(n14611), .ZN(n13081) );
  OAI21_X1 U14864 ( .B1(n13082), .B2(n14631), .A(n13081), .ZN(n13084) );
  NOR2_X1 U14865 ( .A1(n14731), .A2(n14593), .ZN(n13083) );
  AOI211_X1 U14866 ( .C1(n14727), .C2(n14596), .A(n13084), .B(n13083), .ZN(
        n13085) );
  OAI21_X1 U14867 ( .B1(n14598), .B2(n14730), .A(n13085), .ZN(P2_U3250) );
  XNOR2_X1 U14868 ( .A(n13087), .B(n13086), .ZN(n13093) );
  OAI21_X1 U14869 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(n14722) );
  OR2_X1 U14870 ( .A1(n14722), .A2(n14586), .ZN(n13092) );
  AOI22_X1 U14871 ( .A1(n14601), .A2(n14604), .B1(n14600), .B2(n14397), .ZN(
        n13091) );
  OAI211_X1 U14872 ( .C1(n14619), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n14724) );
  INV_X1 U14873 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13094) );
  OAI22_X1 U14874 ( .A1(n16458), .A2(n13094), .B1(n13155), .B2(n16455), .ZN(
        n13095) );
  AOI21_X1 U14875 ( .B1(n14719), .B2(n16463), .A(n13095), .ZN(n13099) );
  NAND2_X1 U14876 ( .A1(n14719), .A2(n13096), .ZN(n13097) );
  AND2_X1 U14877 ( .A1(n14630), .A2(n13097), .ZN(n14720) );
  NAND2_X1 U14878 ( .A1(n14720), .A2(n16452), .ZN(n13098) );
  OAI211_X1 U14879 ( .C1(n14722), .C2(n14593), .A(n13099), .B(n13098), .ZN(
        n13100) );
  AOI21_X1 U14880 ( .B1(n16458), .B2(n14724), .A(n13100), .ZN(n13101) );
  INV_X1 U14881 ( .A(n13101), .ZN(P2_U3249) );
  INV_X1 U14882 ( .A(n13102), .ZN(n13106) );
  INV_X1 U14883 ( .A(n13103), .ZN(n13104) );
  OAI222_X1 U14884 ( .A1(n7555), .A2(n7719), .B1(n15627), .B2(n13106), .C1(
        P1_U3086), .C2(n13104), .ZN(P1_U3330) );
  OAI222_X1 U14885 ( .A1(n14783), .A2(n13107), .B1(n14780), .B2(n13106), .C1(
        P2_U3088), .C2(n13105), .ZN(P2_U3302) );
  INV_X1 U14886 ( .A(n13108), .ZN(n13110) );
  XOR2_X1 U14887 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n13694), .Z(n13124) );
  INV_X1 U14888 ( .A(n13124), .ZN(n13113) );
  XOR2_X1 U14889 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n13694), .Z(n13120) );
  INV_X1 U14890 ( .A(n13120), .ZN(n13112) );
  MUX2_X1 U14891 ( .A(n13113), .B(n13112), .S(n13775), .Z(n13114) );
  OAI211_X1 U14892 ( .C1(n13115), .C2(n13114), .A(n13692), .B(n16272), .ZN(
        n13132) );
  INV_X1 U14893 ( .A(n13116), .ZN(n13118) );
  AOI21_X1 U14894 ( .B1(n13120), .B2(n13119), .A(n13700), .ZN(n13121) );
  NOR2_X1 U14895 ( .A1(n16285), .A2(n13121), .ZN(n13130) );
  AOI21_X1 U14896 ( .B1(n13124), .B2(n13123), .A(n7540), .ZN(n13125) );
  NOR2_X1 U14897 ( .A1(n16280), .A2(n13125), .ZN(n13129) );
  INV_X1 U14898 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13126) );
  NOR2_X1 U14899 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13126), .ZN(n13349) );
  NOR2_X1 U14900 ( .A1(n16292), .A2(n13127), .ZN(n13128) );
  NOR4_X1 U14901 ( .A1(n13130), .A2(n13129), .A3(n13349), .A4(n13128), .ZN(
        n13131) );
  OAI211_X1 U14902 ( .C1(n16278), .C2(n13701), .A(n13132), .B(n13131), .ZN(
        P3_U3194) );
  INV_X1 U14903 ( .A(n13133), .ZN(n13135) );
  NAND2_X1 U14904 ( .A1(n13135), .A2(n13134), .ZN(n13211) );
  NAND2_X1 U14905 ( .A1(n13136), .A2(n13211), .ZN(n13138) );
  XNOR2_X1 U14906 ( .A(n13137), .B(n13309), .ZN(n13213) );
  NAND2_X1 U14907 ( .A1(n13138), .A2(n13213), .ZN(n13346) );
  OAI211_X1 U14908 ( .C1(n13138), .C2(n13213), .A(n13346), .B(n13442), .ZN(
        n13146) );
  INV_X1 U14909 ( .A(n13139), .ZN(n13144) );
  AOI21_X1 U14910 ( .B1(n13658), .B2(n13439), .A(n13140), .ZN(n13141) );
  OAI21_X1 U14911 ( .B1(n13142), .B2(n13406), .A(n13141), .ZN(n13143) );
  AOI21_X1 U14912 ( .B1(n13144), .B2(n13414), .A(n13143), .ZN(n13145) );
  OAI211_X1 U14913 ( .C1(n13453), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        P3_U3176) );
  AND2_X1 U14914 ( .A1(n14396), .A2(n14305), .ZN(n13149) );
  XNOR2_X1 U14915 ( .A(n14719), .B(n14306), .ZN(n13148) );
  NOR2_X1 U14916 ( .A1(n13148), .A2(n13149), .ZN(n14243) );
  AOI21_X1 U14917 ( .B1(n13149), .B2(n13148), .A(n14243), .ZN(n13153) );
  OAI21_X1 U14918 ( .B1(n13153), .B2(n13152), .A(n14245), .ZN(n13154) );
  NAND2_X1 U14919 ( .A1(n13154), .A2(n14382), .ZN(n13162) );
  INV_X1 U14920 ( .A(n13155), .ZN(n13160) );
  OAI22_X1 U14921 ( .A1(n13157), .A2(n14362), .B1(n14387), .B2(n13156), .ZN(
        n13158) );
  AOI211_X1 U14922 ( .C1(n14385), .C2(n13160), .A(n13159), .B(n13158), .ZN(
        n13161) );
  OAI211_X1 U14923 ( .C1(n13163), .C2(n14393), .A(n13162), .B(n13161), .ZN(
        P2_U3198) );
  MUX2_X1 U14924 ( .A(n13164), .B(P2_REG2_REG_7__SCAN_IN), .S(n14598), .Z(
        n13173) );
  NOR2_X1 U14925 ( .A1(n13165), .A2(n14561), .ZN(n13169) );
  OAI22_X1 U14926 ( .A1(n14631), .A2(n13167), .B1(n13166), .B2(n16455), .ZN(
        n13168) );
  NOR2_X1 U14927 ( .A1(n13169), .A2(n13168), .ZN(n13170) );
  OAI21_X1 U14928 ( .B1(n13171), .B2(n14593), .A(n13170), .ZN(n13172) );
  OR2_X1 U14929 ( .A1(n13173), .A2(n13172), .ZN(P2_U3258) );
  OAI222_X1 U14930 ( .A1(n14780), .A2(n13176), .B1(n13175), .B2(P2_U3088), 
        .C1(n13174), .C2(n14783), .ZN(P2_U3307) );
  NAND2_X1 U14931 ( .A1(n13178), .A2(P3_D_REG_0__SCAN_IN), .ZN(n13177) );
  OAI21_X1 U14932 ( .B1(n13179), .B2(n13178), .A(n13177), .ZN(P3_U3376) );
  INV_X1 U14933 ( .A(n14772), .ZN(n13180) );
  INV_X1 U14934 ( .A(n13181), .ZN(n13182) );
  OAI222_X1 U14935 ( .A1(n14783), .A2(n13456), .B1(n13184), .B2(P2_U3088), 
        .C1(n14780), .C2(n15618), .ZN(P2_U3297) );
  AOI22_X1 U14936 ( .A1(n13849), .A2(n16382), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n16348), .ZN(n13187) );
  OAI21_X1 U14937 ( .B1(n13188), .B2(n14075), .A(n13187), .ZN(n13189) );
  AOI21_X1 U14938 ( .B1(n13186), .B2(n14039), .A(n13189), .ZN(n13190) );
  OAI21_X1 U14939 ( .B1(n13185), .B2(n16348), .A(n13190), .ZN(P3_U3204) );
  AOI22_X1 U14940 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n15619), .B1(n13192), 
        .B2(n13191), .ZN(n13193) );
  AOI22_X1 U14941 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13456), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15617), .ZN(n13455) );
  INV_X1 U14942 ( .A(SI_30_), .ZN(n13463) );
  OAI222_X1 U14943 ( .A1(n8523), .A2(P3_U3151), .B1(n13194), .B2(n13461), .C1(
        n13463), .C2(n14237), .ZN(P3_U3265) );
  OAI21_X1 U14944 ( .B1(n13197), .B2(n13196), .A(n13195), .ZN(n13198) );
  NAND2_X1 U14945 ( .A1(n13198), .A2(n13442), .ZN(n13204) );
  INV_X1 U14946 ( .A(n16312), .ZN(n13199) );
  OAI22_X1 U14947 ( .A1(n13200), .A2(n13446), .B1(n13199), .B2(n13406), .ZN(
        n13201) );
  AOI21_X1 U14948 ( .B1(n13418), .B2(n7952), .A(n13201), .ZN(n13203) );
  OAI211_X1 U14949 ( .C1(n13205), .C2(n16325), .A(n13204), .B(n13203), .ZN(
        P3_U3162) );
  XNOR2_X1 U14950 ( .A(n13874), .B(n13309), .ZN(n13317) );
  NOR2_X1 U14951 ( .A1(n13317), .A2(n13879), .ZN(n13312) );
  AOI21_X1 U14952 ( .B1(n13317), .B2(n13879), .A(n13312), .ZN(n13274) );
  NAND2_X1 U14953 ( .A1(n14058), .A2(n13309), .ZN(n13215) );
  OR2_X1 U14954 ( .A1(n13206), .A2(n13215), .ZN(n13208) );
  OR2_X1 U14955 ( .A1(n14076), .A2(n13309), .ZN(n13207) );
  AND2_X1 U14956 ( .A1(n13208), .A2(n13207), .ZN(n13348) );
  INV_X1 U14957 ( .A(n13348), .ZN(n13210) );
  INV_X1 U14958 ( .A(n13213), .ZN(n13209) );
  NAND2_X1 U14959 ( .A1(n13209), .A2(n14079), .ZN(n13345) );
  AND2_X1 U14960 ( .A1(n13210), .A2(n13345), .ZN(n13212) );
  AND2_X1 U14961 ( .A1(n13211), .A2(n13212), .ZN(n13220) );
  INV_X1 U14962 ( .A(n13212), .ZN(n13214) );
  INV_X1 U14963 ( .A(n13548), .ZN(n13216) );
  OAI21_X1 U14964 ( .B1(n13216), .B2(n13309), .A(n13215), .ZN(n13217) );
  XNOR2_X1 U14965 ( .A(n16466), .B(n13309), .ZN(n13222) );
  XNOR2_X1 U14966 ( .A(n13222), .B(n14078), .ZN(n13403) );
  INV_X1 U14967 ( .A(n13222), .ZN(n13223) );
  NAND2_X1 U14968 ( .A1(n13223), .A2(n14078), .ZN(n13224) );
  XNOR2_X1 U14969 ( .A(n14219), .B(n13309), .ZN(n13225) );
  XNOR2_X1 U14970 ( .A(n13225), .B(n14031), .ZN(n13284) );
  INV_X1 U14971 ( .A(n13225), .ZN(n13226) );
  NAND2_X1 U14972 ( .A1(n13226), .A2(n14031), .ZN(n13368) );
  XNOR2_X1 U14973 ( .A(n14026), .B(n7663), .ZN(n13233) );
  XNOR2_X1 U14974 ( .A(n13233), .B(n14032), .ZN(n13372) );
  INV_X1 U14975 ( .A(n13372), .ZN(n13228) );
  XNOR2_X1 U14976 ( .A(n14159), .B(n13309), .ZN(n13230) );
  INV_X1 U14977 ( .A(n13230), .ZN(n13227) );
  NAND2_X1 U14978 ( .A1(n13227), .A2(n14046), .ZN(n13370) );
  OR2_X1 U14979 ( .A1(n13228), .A2(n13370), .ZN(n13229) );
  INV_X1 U14980 ( .A(n13229), .ZN(n13232) );
  XNOR2_X1 U14981 ( .A(n13230), .B(n14046), .ZN(n13444) );
  AND2_X1 U14982 ( .A1(n13444), .A2(n13372), .ZN(n13231) );
  INV_X1 U14983 ( .A(n13233), .ZN(n13234) );
  NAND2_X1 U14984 ( .A1(n13234), .A2(n14032), .ZN(n13235) );
  NAND2_X1 U14985 ( .A1(n13371), .A2(n13235), .ZN(n13381) );
  XNOR2_X1 U14986 ( .A(n14211), .B(n13309), .ZN(n13236) );
  XNOR2_X1 U14987 ( .A(n13236), .B(n14020), .ZN(n13380) );
  NAND2_X1 U14988 ( .A1(n13381), .A2(n13380), .ZN(n13379) );
  INV_X1 U14989 ( .A(n13236), .ZN(n13237) );
  NAND2_X1 U14990 ( .A1(n13237), .A2(n14020), .ZN(n13238) );
  NAND2_X1 U14991 ( .A1(n13379), .A2(n13238), .ZN(n13425) );
  XNOR2_X1 U14992 ( .A(n14141), .B(n7663), .ZN(n13239) );
  XNOR2_X1 U14993 ( .A(n13239), .B(n13981), .ZN(n13424) );
  INV_X1 U14994 ( .A(n13239), .ZN(n13240) );
  NAND2_X1 U14995 ( .A1(n13240), .A2(n13981), .ZN(n13241) );
  XNOR2_X1 U14996 ( .A(n13987), .B(n13309), .ZN(n13242) );
  XNOR2_X1 U14997 ( .A(n13242), .B(n13993), .ZN(n13303) );
  INV_X1 U14998 ( .A(n13242), .ZN(n13243) );
  NAND2_X1 U14999 ( .A1(n13243), .A2(n13426), .ZN(n13244) );
  NAND2_X1 U15000 ( .A1(n13300), .A2(n13244), .ZN(n13395) );
  INV_X1 U15001 ( .A(n13395), .ZN(n13246) );
  XNOR2_X1 U15002 ( .A(n13972), .B(n13309), .ZN(n13247) );
  XNOR2_X1 U15003 ( .A(n13247), .B(n13980), .ZN(n13394) );
  INV_X1 U15004 ( .A(n13394), .ZN(n13245) );
  NAND2_X1 U15005 ( .A1(n13247), .A2(n13980), .ZN(n13248) );
  INV_X1 U15006 ( .A(n13337), .ZN(n13251) );
  MUX2_X1 U15007 ( .A(n13476), .B(n13249), .S(n13309), .Z(n13335) );
  INV_X1 U15008 ( .A(n13335), .ZN(n13250) );
  MUX2_X1 U15009 ( .A(n13577), .B(n13252), .S(n13309), .Z(n13334) );
  INV_X1 U15010 ( .A(n13334), .ZN(n13253) );
  XNOR2_X1 U15011 ( .A(n13419), .B(n7663), .ZN(n13255) );
  XNOR2_X1 U15012 ( .A(n13257), .B(n13309), .ZN(n13258) );
  XNOR2_X1 U15013 ( .A(n14120), .B(n13309), .ZN(n13261) );
  NAND2_X1 U15014 ( .A1(n13261), .A2(n13921), .ZN(n13264) );
  INV_X1 U15015 ( .A(n13261), .ZN(n13262) );
  NAND2_X1 U15016 ( .A1(n13262), .A2(n13895), .ZN(n13263) );
  NAND2_X1 U15017 ( .A1(n13264), .A2(n13263), .ZN(n13386) );
  INV_X1 U15018 ( .A(n13264), .ZN(n13360) );
  XNOR2_X1 U15019 ( .A(n13356), .B(n7663), .ZN(n13266) );
  NAND2_X1 U15020 ( .A1(n13266), .A2(n13911), .ZN(n13269) );
  INV_X1 U15021 ( .A(n13266), .ZN(n13267) );
  NAND2_X1 U15022 ( .A1(n13267), .A2(n13880), .ZN(n13268) );
  XNOR2_X1 U15023 ( .A(n13887), .B(n13309), .ZN(n13270) );
  NOR2_X1 U15024 ( .A1(n13270), .A2(n13896), .ZN(n13271) );
  AOI21_X1 U15025 ( .B1(n13270), .B2(n13896), .A(n13271), .ZN(n13434) );
  INV_X1 U15026 ( .A(n13271), .ZN(n13272) );
  NAND2_X1 U15027 ( .A1(n13432), .A2(n13272), .ZN(n13273) );
  INV_X1 U15028 ( .A(n13873), .ZN(n13277) );
  AOI22_X1 U15029 ( .A1(n13896), .A2(n13450), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13276) );
  OAI21_X1 U15030 ( .B1(n13277), .B2(n13447), .A(n13276), .ZN(n13278) );
  AOI21_X1 U15031 ( .B1(n13656), .B2(n13439), .A(n13278), .ZN(n13279) );
  INV_X1 U15032 ( .A(n13281), .ZN(n13282) );
  OAI222_X1 U15033 ( .A1(P3_U3151), .A2(n13775), .B1(n14237), .B2(n13283), 
        .C1(n13194), .C2(n13282), .ZN(P3_U3268) );
  OAI211_X1 U15034 ( .C1(n13285), .C2(n13284), .A(n13369), .B(n13442), .ZN(
        n13292) );
  INV_X1 U15035 ( .A(n13286), .ZN(n14049) );
  INV_X1 U15036 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13287) );
  NOR2_X1 U15037 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13287), .ZN(n13727) );
  AOI21_X1 U15038 ( .B1(n14046), .B2(n13439), .A(n13727), .ZN(n13288) );
  OAI21_X1 U15039 ( .B1(n13289), .B2(n13406), .A(n13288), .ZN(n13290) );
  AOI21_X1 U15040 ( .B1(n14049), .B2(n13414), .A(n13290), .ZN(n13291) );
  OAI211_X1 U15041 ( .C1(n13453), .C2(n14219), .A(n13292), .B(n13291), .ZN(
        P3_U3155) );
  OAI21_X1 U15042 ( .B1(n13936), .B2(n13294), .A(n13293), .ZN(n13295) );
  NAND2_X1 U15043 ( .A1(n13295), .A2(n13442), .ZN(n13299) );
  AOI22_X1 U15044 ( .A1(n13657), .A2(n13450), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13296) );
  OAI21_X1 U15045 ( .B1(n13921), .B2(n13446), .A(n13296), .ZN(n13297) );
  AOI21_X1 U15046 ( .B1(n13928), .B2(n13414), .A(n13297), .ZN(n13298) );
  OAI211_X1 U15047 ( .C1(n14189), .C2(n13453), .A(n13299), .B(n13298), .ZN(
        P3_U3156) );
  INV_X1 U15048 ( .A(n13300), .ZN(n13301) );
  AOI21_X1 U15049 ( .B1(n13303), .B2(n13302), .A(n13301), .ZN(n13308) );
  NAND2_X1 U15050 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13836)
         );
  OAI21_X1 U15051 ( .B1(n13950), .B2(n13446), .A(n13836), .ZN(n13304) );
  AOI21_X1 U15052 ( .B1(n13450), .B2(n13981), .A(n13304), .ZN(n13305) );
  OAI21_X1 U15053 ( .B1(n13984), .B2(n13447), .A(n13305), .ZN(n13306) );
  AOI21_X1 U15054 ( .B1(n13987), .B2(n13418), .A(n13306), .ZN(n13307) );
  OAI21_X1 U15055 ( .B1(n13308), .B2(n13421), .A(n13307), .ZN(P3_U3159) );
  XNOR2_X1 U15056 ( .A(n13656), .B(n13309), .ZN(n13310) );
  XNOR2_X1 U15057 ( .A(n13866), .B(n13310), .ZN(n13318) );
  INV_X1 U15058 ( .A(n13318), .ZN(n13311) );
  NAND2_X1 U15059 ( .A1(n13311), .A2(n13442), .ZN(n13324) );
  INV_X1 U15060 ( .A(n13312), .ZN(n13313) );
  NAND4_X1 U15061 ( .A1(n13323), .A2(n13442), .A3(n13318), .A4(n13313), .ZN(
        n13322) );
  AOI22_X1 U15062 ( .A1(n13867), .A2(n13414), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13315) );
  NAND2_X1 U15063 ( .A1(n13860), .A2(n13439), .ZN(n13314) );
  OAI211_X1 U15064 ( .C1(n13316), .C2(n13406), .A(n13315), .B(n13314), .ZN(
        n13320) );
  NOR4_X1 U15065 ( .A1(n13318), .A2(n13317), .A3(n13879), .A4(n13421), .ZN(
        n13319) );
  AOI211_X1 U15066 ( .C1(n13418), .C2(n13866), .A(n13320), .B(n13319), .ZN(
        n13321) );
  OAI211_X1 U15067 ( .C1(n13324), .C2(n13323), .A(n13322), .B(n13321), .ZN(
        P3_U3160) );
  OAI211_X1 U15068 ( .C1(n13327), .C2(n13326), .A(n13325), .B(n13442), .ZN(
        n13333) );
  AOI21_X1 U15069 ( .B1(n13659), .B2(n13439), .A(n13328), .ZN(n13332) );
  AOI22_X1 U15070 ( .A1(n13418), .A2(n13526), .B1(n13661), .B2(n13450), .ZN(
        n13331) );
  OR2_X1 U15071 ( .A1(n13447), .A2(n13329), .ZN(n13330) );
  NAND4_X1 U15072 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        P3_U3161) );
  NOR2_X1 U15073 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  XNOR2_X1 U15074 ( .A(n13337), .B(n13336), .ZN(n13344) );
  INV_X1 U15075 ( .A(n13338), .ZN(n13947) );
  NAND2_X1 U15076 ( .A1(n13657), .A2(n13439), .ZN(n13340) );
  AOI22_X1 U15077 ( .A1(n13980), .A2(n13450), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13339) );
  OAI211_X1 U15078 ( .C1(n13447), .C2(n13947), .A(n13340), .B(n13339), .ZN(
        n13341) );
  AOI21_X1 U15079 ( .B1(n13342), .B2(n13418), .A(n13341), .ZN(n13343) );
  OAI21_X1 U15080 ( .B1(n13344), .B2(n13421), .A(n13343), .ZN(P3_U3163) );
  NAND2_X1 U15081 ( .A1(n13346), .A2(n13345), .ZN(n13347) );
  AOI21_X1 U15082 ( .B1(n13348), .B2(n13347), .A(n7535), .ZN(n13355) );
  AOI21_X1 U15083 ( .B1(n14078), .B2(n13439), .A(n13349), .ZN(n13351) );
  NAND2_X1 U15084 ( .A1(n14079), .A2(n13450), .ZN(n13350) );
  OAI211_X1 U15085 ( .C1(n13447), .C2(n14074), .A(n13351), .B(n13350), .ZN(
        n13352) );
  AOI21_X1 U15086 ( .B1(n13353), .B2(n13418), .A(n13352), .ZN(n13354) );
  OAI21_X1 U15087 ( .B1(n13355), .B2(n13421), .A(n13354), .ZN(P3_U3164) );
  INV_X1 U15088 ( .A(n13357), .ZN(n13362) );
  NOR3_X1 U15089 ( .A1(n13358), .A2(n13360), .A3(n13359), .ZN(n13361) );
  OAI21_X1 U15090 ( .B1(n13362), .B2(n13361), .A(n13442), .ZN(n13367) );
  AOI22_X1 U15091 ( .A1(n13895), .A2(n13450), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13363) );
  OAI21_X1 U15092 ( .B1(n13364), .B2(n13446), .A(n13363), .ZN(n13365) );
  AOI21_X1 U15093 ( .B1(n13903), .B2(n13414), .A(n13365), .ZN(n13366) );
  OAI211_X1 U15094 ( .C1(n14179), .C2(n13453), .A(n13367), .B(n13366), .ZN(
        P3_U3165) );
  INV_X1 U15095 ( .A(n14026), .ZN(n14149) );
  NAND2_X1 U15096 ( .A1(n13369), .A2(n13368), .ZN(n13445) );
  NAND2_X1 U15097 ( .A1(n13445), .A2(n13444), .ZN(n13443) );
  NAND2_X1 U15098 ( .A1(n13443), .A2(n13370), .ZN(n13373) );
  OAI211_X1 U15099 ( .C1(n13373), .C2(n13372), .A(n13371), .B(n13442), .ZN(
        n13378) );
  NAND2_X1 U15100 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13769)
         );
  OAI21_X1 U15101 ( .B1(n13374), .B2(n13446), .A(n13769), .ZN(n13376) );
  NOR2_X1 U15102 ( .A1(n13447), .A2(n14023), .ZN(n13375) );
  AOI211_X1 U15103 ( .C1(n13450), .C2(n14046), .A(n13376), .B(n13375), .ZN(
        n13377) );
  OAI211_X1 U15104 ( .C1(n14149), .C2(n13453), .A(n13378), .B(n13377), .ZN(
        P3_U3166) );
  OAI211_X1 U15105 ( .C1(n13381), .C2(n13380), .A(n13379), .B(n13442), .ZN(
        n13385) );
  NAND2_X1 U15106 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13790)
         );
  OAI21_X1 U15107 ( .B1(n14007), .B2(n13446), .A(n13790), .ZN(n13383) );
  NOR2_X1 U15108 ( .A1(n13447), .A2(n14010), .ZN(n13382) );
  AOI211_X1 U15109 ( .C1(n13450), .C2(n14032), .A(n13383), .B(n13382), .ZN(
        n13384) );
  OAI211_X1 U15110 ( .C1(n13453), .C2(n14211), .A(n13385), .B(n13384), .ZN(
        P3_U3168) );
  AND3_X1 U15111 ( .A1(n13293), .A2(n13387), .A3(n13386), .ZN(n13388) );
  OAI21_X1 U15112 ( .B1(n13358), .B2(n13388), .A(n13442), .ZN(n13393) );
  AOI22_X1 U15113 ( .A1(n13389), .A2(n13450), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13390) );
  OAI21_X1 U15114 ( .B1(n13911), .B2(n13446), .A(n13390), .ZN(n13391) );
  AOI21_X1 U15115 ( .B1(n13916), .B2(n13414), .A(n13391), .ZN(n13392) );
  OAI211_X1 U15116 ( .C1(n13453), .C2(n14120), .A(n13393), .B(n13392), .ZN(
        P3_U3169) );
  AOI21_X1 U15117 ( .B1(n13395), .B2(n13394), .A(n13421), .ZN(n13397) );
  NAND2_X1 U15118 ( .A1(n13397), .A2(n13396), .ZN(n13401) );
  AOI22_X1 U15119 ( .A1(n13967), .A2(n13439), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13398) );
  OAI21_X1 U15120 ( .B1(n13426), .B2(n13406), .A(n13398), .ZN(n13399) );
  AOI21_X1 U15121 ( .B1(n13971), .B2(n13414), .A(n13399), .ZN(n13400) );
  OAI211_X1 U15122 ( .C1(n14200), .C2(n13453), .A(n13401), .B(n13400), .ZN(
        P3_U3173) );
  OAI211_X1 U15123 ( .C1(n13404), .C2(n13403), .A(n13402), .B(n13442), .ZN(
        n13410) );
  INV_X1 U15124 ( .A(n14067), .ZN(n13408) );
  NOR2_X1 U15125 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15914), .ZN(n13706) );
  AOI21_X1 U15126 ( .B1(n14031), .B2(n13439), .A(n13706), .ZN(n13405) );
  OAI21_X1 U15127 ( .B1(n14062), .B2(n13406), .A(n13405), .ZN(n13407) );
  AOI21_X1 U15128 ( .B1(n13408), .B2(n13414), .A(n13407), .ZN(n13409) );
  OAI211_X1 U15129 ( .C1(n13453), .C2(n16466), .A(n13410), .B(n13409), .ZN(
        P3_U3174) );
  INV_X1 U15130 ( .A(n13411), .ZN(n13412) );
  AOI21_X1 U15131 ( .B1(n13657), .B2(n13413), .A(n13412), .ZN(n13422) );
  AOI22_X1 U15132 ( .A1(n13967), .A2(n13450), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13416) );
  NAND2_X1 U15133 ( .A1(n13414), .A2(n13941), .ZN(n13415) );
  OAI211_X1 U15134 ( .C1(n13936), .C2(n13446), .A(n13416), .B(n13415), .ZN(
        n13417) );
  AOI21_X1 U15135 ( .B1(n13419), .B2(n13418), .A(n13417), .ZN(n13420) );
  OAI21_X1 U15136 ( .B1(n13422), .B2(n13421), .A(n13420), .ZN(P3_U3175) );
  INV_X1 U15137 ( .A(n14141), .ZN(n13431) );
  OAI211_X1 U15138 ( .C1(n13425), .C2(n13424), .A(n13423), .B(n13442), .ZN(
        n13430) );
  NAND2_X1 U15139 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13811)
         );
  OAI21_X1 U15140 ( .B1(n13426), .B2(n13446), .A(n13811), .ZN(n13428) );
  NOR2_X1 U15141 ( .A1(n13447), .A2(n13995), .ZN(n13427) );
  AOI211_X1 U15142 ( .C1(n13450), .C2(n14020), .A(n13428), .B(n13427), .ZN(
        n13429) );
  OAI211_X1 U15143 ( .C1(n13431), .C2(n13453), .A(n13430), .B(n13429), .ZN(
        P3_U3178) );
  OAI21_X1 U15144 ( .B1(n13434), .B2(n13433), .A(n13432), .ZN(n13435) );
  NAND2_X1 U15145 ( .A1(n13435), .A2(n13442), .ZN(n13441) );
  INV_X1 U15146 ( .A(n13886), .ZN(n13437) );
  AOI22_X1 U15147 ( .A1(n13880), .A2(n13450), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13436) );
  OAI21_X1 U15148 ( .B1(n13437), .B2(n13447), .A(n13436), .ZN(n13438) );
  AOI21_X1 U15149 ( .B1(n13439), .B2(n13879), .A(n13438), .ZN(n13440) );
  OAI211_X1 U15150 ( .C1(n14175), .C2(n13453), .A(n13441), .B(n13440), .ZN(
        P3_U3180) );
  OAI211_X1 U15151 ( .C1(n13445), .C2(n13444), .A(n13443), .B(n13442), .ZN(
        n13452) );
  NAND2_X1 U15152 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13745)
         );
  OAI21_X1 U15153 ( .B1(n14006), .B2(n13446), .A(n13745), .ZN(n13449) );
  NOR2_X1 U15154 ( .A1(n13447), .A2(n14034), .ZN(n13448) );
  AOI211_X1 U15155 ( .C1(n13450), .C2(n14031), .A(n13449), .B(n13448), .ZN(
        n13451) );
  OAI211_X1 U15156 ( .C1(n13453), .C2(n14159), .A(n13452), .B(n13451), .ZN(
        P3_U3181) );
  AOI22_X1 U15157 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n10136), .B2(n10703), .ZN(n13457) );
  NAND2_X1 U15158 ( .A1(n14230), .A2(n13458), .ZN(n13460) );
  INV_X1 U15159 ( .A(SI_31_), .ZN(n14235) );
  OR2_X1 U15160 ( .A1(n8954), .A2(n14235), .ZN(n13459) );
  OR2_X1 U15161 ( .A1(n8954), .A2(n13463), .ZN(n13464) );
  OR2_X1 U15162 ( .A1(n13465), .A2(n16477), .ZN(n13613) );
  NAND2_X1 U15163 ( .A1(n13613), .A2(n13612), .ZN(n13470) );
  INV_X1 U15164 ( .A(n13608), .ZN(n13468) );
  INV_X1 U15165 ( .A(n13465), .ZN(n13655) );
  OAI211_X1 U15166 ( .C1(n14109), .C2(n13612), .A(n13611), .B(n13639), .ZN(
        n13467) );
  XNOR2_X1 U15167 ( .A(n13471), .B(n13837), .ZN(n13647) );
  INV_X1 U15168 ( .A(n13472), .ZN(n13646) );
  MUX2_X1 U15169 ( .A(n13475), .B(n13922), .S(n13605), .Z(n13583) );
  INV_X1 U15170 ( .A(n13933), .ZN(n13939) );
  NOR2_X1 U15171 ( .A1(n13476), .A2(n13577), .ZN(n13949) );
  INV_X1 U15172 ( .A(n13962), .ZN(n13964) );
  INV_X1 U15173 ( .A(n13480), .ZN(n13478) );
  OAI211_X1 U15174 ( .C1(n13478), .C2(n13477), .A(n13960), .B(n13959), .ZN(
        n13482) );
  NAND3_X1 U15175 ( .A1(n13959), .A2(n14020), .A3(n14211), .ZN(n13479) );
  NAND3_X1 U15176 ( .A1(n13569), .A2(n13480), .A3(n13479), .ZN(n13481) );
  MUX2_X1 U15177 ( .A(n13482), .B(n13481), .S(n13605), .Z(n13571) );
  NAND2_X1 U15178 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  NAND2_X1 U15179 ( .A1(n13486), .A2(n13485), .ZN(n13490) );
  OAI21_X1 U15180 ( .B1(n13490), .B2(n13487), .A(n13598), .ZN(n13488) );
  NAND2_X1 U15181 ( .A1(n13489), .A2(n13488), .ZN(n13493) );
  AOI21_X1 U15182 ( .B1(n13491), .B2(n13490), .A(n13598), .ZN(n13492) );
  AOI21_X1 U15183 ( .B1(n13494), .B2(n13493), .A(n13492), .ZN(n13497) );
  AOI21_X1 U15184 ( .B1(n13505), .B2(n13495), .A(n13605), .ZN(n13496) );
  OAI21_X1 U15185 ( .B1(n13497), .B2(n13496), .A(n13499), .ZN(n13502) );
  NAND2_X1 U15186 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  NAND2_X1 U15187 ( .A1(n13500), .A2(n13605), .ZN(n13501) );
  NAND2_X1 U15188 ( .A1(n13502), .A2(n13501), .ZN(n13504) );
  OAI211_X1 U15189 ( .C1(n13505), .C2(n13598), .A(n13504), .B(n13503), .ZN(
        n13510) );
  MUX2_X1 U15190 ( .A(n13507), .B(n13506), .S(n13605), .Z(n13508) );
  NAND3_X1 U15191 ( .A1(n13510), .A2(n13509), .A3(n13508), .ZN(n13514) );
  MUX2_X1 U15192 ( .A(n13512), .B(n13511), .S(n13598), .Z(n13513) );
  NAND3_X1 U15193 ( .A1(n13514), .A2(n13621), .A3(n13513), .ZN(n13519) );
  MUX2_X1 U15194 ( .A(n13516), .B(n13515), .S(n13605), .Z(n13517) );
  NAND3_X1 U15195 ( .A1(n13519), .A2(n13518), .A3(n13517), .ZN(n13524) );
  MUX2_X1 U15196 ( .A(n13521), .B(n13520), .S(n13598), .Z(n13522) );
  NAND3_X1 U15197 ( .A1(n13524), .A2(n13523), .A3(n13522), .ZN(n13531) );
  NOR2_X1 U15198 ( .A1(n13525), .A2(n14088), .ZN(n13627) );
  NAND2_X1 U15199 ( .A1(n13526), .A2(n13598), .ZN(n13529) );
  NAND2_X1 U15200 ( .A1(n13527), .A2(n13605), .ZN(n13528) );
  MUX2_X1 U15201 ( .A(n13529), .B(n13528), .S(n13660), .Z(n13530) );
  NAND3_X1 U15202 ( .A1(n13531), .A2(n13627), .A3(n13530), .ZN(n13539) );
  OAI21_X1 U15203 ( .B1(n14088), .B2(n7942), .A(n13532), .ZN(n13536) );
  OAI21_X1 U15204 ( .B1(n14088), .B2(n13534), .A(n13533), .ZN(n13535) );
  MUX2_X1 U15205 ( .A(n13536), .B(n13535), .S(n13605), .Z(n13537) );
  AND2_X1 U15206 ( .A1(n13537), .A2(n13632), .ZN(n13538) );
  NAND2_X1 U15207 ( .A1(n13539), .A2(n13538), .ZN(n13547) );
  NAND3_X1 U15208 ( .A1(n13547), .A2(n13548), .A3(n13540), .ZN(n13541) );
  NAND3_X1 U15209 ( .A1(n13541), .A2(n13546), .A3(n13598), .ZN(n13543) );
  AND2_X1 U15210 ( .A1(n13552), .A2(n13542), .ZN(n14061) );
  NAND2_X1 U15211 ( .A1(n13543), .A2(n14061), .ZN(n13545) );
  NAND3_X1 U15212 ( .A1(n16466), .A2(n14078), .A3(n13598), .ZN(n13544) );
  NAND2_X1 U15213 ( .A1(n13545), .A2(n13544), .ZN(n13551) );
  OAI211_X1 U15214 ( .C1(n14091), .C2(n16417), .A(n13547), .B(n13546), .ZN(
        n13549) );
  NAND3_X1 U15215 ( .A1(n13549), .A2(n13605), .A3(n13548), .ZN(n13550) );
  NAND3_X1 U15216 ( .A1(n13551), .A2(n14043), .A3(n13550), .ZN(n13559) );
  NAND2_X1 U15217 ( .A1(n13553), .A2(n13552), .ZN(n13554) );
  NAND2_X1 U15218 ( .A1(n13554), .A2(n13555), .ZN(n13556) );
  MUX2_X1 U15219 ( .A(n13556), .B(n13555), .S(n13598), .Z(n13557) );
  NAND3_X1 U15220 ( .A1(n13559), .A2(n13558), .A3(n13557), .ZN(n13564) );
  MUX2_X1 U15221 ( .A(n13561), .B(n13560), .S(n13605), .Z(n13562) );
  NAND3_X1 U15222 ( .A1(n13564), .A2(n13563), .A3(n13562), .ZN(n13568) );
  MUX2_X1 U15223 ( .A(n13566), .B(n13565), .S(n13605), .Z(n13567) );
  MUX2_X1 U15224 ( .A(n13569), .B(n13960), .S(n13605), .Z(n13570) );
  OAI21_X1 U15225 ( .B1(n13571), .B2(n8498), .A(n13570), .ZN(n13572) );
  NAND2_X1 U15226 ( .A1(n13964), .A2(n13572), .ZN(n13576) );
  MUX2_X1 U15227 ( .A(n13574), .B(n13573), .S(n13605), .Z(n13575) );
  NAND3_X1 U15228 ( .A1(n13949), .A2(n13576), .A3(n13575), .ZN(n13581) );
  INV_X1 U15229 ( .A(n13577), .ZN(n13579) );
  MUX2_X1 U15230 ( .A(n13579), .B(n13578), .S(n13605), .Z(n13580) );
  NAND3_X1 U15231 ( .A1(n13939), .A2(n13581), .A3(n13580), .ZN(n13582) );
  NAND3_X1 U15232 ( .A1(n13583), .A2(n13923), .A3(n13582), .ZN(n13587) );
  MUX2_X1 U15233 ( .A(n13585), .B(n13584), .S(n13598), .Z(n13586) );
  NAND3_X1 U15234 ( .A1(n13910), .A2(n13587), .A3(n13586), .ZN(n13604) );
  NAND2_X1 U15235 ( .A1(n14182), .A2(n13921), .ZN(n13589) );
  MUX2_X1 U15236 ( .A(n13589), .B(n13588), .S(n13598), .Z(n13600) );
  NAND2_X1 U15237 ( .A1(n13591), .A2(n13590), .ZN(n13593) );
  NAND2_X1 U15238 ( .A1(n13593), .A2(n13592), .ZN(n13594) );
  NAND2_X1 U15239 ( .A1(n13595), .A2(n13594), .ZN(n13597) );
  NAND2_X1 U15240 ( .A1(n13597), .A2(n13596), .ZN(n13601) );
  NAND2_X1 U15241 ( .A1(n13601), .A2(n13598), .ZN(n13599) );
  INV_X1 U15242 ( .A(n13601), .ZN(n13602) );
  NAND2_X1 U15243 ( .A1(n13602), .A2(n13605), .ZN(n13603) );
  INV_X1 U15244 ( .A(n13611), .ZN(n13614) );
  INV_X1 U15245 ( .A(n13612), .ZN(n13851) );
  NOR2_X1 U15246 ( .A1(n13620), .A2(n13619), .ZN(n13626) );
  NOR4_X1 U15247 ( .A1(n13624), .A2(n13623), .A3(n8666), .A4(n13622), .ZN(
        n13625) );
  NAND4_X1 U15248 ( .A1(n13628), .A2(n13627), .A3(n13626), .A4(n13625), .ZN(
        n13629) );
  NOR4_X1 U15249 ( .A1(n13630), .A2(n8991), .A3(n14076), .A4(n13629), .ZN(
        n13631) );
  NAND4_X1 U15250 ( .A1(n13632), .A2(n14043), .A3(n14061), .A4(n13631), .ZN(
        n13633) );
  NOR4_X1 U15251 ( .A1(n8808), .A2(n14017), .A3(n13991), .A4(n13633), .ZN(
        n13634) );
  AND4_X1 U15252 ( .A1(n14009), .A2(n13964), .A3(n13949), .A4(n13634), .ZN(
        n13635) );
  NAND4_X1 U15253 ( .A1(n13923), .A2(n13975), .A3(n13910), .A4(n13635), .ZN(
        n13636) );
  NAND3_X1 U15254 ( .A1(n13649), .A2(n13648), .A3(n13775), .ZN(n13650) );
  OAI211_X1 U15255 ( .C1(n13651), .C2(n13653), .A(n13650), .B(P3_B_REG_SCAN_IN), .ZN(n13652) );
  OAI21_X1 U15256 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(P3_U3296) );
  MUX2_X1 U15257 ( .A(n13655), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13666), .Z(
        P3_U3521) );
  MUX2_X1 U15258 ( .A(n13860), .B(P3_DATAO_REG_29__SCAN_IN), .S(n13666), .Z(
        P3_U3520) );
  MUX2_X1 U15259 ( .A(n13656), .B(P3_DATAO_REG_28__SCAN_IN), .S(n13666), .Z(
        P3_U3519) );
  MUX2_X1 U15260 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13879), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15261 ( .A(n13896), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13666), .Z(
        P3_U3517) );
  MUX2_X1 U15262 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13880), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15263 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13895), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15264 ( .A(n13657), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13666), .Z(
        P3_U3513) );
  MUX2_X1 U15265 ( .A(n13967), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13666), .Z(
        P3_U3512) );
  MUX2_X1 U15266 ( .A(n13980), .B(P3_DATAO_REG_20__SCAN_IN), .S(n13666), .Z(
        P3_U3511) );
  MUX2_X1 U15267 ( .A(n13993), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13666), .Z(
        P3_U3510) );
  MUX2_X1 U15268 ( .A(n14020), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13666), .Z(
        P3_U3508) );
  MUX2_X1 U15269 ( .A(n14032), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13666), .Z(
        P3_U3507) );
  MUX2_X1 U15270 ( .A(n14031), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13666), .Z(
        P3_U3505) );
  MUX2_X1 U15271 ( .A(n14078), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13666), .Z(
        P3_U3504) );
  MUX2_X1 U15272 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13658), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15273 ( .A(n14079), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13666), .Z(
        P3_U3502) );
  MUX2_X1 U15274 ( .A(n13659), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13666), .Z(
        P3_U3500) );
  MUX2_X1 U15275 ( .A(n13660), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13666), .Z(
        P3_U3499) );
  MUX2_X1 U15276 ( .A(n13661), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13666), .Z(
        P3_U3498) );
  MUX2_X1 U15277 ( .A(n13662), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13666), .Z(
        P3_U3497) );
  MUX2_X1 U15278 ( .A(n13663), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13666), .Z(
        P3_U3496) );
  MUX2_X1 U15279 ( .A(n13664), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13666), .Z(
        P3_U3495) );
  MUX2_X1 U15280 ( .A(n13665), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13666), .Z(
        P3_U3494) );
  MUX2_X1 U15281 ( .A(n16312), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13666), .Z(
        P3_U3491) );
  AND3_X1 U15282 ( .A1(n13669), .A2(n13668), .A3(n13667), .ZN(n13670) );
  OAI21_X1 U15283 ( .B1(n13671), .B2(n13670), .A(n16272), .ZN(n13689) );
  INV_X1 U15284 ( .A(n13672), .ZN(n13674) );
  NAND3_X1 U15285 ( .A1(n13675), .A2(n13674), .A3(n13673), .ZN(n13676) );
  AOI21_X1 U15286 ( .B1(n13677), .B2(n13676), .A(n16285), .ZN(n13678) );
  AOI211_X1 U15287 ( .C1(n16037), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n13679), .B(
        n13678), .ZN(n13688) );
  NAND2_X1 U15288 ( .A1(n13813), .A2(n13680), .ZN(n13687) );
  AND3_X1 U15289 ( .A1(n13683), .A2(n13682), .A3(n13681), .ZN(n13684) );
  OAI21_X1 U15290 ( .B1(n13685), .B2(n13684), .A(n13840), .ZN(n13686) );
  NAND4_X1 U15291 ( .A1(n13689), .A2(n13688), .A3(n13687), .A4(n13686), .ZN(
        P3_U3186) );
  MUX2_X1 U15292 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13775), .Z(n13717) );
  XNOR2_X1 U15293 ( .A(n13717), .B(n13697), .ZN(n13696) );
  MUX2_X1 U15294 ( .A(n13691), .B(n13690), .S(n13775), .Z(n13693) );
  OAI21_X1 U15295 ( .B1(n13694), .B2(n13693), .A(n13692), .ZN(n13695) );
  NOR2_X1 U15296 ( .A1(n13695), .A2(n13696), .ZN(n13718) );
  AOI21_X1 U15297 ( .B1(n13696), .B2(n13695), .A(n13718), .ZN(n13711) );
  NOR2_X1 U15298 ( .A1(n13720), .A2(n13698), .ZN(n13724) );
  INV_X1 U15299 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14068) );
  AOI21_X1 U15300 ( .B1(n13699), .B2(n14068), .A(n13723), .ZN(n13708) );
  AOI21_X1 U15301 ( .B1(n13701), .B2(P3_REG1_REG_12__SCAN_IN), .A(n13700), 
        .ZN(n13702) );
  NOR2_X1 U15302 ( .A1(n13720), .A2(n13702), .ZN(n13713) );
  INV_X1 U15303 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n16472) );
  AOI21_X1 U15304 ( .B1(n13703), .B2(n16472), .A(n13712), .ZN(n13704) );
  NOR2_X1 U15305 ( .A1(n16285), .A2(n13704), .ZN(n13705) );
  AOI211_X1 U15306 ( .C1(n16037), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n13706), 
        .B(n13705), .ZN(n13707) );
  OAI21_X1 U15307 ( .B1(n13708), .B2(n16280), .A(n13707), .ZN(n13709) );
  AOI21_X1 U15308 ( .B1(n13720), .B2(n13813), .A(n13709), .ZN(n13710) );
  OAI21_X1 U15309 ( .B1(n13711), .B2(n16259), .A(n13710), .ZN(P3_U3195) );
  NAND2_X1 U15310 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n13734), .ZN(n13714) );
  OAI21_X1 U15311 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n13734), .A(n13714), 
        .ZN(n13715) );
  AOI21_X1 U15312 ( .B1(n13716), .B2(n13715), .A(n13735), .ZN(n13733) );
  INV_X1 U15313 ( .A(n13717), .ZN(n13719) );
  MUX2_X1 U15314 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13775), .Z(n13748) );
  XOR2_X1 U15315 ( .A(n13734), .B(n13748), .Z(n13721) );
  OAI211_X1 U15316 ( .C1(n13722), .C2(n13721), .A(n13749), .B(n16272), .ZN(
        n13732) );
  INV_X1 U15317 ( .A(n13734), .ZN(n13751) );
  NAND2_X1 U15318 ( .A1(n13734), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13739) );
  OAI21_X1 U15319 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13734), .A(n13739), 
        .ZN(n13726) );
  AOI21_X1 U15320 ( .B1(n13726), .B2(n13725), .A(n13738), .ZN(n13729) );
  AOI21_X1 U15321 ( .B1(n16037), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13727), 
        .ZN(n13728) );
  OAI21_X1 U15322 ( .B1(n16280), .B2(n13729), .A(n13728), .ZN(n13730) );
  AOI21_X1 U15323 ( .B1(n13751), .B2(n13813), .A(n13730), .ZN(n13731) );
  OAI211_X1 U15324 ( .C1(n13733), .C2(n16285), .A(n13732), .B(n13731), .ZN(
        P3_U3196) );
  NAND2_X1 U15325 ( .A1(n13736), .A2(n13773), .ZN(n13761) );
  OAI21_X1 U15326 ( .B1(n13736), .B2(n13773), .A(n13761), .ZN(n13737) );
  NOR2_X1 U15327 ( .A1(n13753), .A2(n13737), .ZN(n13762) );
  AOI21_X1 U15328 ( .B1(n13737), .B2(n13753), .A(n13762), .ZN(n13760) );
  INV_X1 U15329 ( .A(n13773), .ZN(n13758) );
  NAND2_X1 U15330 ( .A1(n13742), .A2(n14035), .ZN(n13743) );
  NAND2_X1 U15331 ( .A1(n13743), .A2(n7503), .ZN(n13744) );
  NAND2_X1 U15332 ( .A1(n13840), .A2(n13744), .ZN(n13746) );
  OAI211_X1 U15333 ( .C1(n13747), .C2(n16292), .A(n13746), .B(n13745), .ZN(
        n13757) );
  INV_X1 U15334 ( .A(n13748), .ZN(n13750) );
  XOR2_X1 U15335 ( .A(n13773), .B(n13752), .Z(n13755) );
  MUX2_X1 U15336 ( .A(n14035), .B(n13753), .S(n13775), .Z(n13754) );
  NOR2_X1 U15337 ( .A1(n13755), .A2(n13754), .ZN(n13772) );
  AOI211_X1 U15338 ( .C1(n13755), .C2(n13754), .A(n16259), .B(n13772), .ZN(
        n13756) );
  AOI211_X1 U15339 ( .C1(n13813), .C2(n13758), .A(n13757), .B(n13756), .ZN(
        n13759) );
  OAI21_X1 U15340 ( .B1(n13760), .B2(n16285), .A(n13759), .ZN(P3_U3197) );
  INV_X1 U15341 ( .A(n13761), .ZN(n13763) );
  AOI22_X1 U15342 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13780), .B1(n13794), 
        .B2(n14154), .ZN(n13764) );
  NOR2_X1 U15343 ( .A1(n13765), .A2(n13764), .ZN(n13783) );
  AOI21_X1 U15344 ( .B1(n13765), .B2(n13764), .A(n13783), .ZN(n13782) );
  AOI22_X1 U15345 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13780), .B1(n13794), 
        .B2(n14024), .ZN(n13767) );
  AND2_X1 U15346 ( .A1(n13767), .A2(n7516), .ZN(n13768) );
  OAI21_X1 U15347 ( .B1(n13785), .B2(n13768), .A(n13840), .ZN(n13770) );
  OAI211_X1 U15348 ( .C1(n13771), .C2(n16292), .A(n13770), .B(n13769), .ZN(
        n13779) );
  AOI21_X1 U15349 ( .B1(n13774), .B2(n13773), .A(n13772), .ZN(n13777) );
  MUX2_X1 U15350 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13775), .Z(n13795) );
  XNOR2_X1 U15351 ( .A(n13795), .B(n13794), .ZN(n13776) );
  NOR2_X1 U15352 ( .A1(n13777), .A2(n13776), .ZN(n13793) );
  AOI211_X1 U15353 ( .C1(n13777), .C2(n13776), .A(n16259), .B(n13793), .ZN(
        n13778) );
  AOI211_X1 U15354 ( .C1(n13813), .C2(n13780), .A(n13779), .B(n13778), .ZN(
        n13781) );
  OAI21_X1 U15355 ( .B1(n13782), .B2(n16285), .A(n13781), .ZN(P3_U3198) );
  AOI21_X1 U15356 ( .B1(n14147), .B2(n13784), .A(n13814), .ZN(n13801) );
  AOI21_X1 U15357 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13794), .A(n13785), 
        .ZN(n13807) );
  XOR2_X1 U15358 ( .A(n13807), .B(n13803), .Z(n13786) );
  INV_X1 U15359 ( .A(n13786), .ZN(n13788) );
  NOR2_X1 U15360 ( .A1(n14011), .A2(n13786), .ZN(n13809) );
  INV_X1 U15361 ( .A(n13809), .ZN(n13787) );
  OAI21_X1 U15362 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13788), .A(n13787), 
        .ZN(n13789) );
  NAND2_X1 U15363 ( .A1(n13840), .A2(n13789), .ZN(n13791) );
  OAI211_X1 U15364 ( .C1(n13792), .C2(n16292), .A(n13791), .B(n13790), .ZN(
        n13799) );
  MUX2_X1 U15365 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13775), .Z(n13804) );
  XNOR2_X1 U15366 ( .A(n13804), .B(n13803), .ZN(n13796) );
  NOR2_X1 U15367 ( .A1(n13797), .A2(n13796), .ZN(n13802) );
  AOI211_X1 U15368 ( .C1(n13797), .C2(n13796), .A(n16259), .B(n13802), .ZN(
        n13798) );
  OAI21_X1 U15369 ( .B1(n13801), .B2(n16285), .A(n13800), .ZN(P3_U3199) );
  MUX2_X1 U15370 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13775), .Z(n13806) );
  XNOR2_X1 U15371 ( .A(n13828), .B(n13827), .ZN(n13805) );
  AOI21_X1 U15372 ( .B1(n13806), .B2(n13805), .A(n13826), .ZN(n13825) );
  NOR2_X1 U15373 ( .A1(n7977), .A2(n13807), .ZN(n13810) );
  INV_X1 U15374 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13996) );
  NOR2_X1 U15375 ( .A1(n13827), .A2(n13996), .ZN(n13831) );
  AOI21_X1 U15376 ( .B1(n13827), .B2(n13996), .A(n13831), .ZN(n13808) );
  OAI21_X1 U15377 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13833) );
  OR2_X1 U15378 ( .A1(n13815), .A2(n7977), .ZN(n13820) );
  NAND2_X1 U15379 ( .A1(n13816), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13841) );
  INV_X1 U15380 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U15381 ( .A1(n13827), .A2(n13817), .ZN(n13818) );
  NAND2_X1 U15382 ( .A1(n13841), .A2(n13818), .ZN(n13819) );
  AND3_X1 U15383 ( .A1(n13821), .A2(n13820), .A3(n13819), .ZN(n13822) );
  OAI21_X1 U15384 ( .B1(n13843), .B2(n13822), .A(n13847), .ZN(n13823) );
  OAI211_X1 U15385 ( .C1(n13825), .C2(n16259), .A(n13824), .B(n13823), .ZN(
        P3_U3200) );
  XNOR2_X1 U15386 ( .A(n13829), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13834) );
  XNOR2_X1 U15387 ( .A(n13837), .B(n14139), .ZN(n13844) );
  MUX2_X1 U15388 ( .A(n13834), .B(n13844), .S(n13775), .Z(n13830) );
  INV_X1 U15389 ( .A(n13831), .ZN(n13832) );
  NAND2_X1 U15390 ( .A1(n13833), .A2(n13832), .ZN(n13835) );
  OAI21_X1 U15391 ( .B1(n16292), .B2(n8359), .A(n13836), .ZN(n13839) );
  NOR2_X1 U15392 ( .A1(n16278), .A2(n13837), .ZN(n13838) );
  INV_X1 U15393 ( .A(n13841), .ZN(n13842) );
  NOR2_X1 U15394 ( .A1(n13843), .A2(n13842), .ZN(n13846) );
  INV_X1 U15395 ( .A(n13844), .ZN(n13845) );
  XNOR2_X1 U15396 ( .A(n13846), .B(n13845), .ZN(n13848) );
  NAND2_X1 U15397 ( .A1(n13849), .A2(n16382), .ZN(n13852) );
  OR2_X1 U15398 ( .A1(n13851), .A2(n13850), .ZN(n16482) );
  NAND3_X1 U15399 ( .A1(n16390), .A2(n13852), .A3(n16482), .ZN(n13854) );
  OAI21_X1 U15400 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n16386), .A(n13854), 
        .ZN(n13853) );
  OAI21_X1 U15401 ( .B1(n14106), .B2(n14075), .A(n13853), .ZN(P3_U3202) );
  OAI21_X1 U15402 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n16386), .A(n13854), 
        .ZN(n13855) );
  OAI21_X1 U15403 ( .B1(n14109), .B2(n14075), .A(n13855), .ZN(P3_U3203) );
  AOI22_X1 U15404 ( .A1(n13860), .A2(n16313), .B1(n16311), .B2(n13879), .ZN(
        n13861) );
  OAI21_X1 U15405 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n14110) );
  INV_X1 U15406 ( .A(n13866), .ZN(n14170) );
  AOI22_X1 U15407 ( .A1(n13867), .A2(n16382), .B1(n16348), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13868) );
  OAI21_X1 U15408 ( .B1(n14170), .B2(n14075), .A(n13868), .ZN(n13869) );
  AOI21_X1 U15409 ( .B1(n14110), .B2(n14039), .A(n13869), .ZN(n13870) );
  OAI21_X1 U15410 ( .B1(n14111), .B2(n16348), .A(n13870), .ZN(P3_U3205) );
  MUX2_X1 U15411 ( .A(P3_REG2_REG_27__SCAN_IN), .B(n13871), .S(n16390), .Z(
        n13872) );
  INV_X1 U15412 ( .A(n13872), .ZN(n13876) );
  AOI22_X1 U15413 ( .A1(n13874), .A2(n16384), .B1(n16382), .B2(n13873), .ZN(
        n13875) );
  OAI211_X1 U15414 ( .C1(n13877), .C2(n14104), .A(n13876), .B(n13875), .ZN(
        P3_U3206) );
  XNOR2_X1 U15415 ( .A(n13878), .B(n13882), .ZN(n13881) );
  AOI222_X1 U15416 ( .A1(n16309), .A2(n13881), .B1(n13880), .B2(n16311), .C1(
        n13879), .C2(n16313), .ZN(n14112) );
  AND2_X1 U15417 ( .A1(n13883), .A2(n13882), .ZN(n13884) );
  OR2_X1 U15418 ( .A1(n13885), .A2(n13884), .ZN(n14113) );
  AOI22_X1 U15419 ( .A1(n13886), .A2(n16382), .B1(n16348), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U15420 ( .A1(n13887), .A2(n16384), .ZN(n13888) );
  OAI211_X1 U15421 ( .C1(n14113), .C2(n14054), .A(n13889), .B(n13888), .ZN(
        n13890) );
  INV_X1 U15422 ( .A(n13890), .ZN(n13891) );
  OAI21_X1 U15423 ( .B1(n14112), .B2(n16348), .A(n13891), .ZN(P3_U3207) );
  INV_X1 U15424 ( .A(n13892), .ZN(n13894) );
  OAI21_X1 U15425 ( .B1(n13894), .B2(n13893), .A(n16309), .ZN(n13899) );
  AOI22_X1 U15426 ( .A1(n13896), .A2(n16313), .B1(n13895), .B2(n16311), .ZN(
        n13897) );
  OAI21_X1 U15427 ( .B1(n13899), .B2(n13898), .A(n13897), .ZN(n14115) );
  INV_X1 U15428 ( .A(n14115), .ZN(n13907) );
  OAI21_X1 U15429 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n14116) );
  AOI22_X1 U15430 ( .A1(n13903), .A2(n16382), .B1(n16348), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U15431 ( .B1(n14179), .B2(n14075), .A(n13904), .ZN(n13905) );
  AOI21_X1 U15432 ( .B1(n14116), .B2(n14039), .A(n13905), .ZN(n13906) );
  OAI21_X1 U15433 ( .B1(n13907), .B2(n16348), .A(n13906), .ZN(P3_U3208) );
  XNOR2_X1 U15434 ( .A(n13908), .B(n13910), .ZN(n14185) );
  INV_X1 U15435 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13915) );
  XNOR2_X1 U15436 ( .A(n13909), .B(n13910), .ZN(n13913) );
  OAI22_X1 U15437 ( .A1(n13911), .A2(n14090), .B1(n13936), .B2(n14092), .ZN(
        n13912) );
  AOI21_X1 U15438 ( .B1(n13913), .B2(n16309), .A(n13912), .ZN(n13914) );
  OAI21_X1 U15439 ( .B1(n14097), .B2(n14185), .A(n13914), .ZN(n14119) );
  INV_X1 U15440 ( .A(n14119), .ZN(n14180) );
  MUX2_X1 U15441 ( .A(n13915), .B(n14180), .S(n16390), .Z(n13918) );
  AOI22_X1 U15442 ( .A1(n14182), .A2(n16384), .B1(n16382), .B2(n13916), .ZN(
        n13917) );
  OAI211_X1 U15443 ( .C1(n14185), .C2(n14104), .A(n13918), .B(n13917), .ZN(
        P3_U3209) );
  XNOR2_X1 U15444 ( .A(n13919), .B(n13923), .ZN(n13920) );
  OAI222_X1 U15445 ( .A1(n14090), .A2(n13921), .B1(n14092), .B2(n13951), .C1(
        n13920), .C2(n14005), .ZN(n14123) );
  NAND2_X1 U15446 ( .A1(n13938), .A2(n13922), .ZN(n13925) );
  INV_X1 U15447 ( .A(n13923), .ZN(n13924) );
  NAND2_X1 U15448 ( .A1(n13925), .A2(n13924), .ZN(n13927) );
  AND2_X1 U15449 ( .A1(n13927), .A2(n13926), .ZN(n14124) );
  NAND2_X1 U15450 ( .A1(n14124), .A2(n14039), .ZN(n13930) );
  AOI22_X1 U15451 ( .A1(n16348), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13928), 
        .B2(n16382), .ZN(n13929) );
  OAI211_X1 U15452 ( .C1(n14189), .C2(n14075), .A(n13930), .B(n13929), .ZN(
        n13931) );
  AOI21_X1 U15453 ( .B1(n14123), .B2(n16386), .A(n13931), .ZN(n13932) );
  INV_X1 U15454 ( .A(n13932), .ZN(P3_U3210) );
  XNOR2_X1 U15455 ( .A(n13934), .B(n13933), .ZN(n13935) );
  OAI222_X1 U15456 ( .A1(n14092), .A2(n13937), .B1(n14090), .B2(n13936), .C1(
        n13935), .C2(n14005), .ZN(n14127) );
  INV_X1 U15457 ( .A(n14127), .ZN(n13945) );
  OAI21_X1 U15458 ( .B1(n13940), .B2(n13939), .A(n13938), .ZN(n14128) );
  AOI22_X1 U15459 ( .A1(n16348), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n16382), 
        .B2(n13941), .ZN(n13942) );
  OAI21_X1 U15460 ( .B1(n14193), .B2(n14075), .A(n13942), .ZN(n13943) );
  AOI21_X1 U15461 ( .B1(n14128), .B2(n14039), .A(n13943), .ZN(n13944) );
  OAI21_X1 U15462 ( .B1(n13945), .B2(n16348), .A(n13944), .ZN(P3_U3211) );
  XOR2_X1 U15463 ( .A(n13949), .B(n13946), .Z(n14196) );
  INV_X1 U15464 ( .A(n14196), .ZN(n13957) );
  OAI22_X1 U15465 ( .A1(n14195), .A2(n14075), .B1(n13947), .B2(n16339), .ZN(
        n13956) );
  XOR2_X1 U15466 ( .A(n13949), .B(n13948), .Z(n13953) );
  OAI22_X1 U15467 ( .A1(n13951), .A2(n14090), .B1(n13950), .B2(n14092), .ZN(
        n13952) );
  AOI21_X1 U15468 ( .B1(n13953), .B2(n16309), .A(n13952), .ZN(n13954) );
  OAI21_X1 U15469 ( .B1(n14097), .B2(n14196), .A(n13954), .ZN(n14194) );
  MUX2_X1 U15470 ( .A(P3_REG2_REG_21__SCAN_IN), .B(n14194), .S(n16390), .Z(
        n13955) );
  AOI211_X1 U15471 ( .C1(n13957), .C2(n14084), .A(n13956), .B(n13955), .ZN(
        n13958) );
  INV_X1 U15472 ( .A(n13958), .ZN(P3_U3212) );
  NAND2_X1 U15473 ( .A1(n14000), .A2(n13999), .ZN(n13998) );
  NAND2_X1 U15474 ( .A1(n13998), .A2(n13959), .ZN(n13976) );
  NAND2_X1 U15475 ( .A1(n13976), .A2(n13975), .ZN(n13961) );
  NAND2_X1 U15476 ( .A1(n13961), .A2(n13960), .ZN(n13963) );
  XNOR2_X1 U15477 ( .A(n13963), .B(n13962), .ZN(n14201) );
  XNOR2_X1 U15478 ( .A(n13965), .B(n13964), .ZN(n13966) );
  NAND2_X1 U15479 ( .A1(n13966), .A2(n16309), .ZN(n13969) );
  AOI22_X1 U15480 ( .A1(n13967), .A2(n16313), .B1(n13993), .B2(n16311), .ZN(
        n13968) );
  OAI211_X1 U15481 ( .C1(n14097), .C2(n14201), .A(n13969), .B(n13968), .ZN(
        n14199) );
  MUX2_X1 U15482 ( .A(P3_REG2_REG_20__SCAN_IN), .B(n14199), .S(n16390), .Z(
        n13970) );
  INV_X1 U15483 ( .A(n13970), .ZN(n13974) );
  AOI22_X1 U15484 ( .A1(n13972), .A2(n16384), .B1(n16382), .B2(n13971), .ZN(
        n13973) );
  OAI211_X1 U15485 ( .C1(n14201), .C2(n14104), .A(n13974), .B(n13973), .ZN(
        P3_U3213) );
  INV_X1 U15486 ( .A(n13975), .ZN(n13977) );
  XNOR2_X1 U15487 ( .A(n13976), .B(n13977), .ZN(n14136) );
  XNOR2_X1 U15488 ( .A(n13978), .B(n13977), .ZN(n13979) );
  NAND2_X1 U15489 ( .A1(n13979), .A2(n16309), .ZN(n13983) );
  AOI22_X1 U15490 ( .A1(n16311), .A2(n13981), .B1(n13980), .B2(n16313), .ZN(
        n13982) );
  NAND2_X1 U15491 ( .A1(n13983), .A2(n13982), .ZN(n14138) );
  NAND2_X1 U15492 ( .A1(n14138), .A2(n16386), .ZN(n13989) );
  INV_X1 U15493 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13985) );
  OAI22_X1 U15494 ( .A1(n16390), .A2(n13985), .B1(n13984), .B2(n16339), .ZN(
        n13986) );
  AOI21_X1 U15495 ( .B1(n13987), .B2(n16384), .A(n13986), .ZN(n13988) );
  OAI211_X1 U15496 ( .C1(n14136), .C2(n14054), .A(n13989), .B(n13988), .ZN(
        P3_U3214) );
  OAI21_X1 U15497 ( .B1(n13992), .B2(n13991), .A(n13990), .ZN(n13994) );
  AOI222_X1 U15498 ( .A1(n16309), .A2(n13994), .B1(n13993), .B2(n16313), .C1(
        n14020), .C2(n16311), .ZN(n14144) );
  OAI22_X1 U15499 ( .A1(n16390), .A2(n13996), .B1(n13995), .B2(n16339), .ZN(
        n13997) );
  AOI21_X1 U15500 ( .B1(n14141), .B2(n16384), .A(n13997), .ZN(n14002) );
  OAI21_X1 U15501 ( .B1(n14000), .B2(n13999), .A(n13998), .ZN(n14142) );
  NAND2_X1 U15502 ( .A1(n14142), .A2(n14039), .ZN(n14001) );
  OAI211_X1 U15503 ( .C1(n14144), .C2(n16348), .A(n14002), .B(n14001), .ZN(
        P3_U3215) );
  XNOR2_X1 U15504 ( .A(n14003), .B(n14009), .ZN(n14004) );
  OAI222_X1 U15505 ( .A1(n14090), .A2(n14007), .B1(n14092), .B2(n14006), .C1(
        n14005), .C2(n14004), .ZN(n14145) );
  INV_X1 U15506 ( .A(n14145), .ZN(n14015) );
  XNOR2_X1 U15507 ( .A(n14008), .B(n14009), .ZN(n14146) );
  NOR2_X1 U15508 ( .A1(n14211), .A2(n14075), .ZN(n14013) );
  OAI22_X1 U15509 ( .A1(n16390), .A2(n14011), .B1(n14010), .B2(n16339), .ZN(
        n14012) );
  AOI211_X1 U15510 ( .C1(n14146), .C2(n14039), .A(n14013), .B(n14012), .ZN(
        n14014) );
  OAI21_X1 U15511 ( .B1(n14015), .B2(n16348), .A(n14014), .ZN(P3_U3216) );
  XNOR2_X1 U15512 ( .A(n14016), .B(n14017), .ZN(n14151) );
  XNOR2_X1 U15513 ( .A(n14018), .B(n14017), .ZN(n14019) );
  NAND2_X1 U15514 ( .A1(n14019), .A2(n16309), .ZN(n14022) );
  AOI22_X1 U15515 ( .A1(n16311), .A2(n14046), .B1(n14020), .B2(n16313), .ZN(
        n14021) );
  NAND2_X1 U15516 ( .A1(n14022), .A2(n14021), .ZN(n14153) );
  NAND2_X1 U15517 ( .A1(n14153), .A2(n16386), .ZN(n14028) );
  OAI22_X1 U15518 ( .A1(n16390), .A2(n14024), .B1(n14023), .B2(n16339), .ZN(
        n14025) );
  AOI21_X1 U15519 ( .B1(n14026), .B2(n16384), .A(n14025), .ZN(n14027) );
  OAI211_X1 U15520 ( .C1(n14151), .C2(n14054), .A(n14028), .B(n14027), .ZN(
        P3_U3217) );
  OAI21_X1 U15521 ( .B1(n14030), .B2(n8808), .A(n14029), .ZN(n14033) );
  AOI222_X1 U15522 ( .A1(n16309), .A2(n14033), .B1(n14032), .B2(n16313), .C1(
        n14031), .C2(n16311), .ZN(n14158) );
  INV_X1 U15523 ( .A(n14159), .ZN(n14037) );
  OAI22_X1 U15524 ( .A1(n16386), .A2(n14035), .B1(n14034), .B2(n16339), .ZN(
        n14036) );
  AOI21_X1 U15525 ( .B1(n14037), .B2(n16384), .A(n14036), .ZN(n14041) );
  XNOR2_X1 U15526 ( .A(n14038), .B(n8808), .ZN(n14156) );
  NAND2_X1 U15527 ( .A1(n14156), .A2(n14039), .ZN(n14040) );
  OAI211_X1 U15528 ( .C1(n14158), .C2(n16348), .A(n14041), .B(n14040), .ZN(
        P3_U3218) );
  XNOR2_X1 U15529 ( .A(n14042), .B(n14043), .ZN(n14161) );
  INV_X1 U15530 ( .A(n14161), .ZN(n14053) );
  INV_X1 U15531 ( .A(n14043), .ZN(n14045) );
  OAI211_X1 U15532 ( .C1(n7537), .C2(n14045), .A(n16309), .B(n14044), .ZN(
        n14048) );
  AOI22_X1 U15533 ( .A1(n16313), .A2(n14046), .B1(n14078), .B2(n16311), .ZN(
        n14047) );
  NAND2_X1 U15534 ( .A1(n14048), .A2(n14047), .ZN(n14160) );
  AOI22_X1 U15535 ( .A1(n16348), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16382), 
        .B2(n14049), .ZN(n14050) );
  OAI21_X1 U15536 ( .B1(n14219), .B2(n14075), .A(n14050), .ZN(n14051) );
  AOI21_X1 U15537 ( .B1(n14160), .B2(n16386), .A(n14051), .ZN(n14052) );
  OAI21_X1 U15538 ( .B1(n14054), .B2(n14053), .A(n14052), .ZN(P3_U3219) );
  XOR2_X1 U15539 ( .A(n14061), .B(n14055), .Z(n16469) );
  NAND2_X1 U15540 ( .A1(n14056), .A2(n14057), .ZN(n14059) );
  NAND2_X1 U15541 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  XOR2_X1 U15542 ( .A(n14061), .B(n14060), .Z(n14065) );
  OAI22_X1 U15543 ( .A1(n14063), .A2(n14090), .B1(n14062), .B2(n14092), .ZN(
        n14064) );
  AOI21_X1 U15544 ( .B1(n14065), .B2(n16309), .A(n14064), .ZN(n14066) );
  OAI21_X1 U15545 ( .B1(n14097), .B2(n16469), .A(n14066), .ZN(n16471) );
  NAND2_X1 U15546 ( .A1(n16471), .A2(n16386), .ZN(n14072) );
  INV_X1 U15547 ( .A(n16466), .ZN(n14070) );
  OAI22_X1 U15548 ( .A1(n16386), .A2(n14068), .B1(n14067), .B2(n16339), .ZN(
        n14069) );
  AOI21_X1 U15549 ( .B1(n14070), .B2(n16384), .A(n14069), .ZN(n14071) );
  OAI211_X1 U15550 ( .C1(n16469), .C2(n14104), .A(n14072), .B(n14071), .ZN(
        P3_U3220) );
  XNOR2_X1 U15551 ( .A(n14073), .B(n14076), .ZN(n14224) );
  INV_X1 U15552 ( .A(n14224), .ZN(n14085) );
  OAI22_X1 U15553 ( .A1(n14075), .A2(n14222), .B1(n14074), .B2(n16339), .ZN(
        n14083) );
  XNOR2_X1 U15554 ( .A(n14056), .B(n14076), .ZN(n14077) );
  NAND2_X1 U15555 ( .A1(n14077), .A2(n16309), .ZN(n14081) );
  AOI22_X1 U15556 ( .A1(n16311), .A2(n14079), .B1(n14078), .B2(n16313), .ZN(
        n14080) );
  OAI211_X1 U15557 ( .C1(n14097), .C2(n14224), .A(n14081), .B(n14080), .ZN(
        n14220) );
  MUX2_X1 U15558 ( .A(P3_REG2_REG_12__SCAN_IN), .B(n14220), .S(n16390), .Z(
        n14082) );
  AOI211_X1 U15559 ( .C1(n14085), .C2(n14084), .A(n14083), .B(n14082), .ZN(
        n14086) );
  INV_X1 U15560 ( .A(n14086), .ZN(P3_U3221) );
  XOR2_X1 U15561 ( .A(n14088), .B(n14087), .Z(n16400) );
  XOR2_X1 U15562 ( .A(n14089), .B(n14088), .Z(n14095) );
  OAI22_X1 U15563 ( .A1(n14093), .A2(n14092), .B1(n14091), .B2(n14090), .ZN(
        n14094) );
  AOI21_X1 U15564 ( .B1(n14095), .B2(n16309), .A(n14094), .ZN(n14096) );
  OAI21_X1 U15565 ( .B1(n14097), .B2(n16400), .A(n14096), .ZN(n16402) );
  NAND2_X1 U15566 ( .A1(n16402), .A2(n16386), .ZN(n14103) );
  OAI22_X1 U15567 ( .A1(n16386), .A2(n14099), .B1(n14098), .B2(n16339), .ZN(
        n14100) );
  AOI21_X1 U15568 ( .B1(n14101), .B2(n16384), .A(n14100), .ZN(n14102) );
  OAI211_X1 U15569 ( .C1(n16400), .C2(n14104), .A(n14103), .B(n14102), .ZN(
        P3_U3223) );
  NOR2_X1 U15570 ( .A1(n10822), .A2(n16482), .ZN(n14107) );
  AOI21_X1 U15571 ( .B1(n10822), .B2(P3_REG1_REG_31__SCAN_IN), .A(n14107), 
        .ZN(n14105) );
  OAI21_X1 U15572 ( .B1(n14106), .B2(n14164), .A(n14105), .ZN(P3_U3490) );
  AOI21_X1 U15573 ( .B1(n10822), .B2(P3_REG1_REG_30__SCAN_IN), .A(n14107), 
        .ZN(n14108) );
  OAI21_X1 U15574 ( .B1(n14109), .B2(n14164), .A(n14108), .ZN(P3_U3489) );
  OAI21_X1 U15575 ( .B1(n14150), .B2(n14113), .A(n14112), .ZN(n14171) );
  OAI21_X1 U15576 ( .B1(n14175), .B2(n14164), .A(n14114), .ZN(P3_U3485) );
  INV_X1 U15577 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14117) );
  AOI21_X1 U15578 ( .B1(n10820), .B2(n14116), .A(n14115), .ZN(n14176) );
  MUX2_X1 U15579 ( .A(n14117), .B(n14176), .S(n16473), .Z(n14118) );
  OAI21_X1 U15580 ( .B1(n14179), .B2(n14164), .A(n14118), .ZN(P3_U3484) );
  MUX2_X1 U15581 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n14119), .S(n16473), .Z(
        n14122) );
  OAI22_X1 U15582 ( .A1(n14185), .A2(n14165), .B1(n14120), .B2(n14164), .ZN(
        n14121) );
  OR2_X1 U15583 ( .A1(n14122), .A2(n14121), .ZN(P3_U3483) );
  INV_X1 U15584 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14125) );
  AOI21_X1 U15585 ( .B1(n14124), .B2(n10820), .A(n14123), .ZN(n14186) );
  MUX2_X1 U15586 ( .A(n14125), .B(n14186), .S(n16473), .Z(n14126) );
  OAI21_X1 U15587 ( .B1(n14189), .B2(n14164), .A(n14126), .ZN(P3_U3482) );
  INV_X1 U15588 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n14129) );
  AOI21_X1 U15589 ( .B1(n10820), .B2(n14128), .A(n14127), .ZN(n14190) );
  MUX2_X1 U15590 ( .A(n14129), .B(n14190), .S(n16473), .Z(n14130) );
  OAI21_X1 U15591 ( .B1(n14193), .B2(n14164), .A(n14130), .ZN(P3_U3481) );
  MUX2_X1 U15592 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n14194), .S(n16473), .Z(
        n14132) );
  OAI22_X1 U15593 ( .A1(n14196), .A2(n14165), .B1(n14195), .B2(n14164), .ZN(
        n14131) );
  OR2_X1 U15594 ( .A1(n14132), .A2(n14131), .ZN(P3_U3480) );
  MUX2_X1 U15595 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14199), .S(n16473), .Z(
        n14134) );
  OAI22_X1 U15596 ( .A1(n14201), .A2(n14165), .B1(n14200), .B2(n14164), .ZN(
        n14133) );
  OR2_X1 U15597 ( .A1(n14134), .A2(n14133), .ZN(P3_U3479) );
  OAI22_X1 U15598 ( .A1(n14136), .A2(n14150), .B1(n14135), .B2(n16467), .ZN(
        n14137) );
  NOR2_X1 U15599 ( .A1(n14138), .A2(n14137), .ZN(n14204) );
  MUX2_X1 U15600 ( .A(n14139), .B(n14204), .S(n16473), .Z(n14140) );
  INV_X1 U15601 ( .A(n14140), .ZN(P3_U3478) );
  AOI22_X1 U15602 ( .A1(n14142), .A2(n10820), .B1(n16418), .B2(n14141), .ZN(
        n14143) );
  NAND2_X1 U15603 ( .A1(n14144), .A2(n14143), .ZN(n14207) );
  MUX2_X1 U15604 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14207), .S(n16473), .Z(
        P3_U3477) );
  AOI21_X1 U15605 ( .B1(n14146), .B2(n10820), .A(n14145), .ZN(n14208) );
  MUX2_X1 U15606 ( .A(n14147), .B(n14208), .S(n16473), .Z(n14148) );
  OAI21_X1 U15607 ( .B1(n14164), .B2(n14211), .A(n14148), .ZN(P3_U3476) );
  OAI22_X1 U15608 ( .A1(n14151), .A2(n14150), .B1(n14149), .B2(n16467), .ZN(
        n14152) );
  NOR2_X1 U15609 ( .A1(n14153), .A2(n14152), .ZN(n14212) );
  MUX2_X1 U15610 ( .A(n14154), .B(n14212), .S(n16473), .Z(n14155) );
  INV_X1 U15611 ( .A(n14155), .ZN(P3_U3475) );
  NAND2_X1 U15612 ( .A1(n14156), .A2(n10820), .ZN(n14157) );
  OAI211_X1 U15613 ( .C1(n14159), .C2(n16467), .A(n14158), .B(n14157), .ZN(
        n14215) );
  MUX2_X1 U15614 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n14215), .S(n16473), .Z(
        P3_U3474) );
  INV_X1 U15615 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14162) );
  AOI21_X1 U15616 ( .B1(n14161), .B2(n10820), .A(n14160), .ZN(n14216) );
  MUX2_X1 U15617 ( .A(n14162), .B(n14216), .S(n16473), .Z(n14163) );
  OAI21_X1 U15618 ( .B1(n14164), .B2(n14219), .A(n14163), .ZN(P3_U3473) );
  MUX2_X1 U15619 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n14220), .S(n16473), .Z(
        n14167) );
  OAI22_X1 U15620 ( .A1(n14224), .A2(n14165), .B1(n14222), .B2(n14164), .ZN(
        n14166) );
  OR2_X1 U15621 ( .A1(n14167), .A2(n14166), .ZN(P3_U3471) );
  OAI21_X1 U15622 ( .B1(n14170), .B2(n14221), .A(n14169), .ZN(P3_U3455) );
  INV_X1 U15623 ( .A(n14171), .ZN(n14172) );
  MUX2_X1 U15624 ( .A(n14173), .B(n14172), .S(n16476), .Z(n14174) );
  OAI21_X1 U15625 ( .B1(n14175), .B2(n14221), .A(n14174), .ZN(P3_U3453) );
  MUX2_X1 U15626 ( .A(n14177), .B(n14176), .S(n16476), .Z(n14178) );
  OAI21_X1 U15627 ( .B1(n14179), .B2(n14221), .A(n14178), .ZN(P3_U3452) );
  MUX2_X1 U15628 ( .A(n14181), .B(n14180), .S(n16476), .Z(n14184) );
  INV_X1 U15629 ( .A(n14221), .ZN(n16479) );
  NAND2_X1 U15630 ( .A1(n14182), .A2(n16479), .ZN(n14183) );
  OAI211_X1 U15631 ( .C1(n14185), .C2(n14223), .A(n14184), .B(n14183), .ZN(
        P3_U3451) );
  INV_X1 U15632 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14187) );
  MUX2_X1 U15633 ( .A(n14187), .B(n14186), .S(n16476), .Z(n14188) );
  OAI21_X1 U15634 ( .B1(n14189), .B2(n14221), .A(n14188), .ZN(P3_U3450) );
  INV_X1 U15635 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14191) );
  MUX2_X1 U15636 ( .A(n14191), .B(n14190), .S(n16476), .Z(n14192) );
  OAI21_X1 U15637 ( .B1(n14193), .B2(n14221), .A(n14192), .ZN(P3_U3449) );
  MUX2_X1 U15638 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n14194), .S(n16476), .Z(
        n14198) );
  OAI22_X1 U15639 ( .A1(n14196), .A2(n14223), .B1(n14195), .B2(n14221), .ZN(
        n14197) );
  OR2_X1 U15640 ( .A1(n14198), .A2(n14197), .ZN(P3_U3448) );
  MUX2_X1 U15641 ( .A(n14199), .B(P3_REG0_REG_20__SCAN_IN), .S(n16483), .Z(
        n14203) );
  OAI22_X1 U15642 ( .A1(n14201), .A2(n14223), .B1(n14200), .B2(n14221), .ZN(
        n14202) );
  OR2_X1 U15643 ( .A1(n14203), .A2(n14202), .ZN(P3_U3447) );
  INV_X1 U15644 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14205) );
  MUX2_X1 U15645 ( .A(n14205), .B(n14204), .S(n16476), .Z(n14206) );
  INV_X1 U15646 ( .A(n14206), .ZN(P3_U3446) );
  MUX2_X1 U15647 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14207), .S(n16476), .Z(
        P3_U3444) );
  INV_X1 U15648 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14209) );
  MUX2_X1 U15649 ( .A(n14209), .B(n14208), .S(n16476), .Z(n14210) );
  OAI21_X1 U15650 ( .B1(n14221), .B2(n14211), .A(n14210), .ZN(P3_U3441) );
  INV_X1 U15651 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14213) );
  MUX2_X1 U15652 ( .A(n14213), .B(n14212), .S(n16476), .Z(n14214) );
  INV_X1 U15653 ( .A(n14214), .ZN(P3_U3438) );
  MUX2_X1 U15654 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n14215), .S(n16476), .Z(
        P3_U3435) );
  MUX2_X1 U15655 ( .A(n14217), .B(n14216), .S(n16476), .Z(n14218) );
  OAI21_X1 U15656 ( .B1(n14221), .B2(n14219), .A(n14218), .ZN(P3_U3432) );
  MUX2_X1 U15657 ( .A(n14220), .B(P3_REG0_REG_12__SCAN_IN), .S(n16483), .Z(
        n14226) );
  OAI22_X1 U15658 ( .A1(n14224), .A2(n14223), .B1(n14222), .B2(n14221), .ZN(
        n14225) );
  OR2_X1 U15659 ( .A1(n14226), .A2(n14225), .ZN(P3_U3426) );
  MUX2_X1 U15660 ( .A(P3_D_REG_1__SCAN_IN), .B(n14228), .S(n14227), .Z(
        P3_U3377) );
  NAND2_X1 U15661 ( .A1(n14230), .A2(n14229), .ZN(n14234) );
  OR4_X1 U15662 ( .A1(n14232), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n14231), .ZN(n14233) );
  OAI211_X1 U15663 ( .C1(n14235), .C2(n14237), .A(n14234), .B(n14233), .ZN(
        P3_U3264) );
  INV_X1 U15664 ( .A(n14236), .ZN(n14238) );
  OAI222_X1 U15665 ( .A1(n13194), .A2(n14238), .B1(n8525), .B2(P3_U3151), .C1(
        n15633), .C2(n14237), .ZN(P3_U3266) );
  MUX2_X1 U15666 ( .A(n14240), .B(n14239), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3271) );
  MUX2_X1 U15667 ( .A(n14241), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15668 ( .A(n14530), .B(n14306), .ZN(n14267) );
  INV_X1 U15669 ( .A(n14243), .ZN(n14244) );
  AND2_X1 U15670 ( .A1(n14601), .A2(n14305), .ZN(n14247) );
  XNOR2_X1 U15671 ( .A(n14714), .B(n14306), .ZN(n14246) );
  NOR2_X1 U15672 ( .A1(n14246), .A2(n14247), .ZN(n14248) );
  AOI21_X1 U15673 ( .B1(n14247), .B2(n14246), .A(n14248), .ZN(n14333) );
  XNOR2_X1 U15674 ( .A(n14709), .B(n14306), .ZN(n14250) );
  NAND2_X1 U15675 ( .A1(n14582), .A2(n14305), .ZN(n14249) );
  XNOR2_X1 U15676 ( .A(n14250), .B(n14249), .ZN(n14368) );
  INV_X1 U15677 ( .A(n14249), .ZN(n14251) );
  NAND2_X1 U15678 ( .A1(n14605), .A2(n14305), .ZN(n14252) );
  XNOR2_X1 U15679 ( .A(n14253), .B(n14252), .ZN(n14293) );
  XNOR2_X1 U15680 ( .A(n14700), .B(n14254), .ZN(n14256) );
  NAND2_X1 U15681 ( .A1(n14584), .A2(n14305), .ZN(n14255) );
  NAND2_X1 U15682 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  OAI21_X1 U15683 ( .B1(n14256), .B2(n14255), .A(n14257), .ZN(n14352) );
  INV_X1 U15684 ( .A(n14257), .ZN(n14258) );
  NOR2_X1 U15685 ( .A1(n14351), .A2(n14258), .ZN(n14317) );
  XNOR2_X1 U15686 ( .A(n14690), .B(n14306), .ZN(n14261) );
  NAND2_X1 U15687 ( .A1(n14538), .A2(n14305), .ZN(n14259) );
  XNOR2_X1 U15688 ( .A(n14261), .B(n14259), .ZN(n14316) );
  INV_X1 U15689 ( .A(n14259), .ZN(n14260) );
  NAND2_X1 U15692 ( .A1(n14552), .A2(n14305), .ZN(n14359) );
  INV_X1 U15693 ( .A(n14305), .ZN(n14266) );
  NOR2_X1 U15694 ( .A1(n14363), .A2(n14266), .ZN(n14284) );
  NAND2_X1 U15695 ( .A1(n14523), .A2(n14305), .ZN(n14269) );
  XNOR2_X1 U15696 ( .A(n14675), .B(n14306), .ZN(n14268) );
  XOR2_X1 U15697 ( .A(n14269), .B(n14268), .Z(n14342) );
  INV_X1 U15698 ( .A(n14268), .ZN(n14270) );
  XNOR2_X1 U15699 ( .A(n14671), .B(n14306), .ZN(n14272) );
  NAND2_X1 U15700 ( .A1(n14474), .A2(n14305), .ZN(n14271) );
  XNOR2_X1 U15701 ( .A(n14272), .B(n14271), .ZN(n14326) );
  INV_X1 U15702 ( .A(n14271), .ZN(n14273) );
  AND2_X1 U15703 ( .A1(n14395), .A2(n14305), .ZN(n14275) );
  XNOR2_X1 U15704 ( .A(n14664), .B(n14306), .ZN(n14274) );
  NOR2_X1 U15705 ( .A1(n14274), .A2(n14275), .ZN(n14276) );
  AOI21_X1 U15706 ( .B1(n14275), .B2(n14274), .A(n14276), .ZN(n14381) );
  NAND2_X1 U15707 ( .A1(n14380), .A2(n14381), .ZN(n14379) );
  INV_X1 U15708 ( .A(n14276), .ZN(n14277) );
  NAND2_X1 U15709 ( .A1(n14475), .A2(n14305), .ZN(n14301) );
  XNOR2_X1 U15710 ( .A(n14658), .B(n14306), .ZN(n14300) );
  XOR2_X1 U15711 ( .A(n14301), .B(n14300), .Z(n14303) );
  XNOR2_X1 U15712 ( .A(n14304), .B(n14303), .ZN(n14283) );
  OAI22_X1 U15713 ( .A1(n14462), .A2(n14373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14278), .ZN(n14280) );
  NOR2_X1 U15714 ( .A1(n14459), .A2(n14362), .ZN(n14279) );
  AOI211_X1 U15715 ( .C1(n14370), .C2(n14457), .A(n14280), .B(n14279), .ZN(
        n14282) );
  NAND2_X1 U15716 ( .A1(n14658), .A2(n14375), .ZN(n14281) );
  OAI211_X1 U15717 ( .C1(n14283), .C2(n14377), .A(n14282), .B(n14281), .ZN(
        P2_U3186) );
  XNOR2_X1 U15718 ( .A(n14285), .B(n14284), .ZN(n14292) );
  INV_X1 U15719 ( .A(n14529), .ZN(n14287) );
  OAI22_X1 U15720 ( .A1(n14287), .A2(n14373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14286), .ZN(n14290) );
  OAI22_X1 U15721 ( .A1(n14288), .A2(n14387), .B1(n14321), .B2(n14362), .ZN(
        n14289) );
  AOI211_X1 U15722 ( .C1(n14530), .C2(n14375), .A(n14290), .B(n14289), .ZN(
        n14291) );
  OAI21_X1 U15723 ( .B1(n14292), .B2(n14377), .A(n14291), .ZN(P2_U3188) );
  XNOR2_X1 U15724 ( .A(n14294), .B(n14293), .ZN(n14299) );
  OAI22_X1 U15725 ( .A1(n14320), .A2(n14387), .B1(n14362), .B2(n14624), .ZN(
        n14295) );
  AOI211_X1 U15726 ( .C1(n14385), .C2(n14591), .A(n14296), .B(n14295), .ZN(
        n14298) );
  NAND2_X1 U15727 ( .A1(n14704), .A2(n14375), .ZN(n14297) );
  OAI211_X1 U15728 ( .C1(n14299), .C2(n14377), .A(n14298), .B(n14297), .ZN(
        P2_U3191) );
  INV_X1 U15729 ( .A(n14300), .ZN(n14302) );
  MUX2_X1 U15730 ( .A(n14655), .B(n14438), .S(n14305), .Z(n14307) );
  XNOR2_X1 U15731 ( .A(n14307), .B(n14306), .ZN(n14308) );
  XNOR2_X1 U15732 ( .A(n14309), .B(n14308), .ZN(n14315) );
  OAI22_X1 U15733 ( .A1(n14443), .A2(n14373), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14310), .ZN(n14313) );
  INV_X1 U15734 ( .A(n14449), .ZN(n14311) );
  OAI22_X1 U15735 ( .A1(n14311), .A2(n14387), .B1(n14388), .B2(n14362), .ZN(
        n14312) );
  AOI211_X1 U15736 ( .C1(n14655), .C2(n14375), .A(n14313), .B(n14312), .ZN(
        n14314) );
  OAI21_X1 U15737 ( .B1(n14315), .B2(n14377), .A(n14314), .ZN(P2_U3192) );
  XNOR2_X1 U15738 ( .A(n14317), .B(n14316), .ZN(n14325) );
  INV_X1 U15739 ( .A(n14318), .ZN(n14557) );
  OAI22_X1 U15740 ( .A1(n14373), .A2(n14557), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14319), .ZN(n14323) );
  OAI22_X1 U15741 ( .A1(n14321), .A2(n14387), .B1(n14362), .B2(n14320), .ZN(
        n14322) );
  AOI211_X1 U15742 ( .C1(n14690), .C2(n14375), .A(n14323), .B(n14322), .ZN(
        n14324) );
  OAI21_X1 U15743 ( .B1(n14325), .B2(n14377), .A(n14324), .ZN(P2_U3195) );
  XNOR2_X1 U15744 ( .A(n14327), .B(n14326), .ZN(n14332) );
  AOI22_X1 U15745 ( .A1(n14395), .A2(n14583), .B1(n14600), .B2(n14523), .ZN(
        n14489) );
  INV_X1 U15746 ( .A(n14328), .ZN(n14347) );
  AOI22_X1 U15747 ( .A1(n14493), .A2(n14385), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14329) );
  OAI21_X1 U15748 ( .B1(n14489), .B2(n14347), .A(n14329), .ZN(n14330) );
  AOI21_X1 U15749 ( .B1(n14671), .B2(n14375), .A(n14330), .ZN(n14331) );
  OAI21_X1 U15750 ( .B1(n14332), .B2(n14377), .A(n14331), .ZN(P2_U3197) );
  NOR2_X1 U15751 ( .A1(n7666), .A2(n14333), .ZN(n14335) );
  OAI21_X1 U15752 ( .B1(n14336), .B2(n14335), .A(n14382), .ZN(n14341) );
  INV_X1 U15753 ( .A(n14632), .ZN(n14339) );
  OAI22_X1 U15754 ( .A1(n14624), .A2(n14387), .B1(n14362), .B2(n14622), .ZN(
        n14337) );
  AOI211_X1 U15755 ( .C1(n14385), .C2(n14339), .A(n14338), .B(n14337), .ZN(
        n14340) );
  OAI211_X1 U15756 ( .C1(n8169), .C2(n14393), .A(n14341), .B(n14340), .ZN(
        P2_U3200) );
  XNOR2_X1 U15757 ( .A(n14343), .B(n14342), .ZN(n14350) );
  AND2_X1 U15758 ( .A1(n14537), .A2(n14600), .ZN(n14344) );
  AOI21_X1 U15759 ( .B1(n14474), .B2(n14583), .A(n14344), .ZN(n14504) );
  INV_X1 U15760 ( .A(n14345), .ZN(n14512) );
  AOI22_X1 U15761 ( .A1(n14512), .A2(n14385), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14346) );
  OAI21_X1 U15762 ( .B1(n14504), .B2(n14347), .A(n14346), .ZN(n14348) );
  AOI21_X1 U15763 ( .B1(n14675), .B2(n14375), .A(n14348), .ZN(n14349) );
  OAI21_X1 U15764 ( .B1(n14350), .B2(n14377), .A(n14349), .ZN(P2_U3201) );
  AOI21_X1 U15765 ( .B1(n14353), .B2(n14352), .A(n14351), .ZN(n14358) );
  OAI22_X1 U15766 ( .A1(n14373), .A2(n14572), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14354), .ZN(n14356) );
  OAI22_X1 U15767 ( .A1(n14568), .A2(n14362), .B1(n14387), .B2(n14569), .ZN(
        n14355) );
  AOI211_X1 U15768 ( .C1(n14700), .C2(n14375), .A(n14356), .B(n14355), .ZN(
        n14357) );
  OAI21_X1 U15769 ( .B1(n14358), .B2(n14377), .A(n14357), .ZN(P2_U3205) );
  XNOR2_X1 U15770 ( .A(n14360), .B(n14359), .ZN(n14367) );
  OAI22_X1 U15771 ( .A1(n14373), .A2(n14542), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14361), .ZN(n14365) );
  OAI22_X1 U15772 ( .A1(n14363), .A2(n14387), .B1(n14569), .B2(n14362), .ZN(
        n14364) );
  AOI211_X1 U15773 ( .C1(n14686), .C2(n14375), .A(n14365), .B(n14364), .ZN(
        n14366) );
  OAI21_X1 U15774 ( .B1(n14367), .B2(n14377), .A(n14366), .ZN(P2_U3207) );
  XNOR2_X1 U15775 ( .A(n14369), .B(n14368), .ZN(n14378) );
  INV_X1 U15776 ( .A(n14612), .ZN(n14372) );
  AOI22_X1 U15777 ( .A1(n14370), .A2(n14605), .B1(n14390), .B2(n14601), .ZN(
        n14371) );
  NAND2_X1 U15778 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n16172)
         );
  OAI211_X1 U15779 ( .C1(n14373), .C2(n14372), .A(n14371), .B(n16172), .ZN(
        n14374) );
  AOI21_X1 U15780 ( .B1(n14709), .B2(n14375), .A(n14374), .ZN(n14376) );
  OAI21_X1 U15781 ( .B1(n14378), .B2(n14377), .A(n14376), .ZN(P2_U3210) );
  INV_X1 U15782 ( .A(n14664), .ZN(n14480) );
  OAI21_X1 U15783 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(n14383) );
  NAND2_X1 U15784 ( .A1(n14383), .A2(n14382), .ZN(n14392) );
  AOI22_X1 U15785 ( .A1(n14478), .A2(n14385), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14386) );
  OAI21_X1 U15786 ( .B1(n14388), .B2(n14387), .A(n14386), .ZN(n14389) );
  AOI21_X1 U15787 ( .B1(n14390), .B2(n14474), .A(n14389), .ZN(n14391) );
  OAI211_X1 U15788 ( .C1(n14480), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P2_U3212) );
  MUX2_X1 U15789 ( .A(n14394), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14410), .Z(
        P2_U3561) );
  MUX2_X1 U15790 ( .A(n14449), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14410), .Z(
        P2_U3560) );
  MUX2_X1 U15791 ( .A(n14457), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14410), .Z(
        P2_U3559) );
  MUX2_X1 U15792 ( .A(n14475), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14410), .Z(
        P2_U3558) );
  MUX2_X1 U15793 ( .A(n14395), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14410), .Z(
        P2_U3557) );
  MUX2_X1 U15794 ( .A(n14474), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14410), .Z(
        P2_U3556) );
  MUX2_X1 U15795 ( .A(n14523), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14410), .Z(
        P2_U3555) );
  MUX2_X1 U15796 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14552), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15797 ( .A(n14538), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14410), .Z(
        P2_U3552) );
  MUX2_X1 U15798 ( .A(n14584), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14410), .Z(
        P2_U3551) );
  MUX2_X1 U15799 ( .A(n14605), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14410), .Z(
        P2_U3550) );
  MUX2_X1 U15800 ( .A(n14582), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14410), .Z(
        P2_U3549) );
  MUX2_X1 U15801 ( .A(n14601), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14410), .Z(
        P2_U3548) );
  INV_X2 U15802 ( .A(P2_U3947), .ZN(n14410) );
  MUX2_X1 U15803 ( .A(n14396), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14410), .Z(
        P2_U3547) );
  MUX2_X1 U15804 ( .A(n14397), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14410), .Z(
        P2_U3546) );
  MUX2_X1 U15805 ( .A(n14398), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14410), .Z(
        P2_U3545) );
  MUX2_X1 U15806 ( .A(n14399), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14410), .Z(
        P2_U3544) );
  MUX2_X1 U15807 ( .A(n14400), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14410), .Z(
        P2_U3543) );
  MUX2_X1 U15808 ( .A(n14401), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14410), .Z(
        P2_U3542) );
  MUX2_X1 U15809 ( .A(n14402), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14410), .Z(
        P2_U3541) );
  MUX2_X1 U15810 ( .A(n14403), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14410), .Z(
        P2_U3540) );
  MUX2_X1 U15811 ( .A(n14404), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14410), .Z(
        P2_U3539) );
  MUX2_X1 U15812 ( .A(n14405), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14410), .Z(
        P2_U3538) );
  MUX2_X1 U15813 ( .A(n14406), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14410), .Z(
        P2_U3537) );
  MUX2_X1 U15814 ( .A(n14407), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14410), .Z(
        P2_U3536) );
  MUX2_X1 U15815 ( .A(n14408), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14410), .Z(
        P2_U3535) );
  MUX2_X1 U15816 ( .A(n14409), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14410), .Z(
        P2_U3534) );
  MUX2_X1 U15817 ( .A(n9929), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14410), .Z(
        P2_U3533) );
  MUX2_X1 U15818 ( .A(n14411), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14410), .Z(
        P2_U3532) );
  MUX2_X1 U15819 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14412), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI211_X1 U15820 ( .C1(n14415), .C2(n14414), .A(n16163), .B(n14413), .ZN(
        n14423) );
  OAI211_X1 U15821 ( .C1(n14418), .C2(n14417), .A(n16171), .B(n14416), .ZN(
        n14422) );
  AOI22_X1 U15822 ( .A1(n16055), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14421) );
  NAND2_X1 U15823 ( .A1(n16188), .A2(n14419), .ZN(n14420) );
  NAND4_X1 U15824 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        P2_U3215) );
  INV_X1 U15825 ( .A(n14645), .ZN(n14432) );
  XNOR2_X1 U15826 ( .A(n10152), .B(n14430), .ZN(n14641) );
  INV_X1 U15827 ( .A(n14424), .ZN(n14425) );
  NOR2_X1 U15828 ( .A1(n14426), .A2(n14425), .ZN(n14644) );
  NAND2_X1 U15829 ( .A1(n16458), .A2(n14644), .ZN(n14433) );
  OAI21_X1 U15830 ( .B1(n16458), .B2(n14427), .A(n14433), .ZN(n14428) );
  AOI21_X1 U15831 ( .B1(n10152), .B2(n16463), .A(n14428), .ZN(n14429) );
  OAI21_X1 U15832 ( .B1(n14641), .B2(n14561), .A(n14429), .ZN(P2_U3234) );
  OAI21_X1 U15833 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14647) );
  INV_X1 U15834 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14434) );
  OAI21_X1 U15835 ( .B1(n16458), .B2(n14434), .A(n14433), .ZN(n14435) );
  AOI21_X1 U15836 ( .B1(n14645), .B2(n16463), .A(n14435), .ZN(n14436) );
  OAI21_X1 U15837 ( .B1(n14647), .B2(n14561), .A(n14436), .ZN(P2_U3235) );
  OAI21_X1 U15838 ( .B1(n14439), .B2(n14438), .A(n14437), .ZN(n14440) );
  INV_X1 U15839 ( .A(n14440), .ZN(n14656) );
  AOI22_X1 U15840 ( .A1(n14655), .A2(n16463), .B1(n14598), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n14454) );
  AOI211_X1 U15841 ( .C1(n14655), .C2(n14442), .A(n14692), .B(n8163), .ZN(
        n14654) );
  INV_X1 U15842 ( .A(n14654), .ZN(n14445) );
  OAI22_X1 U15843 ( .A1(n14445), .A2(n14444), .B1(n16455), .B2(n14443), .ZN(
        n14452) );
  OAI211_X1 U15844 ( .C1(n14448), .C2(n14447), .A(n14446), .B(n14603), .ZN(
        n14451) );
  AOI22_X1 U15845 ( .A1(n14583), .A2(n14449), .B1(n14475), .B2(n14600), .ZN(
        n14450) );
  OAI21_X1 U15846 ( .B1(n14452), .B2(n14653), .A(n16458), .ZN(n14453) );
  OAI211_X1 U15847 ( .C1(n14656), .C2(n14638), .A(n14454), .B(n14453), .ZN(
        P2_U3237) );
  XNOR2_X1 U15848 ( .A(n14456), .B(n14455), .ZN(n14461) );
  NAND2_X1 U15849 ( .A1(n14457), .A2(n14604), .ZN(n14458) );
  OAI21_X1 U15850 ( .B1(n14459), .B2(n14621), .A(n14458), .ZN(n14460) );
  AOI21_X1 U15851 ( .B1(n14461), .B2(n14603), .A(n14460), .ZN(n14661) );
  XNOR2_X1 U15852 ( .A(n14477), .B(n14658), .ZN(n14659) );
  INV_X1 U15853 ( .A(n14462), .ZN(n14463) );
  AOI22_X1 U15854 ( .A1(n14463), .A2(n14611), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14598), .ZN(n14464) );
  OAI21_X1 U15855 ( .B1(n14465), .B2(n14631), .A(n14464), .ZN(n14466) );
  AOI21_X1 U15856 ( .B1(n14659), .B2(n16452), .A(n14466), .ZN(n14471) );
  INV_X1 U15857 ( .A(n14662), .ZN(n14469) );
  OR2_X1 U15858 ( .A1(n14468), .A2(n14467), .ZN(n14657) );
  NAND3_X1 U15859 ( .A1(n14469), .A2(n14617), .A3(n14657), .ZN(n14470) );
  OAI211_X1 U15860 ( .C1(n14661), .C2(n14598), .A(n14471), .B(n14470), .ZN(
        P2_U3238) );
  XNOR2_X1 U15861 ( .A(n14473), .B(n14472), .ZN(n14476) );
  AOI222_X1 U15862 ( .A1(n14476), .A2(n14603), .B1(n14475), .B2(n14583), .C1(
        n14474), .C2(n14600), .ZN(n14667) );
  AOI21_X1 U15863 ( .B1(n14664), .B2(n14491), .A(n14477), .ZN(n14665) );
  AOI22_X1 U15864 ( .A1(n14478), .A2(n14611), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14598), .ZN(n14479) );
  OAI21_X1 U15865 ( .B1(n14480), .B2(n14631), .A(n14479), .ZN(n14484) );
  XNOR2_X1 U15866 ( .A(n14482), .B(n14481), .ZN(n14668) );
  NOR2_X1 U15867 ( .A1(n14668), .A2(n14638), .ZN(n14483) );
  AOI211_X1 U15868 ( .C1(n16452), .C2(n14665), .A(n14484), .B(n14483), .ZN(
        n14485) );
  OAI21_X1 U15869 ( .B1(n14598), .B2(n14667), .A(n14485), .ZN(P2_U3239) );
  XOR2_X1 U15870 ( .A(n14486), .B(n14487), .Z(n14673) );
  XOR2_X1 U15871 ( .A(n14488), .B(n14487), .Z(n14490) );
  OAI21_X1 U15872 ( .B1(n14490), .B2(n14619), .A(n14489), .ZN(n14669) );
  NAND2_X1 U15873 ( .A1(n14669), .A2(n16458), .ZN(n14498) );
  INV_X1 U15874 ( .A(n14491), .ZN(n14492) );
  AOI211_X1 U15875 ( .C1(n14671), .C2(n14499), .A(n14692), .B(n14492), .ZN(
        n14670) );
  INV_X1 U15876 ( .A(n14671), .ZN(n14495) );
  AOI22_X1 U15877 ( .A1(n14493), .A2(n14611), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14598), .ZN(n14494) );
  OAI21_X1 U15878 ( .B1(n14495), .B2(n14631), .A(n14494), .ZN(n14496) );
  AOI21_X1 U15879 ( .B1(n14670), .B2(n14596), .A(n14496), .ZN(n14497) );
  OAI211_X1 U15880 ( .C1(n14638), .C2(n14673), .A(n14498), .B(n14497), .ZN(
        P2_U3240) );
  INV_X1 U15881 ( .A(n14527), .ZN(n14501) );
  INV_X1 U15882 ( .A(n14499), .ZN(n14500) );
  AOI211_X1 U15883 ( .C1(n14675), .C2(n14501), .A(n14692), .B(n14500), .ZN(
        n14674) );
  XNOR2_X1 U15884 ( .A(n14503), .B(n14502), .ZN(n14506) );
  INV_X1 U15885 ( .A(n14504), .ZN(n14505) );
  AOI21_X1 U15886 ( .B1(n14506), .B2(n14603), .A(n14505), .ZN(n14676) );
  INV_X1 U15887 ( .A(n14676), .ZN(n14507) );
  AOI21_X1 U15888 ( .B1(n14674), .B2(n14508), .A(n14507), .ZN(n14518) );
  OAI21_X1 U15889 ( .B1(n14511), .B2(n14510), .A(n14509), .ZN(n14678) );
  INV_X1 U15890 ( .A(n14678), .ZN(n14516) );
  AOI22_X1 U15891 ( .A1(n14512), .A2(n14611), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14598), .ZN(n14513) );
  OAI21_X1 U15892 ( .B1(n14514), .B2(n14631), .A(n14513), .ZN(n14515) );
  AOI21_X1 U15893 ( .B1(n14516), .B2(n14617), .A(n14515), .ZN(n14517) );
  OAI21_X1 U15894 ( .B1(n14518), .B2(n14598), .A(n14517), .ZN(P2_U3241) );
  XNOR2_X1 U15895 ( .A(n14519), .B(n14520), .ZN(n14526) );
  XNOR2_X1 U15896 ( .A(n14521), .B(n14520), .ZN(n14683) );
  NAND2_X1 U15897 ( .A1(n14683), .A2(n14522), .ZN(n14525) );
  AOI22_X1 U15898 ( .A1(n14523), .A2(n14583), .B1(n14600), .B2(n14552), .ZN(
        n14524) );
  OAI211_X1 U15899 ( .C1(n14619), .C2(n14526), .A(n14525), .B(n14524), .ZN(
        n14681) );
  INV_X1 U15900 ( .A(n14681), .ZN(n14535) );
  AND2_X1 U15901 ( .A1(n14530), .A2(n14540), .ZN(n14528) );
  OR2_X1 U15902 ( .A1(n14528), .A2(n14527), .ZN(n14680) );
  AOI22_X1 U15903 ( .A1(n14598), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14529), 
        .B2(n14611), .ZN(n14532) );
  NAND2_X1 U15904 ( .A1(n14530), .A2(n16463), .ZN(n14531) );
  OAI211_X1 U15905 ( .C1(n14680), .C2(n14561), .A(n14532), .B(n14531), .ZN(
        n14533) );
  AOI21_X1 U15906 ( .B1(n14683), .B2(n16453), .A(n14533), .ZN(n14534) );
  OAI21_X1 U15907 ( .B1(n14535), .B2(n14598), .A(n14534), .ZN(P2_U3242) );
  XOR2_X1 U15908 ( .A(n14545), .B(n14536), .Z(n14539) );
  AOI222_X1 U15909 ( .A1(n14539), .A2(n14603), .B1(n14538), .B2(n14600), .C1(
        n14537), .C2(n14583), .ZN(n14688) );
  INV_X1 U15910 ( .A(n14540), .ZN(n14541) );
  AOI211_X1 U15911 ( .C1(n14686), .C2(n14556), .A(n14692), .B(n14541), .ZN(
        n14685) );
  INV_X1 U15912 ( .A(n14542), .ZN(n14543) );
  AOI22_X1 U15913 ( .A1(n14598), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14543), 
        .B2(n14611), .ZN(n14544) );
  OAI21_X1 U15914 ( .B1(n8165), .B2(n14631), .A(n14544), .ZN(n14548) );
  XNOR2_X1 U15915 ( .A(n14546), .B(n14545), .ZN(n14689) );
  NOR2_X1 U15916 ( .A1(n14689), .A2(n14638), .ZN(n14547) );
  AOI211_X1 U15917 ( .C1(n14685), .C2(n14596), .A(n14548), .B(n14547), .ZN(
        n14549) );
  OAI21_X1 U15918 ( .B1(n14598), .B2(n14688), .A(n14549), .ZN(P2_U3243) );
  XOR2_X1 U15919 ( .A(n14550), .B(n14553), .Z(n14551) );
  AOI222_X1 U15920 ( .A1(n14552), .A2(n14583), .B1(n14603), .B2(n14551), .C1(
        n14584), .C2(n14600), .ZN(n14697) );
  XNOR2_X1 U15921 ( .A(n14554), .B(n14553), .ZN(n14695) );
  NAND2_X1 U15922 ( .A1(n14690), .A2(n14570), .ZN(n14555) );
  NAND2_X1 U15923 ( .A1(n14556), .A2(n14555), .ZN(n14693) );
  INV_X1 U15924 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14558) );
  OAI22_X1 U15925 ( .A1(n16458), .A2(n14558), .B1(n14557), .B2(n16455), .ZN(
        n14559) );
  AOI21_X1 U15926 ( .B1(n14690), .B2(n16463), .A(n14559), .ZN(n14560) );
  OAI21_X1 U15927 ( .B1(n14693), .B2(n14561), .A(n14560), .ZN(n14562) );
  AOI21_X1 U15928 ( .B1(n14695), .B2(n14617), .A(n14562), .ZN(n14563) );
  OAI21_X1 U15929 ( .B1(n14697), .B2(n14598), .A(n14563), .ZN(P2_U3244) );
  XNOR2_X1 U15930 ( .A(n14564), .B(n14566), .ZN(n14702) );
  AOI21_X1 U15931 ( .B1(n14566), .B2(n14565), .A(n7477), .ZN(n14567) );
  OAI222_X1 U15932 ( .A1(n14623), .A2(n14569), .B1(n14621), .B2(n14568), .C1(
        n14567), .C2(n14619), .ZN(n14698) );
  AOI21_X1 U15933 ( .B1(n14700), .B2(n14589), .A(n14692), .ZN(n14571) );
  AND2_X1 U15934 ( .A1(n14571), .A2(n14570), .ZN(n14699) );
  NAND2_X1 U15935 ( .A1(n14699), .A2(n14596), .ZN(n14576) );
  INV_X1 U15936 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n14573) );
  OAI22_X1 U15937 ( .A1(n16458), .A2(n14573), .B1(n14572), .B2(n16455), .ZN(
        n14574) );
  AOI21_X1 U15938 ( .B1(n14700), .B2(n16463), .A(n14574), .ZN(n14575) );
  NAND2_X1 U15939 ( .A1(n14576), .A2(n14575), .ZN(n14577) );
  AOI21_X1 U15940 ( .B1(n14698), .B2(n16458), .A(n14577), .ZN(n14578) );
  OAI21_X1 U15941 ( .B1(n14638), .B2(n14702), .A(n14578), .ZN(P2_U3245) );
  XNOR2_X1 U15942 ( .A(n14579), .B(n8066), .ZN(n14588) );
  OAI21_X1 U15943 ( .B1(n14581), .B2(n8066), .A(n14580), .ZN(n14707) );
  AOI22_X1 U15944 ( .A1(n14584), .A2(n14583), .B1(n14600), .B2(n14582), .ZN(
        n14585) );
  OAI21_X1 U15945 ( .B1(n14707), .B2(n14586), .A(n14585), .ZN(n14587) );
  AOI21_X1 U15946 ( .B1(n14588), .B2(n14603), .A(n14587), .ZN(n14706) );
  INV_X1 U15947 ( .A(n14589), .ZN(n14590) );
  AOI211_X1 U15948 ( .C1(n14704), .C2(n14609), .A(n14692), .B(n14590), .ZN(
        n14703) );
  AOI22_X1 U15949 ( .A1(n14598), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14591), 
        .B2(n14611), .ZN(n14592) );
  OAI21_X1 U15950 ( .B1(n8167), .B2(n14631), .A(n14592), .ZN(n14595) );
  NOR2_X1 U15951 ( .A1(n14707), .A2(n14593), .ZN(n14594) );
  AOI211_X1 U15952 ( .C1(n14703), .C2(n14596), .A(n14595), .B(n14594), .ZN(
        n14597) );
  OAI21_X1 U15953 ( .B1(n14598), .B2(n14706), .A(n14597), .ZN(P2_U3246) );
  XNOR2_X1 U15954 ( .A(n14599), .B(n14607), .ZN(n14602) );
  AOI222_X1 U15955 ( .A1(n14605), .A2(n14604), .B1(n14603), .B2(n14602), .C1(
        n14601), .C2(n14600), .ZN(n14712) );
  OAI21_X1 U15956 ( .B1(n14608), .B2(n14607), .A(n7641), .ZN(n14708) );
  INV_X1 U15957 ( .A(n14709), .ZN(n14615) );
  INV_X1 U15958 ( .A(n14609), .ZN(n14610) );
  AOI21_X1 U15959 ( .B1(n14709), .B2(n14628), .A(n14610), .ZN(n14710) );
  NAND2_X1 U15960 ( .A1(n14710), .A2(n16452), .ZN(n14614) );
  AOI22_X1 U15961 ( .A1(n14598), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14612), 
        .B2(n14611), .ZN(n14613) );
  OAI211_X1 U15962 ( .C1(n14615), .C2(n14631), .A(n14614), .B(n14613), .ZN(
        n14616) );
  AOI21_X1 U15963 ( .B1(n14708), .B2(n14617), .A(n14616), .ZN(n14618) );
  OAI21_X1 U15964 ( .B1(n14712), .B2(n14598), .A(n14618), .ZN(P2_U3247) );
  AOI21_X1 U15965 ( .B1(n14620), .B2(n14636), .A(n14619), .ZN(n14627) );
  OAI22_X1 U15966 ( .A1(n14624), .A2(n14623), .B1(n14622), .B2(n14621), .ZN(
        n14625) );
  AOI21_X1 U15967 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14717) );
  INV_X1 U15968 ( .A(n14628), .ZN(n14629) );
  AOI21_X1 U15969 ( .B1(n14714), .B2(n14630), .A(n14629), .ZN(n14715) );
  NOR2_X1 U15970 ( .A1(n8169), .A2(n14631), .ZN(n14635) );
  OAI22_X1 U15971 ( .A1(n16458), .A2(n14633), .B1(n14632), .B2(n16455), .ZN(
        n14634) );
  AOI211_X1 U15972 ( .C1(n14715), .C2(n16452), .A(n14635), .B(n14634), .ZN(
        n14640) );
  XNOR2_X1 U15973 ( .A(n14637), .B(n14636), .ZN(n14718) );
  OR2_X1 U15974 ( .A1(n14718), .A2(n14638), .ZN(n14639) );
  OAI211_X1 U15975 ( .C1(n14717), .C2(n14598), .A(n14640), .B(n14639), .ZN(
        P2_U3248) );
  AOI21_X1 U15976 ( .B1(n10152), .B2(n14733), .A(n14644), .ZN(n14642) );
  NAND2_X1 U15977 ( .A1(n14643), .A2(n14642), .ZN(n14742) );
  MUX2_X1 U15978 ( .A(n14742), .B(P2_REG1_REG_31__SCAN_IN), .S(n16412), .Z(
        P2_U3530) );
  AOI21_X1 U15979 ( .B1(n14645), .B2(n14733), .A(n14644), .ZN(n14646) );
  OAI21_X1 U15980 ( .B1(n14647), .B2(n14692), .A(n14646), .ZN(n14743) );
  MUX2_X1 U15981 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14743), .S(n16413), .Z(
        P2_U3529) );
  AOI21_X1 U15982 ( .B1(n14733), .B2(n14649), .A(n14648), .ZN(n14650) );
  MUX2_X1 U15983 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14744), .S(n16413), .Z(
        P2_U3528) );
  NAND2_X1 U15984 ( .A1(n14657), .A2(n16374), .ZN(n14663) );
  AOI22_X1 U15985 ( .A1(n14659), .A2(n14734), .B1(n14733), .B2(n14658), .ZN(
        n14660) );
  OAI211_X1 U15986 ( .C1(n14663), .C2(n14662), .A(n14661), .B(n14660), .ZN(
        n14746) );
  MUX2_X1 U15987 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14746), .S(n16413), .Z(
        P2_U3526) );
  AOI22_X1 U15988 ( .A1(n14665), .A2(n14734), .B1(n14733), .B2(n14664), .ZN(
        n14666) );
  OAI211_X1 U15989 ( .C1(n14739), .C2(n14668), .A(n14667), .B(n14666), .ZN(
        n14747) );
  MUX2_X1 U15990 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14747), .S(n16413), .Z(
        P2_U3525) );
  AOI211_X1 U15991 ( .C1(n14733), .C2(n14671), .A(n14670), .B(n14669), .ZN(
        n14672) );
  OAI21_X1 U15992 ( .B1(n14739), .B2(n14673), .A(n14672), .ZN(n14748) );
  MUX2_X1 U15993 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14748), .S(n16413), .Z(
        P2_U3524) );
  AOI21_X1 U15994 ( .B1(n14733), .B2(n14675), .A(n14674), .ZN(n14677) );
  OAI211_X1 U15995 ( .C1(n14739), .C2(n14678), .A(n14677), .B(n14676), .ZN(
        n14749) );
  MUX2_X1 U15996 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14749), .S(n16413), .Z(
        P2_U3523) );
  OAI22_X1 U15997 ( .A1(n14680), .A2(n14692), .B1(n14679), .B2(n16407), .ZN(
        n14682) );
  AOI211_X1 U15998 ( .C1(n11199), .C2(n14683), .A(n14682), .B(n14681), .ZN(
        n14684) );
  INV_X1 U15999 ( .A(n14684), .ZN(n14750) );
  MUX2_X1 U16000 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14750), .S(n16413), .Z(
        P2_U3522) );
  AOI21_X1 U16001 ( .B1(n14733), .B2(n14686), .A(n14685), .ZN(n14687) );
  OAI211_X1 U16002 ( .C1(n14739), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        n14751) );
  MUX2_X1 U16003 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14751), .S(n16413), .Z(
        P2_U3521) );
  INV_X1 U16004 ( .A(n14690), .ZN(n14691) );
  OAI22_X1 U16005 ( .A1(n14693), .A2(n14692), .B1(n14691), .B2(n16407), .ZN(
        n14694) );
  AOI21_X1 U16006 ( .B1(n14695), .B2(n16374), .A(n14694), .ZN(n14696) );
  NAND2_X1 U16007 ( .A1(n14697), .A2(n14696), .ZN(n14752) );
  MUX2_X1 U16008 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14752), .S(n16413), .Z(
        P2_U3520) );
  AOI211_X1 U16009 ( .C1(n14733), .C2(n14700), .A(n14699), .B(n14698), .ZN(
        n14701) );
  OAI21_X1 U16010 ( .B1(n14739), .B2(n14702), .A(n14701), .ZN(n14753) );
  MUX2_X1 U16011 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14753), .S(n16413), .Z(
        P2_U3519) );
  AOI21_X1 U16012 ( .B1(n14733), .B2(n14704), .A(n14703), .ZN(n14705) );
  OAI211_X1 U16013 ( .C1(n16299), .C2(n14707), .A(n14706), .B(n14705), .ZN(
        n14754) );
  MUX2_X1 U16014 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14754), .S(n16413), .Z(
        P2_U3518) );
  INV_X1 U16015 ( .A(n14708), .ZN(n14713) );
  AOI22_X1 U16016 ( .A1(n14710), .A2(n14734), .B1(n14733), .B2(n14709), .ZN(
        n14711) );
  OAI211_X1 U16017 ( .C1(n14739), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14755) );
  MUX2_X1 U16018 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14755), .S(n16413), .Z(
        P2_U3517) );
  AOI22_X1 U16019 ( .A1(n14715), .A2(n14734), .B1(n14733), .B2(n14714), .ZN(
        n14716) );
  OAI211_X1 U16020 ( .C1(n14739), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14756) );
  MUX2_X1 U16021 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14756), .S(n16413), .Z(
        P2_U3516) );
  AOI22_X1 U16022 ( .A1(n14720), .A2(n14734), .B1(n14733), .B2(n14719), .ZN(
        n14721) );
  OAI21_X1 U16023 ( .B1(n14722), .B2(n16299), .A(n14721), .ZN(n14723) );
  NOR2_X1 U16024 ( .A1(n14724), .A2(n14723), .ZN(n14757) );
  INV_X1 U16025 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n14725) );
  MUX2_X1 U16026 ( .A(n14757), .B(n14725), .S(n16412), .Z(n14726) );
  INV_X1 U16027 ( .A(n14726), .ZN(P2_U3515) );
  AOI21_X1 U16028 ( .B1(n14733), .B2(n14728), .A(n14727), .ZN(n14729) );
  OAI211_X1 U16029 ( .C1(n14731), .C2(n16299), .A(n14730), .B(n14729), .ZN(
        n14759) );
  MUX2_X1 U16030 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14759), .S(n16413), .Z(
        P2_U3514) );
  AOI22_X1 U16031 ( .A1(n14735), .A2(n14734), .B1(n14733), .B2(n14732), .ZN(
        n14736) );
  OAI211_X1 U16032 ( .C1(n14739), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        n14761) );
  NAND2_X1 U16033 ( .A1(n14761), .A2(n16413), .ZN(n14740) );
  OAI21_X1 U16034 ( .B1(n16413), .B2(n12068), .A(n14740), .ZN(P2_U3513) );
  MUX2_X1 U16035 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n14741), .S(n16413), .Z(
        P2_U3501) );
  MUX2_X1 U16036 ( .A(n14742), .B(P2_REG0_REG_31__SCAN_IN), .S(n16414), .Z(
        P2_U3498) );
  MUX2_X1 U16037 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14743), .S(n14760), .Z(
        P2_U3497) );
  MUX2_X1 U16038 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14744), .S(n14760), .Z(
        P2_U3496) );
  MUX2_X1 U16039 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14745), .S(n14760), .Z(
        P2_U3495) );
  MUX2_X1 U16040 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14746), .S(n14760), .Z(
        P2_U3494) );
  MUX2_X1 U16041 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14747), .S(n14760), .Z(
        P2_U3493) );
  MUX2_X1 U16042 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14748), .S(n14760), .Z(
        P2_U3492) );
  MUX2_X1 U16043 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14749), .S(n14760), .Z(
        P2_U3491) );
  MUX2_X1 U16044 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14750), .S(n14760), .Z(
        P2_U3490) );
  MUX2_X1 U16045 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14751), .S(n14760), .Z(
        P2_U3489) );
  MUX2_X1 U16046 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14752), .S(n14760), .Z(
        P2_U3488) );
  MUX2_X1 U16047 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14753), .S(n14760), .Z(
        P2_U3487) );
  MUX2_X1 U16048 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14754), .S(n14760), .Z(
        P2_U3486) );
  MUX2_X1 U16049 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14755), .S(n14760), .Z(
        P2_U3484) );
  MUX2_X1 U16050 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14756), .S(n14760), .Z(
        P2_U3481) );
  INV_X1 U16051 ( .A(n14757), .ZN(n14758) );
  MUX2_X1 U16052 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14758), .S(n14760), .Z(
        P2_U3478) );
  MUX2_X1 U16053 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14759), .S(n14760), .Z(
        P2_U3475) );
  NAND2_X1 U16054 ( .A1(n14761), .A2(n14760), .ZN(n14762) );
  OAI21_X1 U16055 ( .B1(n14760), .B2(n9600), .A(n14762), .ZN(P2_U3472) );
  NAND3_X1 U16056 ( .A1(n14763), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14764) );
  OAI22_X1 U16057 ( .A1(n14765), .A2(n14764), .B1(n10136), .B2(n14783), .ZN(
        n14766) );
  AOI21_X1 U16058 ( .B1(n10701), .B2(n14771), .A(n14766), .ZN(n14767) );
  INV_X1 U16059 ( .A(n14767), .ZN(P2_U3296) );
  INV_X1 U16060 ( .A(n14768), .ZN(n15620) );
  OAI222_X1 U16061 ( .A1(n14780), .A2(n15620), .B1(n14770), .B2(P2_U3088), 
        .C1(n14769), .C2(n14783), .ZN(P2_U3298) );
  NAND2_X1 U16062 ( .A1(n14772), .A2(n14771), .ZN(n14774) );
  OAI211_X1 U16063 ( .C1(n14783), .C2(n14775), .A(n14774), .B(n14773), .ZN(
        P2_U3299) );
  INV_X1 U16064 ( .A(n14776), .ZN(n15623) );
  OAI222_X1 U16065 ( .A1(n14780), .A2(n15623), .B1(n14778), .B2(P2_U3088), 
        .C1(n14777), .C2(n14783), .ZN(P2_U3300) );
  INV_X1 U16066 ( .A(n14779), .ZN(n15626) );
  OAI222_X1 U16067 ( .A1(n14783), .A2(n14782), .B1(n14781), .B2(P2_U3088), 
        .C1(n14780), .C2(n15626), .ZN(P2_U3301) );
  MUX2_X1 U16068 ( .A(n7554), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16069 ( .A1(n15489), .A2(n11013), .ZN(n14785) );
  NAND2_X1 U16070 ( .A1(n15217), .A2(n14831), .ZN(n14784) );
  NAND2_X1 U16071 ( .A1(n14785), .A2(n14784), .ZN(n14786) );
  XNOR2_X1 U16072 ( .A(n14786), .B(n11130), .ZN(n14790) );
  NAND2_X1 U16073 ( .A1(n15489), .A2(n14831), .ZN(n14788) );
  NAND2_X1 U16074 ( .A1(n15217), .A2(n12699), .ZN(n14787) );
  NAND2_X1 U16075 ( .A1(n14788), .A2(n14787), .ZN(n14789) );
  NOR2_X1 U16076 ( .A1(n14790), .A2(n14789), .ZN(n14929) );
  AOI21_X1 U16077 ( .B1(n14790), .B2(n14789), .A(n14929), .ZN(n14885) );
  AOI22_X1 U16078 ( .A1(n15509), .A2(n14831), .B1(n12699), .B2(n15183), .ZN(
        n14863) );
  INV_X1 U16079 ( .A(n14863), .ZN(n14865) );
  NAND2_X1 U16080 ( .A1(n15509), .A2(n14856), .ZN(n14792) );
  NAND2_X1 U16081 ( .A1(n15183), .A2(n14831), .ZN(n14791) );
  NAND2_X1 U16082 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  XNOR2_X1 U16083 ( .A(n14793), .B(n11130), .ZN(n14864) );
  OAI22_X1 U16084 ( .A1(n15329), .A2(n14935), .B1(n15197), .B2(n14934), .ZN(
        n14855) );
  OAI22_X1 U16085 ( .A1(n15329), .A2(n14932), .B1(n15197), .B2(n14935), .ZN(
        n14794) );
  XNOR2_X1 U16086 ( .A(n14794), .B(n11130), .ZN(n14854) );
  OAI22_X1 U16087 ( .A1(n15360), .A2(n14935), .B1(n15182), .B2(n14934), .ZN(
        n14848) );
  OAI22_X1 U16088 ( .A1(n15360), .A2(n14932), .B1(n15182), .B2(n14935), .ZN(
        n14795) );
  XNOR2_X1 U16089 ( .A(n14795), .B(n11130), .ZN(n14847) );
  NAND2_X1 U16090 ( .A1(n15396), .A2(n11013), .ZN(n14797) );
  NAND2_X1 U16091 ( .A1(n15370), .A2(n14831), .ZN(n14796) );
  NAND2_X1 U16092 ( .A1(n14797), .A2(n14796), .ZN(n14798) );
  XNOR2_X1 U16093 ( .A(n14798), .B(n11130), .ZN(n14839) );
  OAI22_X1 U16094 ( .A1(n15545), .A2(n14935), .B1(n15411), .B2(n14934), .ZN(
        n14838) );
  INV_X1 U16095 ( .A(n14799), .ZN(n14801) );
  NAND2_X1 U16096 ( .A1(n15579), .A2(n14856), .ZN(n14805) );
  NAND2_X1 U16097 ( .A1(n15047), .A2(n14831), .ZN(n14804) );
  NAND2_X1 U16098 ( .A1(n14805), .A2(n14804), .ZN(n14806) );
  XNOR2_X1 U16099 ( .A(n14806), .B(n11130), .ZN(n14810) );
  NAND2_X1 U16100 ( .A1(n15579), .A2(n14831), .ZN(n14808) );
  NAND2_X1 U16101 ( .A1(n15047), .A2(n14817), .ZN(n14807) );
  NAND2_X1 U16102 ( .A1(n14808), .A2(n14807), .ZN(n14809) );
  NOR2_X1 U16103 ( .A1(n14810), .A2(n14809), .ZN(n14811) );
  AOI21_X1 U16104 ( .B1(n14810), .B2(n14809), .A(n14811), .ZN(n14893) );
  INV_X1 U16105 ( .A(n14811), .ZN(n14812) );
  NAND2_X1 U16106 ( .A1(n15571), .A2(n14856), .ZN(n14814) );
  NAND2_X1 U16107 ( .A1(n15175), .A2(n14831), .ZN(n14813) );
  NAND2_X1 U16108 ( .A1(n14814), .A2(n14813), .ZN(n14815) );
  XNOR2_X1 U16109 ( .A(n14815), .B(n11130), .ZN(n14818) );
  AOI22_X1 U16110 ( .A1(n15571), .A2(n14831), .B1(n14817), .B2(n15175), .ZN(
        n15033) );
  NAND2_X1 U16111 ( .A1(n15562), .A2(n14856), .ZN(n14821) );
  NAND2_X1 U16112 ( .A1(n15177), .A2(n14831), .ZN(n14820) );
  NAND2_X1 U16113 ( .A1(n14821), .A2(n14820), .ZN(n14822) );
  XNOR2_X1 U16114 ( .A(n14822), .B(n12183), .ZN(n14825) );
  AND2_X1 U16115 ( .A1(n15177), .A2(n14817), .ZN(n14823) );
  AOI21_X1 U16116 ( .B1(n15562), .B2(n14831), .A(n14823), .ZN(n14824) );
  NAND2_X1 U16117 ( .A1(n14825), .A2(n14824), .ZN(n14826) );
  OAI21_X1 U16118 ( .B1(n14825), .B2(n14824), .A(n14826), .ZN(n14964) );
  INV_X1 U16119 ( .A(n14826), .ZN(n14972) );
  NAND2_X1 U16120 ( .A1(n15555), .A2(n11013), .ZN(n14828) );
  NAND2_X1 U16121 ( .A1(n15385), .A2(n14831), .ZN(n14827) );
  NAND2_X1 U16122 ( .A1(n14828), .A2(n14827), .ZN(n14829) );
  XNOR2_X1 U16123 ( .A(n14829), .B(n12183), .ZN(n14832) );
  AND2_X1 U16124 ( .A1(n15385), .A2(n14817), .ZN(n14830) );
  AOI21_X1 U16125 ( .B1(n15555), .B2(n14831), .A(n14830), .ZN(n14833) );
  NAND2_X1 U16126 ( .A1(n14832), .A2(n14833), .ZN(n14837) );
  INV_X1 U16127 ( .A(n14832), .ZN(n14835) );
  INV_X1 U16128 ( .A(n14833), .ZN(n14834) );
  NAND2_X1 U16129 ( .A1(n14835), .A2(n14834), .ZN(n14836) );
  AND2_X1 U16130 ( .A1(n14837), .A2(n14836), .ZN(n14971) );
  NAND2_X1 U16131 ( .A1(n14970), .A2(n14837), .ZN(n15010) );
  XOR2_X1 U16132 ( .A(n14838), .B(n14839), .Z(n15011) );
  NAND2_X1 U16133 ( .A1(n15010), .A2(n15011), .ZN(n15009) );
  NAND2_X1 U16134 ( .A1(n15538), .A2(n11013), .ZN(n14841) );
  NAND2_X1 U16135 ( .A1(n15387), .A2(n14831), .ZN(n14840) );
  NAND2_X1 U16136 ( .A1(n14841), .A2(n14840), .ZN(n14842) );
  XNOR2_X1 U16137 ( .A(n14842), .B(n11130), .ZN(n14846) );
  NAND2_X1 U16138 ( .A1(n15538), .A2(n11694), .ZN(n14844) );
  NAND2_X1 U16139 ( .A1(n15387), .A2(n12699), .ZN(n14843) );
  NAND2_X1 U16140 ( .A1(n14844), .A2(n14843), .ZN(n14845) );
  NAND2_X1 U16141 ( .A1(n14846), .A2(n14845), .ZN(n14921) );
  NOR2_X1 U16142 ( .A1(n14846), .A2(n14845), .ZN(n14920) );
  XOR2_X1 U16143 ( .A(n14848), .B(n14847), .Z(n14991) );
  AOI22_X1 U16144 ( .A1(n15528), .A2(n11013), .B1(n11694), .B2(n15319), .ZN(
        n14849) );
  XNOR2_X1 U16145 ( .A(n14849), .B(n11130), .ZN(n14850) );
  AOI22_X1 U16146 ( .A1(n15528), .A2(n14831), .B1(n12699), .B2(n15319), .ZN(
        n14851) );
  XNOR2_X1 U16147 ( .A(n14850), .B(n14851), .ZN(n14947) );
  INV_X1 U16148 ( .A(n14850), .ZN(n14853) );
  INV_X1 U16149 ( .A(n14851), .ZN(n14852) );
  XOR2_X1 U16150 ( .A(n14855), .B(n14854), .Z(n15001) );
  NAND2_X1 U16151 ( .A1(n15517), .A2(n14856), .ZN(n14858) );
  NAND2_X1 U16152 ( .A1(n15320), .A2(n14831), .ZN(n14857) );
  NAND2_X1 U16153 ( .A1(n14858), .A2(n14857), .ZN(n14859) );
  XNOR2_X1 U16154 ( .A(n14859), .B(n11130), .ZN(n14861) );
  OAI22_X1 U16155 ( .A1(n15313), .A2(n14935), .B1(n8435), .B2(n14934), .ZN(
        n14860) );
  XNOR2_X1 U16156 ( .A(n14861), .B(n14860), .ZN(n14906) );
  XNOR2_X1 U16157 ( .A(n14864), .B(n14863), .ZN(n14983) );
  NAND2_X1 U16158 ( .A1(n15501), .A2(n11013), .ZN(n14867) );
  NAND2_X1 U16159 ( .A1(n15290), .A2(n11694), .ZN(n14866) );
  NAND2_X1 U16160 ( .A1(n14867), .A2(n14866), .ZN(n14868) );
  XNOR2_X1 U16161 ( .A(n14868), .B(n11130), .ZN(n14869) );
  AOI22_X1 U16162 ( .A1(n15501), .A2(n14831), .B1(n12699), .B2(n15290), .ZN(
        n14870) );
  XNOR2_X1 U16163 ( .A(n14869), .B(n14870), .ZN(n14955) );
  NAND2_X1 U16164 ( .A1(n14954), .A2(n14955), .ZN(n14873) );
  INV_X1 U16165 ( .A(n14869), .ZN(n14871) );
  NAND2_X1 U16166 ( .A1(n14871), .A2(n14870), .ZN(n14872) );
  NAND2_X1 U16167 ( .A1(n14873), .A2(n14872), .ZN(n15023) );
  NAND2_X1 U16168 ( .A1(n15495), .A2(n11013), .ZN(n14875) );
  NAND2_X1 U16169 ( .A1(n15046), .A2(n11694), .ZN(n14874) );
  NAND2_X1 U16170 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  XNOR2_X1 U16171 ( .A(n14876), .B(n11130), .ZN(n14879) );
  NAND2_X1 U16172 ( .A1(n15495), .A2(n14831), .ZN(n14878) );
  NAND2_X1 U16173 ( .A1(n15046), .A2(n12699), .ZN(n14877) );
  NAND2_X1 U16174 ( .A1(n14878), .A2(n14877), .ZN(n14880) );
  NAND2_X1 U16175 ( .A1(n14879), .A2(n14880), .ZN(n15020) );
  NAND2_X1 U16176 ( .A1(n15023), .A2(n15020), .ZN(n14883) );
  INV_X1 U16177 ( .A(n14879), .ZN(n14882) );
  INV_X1 U16178 ( .A(n14880), .ZN(n14881) );
  NAND2_X1 U16179 ( .A1(n14882), .A2(n14881), .ZN(n15021) );
  NAND2_X1 U16180 ( .A1(n14883), .A2(n15021), .ZN(n14884) );
  OAI21_X1 U16181 ( .B1(n14885), .B2(n14884), .A(n14931), .ZN(n14886) );
  NAND2_X1 U16182 ( .A1(n14886), .A2(n15012), .ZN(n14890) );
  NOR2_X1 U16183 ( .A1(n15036), .A2(n15250), .ZN(n14888) );
  OAI22_X1 U16184 ( .A1(n15243), .A2(n15038), .B1(n15037), .B2(n15242), .ZN(
        n14887) );
  AOI211_X1 U16185 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n14888), 
        .B(n14887), .ZN(n14889) );
  OAI211_X1 U16186 ( .C1(n15249), .C2(n15026), .A(n14890), .B(n14889), .ZN(
        P1_U3214) );
  OAI21_X1 U16187 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n14894) );
  NAND2_X1 U16188 ( .A1(n14894), .A2(n15012), .ZN(n14901) );
  INV_X1 U16189 ( .A(n14895), .ZN(n14898) );
  OAI22_X1 U16190 ( .A1(n14896), .A2(n15038), .B1(n15037), .B2(n15186), .ZN(
        n14897) );
  AOI211_X1 U16191 ( .C1(n14899), .C2(n15017), .A(n14898), .B(n14897), .ZN(
        n14900) );
  OAI211_X1 U16192 ( .C1(n14902), .C2(n15026), .A(n14901), .B(n14900), .ZN(
        P1_U3215) );
  INV_X1 U16193 ( .A(n14903), .ZN(n14904) );
  AOI21_X1 U16194 ( .B1(n14906), .B2(n14905), .A(n14904), .ZN(n14911) );
  INV_X1 U16195 ( .A(n15183), .ZN(n15198) );
  OAI22_X1 U16196 ( .A1(n15197), .A2(n15451), .B1(n15198), .B2(n15410), .ZN(
        n15516) );
  INV_X1 U16197 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14907) );
  OAI22_X1 U16198 ( .A1(n15309), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14907), .ZN(n14909) );
  NOR2_X1 U16199 ( .A1(n15313), .A2(n15026), .ZN(n14908) );
  AOI211_X1 U16200 ( .C1(n15029), .C2(n15516), .A(n14909), .B(n14908), .ZN(
        n14910) );
  OAI21_X1 U16201 ( .B1(n14911), .B2(n15044), .A(n14910), .ZN(P1_U3216) );
  OAI211_X1 U16202 ( .C1(n14914), .C2(n14913), .A(n14912), .B(n15012), .ZN(
        n14919) );
  AOI22_X1 U16203 ( .A1(n15017), .A2(n15090), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14918) );
  NAND2_X1 U16204 ( .A1(n15042), .A2(n10314), .ZN(n14917) );
  NAND2_X1 U16205 ( .A1(n14915), .A2(n15029), .ZN(n14916) );
  NAND4_X1 U16206 ( .A1(n14919), .A2(n14918), .A3(n14917), .A4(n14916), .ZN(
        P1_U3218) );
  INV_X1 U16207 ( .A(n14920), .ZN(n14922) );
  NAND2_X1 U16208 ( .A1(n14922), .A2(n14921), .ZN(n14923) );
  XNOR2_X1 U16209 ( .A(n14924), .B(n14923), .ZN(n14928) );
  NAND2_X1 U16210 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15160)
         );
  OAI21_X1 U16211 ( .B1(n15375), .B2(n15036), .A(n15160), .ZN(n14926) );
  OAI22_X1 U16212 ( .A1(n15182), .A2(n15037), .B1(n15411), .B2(n15038), .ZN(
        n14925) );
  AOI211_X1 U16213 ( .C1(n15538), .C2(n15042), .A(n14926), .B(n14925), .ZN(
        n14927) );
  OAI21_X1 U16214 ( .B1(n14928), .B2(n15044), .A(n14927), .ZN(P1_U3219) );
  INV_X1 U16215 ( .A(n14929), .ZN(n14930) );
  NAND2_X1 U16216 ( .A1(n14931), .A2(n14930), .ZN(n14939) );
  OAI22_X1 U16217 ( .A1(n15227), .A2(n14932), .B1(n15242), .B2(n14935), .ZN(
        n14933) );
  XNOR2_X1 U16218 ( .A(n14933), .B(n11130), .ZN(n14937) );
  OAI22_X1 U16219 ( .A1(n15227), .A2(n14935), .B1(n15242), .B2(n14934), .ZN(
        n14936) );
  XNOR2_X1 U16220 ( .A(n14937), .B(n14936), .ZN(n14938) );
  XNOR2_X1 U16221 ( .A(n14939), .B(n14938), .ZN(n14945) );
  INV_X1 U16222 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14940) );
  OAI22_X1 U16223 ( .A1(n15036), .A2(n15228), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14940), .ZN(n14943) );
  OAI22_X1 U16224 ( .A1(n15200), .A2(n15038), .B1(n15037), .B2(n14941), .ZN(
        n14942) );
  AOI211_X1 U16225 ( .C1(n15483), .C2(n15042), .A(n14943), .B(n14942), .ZN(
        n14944) );
  OAI21_X1 U16226 ( .B1(n14945), .B2(n15044), .A(n14944), .ZN(P1_U3220) );
  AOI21_X1 U16227 ( .B1(n14947), .B2(n14946), .A(n7523), .ZN(n14953) );
  NAND2_X1 U16228 ( .A1(n15333), .A2(n15006), .ZN(n14950) );
  INV_X1 U16229 ( .A(n14948), .ZN(n15337) );
  AOI22_X1 U16230 ( .A1(n15337), .A2(n15017), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14949) );
  OAI211_X1 U16231 ( .C1(n15182), .C2(n15038), .A(n14950), .B(n14949), .ZN(
        n14951) );
  AOI21_X1 U16232 ( .B1(n15528), .B2(n15042), .A(n14951), .ZN(n14952) );
  OAI21_X1 U16233 ( .B1(n14953), .B2(n15044), .A(n14952), .ZN(P1_U3223) );
  XOR2_X1 U16234 ( .A(n14955), .B(n14954), .Z(n14962) );
  NAND2_X1 U16235 ( .A1(n15183), .A2(n15386), .ZN(n14957) );
  NAND2_X1 U16236 ( .A1(n15046), .A2(n15448), .ZN(n14956) );
  NAND2_X1 U16237 ( .A1(n14957), .A2(n14956), .ZN(n15500) );
  INV_X1 U16238 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14958) );
  OAI22_X1 U16239 ( .A1(n15036), .A2(n15279), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14958), .ZN(n14960) );
  NOR2_X1 U16240 ( .A1(n8174), .A2(n15026), .ZN(n14959) );
  AOI211_X1 U16241 ( .C1(n15029), .C2(n15500), .A(n14960), .B(n14959), .ZN(
        n14961) );
  OAI21_X1 U16242 ( .B1(n14962), .B2(n15044), .A(n14961), .ZN(P1_U3225) );
  AOI21_X1 U16243 ( .B1(n14964), .B2(n14963), .A(n7442), .ZN(n14969) );
  INV_X1 U16244 ( .A(n15385), .ZN(n15191) );
  OAI22_X1 U16245 ( .A1(n15191), .A2(n15410), .B1(n15186), .B2(n15451), .ZN(
        n15561) );
  NAND2_X1 U16246 ( .A1(n15561), .A2(n15029), .ZN(n14966) );
  OAI211_X1 U16247 ( .C1(n15036), .C2(n15429), .A(n14966), .B(n14965), .ZN(
        n14967) );
  AOI21_X1 U16248 ( .B1(n15562), .B2(n15042), .A(n14967), .ZN(n14968) );
  OAI21_X1 U16249 ( .B1(n14969), .B2(n15044), .A(n14968), .ZN(P1_U3226) );
  INV_X1 U16250 ( .A(n15555), .ZN(n15416) );
  INV_X1 U16251 ( .A(n14970), .ZN(n14974) );
  NOR3_X1 U16252 ( .A1(n7442), .A2(n14972), .A3(n14971), .ZN(n14973) );
  OAI21_X1 U16253 ( .B1(n14974), .B2(n14973), .A(n15012), .ZN(n14980) );
  INV_X1 U16254 ( .A(n14975), .ZN(n15412) );
  INV_X1 U16255 ( .A(n14976), .ZN(n14978) );
  INV_X1 U16256 ( .A(n15177), .ZN(n15409) );
  OAI22_X1 U16257 ( .A1(n15411), .A2(n15037), .B1(n15409), .B2(n15038), .ZN(
        n14977) );
  AOI211_X1 U16258 ( .C1(n15017), .C2(n15412), .A(n14978), .B(n14977), .ZN(
        n14979) );
  OAI211_X1 U16259 ( .C1(n15416), .C2(n15026), .A(n14980), .B(n14979), .ZN(
        P1_U3228) );
  INV_X1 U16260 ( .A(n15509), .ZN(n15295) );
  OAI21_X1 U16261 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n14984) );
  NAND2_X1 U16262 ( .A1(n14984), .A2(n15012), .ZN(n14989) );
  INV_X1 U16263 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14985) );
  OAI22_X1 U16264 ( .A1(n15036), .A2(n15296), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14985), .ZN(n14987) );
  NOR2_X1 U16265 ( .A1(n8435), .A2(n15038), .ZN(n14986) );
  AOI211_X1 U16266 ( .C1(n15006), .C2(n15290), .A(n14987), .B(n14986), .ZN(
        n14988) );
  OAI211_X1 U16267 ( .C1(n15295), .C2(n15026), .A(n14989), .B(n14988), .ZN(
        P1_U3229) );
  OAI211_X1 U16268 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n15012), .ZN(
        n14999) );
  NAND2_X1 U16269 ( .A1(n15319), .A2(n15448), .ZN(n14994) );
  NAND2_X1 U16270 ( .A1(n15387), .A2(n15386), .ZN(n14993) );
  NAND2_X1 U16271 ( .A1(n14994), .A2(n14993), .ZN(n15348) );
  INV_X1 U16272 ( .A(n15357), .ZN(n14996) );
  OAI22_X1 U16273 ( .A1(n14996), .A2(n15036), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14995), .ZN(n14997) );
  AOI21_X1 U16274 ( .B1(n15348), .B2(n15029), .A(n14997), .ZN(n14998) );
  OAI211_X1 U16275 ( .C1(n15360), .C2(n15026), .A(n14999), .B(n14998), .ZN(
        P1_U3233) );
  OAI211_X1 U16276 ( .C1(n15002), .C2(n15001), .A(n15000), .B(n15012), .ZN(
        n15008) );
  INV_X1 U16277 ( .A(n15003), .ZN(n15326) );
  AOI22_X1 U16278 ( .A1(n15326), .A2(n15017), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15004) );
  OAI21_X1 U16279 ( .B1(n8474), .B2(n15038), .A(n15004), .ZN(n15005) );
  AOI21_X1 U16280 ( .B1(n15006), .B2(n15320), .A(n15005), .ZN(n15007) );
  OAI211_X1 U16281 ( .C1(n15026), .C2(n15329), .A(n15008), .B(n15007), .ZN(
        P1_U3235) );
  OAI21_X1 U16282 ( .B1(n15011), .B2(n15010), .A(n15009), .ZN(n15013) );
  NAND2_X1 U16283 ( .A1(n15013), .A2(n15012), .ZN(n15019) );
  INV_X1 U16284 ( .A(n15394), .ZN(n15016) );
  NAND2_X1 U16285 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15134)
         );
  INV_X1 U16286 ( .A(n15134), .ZN(n15015) );
  OAI22_X1 U16287 ( .A1(n15193), .A2(n15037), .B1(n15191), .B2(n15038), .ZN(
        n15014) );
  AOI211_X1 U16288 ( .C1(n15017), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        n15018) );
  OAI211_X1 U16289 ( .C1(n15545), .C2(n15026), .A(n15019), .B(n15018), .ZN(
        P1_U3238) );
  NAND2_X1 U16290 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  XNOR2_X1 U16291 ( .A(n15023), .B(n15022), .ZN(n15031) );
  INV_X1 U16292 ( .A(n15290), .ZN(n15024) );
  OAI22_X1 U16293 ( .A1(n15024), .A2(n15451), .B1(n15200), .B2(n15410), .ZN(
        n15494) );
  INV_X1 U16294 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15025) );
  OAI22_X1 U16295 ( .A1(n15036), .A2(n15262), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15025), .ZN(n15028) );
  INV_X1 U16296 ( .A(n15495), .ZN(n15267) );
  NOR2_X1 U16297 ( .A1(n15267), .A2(n15026), .ZN(n15027) );
  AOI211_X1 U16298 ( .C1(n15029), .C2(n15494), .A(n15028), .B(n15027), .ZN(
        n15030) );
  OAI21_X1 U16299 ( .B1(n15031), .B2(n15044), .A(n15030), .ZN(P1_U3240) );
  XNOR2_X1 U16300 ( .A(n15032), .B(n15033), .ZN(n15045) );
  OAI22_X1 U16301 ( .A1(n15036), .A2(n15035), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15034), .ZN(n15041) );
  OAI22_X1 U16302 ( .A1(n15039), .A2(n15038), .B1(n15037), .B2(n15409), .ZN(
        n15040) );
  AOI211_X1 U16303 ( .C1(n15571), .C2(n15042), .A(n15041), .B(n15040), .ZN(
        n15043) );
  OAI21_X1 U16304 ( .B1(n15045), .B2(n15044), .A(n15043), .ZN(P1_U3241) );
  MUX2_X1 U16305 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15475), .S(n15059), .Z(
        P1_U3590) );
  MUX2_X1 U16306 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15216), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16307 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15201), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16308 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15217), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16309 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15046), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16310 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15290), .S(n15059), .Z(
        P1_U3585) );
  MUX2_X1 U16311 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15183), .S(n15059), .Z(
        P1_U3584) );
  MUX2_X1 U16312 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15333), .S(n15059), .Z(
        P1_U3582) );
  MUX2_X1 U16313 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15319), .S(n15059), .Z(
        P1_U3581) );
  MUX2_X1 U16314 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15369), .S(n15059), .Z(
        P1_U3580) );
  MUX2_X1 U16315 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15387), .S(n15059), .Z(
        P1_U3579) );
  MUX2_X1 U16316 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15370), .S(n15059), .Z(
        P1_U3578) );
  MUX2_X1 U16317 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15385), .S(n15059), .Z(
        P1_U3577) );
  MUX2_X1 U16318 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15177), .S(n15059), .Z(
        P1_U3576) );
  MUX2_X1 U16319 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15175), .S(n15059), .Z(
        P1_U3575) );
  MUX2_X1 U16320 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15047), .S(n15059), .Z(
        P1_U3574) );
  MUX2_X1 U16321 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15048), .S(n15059), .Z(
        P1_U3573) );
  MUX2_X1 U16322 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15049), .S(n15059), .Z(
        P1_U3572) );
  MUX2_X1 U16323 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15050), .S(n15059), .Z(
        P1_U3571) );
  MUX2_X1 U16324 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15051), .S(n15059), .Z(
        P1_U3570) );
  MUX2_X1 U16325 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15052), .S(n15059), .Z(
        P1_U3569) );
  MUX2_X1 U16326 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15053), .S(n15059), .Z(
        P1_U3568) );
  MUX2_X1 U16327 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15054), .S(n15059), .Z(
        P1_U3567) );
  MUX2_X1 U16328 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15055), .S(n15059), .Z(
        P1_U3566) );
  MUX2_X1 U16329 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15056), .S(n15059), .Z(
        P1_U3565) );
  MUX2_X1 U16330 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15057), .S(n15059), .Z(
        P1_U3564) );
  MUX2_X1 U16331 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15058), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16332 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15449), .S(n15059), .Z(
        P1_U3562) );
  MUX2_X1 U16333 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15060), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16334 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15061), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16335 ( .C1(n15075), .C2(n15063), .A(n15154), .B(n15062), .ZN(
        n15072) );
  OAI211_X1 U16336 ( .C1(n15066), .C2(n15065), .A(n15155), .B(n15064), .ZN(
        n15071) );
  AOI22_X1 U16337 ( .A1(n16197), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n15070) );
  INV_X1 U16338 ( .A(n15067), .ZN(n15068) );
  NAND2_X1 U16339 ( .A1(n15118), .A2(n15068), .ZN(n15069) );
  NAND4_X1 U16340 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        P1_U3244) );
  INV_X1 U16341 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15074) );
  AOI21_X1 U16342 ( .B1(n16194), .B2(n15074), .A(n15073), .ZN(n16193) );
  MUX2_X1 U16343 ( .A(n15076), .B(n15075), .S(n16194), .Z(n15078) );
  NAND2_X1 U16344 ( .A1(n15078), .A2(n15077), .ZN(n15079) );
  OAI211_X1 U16345 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n16193), .A(n15079), .B(
        P1_U4016), .ZN(n15125) );
  AOI22_X1 U16346 ( .A1(n16197), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n15089) );
  OAI211_X1 U16347 ( .C1(n15081), .C2(n15080), .A(n15154), .B(n15096), .ZN(
        n15085) );
  OAI211_X1 U16348 ( .C1(n15083), .C2(n15082), .A(n15155), .B(n15101), .ZN(
        n15084) );
  OAI211_X1 U16349 ( .C1(n15149), .C2(n15086), .A(n15085), .B(n15084), .ZN(
        n15087) );
  INV_X1 U16350 ( .A(n15087), .ZN(n15088) );
  NAND3_X1 U16351 ( .A1(n15125), .A2(n15089), .A3(n15088), .ZN(P1_U3245) );
  INV_X1 U16352 ( .A(n15098), .ZN(n15093) );
  OAI22_X1 U16353 ( .A1(n15162), .A2(n15091), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15090), .ZN(n15092) );
  AOI21_X1 U16354 ( .B1(n15093), .B2(n15118), .A(n15092), .ZN(n15105) );
  MUX2_X1 U16355 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10901), .S(n15098), .Z(
        n15094) );
  NAND3_X1 U16356 ( .A1(n15096), .A2(n15095), .A3(n15094), .ZN(n15097) );
  NAND3_X1 U16357 ( .A1(n15154), .A2(n15108), .A3(n15097), .ZN(n15104) );
  MUX2_X1 U16358 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10895), .S(n15098), .Z(
        n15099) );
  NAND3_X1 U16359 ( .A1(n15101), .A2(n15100), .A3(n15099), .ZN(n15102) );
  NAND3_X1 U16360 ( .A1(n15155), .A2(n15114), .A3(n15102), .ZN(n15103) );
  NAND3_X1 U16361 ( .A1(n15105), .A2(n15104), .A3(n15103), .ZN(P1_U3246) );
  NAND2_X1 U16362 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n16197), .ZN(n15124) );
  MUX2_X1 U16363 ( .A(n11529), .B(P1_REG2_REG_4__SCAN_IN), .S(n15117), .Z(
        n15106) );
  NAND3_X1 U16364 ( .A1(n15108), .A2(n15107), .A3(n15106), .ZN(n15109) );
  NAND3_X1 U16365 ( .A1(n15154), .A2(n15110), .A3(n15109), .ZN(n15122) );
  INV_X1 U16366 ( .A(n15111), .ZN(n15116) );
  NAND3_X1 U16367 ( .A1(n15114), .A2(n15113), .A3(n15112), .ZN(n15115) );
  NAND3_X1 U16368 ( .A1(n15155), .A2(n15116), .A3(n15115), .ZN(n15121) );
  NAND2_X1 U16369 ( .A1(n15118), .A2(n15117), .ZN(n15120) );
  AND4_X1 U16370 ( .A1(n15122), .A2(n15121), .A3(n15120), .A4(n15119), .ZN(
        n15123) );
  NAND3_X1 U16371 ( .A1(n15125), .A2(n15124), .A3(n15123), .ZN(P1_U3247) );
  INV_X1 U16372 ( .A(n15145), .ZN(n15138) );
  OAI21_X1 U16373 ( .B1(n15127), .B2(n15130), .A(n15126), .ZN(n15144) );
  XOR2_X1 U16374 ( .A(n15144), .B(n15145), .Z(n15128) );
  NAND2_X1 U16375 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15128), .ZN(n15147) );
  OAI211_X1 U16376 ( .C1(n15128), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15154), 
        .B(n15147), .ZN(n15137) );
  XNOR2_X1 U16377 ( .A(n15139), .B(n15138), .ZN(n15132) );
  NAND2_X1 U16378 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n15132), .ZN(n15141) );
  OAI211_X1 U16379 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n15132), .A(n15155), 
        .B(n15141), .ZN(n15133) );
  NAND2_X1 U16380 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  AOI21_X1 U16381 ( .B1(n16197), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15135), 
        .ZN(n15136) );
  OAI211_X1 U16382 ( .C1(n15149), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        P1_U3261) );
  NAND2_X1 U16383 ( .A1(n15145), .A2(n15139), .ZN(n15140) );
  NAND2_X1 U16384 ( .A1(n15141), .A2(n15140), .ZN(n15143) );
  XNOR2_X1 U16385 ( .A(n15143), .B(n15142), .ZN(n15156) );
  INV_X1 U16386 ( .A(n15156), .ZN(n15152) );
  NAND2_X1 U16387 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  NAND2_X1 U16388 ( .A1(n15147), .A2(n15146), .ZN(n15148) );
  XOR2_X1 U16389 ( .A(n15148), .B(P1_REG2_REG_19__SCAN_IN), .Z(n15153) );
  OAI21_X1 U16390 ( .B1(n15153), .B2(n15150), .A(n15149), .ZN(n15151) );
  AOI21_X1 U16391 ( .B1(n15152), .B2(n15155), .A(n15151), .ZN(n15159) );
  AOI22_X1 U16392 ( .A1(n15156), .A2(n15155), .B1(n15154), .B2(n15153), .ZN(
        n15158) );
  OAI211_X1 U16393 ( .C1(n8565), .C2(n15162), .A(n15161), .B(n15160), .ZN(
        P1_U3262) );
  NAND2_X1 U16394 ( .A1(n15416), .A2(n15426), .ZN(n15406) );
  NAND2_X1 U16395 ( .A1(n15313), .A2(n15325), .ZN(n15306) );
  OR2_X2 U16396 ( .A1(n15246), .A2(n15483), .ZN(n15204) );
  NAND2_X1 U16397 ( .A1(n15226), .A2(n15211), .ZN(n15170) );
  XNOR2_X1 U16398 ( .A(n15169), .B(n15165), .ZN(n15163) );
  NAND2_X1 U16399 ( .A1(n15163), .A2(n16326), .ZN(n15468) );
  AOI21_X1 U16400 ( .B1(n16194), .B2(P1_B_REG_SCAN_IN), .A(n15410), .ZN(n15476) );
  NAND2_X1 U16401 ( .A1(n15164), .A2(n15476), .ZN(n15471) );
  NOR2_X1 U16402 ( .A1(n15356), .A2(n15471), .ZN(n15172) );
  INV_X1 U16403 ( .A(n15165), .ZN(n15469) );
  NOR2_X1 U16404 ( .A1(n15469), .A2(n15434), .ZN(n15166) );
  AOI211_X1 U16405 ( .C1(n15356), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15172), 
        .B(n15166), .ZN(n15167) );
  OAI21_X1 U16406 ( .B1(n15468), .B2(n15168), .A(n15167), .ZN(P1_U3263) );
  INV_X1 U16407 ( .A(n15171), .ZN(n15473) );
  AOI21_X1 U16408 ( .B1(n15171), .B2(n15170), .A(n15169), .ZN(n15470) );
  NAND2_X1 U16409 ( .A1(n15470), .A2(n15463), .ZN(n15174) );
  AOI21_X1 U16410 ( .B1(n15356), .B2(P1_REG2_REG_30__SCAN_IN), .A(n15172), 
        .ZN(n15173) );
  OAI211_X1 U16411 ( .C1(n15473), .C2(n15434), .A(n15174), .B(n15173), .ZN(
        P1_U3264) );
  OR2_X1 U16412 ( .A1(n15562), .A2(n15177), .ZN(n15178) );
  INV_X1 U16413 ( .A(n15405), .ZN(n15179) );
  NAND2_X1 U16414 ( .A1(n15555), .A2(n15385), .ZN(n15180) );
  NAND2_X1 U16415 ( .A1(n15552), .A2(n15180), .ZN(n15381) );
  NAND2_X1 U16416 ( .A1(n15545), .A2(n15411), .ZN(n15181) );
  INV_X1 U16417 ( .A(n15317), .ZN(n15323) );
  INV_X1 U16418 ( .A(n15288), .ZN(n15285) );
  NAND2_X1 U16419 ( .A1(n15562), .A2(n15409), .ZN(n15189) );
  NAND2_X1 U16420 ( .A1(n15555), .A2(n15191), .ZN(n15192) );
  INV_X1 U16421 ( .A(n15365), .ZN(n15194) );
  INV_X1 U16422 ( .A(n15352), .ZN(n15195) );
  NAND2_X1 U16423 ( .A1(n15346), .A2(n15195), .ZN(n15349) );
  NAND2_X1 U16424 ( .A1(n15349), .A2(n15196), .ZN(n15332) );
  AOI22_X2 U16425 ( .A1(n15332), .A2(n15340), .B1(n8181), .B2(n15319), .ZN(
        n15318) );
  INV_X1 U16426 ( .A(n15274), .ZN(n15199) );
  NOR2_X1 U16427 ( .A1(n15479), .A2(n15398), .ZN(n15213) );
  NOR2_X1 U16428 ( .A1(n15242), .A2(n15451), .ZN(n15474) );
  AND3_X1 U16429 ( .A1(n15205), .A2(n15476), .A3(n15475), .ZN(n15209) );
  OAI22_X1 U16430 ( .A1(n15430), .A2(n15207), .B1(n15206), .B2(n15428), .ZN(
        n15208) );
  AOI211_X1 U16431 ( .C1(n15474), .C2(n15430), .A(n15209), .B(n15208), .ZN(
        n15210) );
  OAI21_X1 U16432 ( .B1(n15211), .B2(n15434), .A(n15210), .ZN(n15212) );
  AOI211_X1 U16433 ( .C1(n15481), .C2(n15269), .A(n15213), .B(n15212), .ZN(
        n15214) );
  OAI21_X1 U16434 ( .B1(n15482), .B2(n15342), .A(n15214), .ZN(P1_U3356) );
  NAND2_X1 U16435 ( .A1(n15216), .A2(n15448), .ZN(n15219) );
  NAND2_X1 U16436 ( .A1(n15217), .A2(n15386), .ZN(n15218) );
  OAI21_X1 U16437 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15487) );
  INV_X1 U16438 ( .A(n15487), .ZN(n15225) );
  NAND2_X1 U16439 ( .A1(n15225), .A2(n15224), .ZN(n15233) );
  AOI21_X1 U16440 ( .B1(n15483), .B2(n15246), .A(n15226), .ZN(n15484) );
  NOR2_X1 U16441 ( .A1(n15227), .A2(n15434), .ZN(n15231) );
  OAI22_X1 U16442 ( .A1(n15430), .A2(n15229), .B1(n15228), .B2(n15428), .ZN(
        n15230) );
  AOI211_X1 U16443 ( .C1(n15484), .C2(n15463), .A(n15231), .B(n15230), .ZN(
        n15232) );
  OAI211_X1 U16444 ( .C1(n15486), .C2(n15356), .A(n15233), .B(n15232), .ZN(
        P1_U3265) );
  AOI21_X1 U16445 ( .B1(n15236), .B2(n15235), .A(n15234), .ZN(n15492) );
  INV_X1 U16446 ( .A(n15492), .ZN(n15254) );
  INV_X1 U16447 ( .A(n15237), .ZN(n15241) );
  AOI21_X1 U16448 ( .B1(n15241), .B2(n15240), .A(n15567), .ZN(n15245) );
  OAI22_X1 U16449 ( .A1(n15243), .A2(n15451), .B1(n15242), .B2(n15410), .ZN(
        n15244) );
  INV_X1 U16450 ( .A(n15261), .ZN(n15248) );
  INV_X1 U16451 ( .A(n15246), .ZN(n15247) );
  AOI211_X1 U16452 ( .C1(n15489), .C2(n15248), .A(n16428), .B(n15247), .ZN(
        n15488) );
  NOR2_X1 U16453 ( .A1(n15249), .A2(n15434), .ZN(n15253) );
  OAI22_X1 U16454 ( .A1(n15430), .A2(n15251), .B1(n15250), .B2(n15428), .ZN(
        n15252) );
  AOI211_X1 U16455 ( .C1(n15488), .C2(n15437), .A(n15253), .B(n15252), .ZN(
        n15256) );
  NAND2_X1 U16456 ( .A1(n15254), .A2(n15460), .ZN(n15255) );
  OAI211_X1 U16457 ( .C1(n15491), .C2(n15356), .A(n15256), .B(n15255), .ZN(
        P1_U3266) );
  XNOR2_X1 U16458 ( .A(n15257), .B(n15259), .ZN(n15499) );
  OAI21_X1 U16459 ( .B1(n15260), .B2(n15259), .A(n15258), .ZN(n15496) );
  AOI211_X1 U16460 ( .C1(n15495), .C2(n15276), .A(n16428), .B(n15261), .ZN(
        n15493) );
  NAND2_X1 U16461 ( .A1(n15493), .A2(n15437), .ZN(n15266) );
  OAI22_X1 U16462 ( .A1(n15430), .A2(n15263), .B1(n15262), .B2(n15428), .ZN(
        n15264) );
  AOI21_X1 U16463 ( .B1(n15494), .B2(n15432), .A(n15264), .ZN(n15265) );
  OAI211_X1 U16464 ( .C1(n15267), .C2(n15434), .A(n15266), .B(n15265), .ZN(
        n15268) );
  AOI21_X1 U16465 ( .B1(n15496), .B2(n15269), .A(n15268), .ZN(n15270) );
  OAI21_X1 U16466 ( .B1(n15499), .B2(n15342), .A(n15270), .ZN(P1_U3267) );
  XNOR2_X1 U16467 ( .A(n15271), .B(n15274), .ZN(n15507) );
  AOI21_X1 U16468 ( .B1(n15274), .B2(n15273), .A(n15272), .ZN(n15505) );
  NAND2_X1 U16469 ( .A1(n15294), .A2(n15501), .ZN(n15275) );
  NAND2_X1 U16470 ( .A1(n15276), .A2(n15275), .ZN(n15503) );
  NAND2_X1 U16471 ( .A1(n15356), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U16472 ( .A1(n15500), .A2(n15432), .ZN(n15277) );
  OAI211_X1 U16473 ( .C1(n15428), .C2(n15279), .A(n15278), .B(n15277), .ZN(
        n15280) );
  AOI21_X1 U16474 ( .B1(n15501), .B2(n15459), .A(n15280), .ZN(n15281) );
  OAI21_X1 U16475 ( .B1(n15503), .B2(n15398), .A(n15281), .ZN(n15282) );
  AOI21_X1 U16476 ( .B1(n15505), .B2(n15425), .A(n15282), .ZN(n15283) );
  OAI21_X1 U16477 ( .B1(n15440), .B2(n15507), .A(n15283), .ZN(P1_U3268) );
  OAI21_X1 U16478 ( .B1(n15286), .B2(n15285), .A(n15284), .ZN(n15508) );
  OAI211_X1 U16479 ( .C1(n15289), .C2(n15288), .A(n15287), .B(n15584), .ZN(
        n15292) );
  AOI22_X1 U16480 ( .A1(n15320), .A2(n15386), .B1(n15448), .B2(n15290), .ZN(
        n15291) );
  NAND2_X1 U16481 ( .A1(n15292), .A2(n15291), .ZN(n15293) );
  AOI21_X1 U16482 ( .B1(n15508), .B2(n15445), .A(n15293), .ZN(n15512) );
  AOI21_X1 U16483 ( .B1(n15509), .B2(n15306), .A(n8175), .ZN(n15510) );
  NOR2_X1 U16484 ( .A1(n15295), .A2(n15434), .ZN(n15299) );
  OAI22_X1 U16485 ( .A1(n15430), .A2(n15297), .B1(n15296), .B2(n15428), .ZN(
        n15298) );
  AOI211_X1 U16486 ( .C1(n15510), .C2(n15463), .A(n15299), .B(n15298), .ZN(
        n15301) );
  NAND2_X1 U16487 ( .A1(n15508), .A2(n15460), .ZN(n15300) );
  OAI211_X1 U16488 ( .C1(n15512), .C2(n15356), .A(n15301), .B(n15300), .ZN(
        P1_U3269) );
  AOI21_X1 U16489 ( .B1(n15303), .B2(n15302), .A(n7486), .ZN(n15520) );
  AOI21_X1 U16490 ( .B1(n8428), .B2(n15305), .A(n15304), .ZN(n15514) );
  NAND2_X1 U16491 ( .A1(n15514), .A2(n15425), .ZN(n15316) );
  INV_X1 U16492 ( .A(n15325), .ZN(n15308) );
  INV_X1 U16493 ( .A(n15306), .ZN(n15307) );
  AOI211_X1 U16494 ( .C1(n15517), .C2(n15308), .A(n16428), .B(n15307), .ZN(
        n15515) );
  INV_X1 U16495 ( .A(n15309), .ZN(n15310) );
  AOI22_X1 U16496 ( .A1(n15310), .A2(n15458), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15356), .ZN(n15312) );
  NAND2_X1 U16497 ( .A1(n15516), .A2(n15432), .ZN(n15311) );
  OAI211_X1 U16498 ( .C1(n15313), .C2(n15434), .A(n15312), .B(n15311), .ZN(
        n15314) );
  AOI21_X1 U16499 ( .B1(n15515), .B2(n15437), .A(n15314), .ZN(n15315) );
  OAI211_X1 U16500 ( .C1(n15520), .C2(n15440), .A(n15316), .B(n15315), .ZN(
        P1_U3270) );
  XNOR2_X1 U16501 ( .A(n15318), .B(n15317), .ZN(n15321) );
  AOI222_X1 U16502 ( .A1(n15584), .A2(n15321), .B1(n15320), .B2(n15448), .C1(
        n15319), .C2(n15386), .ZN(n15525) );
  OAI21_X1 U16503 ( .B1(n15324), .B2(n15323), .A(n15322), .ZN(n15521) );
  AOI21_X1 U16504 ( .B1(n15522), .B2(n15336), .A(n15325), .ZN(n15523) );
  NAND2_X1 U16505 ( .A1(n15523), .A2(n15463), .ZN(n15328) );
  AOI22_X1 U16506 ( .A1(n15326), .A2(n15458), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15356), .ZN(n15327) );
  OAI211_X1 U16507 ( .C1(n15434), .C2(n15329), .A(n15328), .B(n15327), .ZN(
        n15330) );
  AOI21_X1 U16508 ( .B1(n15521), .B2(n15425), .A(n15330), .ZN(n15331) );
  OAI21_X1 U16509 ( .B1(n15525), .B2(n15356), .A(n15331), .ZN(P1_U3271) );
  XOR2_X1 U16510 ( .A(n15340), .B(n15332), .Z(n15334) );
  AOI222_X1 U16511 ( .A1(n15584), .A2(n15334), .B1(n15333), .B2(n15448), .C1(
        n15369), .C2(n15386), .ZN(n15530) );
  AOI21_X1 U16512 ( .B1(n15528), .B2(n15354), .A(n16428), .ZN(n15335) );
  AND2_X1 U16513 ( .A1(n15336), .A2(n15335), .ZN(n15527) );
  NAND2_X1 U16514 ( .A1(n15528), .A2(n15459), .ZN(n15339) );
  AOI22_X1 U16515 ( .A1(n15337), .A2(n15458), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15356), .ZN(n15338) );
  NAND2_X1 U16516 ( .A1(n15339), .A2(n15338), .ZN(n15344) );
  XOR2_X1 U16517 ( .A(n15341), .B(n15340), .Z(n15531) );
  NOR2_X1 U16518 ( .A1(n15531), .A2(n15342), .ZN(n15343) );
  AOI211_X1 U16519 ( .C1(n15527), .C2(n15437), .A(n15344), .B(n15343), .ZN(
        n15345) );
  OAI21_X1 U16520 ( .B1(n15356), .B2(n15530), .A(n15345), .ZN(P1_U3272) );
  INV_X1 U16521 ( .A(n15346), .ZN(n15347) );
  AOI21_X1 U16522 ( .B1(n15347), .B2(n15352), .A(n15567), .ZN(n15350) );
  AOI21_X1 U16523 ( .B1(n15350), .B2(n15349), .A(n15348), .ZN(n15535) );
  OAI21_X1 U16524 ( .B1(n15353), .B2(n15352), .A(n15351), .ZN(n15536) );
  INV_X1 U16525 ( .A(n15536), .ZN(n15362) );
  AOI21_X1 U16526 ( .B1(n15533), .B2(n15368), .A(n16428), .ZN(n15355) );
  AND2_X1 U16527 ( .A1(n15355), .A2(n15354), .ZN(n15532) );
  NAND2_X1 U16528 ( .A1(n15532), .A2(n15437), .ZN(n15359) );
  AOI22_X1 U16529 ( .A1(n15357), .A2(n15458), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n15356), .ZN(n15358) );
  OAI211_X1 U16530 ( .C1(n15360), .C2(n15434), .A(n15359), .B(n15358), .ZN(
        n15361) );
  AOI21_X1 U16531 ( .B1(n15362), .B2(n15425), .A(n15361), .ZN(n15363) );
  OAI21_X1 U16532 ( .B1(n15356), .B2(n15535), .A(n15363), .ZN(P1_U3273) );
  XNOR2_X1 U16533 ( .A(n15364), .B(n15365), .ZN(n15544) );
  XNOR2_X1 U16534 ( .A(n15366), .B(n15365), .ZN(n15542) );
  NAND2_X1 U16535 ( .A1(n15538), .A2(n15392), .ZN(n15367) );
  NAND2_X1 U16536 ( .A1(n15368), .A2(n15367), .ZN(n15540) );
  NAND2_X1 U16537 ( .A1(n15369), .A2(n15448), .ZN(n15372) );
  NAND2_X1 U16538 ( .A1(n15370), .A2(n15386), .ZN(n15371) );
  NAND2_X1 U16539 ( .A1(n15372), .A2(n15371), .ZN(n15537) );
  NAND2_X1 U16540 ( .A1(n15537), .A2(n15432), .ZN(n15374) );
  NAND2_X1 U16541 ( .A1(n15356), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n15373) );
  OAI211_X1 U16542 ( .C1(n15428), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        n15376) );
  AOI21_X1 U16543 ( .B1(n15538), .B2(n15459), .A(n15376), .ZN(n15377) );
  OAI21_X1 U16544 ( .B1(n15540), .B2(n15398), .A(n15377), .ZN(n15378) );
  AOI21_X1 U16545 ( .B1(n15542), .B2(n15425), .A(n15378), .ZN(n15379) );
  OAI21_X1 U16546 ( .B1(n15440), .B2(n15544), .A(n15379), .ZN(P1_U3274) );
  INV_X1 U16547 ( .A(n15382), .ZN(n15380) );
  XNOR2_X1 U16548 ( .A(n15381), .B(n15380), .ZN(n15548) );
  NAND2_X1 U16549 ( .A1(n15383), .A2(n15382), .ZN(n15384) );
  NAND2_X1 U16550 ( .A1(n15384), .A2(n15584), .ZN(n15389) );
  AOI22_X1 U16551 ( .A1(n15387), .A2(n15448), .B1(n15386), .B2(n15385), .ZN(
        n15388) );
  OAI21_X1 U16552 ( .B1(n7534), .B2(n15389), .A(n15388), .ZN(n15390) );
  AOI21_X1 U16553 ( .B1(n15548), .B2(n15445), .A(n15390), .ZN(n15550) );
  NAND2_X1 U16554 ( .A1(n15396), .A2(n15406), .ZN(n15391) );
  NAND2_X1 U16555 ( .A1(n15392), .A2(n15391), .ZN(n15546) );
  OAI22_X1 U16556 ( .A1(n15394), .A2(n15428), .B1(n15393), .B2(n15432), .ZN(
        n15395) );
  AOI21_X1 U16557 ( .B1(n15396), .B2(n15459), .A(n15395), .ZN(n15397) );
  OAI21_X1 U16558 ( .B1(n15546), .B2(n15398), .A(n15397), .ZN(n15399) );
  AOI21_X1 U16559 ( .B1(n15548), .B2(n15460), .A(n15399), .ZN(n15400) );
  OAI21_X1 U16560 ( .B1(n15550), .B2(n15356), .A(n15400), .ZN(P1_U3275) );
  OAI21_X1 U16561 ( .B1(n15402), .B2(n15405), .A(n15401), .ZN(n15403) );
  INV_X1 U16562 ( .A(n15403), .ZN(n15558) );
  NAND2_X1 U16563 ( .A1(n15404), .A2(n15405), .ZN(n15551) );
  NAND3_X1 U16564 ( .A1(n15552), .A2(n15551), .A3(n15425), .ZN(n15420) );
  INV_X1 U16565 ( .A(n15426), .ZN(n15408) );
  INV_X1 U16566 ( .A(n15406), .ZN(n15407) );
  AOI211_X1 U16567 ( .C1(n15555), .C2(n15408), .A(n16428), .B(n15407), .ZN(
        n15553) );
  INV_X1 U16568 ( .A(n15553), .ZN(n15415) );
  OAI22_X1 U16569 ( .A1(n15411), .A2(n15410), .B1(n15409), .B2(n15451), .ZN(
        n15554) );
  AOI21_X1 U16570 ( .B1(n15412), .B2(n15458), .A(n15554), .ZN(n15413) );
  OAI21_X1 U16571 ( .B1(n15415), .B2(n15414), .A(n15413), .ZN(n15418) );
  OAI22_X1 U16572 ( .A1(n15416), .A2(n15434), .B1(n15430), .B2(n15127), .ZN(
        n15417) );
  AOI21_X1 U16573 ( .B1(n15418), .B2(n15432), .A(n15417), .ZN(n15419) );
  OAI211_X1 U16574 ( .C1(n15558), .C2(n15440), .A(n15420), .B(n15419), .ZN(
        P1_U3276) );
  XNOR2_X1 U16575 ( .A(n15422), .B(n15421), .ZN(n15566) );
  XNOR2_X1 U16576 ( .A(n15423), .B(n15424), .ZN(n15559) );
  NAND2_X1 U16577 ( .A1(n15559), .A2(n15425), .ZN(n15439) );
  AOI211_X1 U16578 ( .C1(n15562), .C2(n15427), .A(n16428), .B(n15426), .ZN(
        n15560) );
  INV_X1 U16579 ( .A(n15562), .ZN(n15435) );
  OAI22_X1 U16580 ( .A1(n15430), .A2(n12801), .B1(n15429), .B2(n15428), .ZN(
        n15431) );
  AOI21_X1 U16581 ( .B1(n15561), .B2(n15432), .A(n15431), .ZN(n15433) );
  OAI21_X1 U16582 ( .B1(n15435), .B2(n15434), .A(n15433), .ZN(n15436) );
  AOI21_X1 U16583 ( .B1(n15560), .B2(n15437), .A(n15436), .ZN(n15438) );
  OAI211_X1 U16584 ( .C1(n15566), .C2(n15440), .A(n15439), .B(n15438), .ZN(
        P1_U3277) );
  INV_X1 U16585 ( .A(n15441), .ZN(n15442) );
  NAND2_X1 U16586 ( .A1(n11294), .A2(n15442), .ZN(n15443) );
  NAND2_X1 U16587 ( .A1(n15444), .A2(n15443), .ZN(n16334) );
  NAND2_X1 U16588 ( .A1(n16334), .A2(n15445), .ZN(n15456) );
  OAI21_X1 U16589 ( .B1(n15447), .B2(n11294), .A(n15446), .ZN(n15454) );
  NAND2_X1 U16590 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  OAI21_X1 U16591 ( .B1(n15452), .B2(n15451), .A(n15450), .ZN(n15453) );
  AOI21_X1 U16592 ( .B1(n15454), .B2(n15584), .A(n15453), .ZN(n15455) );
  AND2_X1 U16593 ( .A1(n15456), .A2(n15455), .ZN(n16331) );
  MUX2_X1 U16594 ( .A(n16331), .B(n15457), .S(n15356), .Z(n15467) );
  AOI22_X1 U16595 ( .A1(n15459), .A2(n7438), .B1(n15458), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n15466) );
  NAND2_X1 U16596 ( .A1(n16334), .A2(n15460), .ZN(n15465) );
  NAND2_X1 U16597 ( .A1(n15462), .A2(n7438), .ZN(n16327) );
  NAND3_X1 U16598 ( .A1(n15463), .A2(n16328), .A3(n16327), .ZN(n15464) );
  NAND4_X1 U16599 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        P1_U3292) );
  OAI211_X1 U16600 ( .C1(n15469), .C2(n16437), .A(n15468), .B(n15471), .ZN(
        n15590) );
  MUX2_X1 U16601 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15590), .S(n16446), .Z(
        P1_U3559) );
  NAND2_X1 U16602 ( .A1(n15470), .A2(n16326), .ZN(n15472) );
  OAI211_X1 U16603 ( .C1(n15473), .C2(n16437), .A(n15472), .B(n15471), .ZN(
        n15591) );
  MUX2_X1 U16604 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15591), .S(n16446), .Z(
        P1_U3558) );
  AOI21_X1 U16605 ( .B1(n15476), .B2(n15475), .A(n15474), .ZN(n15478) );
  MUX2_X1 U16606 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15592), .S(n16446), .Z(
        P1_U3557) );
  AOI22_X1 U16607 ( .A1(n15484), .A2(n16326), .B1(n16358), .B2(n15483), .ZN(
        n15485) );
  OAI211_X1 U16608 ( .C1(n15487), .C2(n16425), .A(n15486), .B(n15485), .ZN(
        n15593) );
  MUX2_X1 U16609 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15593), .S(n16446), .Z(
        P1_U3556) );
  AOI21_X1 U16610 ( .B1(n15563), .B2(n15489), .A(n15488), .ZN(n15490) );
  MUX2_X1 U16611 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15594), .S(n16446), .Z(
        P1_U3555) );
  AOI211_X1 U16612 ( .C1(n15563), .C2(n15495), .A(n15494), .B(n15493), .ZN(
        n15498) );
  NAND2_X1 U16613 ( .A1(n15496), .A2(n15584), .ZN(n15497) );
  OAI211_X1 U16614 ( .C1(n15499), .C2(n16425), .A(n15498), .B(n15497), .ZN(
        n15595) );
  MUX2_X1 U16615 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15595), .S(n16446), .Z(
        P1_U3554) );
  AOI21_X1 U16616 ( .B1(n15501), .B2(n16358), .A(n15500), .ZN(n15502) );
  OAI21_X1 U16617 ( .B1(n15503), .B2(n16428), .A(n15502), .ZN(n15504) );
  AOI21_X1 U16618 ( .B1(n15505), .B2(n15568), .A(n15504), .ZN(n15506) );
  OAI21_X1 U16619 ( .B1(n15567), .B2(n15507), .A(n15506), .ZN(n15596) );
  MUX2_X1 U16620 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15596), .S(n16446), .Z(
        P1_U3553) );
  INV_X1 U16621 ( .A(n15508), .ZN(n15513) );
  AOI22_X1 U16622 ( .A1(n15510), .A2(n16326), .B1(n15563), .B2(n15509), .ZN(
        n15511) );
  OAI211_X1 U16623 ( .C1(n15513), .C2(n16353), .A(n15512), .B(n15511), .ZN(
        n15597) );
  MUX2_X1 U16624 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15597), .S(n16446), .Z(
        P1_U3552) );
  NAND2_X1 U16625 ( .A1(n15514), .A2(n15568), .ZN(n15519) );
  AOI211_X1 U16626 ( .C1(n15563), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15518) );
  OAI211_X1 U16627 ( .C1(n15567), .C2(n15520), .A(n15519), .B(n15518), .ZN(
        n15598) );
  MUX2_X1 U16628 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15598), .S(n16446), .Z(
        P1_U3551) );
  INV_X1 U16629 ( .A(n15521), .ZN(n15526) );
  AOI22_X1 U16630 ( .A1(n15523), .A2(n16326), .B1(n15522), .B2(n16358), .ZN(
        n15524) );
  OAI211_X1 U16631 ( .C1(n16425), .C2(n15526), .A(n15525), .B(n15524), .ZN(
        n15599) );
  MUX2_X1 U16632 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15599), .S(n16446), .Z(
        P1_U3550) );
  AOI21_X1 U16633 ( .B1(n15563), .B2(n15528), .A(n15527), .ZN(n15529) );
  OAI211_X1 U16634 ( .C1(n16425), .C2(n15531), .A(n15530), .B(n15529), .ZN(
        n15600) );
  MUX2_X1 U16635 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15600), .S(n16446), .Z(
        P1_U3549) );
  AOI21_X1 U16636 ( .B1(n15563), .B2(n15533), .A(n15532), .ZN(n15534) );
  OAI211_X1 U16637 ( .C1(n15536), .C2(n16425), .A(n15535), .B(n15534), .ZN(
        n15601) );
  MUX2_X1 U16638 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15601), .S(n16446), .Z(
        P1_U3548) );
  AOI21_X1 U16639 ( .B1(n15538), .B2(n16358), .A(n15537), .ZN(n15539) );
  OAI21_X1 U16640 ( .B1(n15540), .B2(n16428), .A(n15539), .ZN(n15541) );
  AOI21_X1 U16641 ( .B1(n15542), .B2(n15568), .A(n15541), .ZN(n15543) );
  OAI21_X1 U16642 ( .B1(n15567), .B2(n15544), .A(n15543), .ZN(n15602) );
  MUX2_X1 U16643 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15602), .S(n16446), .Z(
        P1_U3547) );
  INV_X1 U16644 ( .A(n16353), .ZN(n16440) );
  OAI22_X1 U16645 ( .A1(n15546), .A2(n16428), .B1(n15545), .B2(n16437), .ZN(
        n15547) );
  AOI21_X1 U16646 ( .B1(n15548), .B2(n16440), .A(n15547), .ZN(n15549) );
  NAND2_X1 U16647 ( .A1(n15550), .A2(n15549), .ZN(n15603) );
  MUX2_X1 U16648 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15603), .S(n16446), .Z(
        P1_U3546) );
  NAND3_X1 U16649 ( .A1(n15552), .A2(n15568), .A3(n15551), .ZN(n15557) );
  AOI211_X1 U16650 ( .C1(n15563), .C2(n15555), .A(n15554), .B(n15553), .ZN(
        n15556) );
  OAI211_X1 U16651 ( .C1(n15567), .C2(n15558), .A(n15557), .B(n15556), .ZN(
        n15604) );
  MUX2_X1 U16652 ( .A(n15604), .B(P1_REG1_REG_17__SCAN_IN), .S(n16444), .Z(
        P1_U3545) );
  NAND2_X1 U16653 ( .A1(n15559), .A2(n15568), .ZN(n15565) );
  AOI211_X1 U16654 ( .C1(n15563), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15564) );
  OAI211_X1 U16655 ( .C1(n15567), .C2(n15566), .A(n15565), .B(n15564), .ZN(
        n15605) );
  MUX2_X1 U16656 ( .A(n15605), .B(P1_REG1_REG_16__SCAN_IN), .S(n16444), .Z(
        P1_U3544) );
  NAND2_X1 U16657 ( .A1(n15569), .A2(n15568), .ZN(n15577) );
  AOI21_X1 U16658 ( .B1(n15571), .B2(n16358), .A(n15570), .ZN(n15572) );
  NAND2_X1 U16659 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  AOI21_X1 U16660 ( .B1(n15575), .B2(n15584), .A(n15574), .ZN(n15576) );
  NAND2_X1 U16661 ( .A1(n15577), .A2(n15576), .ZN(n15606) );
  MUX2_X1 U16662 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15606), .S(n16446), .Z(
        P1_U3543) );
  OR2_X1 U16663 ( .A1(n15578), .A2(n16425), .ZN(n15587) );
  NAND2_X1 U16664 ( .A1(n15579), .A2(n16358), .ZN(n15580) );
  OAI211_X1 U16665 ( .C1(n15582), .C2(n16428), .A(n15581), .B(n15580), .ZN(
        n15583) );
  AOI21_X1 U16666 ( .B1(n15585), .B2(n15584), .A(n15583), .ZN(n15586) );
  NAND2_X1 U16667 ( .A1(n15587), .A2(n15586), .ZN(n15607) );
  MUX2_X1 U16668 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15607), .S(n16446), .Z(
        P1_U3542) );
  MUX2_X1 U16669 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15588), .S(n16446), .Z(
        P1_U3534) );
  MUX2_X1 U16670 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15589), .S(n16446), .Z(
        P1_U3533) );
  MUX2_X1 U16671 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15590), .S(n16338), .Z(
        P1_U3527) );
  MUX2_X1 U16672 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15591), .S(n16338), .Z(
        P1_U3526) );
  MUX2_X1 U16673 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15593), .S(n16338), .Z(
        P1_U3524) );
  MUX2_X1 U16674 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15594), .S(n16338), .Z(
        P1_U3523) );
  MUX2_X1 U16675 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15595), .S(n16338), .Z(
        P1_U3522) );
  MUX2_X1 U16676 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15596), .S(n16338), .Z(
        P1_U3521) );
  MUX2_X1 U16677 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15597), .S(n16338), .Z(
        P1_U3520) );
  MUX2_X1 U16678 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15598), .S(n16338), .Z(
        P1_U3519) );
  MUX2_X1 U16679 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15599), .S(n16338), .Z(
        P1_U3518) );
  MUX2_X1 U16680 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15600), .S(n16338), .Z(
        P1_U3517) );
  MUX2_X1 U16681 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15601), .S(n16338), .Z(
        P1_U3516) );
  MUX2_X1 U16682 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15602), .S(n16338), .Z(
        P1_U3515) );
  MUX2_X1 U16683 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15603), .S(n16338), .Z(
        P1_U3513) );
  MUX2_X1 U16684 ( .A(n15604), .B(P1_REG0_REG_17__SCAN_IN), .S(n16447), .Z(
        P1_U3510) );
  MUX2_X1 U16685 ( .A(n15605), .B(P1_REG0_REG_16__SCAN_IN), .S(n16447), .Z(
        P1_U3507) );
  MUX2_X1 U16686 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15606), .S(n16338), .Z(
        P1_U3504) );
  MUX2_X1 U16687 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15607), .S(n16338), .Z(
        P1_U3501) );
  MUX2_X1 U16689 ( .A(n15610), .B(P1_D_REG_1__SCAN_IN), .S(n7430), .Z(P1_U3446) );
  MUX2_X1 U16690 ( .A(n15611), .B(P1_D_REG_0__SCAN_IN), .S(n7430), .Z(P1_U3445) );
  NAND2_X1 U16691 ( .A1(n10701), .A2(n15612), .ZN(n15615) );
  OR4_X1 U16692 ( .A1(n15613), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10291), .A4(
        P1_U3086), .ZN(n15614) );
  OAI211_X1 U16693 ( .C1(n10703), .C2(n7555), .A(n15615), .B(n15614), .ZN(
        P1_U3324) );
  OAI222_X1 U16694 ( .A1(P1_U3086), .A2(n15621), .B1(n15627), .B2(n15620), 
        .C1(n15619), .C2(n7555), .ZN(P1_U3326) );
  OAI222_X1 U16695 ( .A1(P1_U3086), .A2(n15628), .B1(n15627), .B2(n15626), 
        .C1(n7735), .C2(n7555), .ZN(P1_U3329) );
  MUX2_X1 U16696 ( .A(n15630), .B(n15629), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16697 ( .A(n15631), .ZN(n15632) );
  MUX2_X1 U16698 ( .A(n15632), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16699 ( .A(SI_31_), .B(keyinput_129), .ZN(n15636) );
  XNOR2_X1 U16700 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n15635) );
  OAI21_X1 U16701 ( .B1(n15636), .B2(n15635), .A(n15634), .ZN(n15640) );
  XOR2_X1 U16702 ( .A(SI_30_), .B(keyinput_130), .Z(n15639) );
  XNOR2_X1 U16703 ( .A(n15637), .B(keyinput_132), .ZN(n15638) );
  XOR2_X1 U16704 ( .A(SI_27_), .B(keyinput_133), .Z(n15642) );
  XNOR2_X1 U16705 ( .A(SI_26_), .B(keyinput_134), .ZN(n15641) );
  NOR3_X1 U16706 ( .A1(n15643), .A2(n15642), .A3(n15641), .ZN(n15647) );
  XNOR2_X1 U16707 ( .A(n15644), .B(keyinput_135), .ZN(n15646) );
  XOR2_X1 U16708 ( .A(SI_24_), .B(keyinput_136), .Z(n15645) );
  XNOR2_X1 U16709 ( .A(SI_23_), .B(keyinput_137), .ZN(n15649) );
  XNOR2_X1 U16710 ( .A(SI_22_), .B(keyinput_138), .ZN(n15648) );
  OAI21_X1 U16711 ( .B1(n15650), .B2(n15649), .A(n15648), .ZN(n15653) );
  XNOR2_X1 U16712 ( .A(n15839), .B(keyinput_140), .ZN(n15652) );
  XNOR2_X1 U16713 ( .A(SI_21_), .B(keyinput_139), .ZN(n15651) );
  NAND3_X1 U16714 ( .A1(n15653), .A2(n15652), .A3(n15651), .ZN(n15656) );
  XNOR2_X1 U16715 ( .A(SI_19_), .B(keyinput_141), .ZN(n15655) );
  XNOR2_X1 U16716 ( .A(n15843), .B(keyinput_142), .ZN(n15654) );
  AOI21_X1 U16717 ( .B1(n15656), .B2(n15655), .A(n15654), .ZN(n15660) );
  XNOR2_X1 U16718 ( .A(n15657), .B(keyinput_143), .ZN(n15659) );
  XNOR2_X1 U16719 ( .A(SI_16_), .B(keyinput_144), .ZN(n15658) );
  XNOR2_X1 U16720 ( .A(SI_15_), .B(keyinput_145), .ZN(n15662) );
  XNOR2_X1 U16721 ( .A(n15851), .B(keyinput_146), .ZN(n15661) );
  AOI21_X1 U16722 ( .B1(n15663), .B2(n15662), .A(n15661), .ZN(n15667) );
  XNOR2_X1 U16723 ( .A(n15857), .B(keyinput_149), .ZN(n15666) );
  XNOR2_X1 U16724 ( .A(SI_12_), .B(keyinput_148), .ZN(n15665) );
  XNOR2_X1 U16725 ( .A(SI_13_), .B(keyinput_147), .ZN(n15664) );
  XOR2_X1 U16726 ( .A(SI_8_), .B(keyinput_152), .Z(n15670) );
  XOR2_X1 U16727 ( .A(SI_9_), .B(keyinput_151), .Z(n15669) );
  XNOR2_X1 U16728 ( .A(SI_10_), .B(keyinput_150), .ZN(n15668) );
  NOR4_X1 U16729 ( .A1(n15671), .A2(n15670), .A3(n15669), .A4(n15668), .ZN(
        n15675) );
  XOR2_X1 U16730 ( .A(SI_6_), .B(keyinput_154), .Z(n15674) );
  XOR2_X1 U16731 ( .A(SI_7_), .B(keyinput_153), .Z(n15673) );
  XNOR2_X1 U16732 ( .A(SI_5_), .B(keyinput_155), .ZN(n15672) );
  XOR2_X1 U16733 ( .A(SI_4_), .B(keyinput_156), .Z(n15677) );
  XOR2_X1 U16734 ( .A(SI_3_), .B(keyinput_157), .Z(n15676) );
  OAI21_X1 U16735 ( .B1(n15678), .B2(n15677), .A(n15676), .ZN(n15681) );
  XNOR2_X1 U16736 ( .A(SI_2_), .B(keyinput_158), .ZN(n15680) );
  XOR2_X1 U16737 ( .A(SI_1_), .B(keyinput_159), .Z(n15679) );
  AOI21_X1 U16738 ( .B1(n15681), .B2(n15680), .A(n15679), .ZN(n15684) );
  INV_X1 U16739 ( .A(P3_RD_REG_SCAN_IN), .ZN(n16293) );
  XNOR2_X1 U16740 ( .A(n16293), .B(keyinput_161), .ZN(n15683) );
  XNOR2_X1 U16741 ( .A(SI_0_), .B(keyinput_160), .ZN(n15682) );
  NOR3_X1 U16742 ( .A1(n15684), .A2(n15683), .A3(n15682), .ZN(n15688) );
  XNOR2_X1 U16743 ( .A(P3_U3151), .B(keyinput_162), .ZN(n15687) );
  XOR2_X1 U16744 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .Z(n15686) );
  XNOR2_X1 U16745 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n15685)
         );
  XOR2_X1 U16746 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n15690)
         );
  XOR2_X1 U16747 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n15689)
         );
  OAI21_X1 U16748 ( .B1(n15691), .B2(n15690), .A(n15689), .ZN(n15700) );
  XOR2_X1 U16749 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n15699)
         );
  XOR2_X1 U16750 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .Z(n15694)
         );
  XNOR2_X1 U16751 ( .A(n15892), .B(keyinput_171), .ZN(n15693) );
  XNOR2_X1 U16752 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n15692)
         );
  NOR3_X1 U16753 ( .A1(n15694), .A2(n15693), .A3(n15692), .ZN(n15697) );
  XNOR2_X1 U16754 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n15696)
         );
  XNOR2_X1 U16755 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n15695)
         );
  NAND3_X1 U16756 ( .A1(n15697), .A2(n15696), .A3(n15695), .ZN(n15698) );
  AOI21_X1 U16757 ( .B1(n15700), .B2(n15699), .A(n15698), .ZN(n15705) );
  XNOR2_X1 U16758 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n15704)
         );
  XNOR2_X1 U16759 ( .A(n15701), .B(keyinput_175), .ZN(n15703) );
  XNOR2_X1 U16760 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n15702)
         );
  OAI211_X1 U16761 ( .C1(n15705), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        n15709) );
  XNOR2_X1 U16762 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n15708)
         );
  XNOR2_X1 U16763 ( .A(n15902), .B(keyinput_177), .ZN(n15707) );
  XNOR2_X1 U16764 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n15706)
         );
  XNOR2_X1 U16765 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_179), .ZN(n15711)
         );
  XNOR2_X1 U16766 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n15710)
         );
  NOR3_X1 U16767 ( .A1(n15712), .A2(n15711), .A3(n15710), .ZN(n15716) );
  XNOR2_X1 U16768 ( .A(n15713), .B(keyinput_181), .ZN(n15715) );
  XNOR2_X1 U16769 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n15714)
         );
  XNOR2_X1 U16770 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_183), .ZN(n15718)
         );
  XNOR2_X1 U16771 ( .A(P3_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n15717)
         );
  NOR3_X1 U16772 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(n15722) );
  XOR2_X1 U16773 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n15721)
         );
  XNOR2_X1 U16774 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n15720)
         );
  XNOR2_X1 U16775 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n15725)
         );
  XOR2_X1 U16776 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .Z(n15724) );
  XOR2_X1 U16777 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .Z(n15723)
         );
  OAI211_X1 U16778 ( .C1(n15726), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15730) );
  XNOR2_X1 U16779 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_190), .ZN(n15729)
         );
  XOR2_X1 U16780 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .Z(n15728)
         );
  XOR2_X1 U16781 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_192), .Z(n15727) );
  XNOR2_X1 U16782 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n15732) );
  XOR2_X1 U16783 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .Z(n15731)
         );
  OAI21_X1 U16784 ( .B1(n15733), .B2(n15732), .A(n15731), .ZN(n15736) );
  XNOR2_X1 U16785 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n15735) );
  XNOR2_X1 U16786 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n15734) );
  XOR2_X1 U16787 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .Z(n15738)
         );
  XOR2_X1 U16788 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n15737)
         );
  NOR3_X1 U16789 ( .A1(n15739), .A2(n15738), .A3(n15737), .ZN(n15743) );
  XNOR2_X1 U16790 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n15742) );
  XNOR2_X1 U16791 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .ZN(n15741) );
  XNOR2_X1 U16792 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n15740) );
  XOR2_X1 U16793 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .Z(n15748)
         );
  XOR2_X1 U16794 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n15747)
         );
  OAI22_X1 U16795 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_203), .B1(
        P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_204), .ZN(n15745) );
  AND2_X1 U16796 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_203), .ZN(
        n15744) );
  AOI211_X1 U16797 ( .C1(keyinput_204), .C2(P3_DATAO_REG_20__SCAN_IN), .A(
        n15745), .B(n15744), .ZN(n15746) );
  OAI211_X1 U16798 ( .C1(n15749), .C2(n15748), .A(n15747), .B(n15746), .ZN(
        n15752) );
  XOR2_X1 U16799 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n15751)
         );
  XOR2_X1 U16800 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .Z(n15750)
         );
  NAND3_X1 U16801 ( .A1(n15752), .A2(n15751), .A3(n15750), .ZN(n15755) );
  XOR2_X1 U16802 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .Z(n15754)
         );
  XOR2_X1 U16803 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n15753)
         );
  NAND3_X1 U16804 ( .A1(n15755), .A2(n15754), .A3(n15753), .ZN(n15759) );
  XOR2_X1 U16805 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n15758)
         );
  XOR2_X1 U16806 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n15757)
         );
  XOR2_X1 U16807 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n15756)
         );
  INV_X1 U16808 ( .A(keyinput_214), .ZN(n15760) );
  XNOR2_X1 U16809 ( .A(n15760), .B(P3_DATAO_REG_10__SCAN_IN), .ZN(n15764) );
  XNOR2_X1 U16810 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n15763)
         );
  XNOR2_X1 U16811 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n15762)
         );
  XNOR2_X1 U16812 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n15761) );
  NAND4_X1 U16813 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15766) );
  XNOR2_X1 U16814 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n15765)
         );
  OAI21_X1 U16815 ( .B1(n15767), .B2(n15766), .A(n15765), .ZN(n15770) );
  XNOR2_X1 U16816 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n15769)
         );
  XNOR2_X1 U16817 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_219), .ZN(n15768)
         );
  XOR2_X1 U16818 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_220), .Z(n15772)
         );
  XNOR2_X1 U16819 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n15771)
         );
  XOR2_X1 U16820 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_222), .Z(n15774)
         );
  XOR2_X1 U16821 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_223), .Z(n15773)
         );
  NAND3_X1 U16822 ( .A1(n15775), .A2(n15774), .A3(n15773), .ZN(n15779) );
  XNOR2_X1 U16823 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_224), .ZN(n15778)
         );
  XOR2_X1 U16824 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_225), .Z(n15777) );
  XNOR2_X1 U16825 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_226), .ZN(n15776)
         );
  AOI211_X1 U16826 ( .C1(n15779), .C2(n15778), .A(n15777), .B(n15776), .ZN(
        n15782) );
  XOR2_X1 U16827 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_227), .Z(n15781) );
  XNOR2_X1 U16828 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_228), .ZN(n15780)
         );
  XOR2_X1 U16829 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_229), .Z(n15785) );
  XNOR2_X1 U16830 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .ZN(n15784)
         );
  XNOR2_X1 U16831 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_230), .ZN(n15783)
         );
  AOI211_X1 U16832 ( .C1(n15786), .C2(n15785), .A(n15784), .B(n15783), .ZN(
        n15789) );
  XOR2_X1 U16833 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_232), .Z(n15788) );
  XNOR2_X1 U16834 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_233), .ZN(n15787)
         );
  OAI21_X1 U16835 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n15797) );
  XNOR2_X1 U16836 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .ZN(n15792) );
  XNOR2_X1 U16837 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n15791)
         );
  XNOR2_X1 U16838 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .ZN(n15790) );
  NOR3_X1 U16839 ( .A1(n15792), .A2(n15791), .A3(n15790), .ZN(n15796) );
  XNOR2_X1 U16840 ( .A(n7858), .B(keyinput_238), .ZN(n15795) );
  XNOR2_X1 U16841 ( .A(n15793), .B(keyinput_237), .ZN(n15794) );
  XOR2_X1 U16842 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .Z(n15801) );
  XNOR2_X1 U16843 ( .A(n15995), .B(keyinput_241), .ZN(n15800) );
  XNOR2_X1 U16844 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_240), .ZN(n15799) );
  XNOR2_X1 U16845 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n15798) );
  NAND4_X1 U16846 ( .A1(n15801), .A2(n15800), .A3(n15799), .A4(n15798), .ZN(
        n15803) );
  XNOR2_X1 U16847 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_243), .ZN(n15802) );
  OAI21_X1 U16848 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n15809) );
  XNOR2_X1 U16849 ( .A(n15805), .B(keyinput_245), .ZN(n15808) );
  XNOR2_X1 U16850 ( .A(n15806), .B(keyinput_244), .ZN(n15807) );
  NAND3_X1 U16851 ( .A1(n15809), .A2(n15808), .A3(n15807), .ZN(n15816) );
  XOR2_X1 U16852 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .Z(n15812) );
  XNOR2_X1 U16853 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_248), .ZN(n15811)
         );
  XNOR2_X1 U16854 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_247), .ZN(n15810)
         );
  NOR3_X1 U16855 ( .A1(n15812), .A2(n15811), .A3(n15810), .ZN(n15815) );
  XNOR2_X1 U16856 ( .A(n16013), .B(keyinput_249), .ZN(n15814) );
  XNOR2_X1 U16857 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n15813)
         );
  AOI211_X1 U16858 ( .C1(n15816), .C2(n15815), .A(n15814), .B(n15813), .ZN(
        n15820) );
  XNOR2_X1 U16859 ( .A(n16017), .B(keyinput_251), .ZN(n15819) );
  XNOR2_X1 U16860 ( .A(n16018), .B(keyinput_252), .ZN(n15818) );
  XNOR2_X1 U16861 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_253), .ZN(n15817)
         );
  OAI211_X1 U16862 ( .C1(n15820), .C2(n15819), .A(n15818), .B(n15817), .ZN(
        n15823) );
  XNOR2_X1 U16863 ( .A(n16023), .B(keyinput_254), .ZN(n15822) );
  XNOR2_X1 U16864 ( .A(keyinput_127), .B(keyinput_255), .ZN(n15821) );
  AOI21_X1 U16865 ( .B1(n15823), .B2(n15822), .A(n15821), .ZN(n16029) );
  XOR2_X1 U16866 ( .A(SI_31_), .B(keyinput_1), .Z(n15826) );
  XOR2_X1 U16867 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n15825) );
  XNOR2_X1 U16868 ( .A(SI_29_), .B(keyinput_3), .ZN(n15824) );
  AOI21_X1 U16869 ( .B1(n15826), .B2(n15825), .A(n15824), .ZN(n15829) );
  XOR2_X1 U16870 ( .A(SI_30_), .B(keyinput_2), .Z(n15828) );
  XNOR2_X1 U16871 ( .A(SI_28_), .B(keyinput_4), .ZN(n15827) );
  NAND3_X1 U16872 ( .A1(n15829), .A2(n15828), .A3(n15827), .ZN(n15832) );
  XNOR2_X1 U16873 ( .A(SI_26_), .B(keyinput_6), .ZN(n15831) );
  XNOR2_X1 U16874 ( .A(SI_27_), .B(keyinput_5), .ZN(n15830) );
  NAND3_X1 U16875 ( .A1(n15832), .A2(n15831), .A3(n15830), .ZN(n15835) );
  XNOR2_X1 U16876 ( .A(SI_25_), .B(keyinput_7), .ZN(n15834) );
  XNOR2_X1 U16877 ( .A(SI_24_), .B(keyinput_8), .ZN(n15833) );
  NAND3_X1 U16878 ( .A1(n15835), .A2(n15834), .A3(n15833), .ZN(n15838) );
  XNOR2_X1 U16879 ( .A(SI_23_), .B(keyinput_9), .ZN(n15837) );
  XNOR2_X1 U16880 ( .A(SI_22_), .B(keyinput_10), .ZN(n15836) );
  AOI21_X1 U16881 ( .B1(n15838), .B2(n15837), .A(n15836), .ZN(n15842) );
  XOR2_X1 U16882 ( .A(SI_21_), .B(keyinput_11), .Z(n15841) );
  XNOR2_X1 U16883 ( .A(n15839), .B(keyinput_12), .ZN(n15840) );
  NOR3_X1 U16884 ( .A1(n15842), .A2(n15841), .A3(n15840), .ZN(n15846) );
  XNOR2_X1 U16885 ( .A(SI_19_), .B(keyinput_13), .ZN(n15845) );
  XNOR2_X1 U16886 ( .A(n15843), .B(keyinput_14), .ZN(n15844) );
  OAI21_X1 U16887 ( .B1(n15846), .B2(n15845), .A(n15844), .ZN(n15849) );
  XNOR2_X1 U16888 ( .A(SI_17_), .B(keyinput_15), .ZN(n15848) );
  XNOR2_X1 U16889 ( .A(SI_16_), .B(keyinput_16), .ZN(n15847) );
  AOI21_X1 U16890 ( .B1(n15849), .B2(n15848), .A(n15847), .ZN(n15854) );
  XNOR2_X1 U16891 ( .A(n15850), .B(keyinput_17), .ZN(n15853) );
  XNOR2_X1 U16892 ( .A(n15851), .B(keyinput_18), .ZN(n15852) );
  OAI21_X1 U16893 ( .B1(n15854), .B2(n15853), .A(n15852), .ZN(n15861) );
  XNOR2_X1 U16894 ( .A(n15855), .B(keyinput_19), .ZN(n15860) );
  XNOR2_X1 U16895 ( .A(n15856), .B(keyinput_20), .ZN(n15859) );
  XNOR2_X1 U16896 ( .A(n15857), .B(keyinput_21), .ZN(n15858) );
  NAND4_X1 U16897 ( .A1(n15861), .A2(n15860), .A3(n15859), .A4(n15858), .ZN(
        n15865) );
  XOR2_X1 U16898 ( .A(SI_8_), .B(keyinput_24), .Z(n15864) );
  XNOR2_X1 U16899 ( .A(SI_9_), .B(keyinput_23), .ZN(n15863) );
  XNOR2_X1 U16900 ( .A(SI_10_), .B(keyinput_22), .ZN(n15862) );
  NAND4_X1 U16901 ( .A1(n15865), .A2(n15864), .A3(n15863), .A4(n15862), .ZN(
        n15869) );
  XOR2_X1 U16902 ( .A(SI_5_), .B(keyinput_27), .Z(n15868) );
  XOR2_X1 U16903 ( .A(SI_7_), .B(keyinput_25), .Z(n15867) );
  XNOR2_X1 U16904 ( .A(SI_6_), .B(keyinput_26), .ZN(n15866) );
  NAND4_X1 U16905 ( .A1(n15869), .A2(n15868), .A3(n15867), .A4(n15866), .ZN(
        n15872) );
  XOR2_X1 U16906 ( .A(SI_4_), .B(keyinput_28), .Z(n15871) );
  XNOR2_X1 U16907 ( .A(SI_3_), .B(keyinput_29), .ZN(n15870) );
  AOI21_X1 U16908 ( .B1(n15872), .B2(n15871), .A(n15870), .ZN(n15876) );
  XNOR2_X1 U16909 ( .A(n15873), .B(keyinput_30), .ZN(n15875) );
  XNOR2_X1 U16910 ( .A(SI_1_), .B(keyinput_31), .ZN(n15874) );
  OAI21_X1 U16911 ( .B1(n15876), .B2(n15875), .A(n15874), .ZN(n15879) );
  XNOR2_X1 U16912 ( .A(n16293), .B(keyinput_33), .ZN(n15878) );
  XOR2_X1 U16913 ( .A(SI_0_), .B(keyinput_32), .Z(n15877) );
  NAND3_X1 U16914 ( .A1(n15879), .A2(n15878), .A3(n15877), .ZN(n15883) );
  XOR2_X1 U16915 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n15882) );
  XNOR2_X1 U16916 ( .A(P3_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n15881) );
  XNOR2_X1 U16917 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n15880)
         );
  NAND4_X1 U16918 ( .A1(n15883), .A2(n15882), .A3(n15881), .A4(n15880), .ZN(
        n15886) );
  XNOR2_X1 U16919 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n15885)
         );
  XNOR2_X1 U16920 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n15884)
         );
  AOI21_X1 U16921 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n15888) );
  XNOR2_X1 U16922 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n15887)
         );
  NOR2_X1 U16923 ( .A1(n15888), .A2(n15887), .ZN(n15896) );
  INV_X1 U16924 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15890) );
  AOI22_X1 U16925 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_42), .B1(n15890), .B2(keyinput_41), .ZN(n15889) );
  OAI221_X1 U16926 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .C1(
        n15890), .C2(keyinput_41), .A(n15889), .ZN(n15895) );
  AOI22_X1 U16927 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(n15892), 
        .B2(keyinput_43), .ZN(n15891) );
  OAI221_X1 U16928 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n15892), .C2(keyinput_43), .A(n15891), .ZN(n15894) );
  XNOR2_X1 U16929 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n15893)
         );
  NOR4_X1 U16930 ( .A1(n15896), .A2(n15895), .A3(n15894), .A4(n15893), .ZN(
        n15901) );
  XNOR2_X1 U16931 ( .A(n15897), .B(keyinput_45), .ZN(n15900) );
  XOR2_X1 U16932 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .Z(n15899) );
  XNOR2_X1 U16933 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n15898)
         );
  OAI211_X1 U16934 ( .C1(n15901), .C2(n15900), .A(n15899), .B(n15898), .ZN(
        n15906) );
  XNOR2_X1 U16935 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n15905)
         );
  XNOR2_X1 U16936 ( .A(n15902), .B(keyinput_49), .ZN(n15904) );
  XNOR2_X1 U16937 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n15903)
         );
  AOI211_X1 U16938 ( .C1(n15906), .C2(n15905), .A(n15904), .B(n15903), .ZN(
        n15909) );
  XOR2_X1 U16939 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n15908) );
  XNOR2_X1 U16940 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n15907)
         );
  NOR3_X1 U16941 ( .A1(n15909), .A2(n15908), .A3(n15907), .ZN(n15912) );
  XNOR2_X1 U16942 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n15911)
         );
  XNOR2_X1 U16943 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n15910)
         );
  NOR3_X1 U16944 ( .A1(n15912), .A2(n15911), .A3(n15910), .ZN(n15917) );
  XNOR2_X1 U16945 ( .A(n15913), .B(keyinput_55), .ZN(n15916) );
  XNOR2_X1 U16946 ( .A(n15914), .B(keyinput_56), .ZN(n15915) );
  NOR3_X1 U16947 ( .A1(n15917), .A2(n15916), .A3(n15915), .ZN(n15920) );
  XNOR2_X1 U16948 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n15919)
         );
  XNOR2_X1 U16949 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n15918)
         );
  NOR3_X1 U16950 ( .A1(n15920), .A2(n15919), .A3(n15918), .ZN(n15924) );
  XNOR2_X1 U16951 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n15923)
         );
  XOR2_X1 U16952 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .Z(n15922) );
  XNOR2_X1 U16953 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n15921)
         );
  OAI211_X1 U16954 ( .C1(n15924), .C2(n15923), .A(n15922), .B(n15921), .ZN(
        n15928) );
  XNOR2_X1 U16955 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n15927)
         );
  XOR2_X1 U16956 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_63), .Z(n15926) );
  XOR2_X1 U16957 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .Z(n15925) );
  AOI211_X1 U16958 ( .C1(n15928), .C2(n15927), .A(n15926), .B(n15925), .ZN(
        n15931) );
  XNOR2_X1 U16959 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .ZN(n15930)
         );
  XOR2_X1 U16960 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n15929)
         );
  OAI21_X1 U16961 ( .B1(n15931), .B2(n15930), .A(n15929), .ZN(n15934) );
  XNOR2_X1 U16962 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n15933)
         );
  XOR2_X1 U16963 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n15932)
         );
  AOI21_X1 U16964 ( .B1(n15934), .B2(n15933), .A(n15932), .ZN(n15937) );
  XOR2_X1 U16965 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .Z(n15936)
         );
  XNOR2_X1 U16966 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n15935)
         );
  NOR3_X1 U16967 ( .A1(n15937), .A2(n15936), .A3(n15935), .ZN(n15941) );
  XOR2_X1 U16968 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n15940)
         );
  XOR2_X1 U16969 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n15939)
         );
  XNOR2_X1 U16970 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n15938)
         );
  NOR4_X1 U16971 ( .A1(n15941), .A2(n15940), .A3(n15939), .A4(n15938), .ZN(
        n15947) );
  XNOR2_X1 U16972 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n15946)
         );
  XOR2_X1 U16973 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n15944)
         );
  XOR2_X1 U16974 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n15943)
         );
  XOR2_X1 U16975 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .Z(n15942)
         );
  NOR3_X1 U16976 ( .A1(n15944), .A2(n15943), .A3(n15942), .ZN(n15945) );
  OAI21_X1 U16977 ( .B1(n15947), .B2(n15946), .A(n15945), .ZN(n15950) );
  XOR2_X1 U16978 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n15949)
         );
  XNOR2_X1 U16979 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n15948)
         );
  NAND3_X1 U16980 ( .A1(n15950), .A2(n15949), .A3(n15948), .ZN(n15953) );
  XOR2_X1 U16981 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n15952)
         );
  XNOR2_X1 U16982 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n15951)
         );
  NAND3_X1 U16983 ( .A1(n15953), .A2(n15952), .A3(n15951), .ZN(n15957) );
  XNOR2_X1 U16984 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n15956)
         );
  XOR2_X1 U16985 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .Z(n15955)
         );
  XOR2_X1 U16986 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n15954)
         );
  AOI211_X1 U16987 ( .C1(n15957), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        n15964) );
  XOR2_X1 U16988 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n15961) );
  XOR2_X1 U16989 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n15960)
         );
  XOR2_X1 U16990 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n15959) );
  XNOR2_X1 U16991 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n15958)
         );
  NAND4_X1 U16992 ( .A1(n15961), .A2(n15960), .A3(n15959), .A4(n15958), .ZN(
        n15963) );
  XNOR2_X1 U16993 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n15962)
         );
  OAI21_X1 U16994 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(n15967) );
  XNOR2_X1 U16995 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n15966)
         );
  XOR2_X1 U16996 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .Z(n15965) );
  AOI21_X1 U16997 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(n15970) );
  XOR2_X1 U16998 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .Z(n15969) );
  XNOR2_X1 U16999 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n15968)
         );
  OAI21_X1 U17000 ( .B1(n15970), .B2(n15969), .A(n15968), .ZN(n15973) );
  XOR2_X1 U17001 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .Z(n15972) );
  XOR2_X1 U17002 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .Z(n15971) );
  NAND3_X1 U17003 ( .A1(n15973), .A2(n15972), .A3(n15971), .ZN(n15977) );
  XNOR2_X1 U17004 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n15976)
         );
  XNOR2_X1 U17005 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .ZN(n15975)
         );
  XNOR2_X1 U17006 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .ZN(n15974)
         );
  AOI211_X1 U17007 ( .C1(n15977), .C2(n15976), .A(n15975), .B(n15974), .ZN(
        n15980) );
  XNOR2_X1 U17008 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .ZN(n15979)
         );
  XNOR2_X1 U17009 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .ZN(n15978)
         );
  NOR3_X1 U17010 ( .A1(n15980), .A2(n15979), .A3(n15978), .ZN(n15984) );
  XNOR2_X1 U17011 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .ZN(n15983)
         );
  XOR2_X1 U17012 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .Z(n15982) );
  XNOR2_X1 U17013 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .ZN(n15981)
         );
  OAI211_X1 U17014 ( .C1(n15984), .C2(n15983), .A(n15982), .B(n15981), .ZN(
        n15987) );
  XNOR2_X1 U17015 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .ZN(n15986)
         );
  XNOR2_X1 U17016 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n15985)
         );
  AOI21_X1 U17017 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n15991) );
  XNOR2_X1 U17018 ( .A(n16195), .B(keyinput_107), .ZN(n15990) );
  XNOR2_X1 U17019 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n15989)
         );
  XNOR2_X1 U17020 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n15988) );
  NOR4_X1 U17021 ( .A1(n15991), .A2(n15990), .A3(n15989), .A4(n15988), .ZN(
        n15994) );
  XNOR2_X1 U17022 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .ZN(n15993) );
  XNOR2_X1 U17023 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_109), .ZN(n15992) );
  NOR3_X1 U17024 ( .A1(n15994), .A2(n15993), .A3(n15992), .ZN(n16002) );
  XNOR2_X1 U17025 ( .A(n15995), .B(keyinput_113), .ZN(n15999) );
  XNOR2_X1 U17026 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .ZN(n15998) );
  XNOR2_X1 U17027 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_112), .ZN(n15997) );
  XNOR2_X1 U17028 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15996) );
  NAND4_X1 U17029 ( .A1(n15999), .A2(n15998), .A3(n15997), .A4(n15996), .ZN(
        n16001) );
  XNOR2_X1 U17030 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_115), .ZN(n16000) );
  OAI21_X1 U17031 ( .B1(n16002), .B2(n16001), .A(n16000), .ZN(n16005) );
  XNOR2_X1 U17032 ( .A(n15805), .B(keyinput_117), .ZN(n16004) );
  XNOR2_X1 U17033 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_116), .ZN(n16003) );
  NAND3_X1 U17034 ( .A1(n16005), .A2(n16004), .A3(n16003), .ZN(n16011) );
  XOR2_X1 U17035 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_118), .Z(n16010) );
  XNOR2_X1 U17036 ( .A(n16006), .B(keyinput_119), .ZN(n16009) );
  XNOR2_X1 U17037 ( .A(n16007), .B(keyinput_120), .ZN(n16008) );
  NAND4_X1 U17038 ( .A1(n16011), .A2(n16010), .A3(n16009), .A4(n16008), .ZN(
        n16016) );
  XNOR2_X1 U17039 ( .A(n16012), .B(keyinput_122), .ZN(n16015) );
  XNOR2_X1 U17040 ( .A(n16013), .B(keyinput_121), .ZN(n16014) );
  NAND3_X1 U17041 ( .A1(n16016), .A2(n16015), .A3(n16014), .ZN(n16022) );
  XNOR2_X1 U17042 ( .A(n16017), .B(keyinput_123), .ZN(n16021) );
  XNOR2_X1 U17043 ( .A(n16018), .B(keyinput_124), .ZN(n16020) );
  XNOR2_X1 U17044 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n16019)
         );
  AOI211_X1 U17045 ( .C1(n16022), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        n16027) );
  XNOR2_X1 U17046 ( .A(n16023), .B(keyinput_126), .ZN(n16026) );
  XNOR2_X1 U17047 ( .A(n16024), .B(keyinput_127), .ZN(n16025) );
  OAI21_X1 U17048 ( .B1(n16027), .B2(n16026), .A(n16025), .ZN(n16028) );
  AND2_X1 U17049 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n7430), .ZN(P1_U3323) );
  AND2_X1 U17050 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n7430), .ZN(P1_U3322) );
  AND2_X1 U17051 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n7430), .ZN(P1_U3321) );
  AND2_X1 U17052 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n7430), .ZN(P1_U3320) );
  AND2_X1 U17053 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n7430), .ZN(P1_U3319) );
  AND2_X1 U17054 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n7430), .ZN(P1_U3318) );
  AND2_X1 U17055 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n7430), .ZN(P1_U3317) );
  AND2_X1 U17056 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n7430), .ZN(P1_U3316) );
  AND2_X1 U17057 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n7430), .ZN(P1_U3315) );
  AND2_X1 U17058 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n7430), .ZN(P1_U3314) );
  AND2_X1 U17059 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n7430), .ZN(P1_U3313) );
  AND2_X1 U17060 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n7430), .ZN(P1_U3312) );
  AND2_X1 U17061 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n7430), .ZN(P1_U3311) );
  AND2_X1 U17062 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n7430), .ZN(P1_U3310) );
  AND2_X1 U17063 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n7430), .ZN(P1_U3309) );
  AND2_X1 U17064 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n7430), .ZN(P1_U3308) );
  AND2_X1 U17065 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n7430), .ZN(P1_U3307) );
  AND2_X1 U17066 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n7430), .ZN(P1_U3306) );
  AND2_X1 U17067 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n7430), .ZN(P1_U3305) );
  AND2_X1 U17068 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n7430), .ZN(P1_U3304) );
  AND2_X1 U17069 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n7430), .ZN(P1_U3303) );
  AND2_X1 U17070 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n7430), .ZN(P1_U3302) );
  AND2_X1 U17071 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n7430), .ZN(P1_U3301) );
  AND2_X1 U17072 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n7430), .ZN(P1_U3300) );
  AND2_X1 U17073 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n7430), .ZN(P1_U3299) );
  AND2_X1 U17074 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n7430), .ZN(P1_U3298) );
  AND2_X1 U17075 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n7430), .ZN(P1_U3297) );
  AND2_X1 U17076 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n7430), .ZN(P1_U3296) );
  AND2_X1 U17077 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n7430), .ZN(P1_U3295) );
  AND2_X1 U17078 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n7430), .ZN(P1_U3294) );
  INV_X1 U17079 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16034) );
  AOI21_X1 U17080 ( .B1(n16034), .B2(n16038), .A(n16033), .ZN(P2_U3417) );
  AND2_X1 U17081 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n16036), .ZN(P2_U3295) );
  AND2_X1 U17082 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n16036), .ZN(P2_U3294) );
  AND2_X1 U17083 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n16036), .ZN(P2_U3293) );
  AND2_X1 U17084 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n16036), .ZN(P2_U3292) );
  AND2_X1 U17085 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n16036), .ZN(P2_U3291) );
  AND2_X1 U17086 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n16036), .ZN(P2_U3290) );
  AND2_X1 U17087 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n16036), .ZN(P2_U3289) );
  AND2_X1 U17088 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n16036), .ZN(P2_U3288) );
  AND2_X1 U17089 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n16036), .ZN(P2_U3287) );
  AND2_X1 U17090 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n16036), .ZN(P2_U3286) );
  AND2_X1 U17091 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n16036), .ZN(P2_U3285) );
  AND2_X1 U17092 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n16036), .ZN(P2_U3284) );
  AND2_X1 U17093 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n16036), .ZN(P2_U3283) );
  AND2_X1 U17094 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n16036), .ZN(P2_U3282) );
  AND2_X1 U17095 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n16036), .ZN(P2_U3281) );
  AND2_X1 U17096 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n16036), .ZN(P2_U3280) );
  AND2_X1 U17097 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n16036), .ZN(P2_U3279) );
  AND2_X1 U17098 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n16036), .ZN(P2_U3278) );
  AND2_X1 U17099 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n16036), .ZN(P2_U3277) );
  AND2_X1 U17100 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n16036), .ZN(P2_U3276) );
  AND2_X1 U17101 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n16036), .ZN(P2_U3275) );
  AND2_X1 U17102 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n16036), .ZN(P2_U3274) );
  AND2_X1 U17103 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n16036), .ZN(P2_U3273) );
  AND2_X1 U17104 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n16036), .ZN(P2_U3272) );
  AND2_X1 U17105 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n16036), .ZN(P2_U3271) );
  AND2_X1 U17106 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n16036), .ZN(P2_U3270) );
  AND2_X1 U17107 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n16036), .ZN(P2_U3269) );
  AND2_X1 U17108 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n16036), .ZN(P2_U3268) );
  AND2_X1 U17109 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n16036), .ZN(P2_U3267) );
  AND2_X1 U17110 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n16036), .ZN(P2_U3266) );
  NOR2_X1 U17111 ( .A1(n16055), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17112 ( .A1(P3_U3897), .A2(n16037), .ZN(P3_U3150) );
  INV_X1 U17113 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U17114 ( .A1(n16041), .A2(n16040), .B1(n16039), .B2(n16038), .ZN(
        P2_U3416) );
  OAI21_X1 U17115 ( .B1(n16043), .B2(n16042), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n16044) );
  OAI21_X1 U17116 ( .B1(P2_STATE_REG_SCAN_IN), .B2(P2_REG3_REG_2__SCAN_IN), 
        .A(n16044), .ZN(n16057) );
  OAI211_X1 U17117 ( .C1(n16047), .C2(n16046), .A(n16171), .B(n16045), .ZN(
        n16048) );
  INV_X1 U17118 ( .A(n16048), .ZN(n16054) );
  OAI211_X1 U17119 ( .C1(n16051), .C2(n16050), .A(n16163), .B(n16049), .ZN(
        n16052) );
  INV_X1 U17120 ( .A(n16052), .ZN(n16053) );
  AOI211_X1 U17121 ( .C1(n16055), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n16054), .B(
        n16053), .ZN(n16056) );
  NAND2_X1 U17122 ( .A1(n16057), .A2(n16056), .ZN(P2_U3216) );
  INV_X1 U17123 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n16071) );
  OAI211_X1 U17124 ( .C1(n16060), .C2(n16059), .A(n16163), .B(n16058), .ZN(
        n16066) );
  OAI21_X1 U17125 ( .B1(n16063), .B2(n16062), .A(n16061), .ZN(n16064) );
  OR2_X1 U17126 ( .A1(n16182), .A2(n16064), .ZN(n16065) );
  OAI211_X1 U17127 ( .C1(n16168), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        n16068) );
  INV_X1 U17128 ( .A(n16068), .ZN(n16070) );
  NAND2_X1 U17129 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n16069) );
  OAI211_X1 U17130 ( .C1(n16191), .C2(n16071), .A(n16070), .B(n16069), .ZN(
        P2_U3217) );
  OAI21_X1 U17131 ( .B1(n16074), .B2(n16073), .A(n16072), .ZN(n16081) );
  OAI211_X1 U17132 ( .C1(n16077), .C2(n16076), .A(n16163), .B(n16075), .ZN(
        n16080) );
  NAND2_X1 U17133 ( .A1(n16188), .A2(n16078), .ZN(n16079) );
  OAI211_X1 U17134 ( .C1(n16182), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16082) );
  INV_X1 U17135 ( .A(n16082), .ZN(n16084) );
  OAI211_X1 U17136 ( .C1(n16191), .C2(n16085), .A(n16084), .B(n16083), .ZN(
        P2_U3218) );
  OAI211_X1 U17137 ( .C1(n16088), .C2(n16087), .A(n16171), .B(n16086), .ZN(
        n16093) );
  OAI211_X1 U17138 ( .C1(n16091), .C2(n16090), .A(n16163), .B(n16089), .ZN(
        n16092) );
  OAI211_X1 U17139 ( .C1(n16168), .C2(n16094), .A(n16093), .B(n16092), .ZN(
        n16095) );
  INV_X1 U17140 ( .A(n16095), .ZN(n16097) );
  OAI211_X1 U17141 ( .C1(n16191), .C2(n16212), .A(n16097), .B(n16096), .ZN(
        P2_U3219) );
  INV_X1 U17142 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n16251) );
  OAI211_X1 U17143 ( .C1(n16100), .C2(n16099), .A(n16171), .B(n16098), .ZN(
        n16105) );
  OAI211_X1 U17144 ( .C1(n16103), .C2(n16102), .A(n16163), .B(n16101), .ZN(
        n16104) );
  OAI211_X1 U17145 ( .C1(n16168), .C2(n16106), .A(n16105), .B(n16104), .ZN(
        n16107) );
  INV_X1 U17146 ( .A(n16107), .ZN(n16109) );
  OAI211_X1 U17147 ( .C1(n16191), .C2(n16251), .A(n16109), .B(n16108), .ZN(
        P2_U3220) );
  INV_X1 U17148 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n16122) );
  OAI211_X1 U17149 ( .C1(n16112), .C2(n16111), .A(n16171), .B(n16110), .ZN(
        n16117) );
  OAI211_X1 U17150 ( .C1(n16115), .C2(n16114), .A(n16163), .B(n16113), .ZN(
        n16116) );
  OAI211_X1 U17151 ( .C1(n16168), .C2(n16118), .A(n16117), .B(n16116), .ZN(
        n16119) );
  INV_X1 U17152 ( .A(n16119), .ZN(n16121) );
  OAI211_X1 U17153 ( .C1(n16191), .C2(n16122), .A(n16121), .B(n16120), .ZN(
        P2_U3221) );
  INV_X1 U17154 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n16135) );
  OAI211_X1 U17155 ( .C1(n16125), .C2(n16124), .A(n16123), .B(n16171), .ZN(
        n16130) );
  OAI211_X1 U17156 ( .C1(n16128), .C2(n16127), .A(n16126), .B(n16163), .ZN(
        n16129) );
  OAI211_X1 U17157 ( .C1(n16168), .C2(n16131), .A(n16130), .B(n16129), .ZN(
        n16132) );
  INV_X1 U17158 ( .A(n16132), .ZN(n16134) );
  OAI211_X1 U17159 ( .C1(n16191), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        P2_U3222) );
  OAI21_X1 U17160 ( .B1(n16138), .B2(n16137), .A(n16136), .ZN(n16139) );
  NAND2_X1 U17161 ( .A1(n16139), .A2(n16171), .ZN(n16144) );
  OAI211_X1 U17162 ( .C1(n16142), .C2(n16141), .A(n16140), .B(n16163), .ZN(
        n16143) );
  OAI211_X1 U17163 ( .C1(n16168), .C2(n16145), .A(n16144), .B(n16143), .ZN(
        n16146) );
  INV_X1 U17164 ( .A(n16146), .ZN(n16148) );
  NAND2_X1 U17165 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n16147)
         );
  OAI211_X1 U17166 ( .C1(n16225), .C2(n16191), .A(n16148), .B(n16147), .ZN(
        P2_U3225) );
  INV_X1 U17167 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n16161) );
  OAI21_X1 U17168 ( .B1(n16150), .B2(n16149), .A(n16171), .ZN(n16152) );
  NOR2_X1 U17169 ( .A1(n16152), .A2(n16151), .ZN(n16157) );
  AOI211_X1 U17170 ( .C1(n16155), .C2(n16154), .A(n16177), .B(n16153), .ZN(
        n16156) );
  AOI211_X1 U17171 ( .C1(n16188), .C2(n16158), .A(n16157), .B(n16156), .ZN(
        n16160) );
  OAI211_X1 U17172 ( .C1(n16161), .C2(n16191), .A(n16160), .B(n16159), .ZN(
        P2_U3228) );
  INV_X1 U17173 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n16174) );
  XNOR2_X1 U17174 ( .A(n16162), .B(n9664), .ZN(n16170) );
  OAI211_X1 U17175 ( .C1(n16165), .C2(P2_REG1_REG_18__SCAN_IN), .A(n16164), 
        .B(n16163), .ZN(n16166) );
  OAI21_X1 U17176 ( .B1(n16168), .B2(n16167), .A(n16166), .ZN(n16169) );
  AOI21_X1 U17177 ( .B1(n16171), .B2(n16170), .A(n16169), .ZN(n16173) );
  OAI211_X1 U17178 ( .C1(n16174), .C2(n16191), .A(n16173), .B(n16172), .ZN(
        P2_U3232) );
  INV_X1 U17179 ( .A(n16175), .ZN(n16176) );
  AOI211_X1 U17180 ( .C1(n16179), .C2(n16178), .A(n16177), .B(n16176), .ZN(
        n16186) );
  INV_X1 U17181 ( .A(n16180), .ZN(n16181) );
  AOI211_X1 U17182 ( .C1(n16184), .C2(n16183), .A(n16182), .B(n16181), .ZN(
        n16185) );
  AOI211_X1 U17183 ( .C1(n16188), .C2(n16187), .A(n16186), .B(n16185), .ZN(
        n16190) );
  OAI211_X1 U17184 ( .C1(n16192), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        P2_U3224) );
  OAI21_X1 U17185 ( .B1(n16194), .B2(P1_REG1_REG_0__SCAN_IN), .A(n16193), .ZN(
        n16196) );
  XNOR2_X1 U17186 ( .A(n16196), .B(n16195), .ZN(n16200) );
  AOI22_X1 U17187 ( .A1(n16197), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n16198) );
  OAI21_X1 U17188 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(P1_U3243) );
  AOI21_X1 U17189 ( .B1(n16202), .B2(n16201), .A(n16254), .ZN(SUB_1596_U53) );
  NOR2_X1 U17190 ( .A1(n16204), .A2(n16203), .ZN(n16205) );
  XOR2_X1 U17191 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n16205), .Z(SUB_1596_U61) );
  XNOR2_X1 U17192 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n16206), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17193 ( .A(n16208), .B(n16207), .Z(SUB_1596_U59) );
  AOI21_X1 U17194 ( .B1(n16211), .B2(n16210), .A(n16209), .ZN(n16213) );
  XNOR2_X1 U17195 ( .A(n16213), .B(n16212), .ZN(SUB_1596_U58) );
  XNOR2_X1 U17196 ( .A(n16215), .B(n16214), .ZN(SUB_1596_U56) );
  XOR2_X1 U17197 ( .A(n16216), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  XOR2_X1 U17198 ( .A(n16217), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI21_X1 U17199 ( .B1(n16220), .B2(n16219), .A(n16218), .ZN(n16221) );
  XNOR2_X1 U17200 ( .A(n16221), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  AOI21_X1 U17201 ( .B1(n16224), .B2(n16223), .A(n16222), .ZN(n16226) );
  XNOR2_X1 U17202 ( .A(n16226), .B(n16225), .ZN(SUB_1596_U69) );
  AOI21_X1 U17203 ( .B1(n16229), .B2(n16228), .A(n16227), .ZN(n16231) );
  XNOR2_X1 U17204 ( .A(n16231), .B(n16230), .ZN(SUB_1596_U68) );
  AOI21_X1 U17205 ( .B1(n16234), .B2(n16233), .A(n16232), .ZN(n16235) );
  XOR2_X1 U17206 ( .A(n16235), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  NOR2_X1 U17207 ( .A1(n16237), .A2(n16236), .ZN(n16238) );
  XOR2_X1 U17208 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n16238), .Z(SUB_1596_U66)
         );
  NOR2_X1 U17209 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  XOR2_X1 U17210 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n16241), .Z(SUB_1596_U65)
         );
  XNOR2_X1 U17211 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n16242), .ZN(n16244) );
  XNOR2_X1 U17212 ( .A(n16244), .B(n16243), .ZN(SUB_1596_U63) );
  AOI21_X1 U17213 ( .B1(n16247), .B2(n16246), .A(n16245), .ZN(n16248) );
  XOR2_X1 U17214 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n16248), .Z(SUB_1596_U62)
         );
  NOR2_X1 U17215 ( .A1(n16250), .A2(n16249), .ZN(n16252) );
  XNOR2_X1 U17216 ( .A(n16252), .B(n16251), .ZN(SUB_1596_U57) );
  OAI21_X1 U17217 ( .B1(n16255), .B2(n16254), .A(n16253), .ZN(n16256) );
  XNOR2_X1 U17218 ( .A(n16256), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(SUB_1596_U5)
         );
  INV_X1 U17219 ( .A(n16257), .ZN(n16258) );
  NOR2_X1 U17220 ( .A1(n16258), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n16261) );
  NAND3_X1 U17221 ( .A1(n16285), .A2(n16280), .A3(n16259), .ZN(n16260) );
  OAI21_X1 U17222 ( .B1(n16262), .B2(n16261), .A(n16260), .ZN(n16267) );
  OAI22_X1 U17223 ( .A1(n16278), .A2(n16264), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16263), .ZN(n16265) );
  INV_X1 U17224 ( .A(n16265), .ZN(n16266) );
  OAI211_X1 U17225 ( .C1(n16292), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        P3_U3182) );
  AOI21_X1 U17226 ( .B1(n16271), .B2(n16270), .A(n16269), .ZN(n16286) );
  OAI211_X1 U17227 ( .C1(n16275), .C2(n16274), .A(n16273), .B(n16272), .ZN(
        n16284) );
  AOI21_X1 U17228 ( .B1(n16277), .B2(n16389), .A(n16276), .ZN(n16281) );
  OAI22_X1 U17229 ( .A1(n16281), .A2(n16280), .B1(n16279), .B2(n16278), .ZN(
        n16282) );
  INV_X1 U17230 ( .A(n16282), .ZN(n16283) );
  OAI211_X1 U17231 ( .C1(n16286), .C2(n16285), .A(n16284), .B(n16283), .ZN(
        n16287) );
  INV_X1 U17232 ( .A(n16287), .ZN(n16290) );
  INV_X1 U17233 ( .A(n16288), .ZN(n16289) );
  OAI211_X1 U17234 ( .C1(n16292), .C2(n16291), .A(n16290), .B(n16289), .ZN(
        P3_U3191) );
  INV_X1 U17235 ( .A(P2_RD_REG_SCAN_IN), .ZN(n16295) );
  OAI221_X1 U17236 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n16295), .C2(n16294), .A(n16293), .ZN(U29) );
  INV_X1 U17237 ( .A(n16296), .ZN(n16302) );
  OAI22_X1 U17238 ( .A1(n16300), .A2(n16299), .B1(n16298), .B2(n16297), .ZN(
        n16301) );
  NOR2_X1 U17239 ( .A1(n16302), .A2(n16301), .ZN(n16304) );
  AOI22_X1 U17240 ( .A1(n16413), .A2(n16304), .B1(n11075), .B2(n16412), .ZN(
        P2_U3499) );
  INV_X1 U17241 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n16303) );
  AOI22_X1 U17242 ( .A1(n14760), .A2(n16304), .B1(n16303), .B2(n16414), .ZN(
        P2_U3430) );
  OAI21_X1 U17243 ( .B1(n16307), .B2(n16306), .A(n16305), .ZN(n16320) );
  NOR2_X1 U17244 ( .A1(n13483), .A2(n16467), .ZN(n16316) );
  XNOR2_X1 U17245 ( .A(n8991), .B(n16308), .ZN(n16310) );
  NAND2_X1 U17246 ( .A1(n16310), .A2(n16309), .ZN(n16315) );
  AOI22_X1 U17247 ( .A1(n16313), .A2(n8598), .B1(n16312), .B2(n16311), .ZN(
        n16314) );
  NAND2_X1 U17248 ( .A1(n16315), .A2(n16314), .ZN(n16322) );
  AOI211_X1 U17249 ( .C1(n10820), .C2(n16320), .A(n16316), .B(n16322), .ZN(
        n16318) );
  AOI22_X1 U17250 ( .A1(n16473), .A2(n16318), .B1(n8568), .B2(n10822), .ZN(
        P3_U3460) );
  INV_X1 U17251 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16317) );
  AOI22_X1 U17252 ( .A1(n16476), .A2(n16318), .B1(n16317), .B2(n16483), .ZN(
        P3_U3393) );
  INV_X1 U17253 ( .A(n16319), .ZN(n16341) );
  NAND2_X1 U17254 ( .A1(n16320), .A2(n16377), .ZN(n16321) );
  OAI211_X1 U17255 ( .C1(n13483), .C2(n16341), .A(n16321), .B(n16386), .ZN(
        n16323) );
  OAI22_X1 U17256 ( .A1(n16323), .A2(n16322), .B1(P3_REG2_REG_1__SCAN_IN), 
        .B2(n16386), .ZN(n16324) );
  OAI21_X1 U17257 ( .B1(n16325), .B2(n16339), .A(n16324), .ZN(P3_U3232) );
  NAND3_X1 U17258 ( .A1(n16328), .A2(n16327), .A3(n16326), .ZN(n16329) );
  OAI21_X1 U17259 ( .B1(n16330), .B2(n16437), .A(n16329), .ZN(n16333) );
  INV_X1 U17260 ( .A(n16331), .ZN(n16332) );
  AOI211_X1 U17261 ( .C1(n16440), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16337) );
  AOI22_X1 U17262 ( .A1(n16446), .A2(n16337), .B1(n16335), .B2(n16444), .ZN(
        P1_U3529) );
  INV_X1 U17263 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n16336) );
  AOI22_X1 U17264 ( .A1(n16338), .A2(n16337), .B1(n16336), .B2(n16447), .ZN(
        P1_U3462) );
  OAI22_X1 U17265 ( .A1(n16342), .A2(n16341), .B1(n16340), .B2(n16339), .ZN(
        n16344) );
  AOI211_X1 U17266 ( .C1(n16346), .C2(n16345), .A(n16344), .B(n16343), .ZN(
        n16347) );
  AOI22_X1 U17267 ( .A1(n16348), .A2(n11657), .B1(n16347), .B2(n16390), .ZN(
        P3_U3231) );
  AOI21_X1 U17268 ( .B1(n16358), .B2(n16350), .A(n16349), .ZN(n16351) );
  OAI211_X1 U17269 ( .C1(n16354), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        n16355) );
  INV_X1 U17270 ( .A(n16355), .ZN(n16357) );
  AOI22_X1 U17271 ( .A1(n16446), .A2(n16357), .B1(n10365), .B2(n16444), .ZN(
        P1_U3535) );
  INV_X1 U17272 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U17273 ( .A1(n16338), .A2(n16357), .B1(n16356), .B2(n16447), .ZN(
        P1_U3480) );
  AND2_X1 U17274 ( .A1(n16359), .A2(n16358), .ZN(n16360) );
  OR2_X1 U17275 ( .A1(n16361), .A2(n16360), .ZN(n16362) );
  AOI21_X1 U17276 ( .B1(n16363), .B2(n16440), .A(n16362), .ZN(n16364) );
  AND2_X1 U17277 ( .A1(n16365), .A2(n16364), .ZN(n16368) );
  AOI22_X1 U17278 ( .A1(n16446), .A2(n16368), .B1(n16366), .B2(n16444), .ZN(
        P1_U3536) );
  INV_X1 U17279 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U17280 ( .A1(n16338), .A2(n16368), .B1(n16367), .B2(n16447), .ZN(
        P1_U3483) );
  OAI21_X1 U17281 ( .B1(n16370), .B2(n16407), .A(n16369), .ZN(n16372) );
  AOI211_X1 U17282 ( .C1(n16374), .C2(n16373), .A(n16372), .B(n16371), .ZN(
        n16376) );
  AOI22_X1 U17283 ( .A1(n16413), .A2(n16376), .B1(n11118), .B2(n16412), .ZN(
        P2_U3507) );
  INV_X1 U17284 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U17285 ( .A1(n14760), .A2(n16376), .B1(n16375), .B2(n16414), .ZN(
        P2_U3454) );
  INV_X1 U17286 ( .A(n16377), .ZN(n16380) );
  OAI21_X1 U17287 ( .B1(n16380), .B2(n16379), .A(n16378), .ZN(n16387) );
  INV_X1 U17288 ( .A(n16381), .ZN(n16383) );
  AOI222_X1 U17289 ( .A1(n16387), .A2(n16386), .B1(n16385), .B2(n16384), .C1(
        n16383), .C2(n16382), .ZN(n16388) );
  OAI21_X1 U17290 ( .B1(n16390), .B2(n16389), .A(n16388), .ZN(P3_U3224) );
  OAI22_X1 U17291 ( .A1(n16392), .A2(n16428), .B1(n16391), .B2(n16437), .ZN(
        n16393) );
  AOI21_X1 U17292 ( .B1(n16394), .B2(n16440), .A(n16393), .ZN(n16395) );
  AND2_X1 U17293 ( .A1(n16396), .A2(n16395), .ZN(n16398) );
  AOI22_X1 U17294 ( .A1(n16446), .A2(n16398), .B1(n10402), .B2(n16444), .ZN(
        P1_U3537) );
  INV_X1 U17295 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16397) );
  AOI22_X1 U17296 ( .A1(n16338), .A2(n16398), .B1(n16397), .B2(n16447), .ZN(
        P1_U3486) );
  OAI22_X1 U17297 ( .A1(n16400), .A2(n16468), .B1(n16467), .B2(n16399), .ZN(
        n16401) );
  NOR2_X1 U17298 ( .A1(n16402), .A2(n16401), .ZN(n16405) );
  AOI22_X1 U17299 ( .A1(n16473), .A2(n16405), .B1(n16403), .B2(n10822), .ZN(
        P3_U3469) );
  INV_X1 U17300 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16404) );
  AOI22_X1 U17301 ( .A1(n16476), .A2(n16405), .B1(n16404), .B2(n16483), .ZN(
        P3_U3420) );
  OAI21_X1 U17302 ( .B1(n16408), .B2(n16407), .A(n16406), .ZN(n16410) );
  AOI211_X1 U17303 ( .C1(n11199), .C2(n16411), .A(n16410), .B(n16409), .ZN(
        n16416) );
  AOI22_X1 U17304 ( .A1(n16413), .A2(n16416), .B1(n11234), .B2(n16412), .ZN(
        P2_U3509) );
  INV_X1 U17305 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U17306 ( .A1(n14760), .A2(n16416), .B1(n16415), .B2(n16414), .ZN(
        P2_U3460) );
  AOI22_X1 U17307 ( .A1(n16419), .A2(n10820), .B1(n16418), .B2(n16417), .ZN(
        n16420) );
  AND2_X1 U17308 ( .A1(n16421), .A2(n16420), .ZN(n16424) );
  AOI22_X1 U17309 ( .A1(n16473), .A2(n16424), .B1(n16422), .B2(n10822), .ZN(
        P3_U3470) );
  INV_X1 U17310 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16423) );
  AOI22_X1 U17311 ( .A1(n16476), .A2(n16424), .B1(n16423), .B2(n16483), .ZN(
        P3_U3423) );
  NOR2_X1 U17312 ( .A1(n16426), .A2(n16425), .ZN(n16432) );
  OAI22_X1 U17313 ( .A1(n16429), .A2(n16428), .B1(n16427), .B2(n16437), .ZN(
        n16431) );
  AOI211_X1 U17314 ( .C1(n16432), .C2(n12600), .A(n16431), .B(n16430), .ZN(
        n16435) );
  AOI22_X1 U17315 ( .A1(n16446), .A2(n16435), .B1(n16433), .B2(n16444), .ZN(
        P1_U3539) );
  INV_X1 U17316 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U17317 ( .A1(n16338), .A2(n16435), .B1(n16434), .B2(n16447), .ZN(
        P1_U3492) );
  OAI21_X1 U17318 ( .B1(n16438), .B2(n16437), .A(n16436), .ZN(n16439) );
  AOI21_X1 U17319 ( .B1(n16441), .B2(n16440), .A(n16439), .ZN(n16442) );
  AND2_X1 U17320 ( .A1(n16443), .A2(n16442), .ZN(n16449) );
  AOI22_X1 U17321 ( .A1(n16446), .A2(n16449), .B1(n16445), .B2(n16444), .ZN(
        P1_U3540) );
  INV_X1 U17322 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U17323 ( .A1(n16338), .A2(n16449), .B1(n16448), .B2(n16447), .ZN(
        P1_U3495) );
  INV_X1 U17324 ( .A(n16450), .ZN(n16454) );
  AOI22_X1 U17325 ( .A1(n16454), .A2(n16453), .B1(n16452), .B2(n16451), .ZN(
        n16465) );
  OAI22_X1 U17326 ( .A1(n16458), .A2(n16457), .B1(n16456), .B2(n16455), .ZN(
        n16461) );
  NOR2_X1 U17327 ( .A1(n16459), .A2(n14598), .ZN(n16460) );
  AOI211_X1 U17328 ( .C1(n16463), .C2(n16462), .A(n16461), .B(n16460), .ZN(
        n16464) );
  NAND2_X1 U17329 ( .A1(n16465), .A2(n16464), .ZN(P2_U3253) );
  OAI22_X1 U17330 ( .A1(n16469), .A2(n16468), .B1(n16467), .B2(n16466), .ZN(
        n16470) );
  NOR2_X1 U17331 ( .A1(n16471), .A2(n16470), .ZN(n16475) );
  AOI22_X1 U17332 ( .A1(n16473), .A2(n16475), .B1(n16472), .B2(n10822), .ZN(
        P3_U3472) );
  INV_X1 U17333 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16474) );
  AOI22_X1 U17334 ( .A1(n16476), .A2(n16475), .B1(n16474), .B2(n16483), .ZN(
        P3_U3429) );
  AOI22_X1 U17335 ( .A1(n16479), .A2(n16477), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16483), .ZN(n16478) );
  OAI21_X1 U17336 ( .B1(n16483), .B2(n16482), .A(n16478), .ZN(P3_U3457) );
  AOI22_X1 U17337 ( .A1(n16480), .A2(n16479), .B1(P3_REG0_REG_31__SCAN_IN), 
        .B2(n16483), .ZN(n16481) );
  OAI21_X1 U17338 ( .B1(n16483), .B2(n16482), .A(n16481), .ZN(P3_U3458) );
  AOI21_X1 U17339 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16484) );
  OAI21_X1 U17340 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16484), 
        .ZN(U28) );
  XNOR2_X1 U7810 ( .A(n9343), .B(n9342), .ZN(n9910) );
  NAND2_X1 U9850 ( .A1(n9910), .A2(n9904), .ZN(n11067) );
  OR2_X1 U11214 ( .A1(n9401), .A2(n10847), .ZN(n9377) );
  INV_X1 U12133 ( .A(n10322), .ZN(n10560) );
  INV_X1 U7540 ( .A(n11694), .ZN(n14935) );
  BUF_X2 U7545 ( .A(n15461), .Z(n7438) );
  NAND2_X1 U7553 ( .A1(n11067), .A2(n10838), .ZN(n9401) );
  CLKBUF_X2 U7564 ( .A(n9401), .Z(n10137) );
  CLKBUF_X1 U7567 ( .A(n9388), .Z(n9685) );
  CLKBUF_X2 U7572 ( .A(n12699), .Z(n14817) );
  CLKBUF_X1 U7678 ( .A(n10331), .Z(n7433) );
  CLKBUF_X1 U7687 ( .A(n9391), .Z(n10118) );
  XOR2_X1 U9546 ( .A(n14686), .B(n14306), .Z(n16491) );
  AND2_X1 U9851 ( .A1(n15609), .A2(n15608), .ZN(n16492) );
endmodule

