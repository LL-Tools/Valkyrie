

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4864, n4866, n4867, n4868, n4869, n4870, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659;

  AOI21_X1 U4928 ( .B1(n8541), .B2(n5286), .A(n4891), .ZN(n9392) );
  NAND4_X1 U4929 ( .A1(n6301), .A2(n6300), .A3(n6299), .A4(n6298), .ZN(n8662)
         );
  NAND2_X2 U4931 ( .A1(n6253), .A2(n6251), .ZN(n6309) );
  INV_X4 U4932 ( .A(n6220), .ZN(n7284) );
  INV_X1 U4933 ( .A(n6302), .ZN(n6715) );
  INV_X1 U4934 ( .A(n6279), .ZN(n6640) );
  INV_X1 U4935 ( .A(n5907), .ZN(n5713) );
  INV_X1 U4936 ( .A(n6112), .ZN(n6141) );
  INV_X1 U4937 ( .A(n5548), .ZN(n5915) );
  BUF_X1 U4938 ( .A(n6309), .Z(n4870) );
  INV_X1 U4940 ( .A(n7613), .ZN(n6847) );
  INV_X2 U4941 ( .A(n5907), .ZN(n6000) );
  NAND2_X1 U4942 ( .A1(n8545), .A2(n8547), .ZN(n8541) );
  AND2_X1 U4944 ( .A1(n5153), .A2(n5151), .ZN(n4933) );
  XNOR2_X1 U4945 ( .A(n5439), .B(n5438), .ZN(n8436) );
  INV_X1 U4946 ( .A(n5681), .ZN(n4866) );
  OR2_X2 U4947 ( .A1(n5770), .A2(SI_12_), .ZN(n5796) );
  OAI21_X2 U4948 ( .B1(n9972), .B2(n4906), .A(n5193), .ZN(n9936) );
  NAND2_X2 U4949 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  NAND4_X2 U4950 ( .A1(n6331), .A2(n6330), .A3(n6329), .A4(n6328), .ZN(n8663)
         );
  OAI21_X2 U4951 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8839), .A(n8835), .ZN(
        n8837) );
  NAND2_X2 U4952 ( .A1(n5442), .A2(n6146), .ZN(n7069) );
  NAND2_X1 U4953 ( .A1(n6751), .A2(n6750), .ZN(n4864) );
  NAND2_X1 U4954 ( .A1(n6751), .A2(n6750), .ZN(n10613) );
  NAND2_X2 U4955 ( .A1(n6324), .A2(n6323), .ZN(n7515) );
  OAI21_X2 U4956 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8851), .A(n8850), .ZN(
        n8873) );
  OAI21_X2 U4957 ( .B1(n8984), .B2(n8986), .A(n6803), .ZN(n8968) );
  AOI21_X2 U4958 ( .B1(n8999), .B2(n5081), .A(n6802), .ZN(n8984) );
  OAI211_X4 U4959 ( .C1(n7297), .C2(n6288), .A(n6278), .B(n5231), .ZN(n7613)
         );
  AOI21_X2 U4960 ( .B1(n8884), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8883), .ZN(
        n8885) );
  MUX2_X1 U4961 ( .A(n9615), .B(n9614), .S(n9900), .Z(n9663) );
  XNOR2_X1 U4962 ( .A(n6637), .B(n6635), .ZN(n8652) );
  AND2_X1 U4963 ( .A1(n8542), .A2(n5287), .ZN(n5286) );
  AND2_X1 U4964 ( .A1(n6974), .A2(n6973), .ZN(n6831) );
  INV_X2 U4965 ( .A(n8370), .ZN(P2_U3966) );
  AND2_X1 U4966 ( .A1(n6901), .A2(n6900), .ZN(n8086) );
  OR2_X1 U4967 ( .A1(n7669), .A2(n6790), .ZN(n5262) );
  INV_X1 U4968 ( .A(n10490), .ZN(n7851) );
  NAND2_X1 U4969 ( .A1(n6922), .A2(n6921), .ZN(n6818) );
  OAI21_X1 U4970 ( .B1(n5158), .B2(n7720), .A(n7746), .ZN(n5160) );
  INV_X2 U4971 ( .A(n8662), .ZN(n6779) );
  NAND2_X1 U4972 ( .A1(n7713), .A2(n4879), .ZN(n7746) );
  INV_X1 U4973 ( .A(n7712), .ZN(n7736) );
  INV_X1 U4974 ( .A(n10418), .ZN(n7760) );
  INV_X1 U4975 ( .A(n7773), .ZN(n7846) );
  INV_X2 U4976 ( .A(n5973), .ZN(n5566) );
  INV_X4 U4977 ( .A(n6295), .ZN(n6561) );
  CLKBUF_X2 U4978 ( .A(n5681), .Z(n4875) );
  AND2_X1 U4979 ( .A1(n10192), .A2(n8582), .ZN(n5568) );
  INV_X2 U4980 ( .A(n5992), .ZN(n4867) );
  OAI21_X1 U4981 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5466) );
  NOR2_X1 U4982 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6201) );
  AND2_X1 U4983 ( .A1(n5130), .A2(n5133), .ZN(n4983) );
  AOI21_X1 U4984 ( .B1(n5089), .B2(n10453), .A(n6846), .ZN(n8947) );
  AOI22_X1 U4985 ( .A1(n7033), .A2(n7032), .B1(n7031), .B2(n7030), .ZN(n7035)
         );
  NOR2_X1 U4986 ( .A1(n9797), .A2(n9796), .ZN(n9798) );
  OR2_X1 U4987 ( .A1(n9794), .A2(n9793), .ZN(n10069) );
  NAND2_X1 U4988 ( .A1(n9300), .A2(n9301), .ZN(n9299) );
  OAI21_X1 U4989 ( .B1(n4963), .B2(n4962), .A(n4961), .ZN(n9478) );
  CLKBUF_X1 U4990 ( .A(n9850), .Z(n10096) );
  NAND2_X1 U4991 ( .A1(n9029), .A2(n6990), .ZN(n9013) );
  NAND2_X1 U4992 ( .A1(n9054), .A2(n9055), .ZN(n9053) );
  AOI22_X1 U4993 ( .A1(n9046), .A2(n7046), .B1(n9052), .B2(n9069), .ZN(n9042)
         );
  OAI211_X1 U4994 ( .C1(n9958), .C2(n5184), .A(n4982), .B(n9935), .ZN(n9926)
         );
  AOI21_X1 U4995 ( .B1(n9456), .B2(n4967), .A(n4966), .ZN(n9460) );
  NAND2_X1 U4996 ( .A1(n5253), .A2(n5252), .ZN(n9117) );
  NAND2_X1 U4997 ( .A1(n8595), .A2(n4917), .ZN(n10015) );
  AOI21_X1 U4998 ( .B1(n5006), .B2(n5387), .A(n5005), .ZN(n5004) );
  NAND2_X1 U4999 ( .A1(n8396), .A2(n9525), .ZN(n8595) );
  AND2_X1 U5000 ( .A1(n9598), .A2(n9543), .ZN(n9855) );
  NOR2_X1 U5001 ( .A1(n8673), .A2(n5007), .ZN(n5006) );
  NAND2_X1 U5002 ( .A1(n6059), .A2(n6058), .ZN(n10084) );
  XNOR2_X1 U5003 ( .A(n6120), .B(n6119), .ZN(n10200) );
  NAND2_X1 U5004 ( .A1(n6038), .A2(n6037), .ZN(n10090) );
  NAND2_X1 U5005 ( .A1(n6102), .A2(n6101), .ZN(n6120) );
  NAND2_X1 U5006 ( .A1(n8120), .A2(n8119), .ZN(n8118) );
  OR2_X1 U5007 ( .A1(n6796), .A2(n8718), .ZN(n6974) );
  NAND2_X1 U5008 ( .A1(n6591), .A2(n6590), .ZN(n9216) );
  NAND2_X1 U5009 ( .A1(n8351), .A2(n5208), .ZN(n8373) );
  NAND2_X1 U5010 ( .A1(n5178), .A2(n9522), .ZN(n8374) );
  NAND2_X1 U5011 ( .A1(n8070), .A2(n9520), .ZN(n8351) );
  NAND2_X1 U5012 ( .A1(n5896), .A2(n5895), .ZN(n10123) );
  OAI21_X1 U5013 ( .B1(n8042), .B2(n5176), .A(n5174), .ZN(n8376) );
  NAND2_X1 U5014 ( .A1(n6531), .A2(n6530), .ZN(n9237) );
  OAI21_X1 U5015 ( .B1(n5940), .B2(n5932), .A(n5913), .ZN(n8531) );
  AND2_X1 U5016 ( .A1(n7688), .A2(n6793), .ZN(n7817) );
  NAND2_X1 U5017 ( .A1(n5876), .A2(n5875), .ZN(n10128) );
  OAI211_X1 U5018 ( .C1(n9430), .C2(n10046), .A(n9517), .B(n9429), .ZN(n9433)
         );
  OR2_X1 U5019 ( .A1(n10135), .A2(n10016), .ZN(n9576) );
  NOR2_X1 U5020 ( .A1(n8086), .A2(n5345), .ZN(n5344) );
  AOI21_X1 U5021 ( .B1(n8820), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8819), .ZN(
        n8823) );
  AOI21_X1 U5022 ( .B1(n5192), .B2(n5191), .A(n5188), .ZN(n10047) );
  NAND2_X1 U5023 ( .A1(n6494), .A2(n6493), .ZN(n8093) );
  NAND2_X1 U5024 ( .A1(n6475), .A2(n6474), .ZN(n8128) );
  AND2_X1 U5025 ( .A1(n5841), .A2(n5861), .ZN(n5310) );
  NAND2_X1 U5026 ( .A1(n5777), .A2(n5776), .ZN(n8409) );
  NAND2_X1 U5027 ( .A1(n5754), .A2(n5753), .ZN(n10159) );
  NAND2_X1 U5028 ( .A1(n5658), .A2(n5657), .ZN(n10560) );
  OAI21_X2 U5029 ( .B1(n6768), .B2(n6758), .A(n10470), .ZN(n6759) );
  INV_X1 U5030 ( .A(n6781), .ZN(n10402) );
  NAND2_X1 U5031 ( .A1(n5628), .A2(n5627), .ZN(n5633) );
  NAND2_X1 U5032 ( .A1(n7736), .A2(n7711), .ZN(n9622) );
  AND3_X1 U5033 ( .A1(n5398), .A2(n6281), .A3(n6282), .ZN(n4880) );
  AND2_X1 U5034 ( .A1(n6308), .A2(n6307), .ZN(n6781) );
  NAND2_X1 U5035 ( .A1(n6550), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6300) );
  XNOR2_X1 U5036 ( .A(n6280), .B(n6847), .ZN(n6284) );
  BUF_X1 U5037 ( .A(n7711), .Z(n9680) );
  AND2_X1 U5038 ( .A1(n5525), .A2(n5524), .ZN(n10418) );
  AND2_X2 U5039 ( .A1(n7313), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X2 U5040 ( .A1(n7428), .A2(n5478), .ZN(n10519) );
  AND2_X2 U5041 ( .A1(n5539), .A2(n5481), .ZN(n6112) );
  NAND2_X1 U5042 ( .A1(n7725), .A2(n7724), .ZN(n10511) );
  INV_X1 U5043 ( .A(n4866), .ZN(n4876) );
  OR2_X1 U5044 ( .A1(n5536), .A2(n7298), .ZN(n5495) );
  INV_X1 U5045 ( .A(n9273), .ZN(n6251) );
  NAND2_X4 U5046 ( .A1(n6252), .A2(n9273), .ZN(n6295) );
  BUF_X2 U5047 ( .A(n5568), .Z(n4874) );
  BUF_X2 U5048 ( .A(n5568), .Z(n4873) );
  BUF_X1 U5049 ( .A(n6249), .Z(n6253) );
  INV_X1 U5050 ( .A(n6249), .ZN(n6252) );
  NAND2_X1 U5051 ( .A1(n6248), .A2(n9267), .ZN(n9273) );
  NAND2_X1 U5052 ( .A1(n5466), .A2(n5465), .ZN(n10192) );
  NAND2_X1 U5053 ( .A1(n5440), .A2(n5436), .ZN(n8458) );
  MUX2_X1 U5054 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6247), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6248) );
  NAND2_X1 U5055 ( .A1(n6219), .A2(n5264), .ZN(n6841) );
  XNOR2_X1 U5056 ( .A(n6245), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U5057 ( .A1(n9267), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6245) );
  MUX2_X1 U5058 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6217), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6219) );
  XNOR2_X1 U5059 ( .A(n6232), .B(n6205), .ZN(n6750) );
  AOI21_X1 U5060 ( .B1(n10641), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10637), .ZN(
        n10626) );
  NAND2_X1 U5061 ( .A1(n6218), .A2(n5100), .ZN(n9267) );
  NAND2_X1 U5062 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  INV_X2 U5063 ( .A(n9265), .ZN(n8529) );
  XNOR2_X1 U5064 ( .A(n6734), .B(n6733), .ZN(n6259) );
  NAND2_X2 U5065 ( .A1(n7285), .A2(P2_U3152), .ZN(n9280) );
  OAI21_X1 U5066 ( .B1(n6238), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U5067 ( .A1(n5411), .A2(n5410), .ZN(n5211) );
  NOR2_X1 U5068 ( .A1(n6223), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U5069 ( .A1(n4901), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5070 ( .A1(n5461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  MUX2_X1 U5071 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6274), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6277) );
  AND4_X1 U5072 ( .A1(n6229), .A2(n6228), .A3(n6508), .A4(n5012), .ZN(n6208)
         );
  INV_X1 U5073 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5434) );
  NOR2_X1 U5074 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5445) );
  INV_X1 U5075 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6747) );
  INV_X1 U5076 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6228) );
  INV_X1 U5077 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6222) );
  NOR2_X1 U5078 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5406) );
  NOR2_X1 U5079 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5407) );
  INV_X1 U5080 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6508) );
  INV_X1 U5081 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6490) );
  NOR2_X1 U5082 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6199) );
  NOR2_X1 U5083 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6200) );
  INV_X1 U5084 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5869) );
  INV_X1 U5085 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5404) );
  INV_X1 U5086 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5872) );
  NOR2_X1 U5087 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5403) );
  INV_X4 U5088 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5089 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5558) );
  NOR2_X1 U5090 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5430) );
  NOR2_X1 U5091 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n6203) );
  NAND2_X4 U5092 ( .A1(n6242), .A2(n5391), .ZN(n6325) );
  CLKBUF_X2 U5093 ( .A(n6815), .Z(n4868) );
  NAND2_X1 U5094 ( .A1(n4880), .A2(n6283), .ZN(n6815) );
  NAND2_X2 U5095 ( .A1(n8744), .A2(n6623), .ZN(n6637) );
  INV_X4 U5096 ( .A(n5973), .ZN(n4869) );
  BUF_X4 U5097 ( .A(n10289), .Z(n4872) );
  NAND2_X1 U5098 ( .A1(n7315), .A2(n6180), .ZN(n10289) );
  INV_X1 U5099 ( .A(n4866), .ZN(n4877) );
  AND2_X1 U5100 ( .A1(n10192), .A2(n5468), .ZN(n5681) );
  NAND2_X1 U5101 ( .A1(n4872), .A2(n6220), .ZN(n4878) );
  CLKBUF_X2 U5102 ( .A(n7712), .Z(n4879) );
  OAI211_X1 U5103 ( .C1(n4872), .C2(n7368), .A(n5495), .B(n5494), .ZN(n7712)
         );
  OAI21_X1 U5104 ( .B1(n7002), .B2(n7021), .A(n5104), .ZN(n5103) );
  INV_X1 U5105 ( .A(n5105), .ZN(n5104) );
  OR2_X1 U5106 ( .A1(n8932), .A2(n8057), .ZN(n5360) );
  AND2_X1 U5107 ( .A1(n6887), .A2(n7025), .ZN(n7051) );
  OR2_X1 U5108 ( .A1(n9197), .A2(n9033), .ZN(n6995) );
  OR2_X1 U5109 ( .A1(n9222), .A2(n9067), .ZN(n6980) );
  INV_X1 U5110 ( .A(n6297), .ZN(n6871) );
  OR2_X1 U5111 ( .A1(n9210), .A2(n9069), .ZN(n6988) );
  INV_X1 U5112 ( .A(n5536), .ZN(n9493) );
  OAI211_X1 U5113 ( .C1(n5889), .C2(n4946), .A(n4974), .B(n4973), .ZN(n7970)
         );
  OAI22_X1 U5114 ( .A1(n4975), .A2(n4945), .B1(n4978), .B2(n5936), .ZN(n4974)
         );
  NAND2_X1 U5115 ( .A1(n5889), .A2(n4944), .ZN(n4973) );
  NAND2_X1 U5116 ( .A1(n6928), .A2(n5099), .ZN(n5098) );
  OR2_X1 U5117 ( .A1(n6987), .A2(n9041), .ZN(n6998) );
  AOI21_X1 U5118 ( .B1(n5091), .B2(n7044), .A(n5090), .ZN(n6986) );
  INV_X1 U5119 ( .A(n6985), .ZN(n5090) );
  INV_X1 U5120 ( .A(n6056), .ZN(n5316) );
  OR2_X1 U5121 ( .A1(n9181), .A2(n8765), .ZN(n7013) );
  AND2_X1 U5122 ( .A1(n9110), .A2(n5076), .ZN(n5075) );
  NAND2_X1 U5123 ( .A1(n9116), .A2(n6974), .ZN(n5076) );
  OR2_X1 U5124 ( .A1(n9122), .A2(n5077), .ZN(n5074) );
  INV_X1 U5125 ( .A(n6974), .ZN(n5077) );
  OR2_X1 U5126 ( .A1(n9237), .A2(n8345), .ZN(n6896) );
  AND2_X1 U5127 ( .A1(n6778), .A2(n6777), .ZN(n9151) );
  AND2_X1 U5128 ( .A1(n10343), .A2(n6746), .ZN(n8148) );
  AND2_X1 U5129 ( .A1(n10342), .A2(n10241), .ZN(n6746) );
  OR2_X1 U5131 ( .A1(n10060), .A2(n9508), .ZN(n9651) );
  NAND2_X1 U5132 ( .A1(n5121), .A2(n5120), .ZN(n5119) );
  INV_X1 U5133 ( .A(n10066), .ZN(n5121) );
  NAND2_X1 U5134 ( .A1(n8613), .A2(n8615), .ZN(n5207) );
  INV_X1 U5135 ( .A(n8603), .ZN(n5195) );
  OR2_X1 U5136 ( .A1(n10139), .A2(n9996), .ZN(n9575) );
  INV_X1 U5137 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5138 ( .A1(n5302), .A2(n5796), .ZN(n5305) );
  AND2_X1 U5139 ( .A1(n5795), .A2(n4943), .ZN(n5302) );
  AND2_X1 U5140 ( .A1(n5791), .A2(n5792), .ZN(n5795) );
  OAI21_X1 U5141 ( .B1(n5324), .B2(n5633), .A(n4970), .ZN(n5721) );
  AOI21_X1 U5142 ( .B1(n5323), .B2(n4889), .A(n4926), .ZN(n4970) );
  OAI21_X1 U5143 ( .B1(n7284), .B2(n4965), .A(n4964), .ZN(n5552) );
  NAND2_X1 U5144 ( .A1(n7284), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4964) );
  OAI21_X1 U5145 ( .B1(n9176), .B2(n5380), .A(n5375), .ZN(n5374) );
  NAND2_X1 U5146 ( .A1(n6760), .A2(n5380), .ZN(n5375) );
  NAND2_X1 U5147 ( .A1(n4988), .A2(n4986), .ZN(n8017) );
  OAI21_X1 U5148 ( .B1(n4992), .B2(n4990), .A(n8019), .ZN(n4987) );
  AOI21_X1 U5149 ( .B1(n4928), .B2(n5360), .A(n5357), .ZN(n5356) );
  XNOR2_X1 U5150 ( .A(n7035), .B(n5321), .ZN(n5320) );
  INV_X1 U5151 ( .A(n7034), .ZN(n5321) );
  NAND2_X1 U5152 ( .A1(n8951), .A2(n6837), .ZN(n6861) );
  AND2_X1 U5153 ( .A1(n5239), .A2(n5243), .ZN(n5238) );
  NAND2_X1 U5154 ( .A1(n8972), .A2(n8765), .ZN(n5243) );
  NAND2_X1 U5155 ( .A1(n8973), .A2(n5240), .ZN(n5239) );
  INV_X1 U5156 ( .A(n6803), .ZN(n5240) );
  AND2_X1 U5157 ( .A1(n6708), .A2(n6707), .ZN(n8962) );
  OAI21_X1 U5158 ( .B1(n9017), .B2(n5081), .A(n5078), .ZN(n8985) );
  AND2_X1 U5159 ( .A1(n5082), .A2(n5079), .ZN(n5078) );
  AND2_X1 U5160 ( .A1(n7004), .A2(n8986), .ZN(n5082) );
  NAND2_X1 U5161 ( .A1(n9001), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U5162 ( .A1(n9017), .A2(n6995), .ZN(n9002) );
  NAND2_X1 U5163 ( .A1(n6995), .A2(n6999), .ZN(n9020) );
  NAND2_X1 U5164 ( .A1(n9053), .A2(n5346), .ZN(n9029) );
  AND2_X1 U5165 ( .A1(n6833), .A2(n6988), .ZN(n5346) );
  NAND2_X1 U5166 ( .A1(n5246), .A2(n5244), .ZN(n9046) );
  AOI21_X1 U5167 ( .B1(n4882), .B2(n9091), .A(n5245), .ZN(n5244) );
  INV_X1 U5168 ( .A(n6799), .ZN(n5245) );
  OR2_X1 U5169 ( .A1(n6797), .A2(n8736), .ZN(n6894) );
  AOI21_X1 U5170 ( .B1(n9117), .B2(n9116), .A(n5399), .ZN(n9102) );
  NAND2_X1 U5171 ( .A1(n6965), .A2(n5341), .ZN(n5340) );
  NOR2_X1 U5172 ( .A1(n5344), .A2(n6901), .ZN(n5341) );
  AOI21_X1 U5173 ( .B1(n5069), .B2(n6947), .A(n5067), .ZN(n5066) );
  OR2_X1 U5174 ( .A1(n10598), .A2(n8460), .ZN(n5397) );
  OR2_X1 U5175 ( .A1(n8156), .A2(n9275), .ZN(n9066) );
  INV_X1 U5176 ( .A(n10453), .ZN(n9064) );
  INV_X1 U5177 ( .A(n10448), .ZN(n9068) );
  NAND2_X1 U5178 ( .A1(n4925), .A2(n6922), .ZN(n5086) );
  AND2_X2 U5179 ( .A1(n6915), .A2(n5233), .ZN(n9159) );
  NAND2_X1 U5180 ( .A1(n6575), .A2(n6574), .ZN(n9222) );
  OR2_X1 U5181 ( .A1(n6288), .A2(n6573), .ZN(n6574) );
  AND2_X1 U5182 ( .A1(n7892), .A2(n10596), .ZN(n9245) );
  INV_X1 U5183 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5263) );
  AOI21_X1 U5184 ( .B1(n4907), .B2(n6074), .A(n5057), .ZN(n5056) );
  INV_X1 U5185 ( .A(n9400), .ZN(n5057) );
  XNOR2_X1 U5186 ( .A(n5464), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6180) );
  INV_X1 U5187 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U5188 ( .A1(n5186), .A2(n9586), .ZN(n4982) );
  NAND2_X1 U5189 ( .A1(n9489), .A2(n9488), .ZN(n10056) );
  NAND2_X1 U5190 ( .A1(n5986), .A2(n5985), .ZN(n10102) );
  NOR2_X1 U5191 ( .A1(n8458), .A2(n8436), .ZN(n5442) );
  OAI21_X1 U5192 ( .B1(n5963), .B2(n5329), .A(n5328), .ZN(n6027) );
  AOI21_X1 U5193 ( .B1(n5330), .B2(n5964), .A(n4956), .ZN(n5328) );
  INV_X1 U5194 ( .A(n5330), .ZN(n5329) );
  AND2_X1 U5195 ( .A1(n5475), .A2(n5456), .ZN(n7723) );
  OR2_X1 U5196 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  XNOR2_X1 U5197 ( .A(n5457), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9659) );
  NAND2_X2 U5198 ( .A1(n5865), .A2(n5864), .ZN(n5889) );
  NAND2_X1 U5199 ( .A1(n5146), .A2(n5841), .ZN(n5842) );
  AND2_X1 U5200 ( .A1(n5308), .A2(SI_15_), .ZN(n5146) );
  AND2_X1 U5201 ( .A1(n6650), .A2(n6649), .ZN(n9033) );
  AND2_X1 U5202 ( .A1(n6616), .A2(n6615), .ZN(n9069) );
  NAND2_X1 U5203 ( .A1(n6909), .A2(n5095), .ZN(n6913) );
  INV_X1 U5204 ( .A(n5233), .ZN(n6917) );
  AND2_X1 U5205 ( .A1(n6948), .A2(n6949), .ZN(n5111) );
  MUX2_X1 U5206 ( .A(n9426), .B(n9425), .S(n9485), .Z(n9430) );
  NAND2_X1 U5207 ( .A1(n5092), .A2(n6982), .ZN(n5091) );
  NAND2_X1 U5208 ( .A1(n6993), .A2(n9033), .ZN(n6991) );
  OAI21_X1 U5209 ( .B1(n7001), .B2(n7028), .A(n9001), .ZN(n5105) );
  NOR2_X1 U5210 ( .A1(n9474), .A2(n9475), .ZN(n4963) );
  OAI21_X1 U5211 ( .B1(n5102), .B2(n8973), .A(n5101), .ZN(n7018) );
  AND2_X1 U5212 ( .A1(n8952), .A2(n7015), .ZN(n5101) );
  AOI21_X1 U5213 ( .B1(n5103), .B2(n7012), .A(n7011), .ZN(n5102) );
  NOR2_X1 U5214 ( .A1(n5279), .A2(n7642), .ZN(n5275) );
  INV_X1 U5215 ( .A(n7907), .ZN(n5279) );
  NAND2_X1 U5216 ( .A1(n7907), .A2(n5278), .ZN(n5277) );
  INV_X1 U5217 ( .A(n5626), .ZN(n5278) );
  OR2_X1 U5218 ( .A1(n10063), .A2(n8592), .ZN(n9483) );
  NAND2_X1 U5219 ( .A1(n5888), .A2(n5887), .ZN(n5142) );
  NAND2_X1 U5220 ( .A1(n5797), .A2(SI_14_), .ZN(n5819) );
  INV_X1 U5221 ( .A(SI_9_), .ZN(n7221) );
  NOR2_X1 U5222 ( .A1(n5358), .A2(n5355), .ZN(n5354) );
  INV_X1 U5223 ( .A(n7023), .ZN(n5355) );
  NAND2_X1 U5224 ( .A1(n8952), .A2(n5333), .ZN(n5332) );
  NOR2_X1 U5225 ( .A1(n7048), .A2(n8973), .ZN(n5333) );
  OR2_X1 U5226 ( .A1(n8941), .A2(n8368), .ZN(n7022) );
  NOR2_X1 U5227 ( .A1(n9187), .A2(n9181), .ZN(n5218) );
  OR2_X1 U5228 ( .A1(n6394), .A2(n6393), .ZN(n6411) );
  NAND2_X1 U5229 ( .A1(n7662), .A2(n5227), .ZN(n5226) );
  OR2_X1 U5230 ( .A1(n7792), .A2(n5226), .ZN(n5225) );
  AND2_X1 U5231 ( .A1(n7058), .A2(n5392), .ZN(n8150) );
  NOR2_X1 U5232 ( .A1(n9154), .A2(n10402), .ZN(n10443) );
  INV_X1 U5233 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6212) );
  INV_X1 U5234 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6206) );
  INV_X1 U5235 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6230) );
  AND4_X1 U5236 ( .A1(n5094), .A2(n5013), .A3(n6338), .A4(n5011), .ZN(n6235)
         );
  AND2_X1 U5237 ( .A1(n5012), .A2(n6228), .ZN(n5011) );
  OR2_X1 U5238 ( .A1(n6340), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6371) );
  OR2_X1 U5239 ( .A1(n6025), .A2(n5045), .ZN(n5044) );
  INV_X1 U5240 ( .A(n9303), .ZN(n5045) );
  INV_X1 U5241 ( .A(n6004), .ZN(n5043) );
  NOR2_X1 U5242 ( .A1(n5047), .A2(n9303), .ZN(n5046) );
  NOR2_X1 U5243 ( .A1(n5058), .A2(n5395), .ZN(n5063) );
  INV_X1 U5244 ( .A(n5266), .ZN(n5058) );
  INV_X1 U5245 ( .A(n8616), .ZN(n5205) );
  NAND2_X1 U5246 ( .A1(n5167), .A2(n9542), .ZN(n5166) );
  INV_X1 U5247 ( .A(n9868), .ZN(n5167) );
  INV_X1 U5248 ( .A(n9543), .ZN(n5164) );
  AND2_X1 U5249 ( .A1(n9954), .A2(n8602), .ZN(n5196) );
  NOR2_X1 U5250 ( .A1(n9991), .A2(n8596), .ZN(n5170) );
  INV_X1 U5251 ( .A(n9576), .ZN(n5172) );
  OR2_X1 U5252 ( .A1(n10146), .A2(n10017), .ZN(n9570) );
  OR2_X1 U5253 ( .A1(n8409), .A2(n9292), .ZN(n9569) );
  OR2_X1 U5254 ( .A1(n5679), .A2(n7394), .ZN(n5707) );
  NAND2_X1 U5255 ( .A1(n10565), .A2(n7915), .ZN(n8035) );
  INV_X1 U5256 ( .A(n7854), .ZN(n5190) );
  INV_X1 U5257 ( .A(n10509), .ZN(n7853) );
  XNOR2_X1 U5258 ( .A(n9678), .B(n10434), .ZN(n10413) );
  INV_X1 U5259 ( .A(n5182), .ZN(n5181) );
  OR2_X1 U5260 ( .A1(n10123), .A2(n9975), .ZN(n9583) );
  NAND2_X1 U5261 ( .A1(n5480), .A2(n10494), .ZN(n9485) );
  NAND2_X1 U5262 ( .A1(n5311), .A2(n5312), .ZN(n6098) );
  AND2_X1 U5263 ( .A1(n5313), .A2(n6077), .ZN(n5312) );
  NAND2_X1 U5264 ( .A1(n5453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5455) );
  INV_X1 U5265 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5452) );
  INV_X1 U5266 ( .A(n5771), .ZN(n5150) );
  INV_X1 U5267 ( .A(SI_10_), .ZN(n5723) );
  NAND2_X1 U5268 ( .A1(n5404), .A2(n5285), .ZN(n5284) );
  INV_X1 U5269 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5285) );
  NOR2_X1 U5270 ( .A1(n5671), .A2(n5327), .ZN(n5326) );
  INV_X1 U5271 ( .A(SI_7_), .ZN(n7220) );
  INV_X1 U5272 ( .A(SI_6_), .ZN(n7227) );
  INV_X1 U5273 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5301) );
  OR2_X1 U5274 ( .A1(n8533), .A2(n5386), .ZN(n5385) );
  INV_X1 U5275 ( .A(n8532), .ZN(n5386) );
  NAND2_X1 U5276 ( .A1(n5010), .A2(n5009), .ZN(n5008) );
  AOI22_X1 U5277 ( .A1(n6760), .A2(n8759), .B1(n6761), .B2(n8759), .ZN(n5379)
         );
  NAND2_X1 U5278 ( .A1(n5374), .A2(n5002), .ZN(n5000) );
  INV_X1 U5279 ( .A(n6459), .ZN(n4993) );
  NAND2_X1 U5280 ( .A1(n6431), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6464) );
  AND2_X1 U5281 ( .A1(n6443), .A2(n6422), .ZN(n5390) );
  OR2_X1 U5282 ( .A1(n8531), .A2(n6640), .ZN(n6545) );
  OR2_X1 U5283 ( .A1(n6311), .A2(n7627), .ZN(n6281) );
  OR2_X1 U5284 ( .A1(n6297), .A2(n10643), .ZN(n6270) );
  OR2_X1 U5285 ( .A1(n6309), .A2(n7494), .ZN(n6269) );
  NOR4_X1 U5286 ( .A1(n7281), .A2(n7280), .A3(n7279), .A4(n7278), .ZN(n7282)
         );
  NAND2_X1 U5287 ( .A1(n7023), .A2(n7022), .ZN(n7049) );
  AND2_X1 U5288 ( .A1(n8990), .A2(n5214), .ZN(n8935) );
  NOR2_X1 U5289 ( .A1(n5215), .A2(n8941), .ZN(n5214) );
  INV_X1 U5290 ( .A(n5216), .ZN(n5215) );
  NAND2_X1 U5291 ( .A1(n8983), .A2(n8973), .ZN(n5241) );
  NAND2_X1 U5292 ( .A1(n8985), .A2(n5364), .ZN(n8978) );
  AND2_X1 U5293 ( .A1(n6836), .A2(n7007), .ZN(n5364) );
  INV_X1 U5294 ( .A(n8973), .ZN(n6836) );
  NAND2_X1 U5295 ( .A1(n8990), .A2(n6848), .ZN(n8991) );
  OR2_X1 U5296 ( .A1(n9187), .A2(n8699), .ZN(n6803) );
  NAND2_X1 U5297 ( .A1(n7013), .A2(n7014), .ZN(n8973) );
  NAND2_X1 U5298 ( .A1(n9002), .A2(n9001), .ZN(n9000) );
  INV_X1 U5299 ( .A(n5259), .ZN(n5258) );
  AOI21_X1 U5300 ( .B1(n5259), .B2(n6833), .A(n4924), .ZN(n5257) );
  AND2_X1 U5301 ( .A1(n9020), .A2(n5260), .ZN(n5259) );
  INV_X1 U5302 ( .A(n6800), .ZN(n5260) );
  INV_X1 U5303 ( .A(n9020), .ZN(n6834) );
  NAND2_X1 U5304 ( .A1(n9042), .A2(n9041), .ZN(n5261) );
  NAND2_X1 U5305 ( .A1(n5072), .A2(n5336), .ZN(n9063) );
  AOI21_X1 U5306 ( .B1(n9091), .B2(n5338), .A(n5337), .ZN(n5336) );
  INV_X1 U5307 ( .A(n6894), .ZN(n5338) );
  INV_X1 U5308 ( .A(n7044), .ZN(n9074) );
  OR2_X1 U5309 ( .A1(n6576), .A2(n7270), .ZN(n6592) );
  OR2_X1 U5310 ( .A1(n9090), .A2(n9091), .ZN(n5247) );
  NAND2_X1 U5311 ( .A1(n5074), .A2(n5075), .ZN(n9108) );
  AND2_X1 U5312 ( .A1(n6894), .A2(n6895), .ZN(n9110) );
  NAND2_X1 U5313 ( .A1(n9122), .A2(n6831), .ZN(n9123) );
  INV_X1 U5314 ( .A(n9133), .ZN(n9137) );
  AND2_X1 U5315 ( .A1(n6896), .A2(n6897), .ZN(n9133) );
  AND2_X1 U5316 ( .A1(n6898), .A2(n6899), .ZN(n8443) );
  OR2_X1 U5317 ( .A1(n8442), .A2(n8443), .ZN(n5254) );
  AND2_X1 U5318 ( .A1(n6964), .A2(n6965), .ZN(n8299) );
  AOI21_X1 U5319 ( .B1(n8121), .B2(n8122), .A(n6828), .ZN(n8087) );
  NAND2_X1 U5320 ( .A1(n8087), .A2(n8086), .ZN(n8085) );
  NAND2_X1 U5321 ( .A1(n5249), .A2(n4920), .ZN(n5248) );
  NAND2_X1 U5322 ( .A1(n7816), .A2(n4897), .ZN(n7882) );
  OR2_X1 U5323 ( .A1(n7822), .A2(n8476), .ZN(n7895) );
  INV_X1 U5324 ( .A(n5351), .ZN(n5350) );
  OAI21_X1 U5325 ( .B1(n6790), .B2(n5352), .A(n7691), .ZN(n5351) );
  AND2_X1 U5326 ( .A1(n6944), .A2(n6945), .ZN(n7691) );
  NAND2_X1 U5327 ( .A1(n7670), .A2(n6790), .ZN(n7671) );
  AND2_X1 U5328 ( .A1(n6931), .A2(n6930), .ZN(n7527) );
  INV_X1 U5329 ( .A(n5086), .ZN(n5087) );
  NAND2_X1 U5330 ( .A1(n6780), .A2(n10402), .ZN(n6922) );
  NAND2_X1 U5331 ( .A1(n6909), .A2(n9159), .ZN(n9158) );
  INV_X1 U5332 ( .A(n9066), .ZN(n10450) );
  NAND2_X1 U5333 ( .A1(n6890), .A2(n7034), .ZN(n10453) );
  NAND2_X1 U5334 ( .A1(n6755), .A2(n6754), .ZN(n9176) );
  OR2_X1 U5335 ( .A1(n5251), .A2(n9276), .ZN(n6754) );
  OR2_X1 U5336 ( .A1(n5251), .A2(n8455), .ZN(n6656) );
  OR2_X1 U5337 ( .A1(n6756), .A2(n6757), .ZN(n10596) );
  NAND2_X1 U5338 ( .A1(n10342), .A2(n6739), .ZN(n10243) );
  OR2_X1 U5339 ( .A1(n10241), .A2(n6738), .ZN(n6739) );
  OR2_X1 U5340 ( .A1(n8148), .A2(n6749), .ZN(n10242) );
  NAND2_X1 U5341 ( .A1(n5264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5342 ( .A1(n6213), .A2(n6212), .ZN(n6729) );
  NAND2_X1 U5343 ( .A1(n5382), .A2(n5381), .ZN(n6231) );
  AOI21_X1 U5344 ( .B1(n5383), .B2(n6214), .A(n6214), .ZN(n5381) );
  INV_X1 U5345 ( .A(n5384), .ZN(n5383) );
  NAND2_X1 U5346 ( .A1(n5055), .A2(n4881), .ZN(n5054) );
  INV_X1 U5347 ( .A(n5056), .ZN(n5055) );
  AND3_X1 U5348 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U5349 ( .A1(n7977), .A2(n7980), .ZN(n7937) );
  OR2_X1 U5350 ( .A1(n5693), .A2(n5692), .ZN(n7978) );
  NOR2_X1 U5351 ( .A1(n5718), .A2(n5061), .ZN(n5060) );
  INV_X1 U5352 ( .A(n8025), .ZN(n5061) );
  NOR2_X1 U5353 ( .A1(n5719), .A2(n8025), .ZN(n5062) );
  NAND2_X1 U5354 ( .A1(n5063), .A2(n5718), .ZN(n8024) );
  OR2_X1 U5355 ( .A1(n7416), .A2(n7415), .ZN(n5015) );
  NOR2_X1 U5356 ( .A1(n7340), .A2(n4942), .ZN(n7343) );
  NAND2_X1 U5357 ( .A1(n7343), .A2(n7342), .ZN(n7398) );
  NAND2_X1 U5358 ( .A1(n9702), .A2(n9703), .ZN(n9701) );
  OR2_X1 U5359 ( .A1(n7403), .A2(n7402), .ZN(n5027) );
  AND2_X1 U5360 ( .A1(n5027), .A2(n5026), .ZN(n10308) );
  NAND2_X1 U5361 ( .A1(n7545), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5026) );
  OR2_X1 U5362 ( .A1(n10308), .A2(n10307), .ZN(n5025) );
  NOR2_X1 U5363 ( .A1(n7776), .A2(n4955), .ZN(n7779) );
  NOR2_X1 U5364 ( .A1(n7779), .A2(n7778), .ZN(n7800) );
  OR2_X1 U5365 ( .A1(n5803), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5843) );
  NOR2_X1 U5366 ( .A1(n5119), .A2(n10079), .ZN(n5116) );
  AND2_X1 U5367 ( .A1(n9846), .A2(n5117), .ZN(n9786) );
  NOR2_X1 U5368 ( .A1(n10063), .A2(n5118), .ZN(n5117) );
  OR2_X1 U5369 ( .A1(n5119), .A2(n10079), .ZN(n5118) );
  INV_X1 U5370 ( .A(n5154), .ZN(n8613) );
  OAI21_X1 U5371 ( .B1(n9855), .B2(n9852), .A(n4929), .ZN(n5154) );
  NAND2_X1 U5372 ( .A1(n8614), .A2(n5206), .ZN(n9838) );
  INV_X1 U5373 ( .A(n5207), .ZN(n5206) );
  AND2_X1 U5374 ( .A1(n9599), .A2(n9537), .ZN(n9837) );
  NAND2_X1 U5375 ( .A1(n9887), .A2(n8632), .ZN(n9889) );
  INV_X1 U5376 ( .A(n10094), .ZN(n8632) );
  NAND2_X1 U5377 ( .A1(n9895), .A2(n9901), .ZN(n9896) );
  AND2_X1 U5378 ( .A1(n9412), .A2(n9413), .ZN(n9935) );
  NAND2_X1 U5379 ( .A1(n9958), .A2(n5185), .ZN(n9942) );
  INV_X1 U5380 ( .A(n5186), .ZN(n5185) );
  NAND2_X1 U5381 ( .A1(n9583), .A2(n9582), .ZN(n9954) );
  NOR2_X1 U5382 ( .A1(n5898), .A2(n5897), .ZN(n5918) );
  AND2_X1 U5383 ( .A1(n5831), .A2(n5830), .ZN(n9996) );
  NAND2_X1 U5384 ( .A1(n10018), .A2(n9575), .ZN(n9995) );
  NAND2_X1 U5385 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  AOI21_X1 U5386 ( .B1(n9549), .B2(n8037), .A(n5175), .ZN(n5174) );
  AND2_X1 U5387 ( .A1(n8377), .A2(n8350), .ZN(n5208) );
  NOR2_X1 U5388 ( .A1(n5736), .A2(n5735), .ZN(n5755) );
  NAND2_X1 U5389 ( .A1(n8034), .A2(n10039), .ZN(n5201) );
  NAND2_X1 U5390 ( .A1(n8035), .A2(n5202), .ZN(n5200) );
  OR2_X1 U5391 ( .A1(n8034), .A2(n10039), .ZN(n5202) );
  NAND2_X1 U5392 ( .A1(n5200), .A2(n5198), .ZN(n8069) );
  NOR2_X1 U5393 ( .A1(n9518), .A2(n5199), .ZN(n5198) );
  INV_X1 U5394 ( .A(n5201), .ZN(n5199) );
  OR2_X1 U5395 ( .A1(n10560), .A2(n7919), .ZN(n10033) );
  NAND2_X1 U5396 ( .A1(n5192), .A2(n7853), .ZN(n10503) );
  AND2_X1 U5397 ( .A1(n5604), .A2(n5603), .ZN(n10483) );
  NAND2_X1 U5398 ( .A1(n5160), .A2(n7748), .ZN(n7763) );
  INV_X1 U5399 ( .A(n9622), .ZN(n5158) );
  OR2_X1 U5400 ( .A1(n10550), .A2(n7723), .ZN(n7432) );
  AND2_X1 U5401 ( .A1(n6181), .A2(n7717), .ZN(n10514) );
  OR2_X1 U5402 ( .A1(n6163), .A2(n6162), .ZN(n7428) );
  OAI21_X1 U5403 ( .B1(n10065), .B2(n10550), .A(n5132), .ZN(n5131) );
  NAND2_X1 U5404 ( .A1(n10063), .A2(n10561), .ZN(n5132) );
  AND2_X1 U5405 ( .A1(n7728), .A2(n8016), .ZN(n10562) );
  INV_X1 U5406 ( .A(n7862), .ZN(n10529) );
  INV_X1 U5407 ( .A(n6164), .ZN(n6165) );
  AND2_X1 U5408 ( .A1(n5291), .A2(n5412), .ZN(n5290) );
  NOR2_X1 U5409 ( .A1(n5414), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U5410 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5441) );
  OR2_X1 U5411 ( .A1(n6035), .A2(n6034), .ZN(n6057) );
  NAND2_X1 U5412 ( .A1(n5984), .A2(n5983), .ZN(n6009) );
  OAI22_X1 U5413 ( .A1(n5889), .A2(n5134), .B1(n5956), .B2(n5136), .ZN(n5963)
         );
  NAND2_X1 U5414 ( .A1(n5139), .A2(n5143), .ZN(n5134) );
  AOI21_X1 U5415 ( .B1(n5138), .B2(n5139), .A(n5137), .ZN(n5136) );
  NAND2_X1 U5416 ( .A1(n5135), .A2(n5139), .ZN(n5958) );
  NAND2_X1 U5417 ( .A1(n5889), .A2(n5140), .ZN(n5135) );
  AOI21_X1 U5418 ( .B1(n5888), .B2(n5887), .A(n4981), .ZN(n4980) );
  INV_X1 U5419 ( .A(n5932), .ZN(n4981) );
  NAND2_X1 U5420 ( .A1(n5305), .A2(n5303), .ZN(n5308) );
  NOR2_X1 U5421 ( .A1(n5304), .A2(n5821), .ZN(n5303) );
  INV_X1 U5422 ( .A(n5306), .ZN(n5304) );
  NAND2_X1 U5423 ( .A1(n5305), .A2(n5306), .ZN(n4971) );
  NAND2_X1 U5424 ( .A1(n5726), .A2(n5309), .ZN(n5748) );
  AND2_X1 U5425 ( .A1(n5728), .A2(n5725), .ZN(n5309) );
  INV_X1 U5426 ( .A(n5730), .ZN(n5728) );
  INV_X1 U5427 ( .A(n5589), .ZN(n5155) );
  AND2_X1 U5428 ( .A1(n5587), .A2(n5554), .ZN(n5555) );
  NAND2_X1 U5429 ( .A1(n5428), .A2(n5427), .ZN(n5531) );
  NAND2_X1 U5430 ( .A1(n6625), .A2(n6624), .ZN(n9204) );
  OR2_X1 U5431 ( .A1(n5251), .A2(n8332), .ZN(n6624) );
  OR2_X1 U5432 ( .A1(n6311), .A2(n6296), .ZN(n6299) );
  OR2_X1 U5433 ( .A1(n6295), .A2(n6294), .ZN(n6301) );
  OR2_X1 U5434 ( .A1(n6297), .A2(n8166), .ZN(n6298) );
  NOR2_X1 U5435 ( .A1(n4999), .A2(n5001), .ZN(n4995) );
  NOR2_X1 U5436 ( .A1(n5376), .A2(n5002), .ZN(n5001) );
  INV_X1 U5437 ( .A(n5377), .ZN(n5376) );
  OAI21_X1 U5438 ( .B1(n9176), .B2(n6717), .A(n5378), .ZN(n5377) );
  INV_X1 U5439 ( .A(n5374), .ZN(n4998) );
  NAND2_X1 U5440 ( .A1(n5368), .A2(n8760), .ZN(n5366) );
  AND2_X1 U5441 ( .A1(n7490), .A2(n6273), .ZN(n7423) );
  OR2_X1 U5442 ( .A1(n6288), .A2(n8058), .ZN(n6590) );
  OR2_X1 U5443 ( .A1(n8056), .A2(n6640), .ZN(n6591) );
  INV_X1 U5444 ( .A(n9026), .ZN(n9197) );
  NAND2_X1 U5445 ( .A1(n6513), .A2(n6512), .ZN(n8785) );
  INV_X1 U5446 ( .A(n6259), .ZN(n7058) );
  OAI21_X1 U5447 ( .B1(n7035), .B2(n6756), .A(n5317), .ZN(n5107) );
  NAND2_X1 U5448 ( .A1(n5320), .A2(n5319), .ZN(n5108) );
  NAND2_X1 U5449 ( .A1(n6714), .A2(n6713), .ZN(n8392) );
  AND2_X1 U5450 ( .A1(n6697), .A2(n6696), .ZN(n8765) );
  AND2_X1 U5451 ( .A1(n6681), .A2(n6680), .ZN(n8975) );
  AND2_X1 U5452 ( .A1(n6665), .A2(n6664), .ZN(n9015) );
  INV_X1 U5453 ( .A(n9014), .ZN(n9057) );
  AND2_X1 U5454 ( .A1(n6567), .A2(n6566), .ZN(n8736) );
  AND3_X1 U5455 ( .A1(n6553), .A2(n6552), .A3(n6551), .ZN(n8718) );
  AND3_X1 U5456 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(n8345) );
  INV_X1 U5457 ( .A(n6795), .ZN(n8777) );
  AND4_X1 U5458 ( .A1(n6501), .A2(n6500), .A3(n6499), .A4(n6498), .ZN(n8781)
         );
  AND4_X1 U5459 ( .A1(n6438), .A2(n6437), .A3(n6436), .A4(n6435), .ZN(n8460)
         );
  AND4_X1 U5460 ( .A1(n6416), .A2(n6415), .A3(n6414), .A4(n6413), .ZN(n8315)
         );
  AND4_X1 U5461 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n8556)
         );
  AND3_X1 U5462 ( .A1(n6314), .A2(n6313), .A3(n6312), .ZN(n6315) );
  AND2_X1 U5463 ( .A1(n6885), .A2(n6884), .ZN(n9170) );
  OR2_X1 U5464 ( .A1(n5251), .A2(n9270), .ZN(n6884) );
  XNOR2_X1 U5465 ( .A(n9171), .B(n9170), .ZN(n9169) );
  INV_X1 U5466 ( .A(n5261), .ZN(n9202) );
  NAND2_X1 U5467 ( .A1(n9053), .A2(n6988), .ZN(n9031) );
  NAND2_X1 U5468 ( .A1(n6279), .A2(n5232), .ZN(n5231) );
  INV_X1 U5469 ( .A(n7298), .ZN(n5232) );
  INV_X1 U5470 ( .A(n10460), .ZN(n9100) );
  AOI21_X1 U5471 ( .B1(n9169), .B2(n10404), .A(n5222), .ZN(n5221) );
  OAI21_X1 U5472 ( .B1(n9170), .B2(n10611), .A(n9173), .ZN(n5222) );
  NOR2_X1 U5473 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5100) );
  INV_X1 U5474 ( .A(n5400), .ZN(n5270) );
  INV_X1 U5475 ( .A(n5272), .ZN(n5271) );
  OAI21_X1 U5476 ( .B1(n4881), .B2(n5273), .A(n9381), .ZN(n5272) );
  INV_X1 U5477 ( .A(n4900), .ZN(n5273) );
  NAND2_X1 U5478 ( .A1(n5053), .A2(n5056), .ZN(n6096) );
  NAND2_X1 U5479 ( .A1(n5706), .A2(n5705), .ZN(n8109) );
  NAND2_X1 U5480 ( .A1(n5917), .A2(n5916), .ZN(n10117) );
  AND2_X1 U5481 ( .A1(n5880), .A2(n5879), .ZN(n9999) );
  OAI211_X1 U5482 ( .C1(n4872), .C2(n7286), .A(n5595), .B(n5594), .ZN(n10490)
         );
  OR2_X1 U5483 ( .A1(n7305), .A2(n5536), .ZN(n5595) );
  NAND2_X1 U5484 ( .A1(n6172), .A2(n10531), .ZN(n9408) );
  NAND2_X1 U5485 ( .A1(n9619), .A2(n9659), .ZN(n9662) );
  NAND2_X1 U5486 ( .A1(n9660), .A2(n8016), .ZN(n9661) );
  CLKBUF_X1 U5487 ( .A(n6180), .Z(n6181) );
  XNOR2_X1 U5488 ( .A(n7368), .B(n5028), .ZN(n7364) );
  INV_X1 U5489 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5028) );
  AND2_X1 U5490 ( .A1(n5017), .A2(n5016), .ZN(n7416) );
  NAND2_X1 U5491 ( .A1(n7324), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5016) );
  INV_X1 U5492 ( .A(n9777), .ZN(n5020) );
  NOR2_X1 U5493 ( .A1(n4886), .A2(n5152), .ZN(n5151) );
  INV_X1 U5494 ( .A(n8629), .ZN(n5153) );
  OAI21_X1 U5495 ( .B1(n9798), .B2(n5157), .A(n4922), .ZN(n5152) );
  NAND2_X1 U5496 ( .A1(n5968), .A2(n5967), .ZN(n10108) );
  OR2_X1 U5497 ( .A1(n8056), .A2(n5536), .ZN(n5968) );
  XNOR2_X1 U5498 ( .A(n5041), .B(n5040), .ZN(n5480) );
  INV_X1 U5499 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U5500 ( .A1(n5475), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5041) );
  INV_X1 U5501 ( .A(n9659), .ZN(n8016) );
  INV_X1 U5502 ( .A(n10494), .ZN(n9900) );
  NOR2_X1 U5503 ( .A1(n8514), .A2(n8513), .ZN(n10274) );
  NOR2_X1 U5504 ( .A1(n10272), .A2(n10271), .ZN(n8513) );
  NAND2_X1 U5505 ( .A1(n5096), .A2(n5392), .ZN(n5095) );
  INV_X1 U5506 ( .A(n6910), .ZN(n5096) );
  OAI22_X1 U5507 ( .A1(n4884), .A2(n5097), .B1(n6928), .B2(n6927), .ZN(n6929)
         );
  NAND2_X1 U5508 ( .A1(n6926), .A2(n5098), .ZN(n5097) );
  NAND2_X1 U5509 ( .A1(n5110), .A2(n5109), .ZN(n6957) );
  NOR2_X1 U5510 ( .A1(n7961), .A2(n6956), .ZN(n5109) );
  NAND2_X1 U5511 ( .A1(n5112), .A2(n5111), .ZN(n5110) );
  AND2_X1 U5512 ( .A1(n9959), .A2(n9457), .ZN(n4967) );
  INV_X1 U5513 ( .A(n9458), .ZN(n4966) );
  OAI21_X1 U5514 ( .B1(n6998), .B2(n6989), .A(n6990), .ZN(n6993) );
  AND2_X1 U5515 ( .A1(n9477), .A2(n9476), .ZN(n4961) );
  AND2_X1 U5516 ( .A1(n6607), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6626) );
  NOR2_X1 U5517 ( .A1(n5183), .A2(n5180), .ZN(n5179) );
  INV_X1 U5518 ( .A(n9416), .ZN(n5180) );
  OAI21_X1 U5519 ( .B1(n9901), .B2(n5183), .A(n9876), .ZN(n5182) );
  INV_X1 U5520 ( .A(SI_28_), .ZN(n7191) );
  INV_X1 U5521 ( .A(SI_25_), .ZN(n7092) );
  OR2_X1 U5522 ( .A1(n6033), .A2(n5314), .ZN(n5313) );
  INV_X1 U5523 ( .A(SI_14_), .ZN(n7114) );
  INV_X1 U5524 ( .A(SI_13_), .ZN(n7215) );
  INV_X1 U5525 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5299) );
  NOR2_X1 U5526 ( .A1(n6411), .A2(n6410), .ZN(n6409) );
  AND2_X1 U5527 ( .A1(n9176), .A2(n8743), .ZN(n6760) );
  NOR2_X1 U5528 ( .A1(n6592), .A2(n8690), .ZN(n6607) );
  NOR2_X1 U5529 ( .A1(n6496), .A2(n8102), .ZN(n6495) );
  NOR2_X1 U5530 ( .A1(n6533), .A2(n6532), .ZN(n6546) );
  NOR2_X1 U5531 ( .A1(n4990), .A2(n4991), .ZN(n4989) );
  AND2_X1 U5532 ( .A1(n6409), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6431) );
  INV_X1 U5533 ( .A(n7022), .ZN(n5359) );
  NOR2_X1 U5534 ( .A1(n8937), .A2(n7022), .ZN(n5357) );
  AOI221_X1 U5535 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7275), .C1(n10383), .C2(
        keyinput_123), .A(n7274), .ZN(n7280) );
  AOI21_X1 U5536 ( .B1(keyinput_122), .B2(n8792), .A(n7273), .ZN(n7274) );
  AOI211_X1 U5537 ( .C1(n7175), .C2(n7174), .A(n7173), .B(n7172), .ZN(n7281)
         );
  AND2_X1 U5538 ( .A1(n6689), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6704) );
  NOR2_X1 U5539 ( .A1(n9176), .A2(n5217), .ZN(n5216) );
  INV_X1 U5540 ( .A(n5218), .ZN(n5217) );
  INV_X1 U5541 ( .A(n6995), .ZN(n5080) );
  NOR2_X1 U5542 ( .A1(n6674), .A2(n6673), .ZN(n6689) );
  OR2_X1 U5543 ( .A1(n9216), .A2(n9056), .ZN(n6799) );
  INV_X1 U5544 ( .A(n6980), .ZN(n5337) );
  AND2_X1 U5545 ( .A1(n6546), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6558) );
  INV_X1 U5546 ( .A(n5344), .ZN(n5343) );
  NOR2_X1 U5547 ( .A1(n8305), .A2(n8785), .ZN(n5230) );
  INV_X1 U5548 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8775) );
  OR2_X1 U5549 ( .A1(n8127), .A2(n8128), .ZN(n8090) );
  NAND2_X1 U5550 ( .A1(n5067), .A2(n5250), .ZN(n5249) );
  INV_X1 U5551 ( .A(n5397), .ZN(n5250) );
  INV_X1 U5552 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6410) );
  INV_X1 U5553 ( .A(n6940), .ZN(n5352) );
  NOR2_X1 U5554 ( .A1(n5352), .A2(n5349), .ZN(n5348) );
  NAND2_X1 U5555 ( .A1(n5230), .A2(n5229), .ZN(n9143) );
  AND2_X1 U5556 ( .A1(n6204), .A2(n6211), .ZN(n5093) );
  OAI21_X1 U5557 ( .B1(n6214), .B2(n6228), .A(n6229), .ZN(n5384) );
  OR2_X1 U5558 ( .A1(n6405), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6406) );
  AND2_X1 U5559 ( .A1(n5277), .A2(n5654), .ZN(n5276) );
  INV_X1 U5560 ( .A(n5508), .ZN(n5618) );
  NOR2_X1 U5561 ( .A1(n5035), .A2(n5031), .ZN(n5030) );
  NOR2_X1 U5562 ( .A1(n5818), .A2(n9289), .ZN(n5035) );
  OR2_X1 U5563 ( .A1(n10074), .A2(n8588), .ZN(n9603) );
  NAND2_X1 U5564 ( .A1(n8585), .A2(n9583), .ZN(n5186) );
  NOR2_X1 U5565 ( .A1(n10024), .A2(n10139), .ZN(n10000) );
  OR2_X1 U5566 ( .A1(n10128), .A2(n9999), .ZN(n9580) );
  NOR2_X1 U5567 ( .A1(n5127), .A2(n8409), .ZN(n5126) );
  INV_X1 U5568 ( .A(n5128), .ZN(n5127) );
  INV_X1 U5569 ( .A(n9563), .ZN(n5175) );
  NOR2_X1 U5570 ( .A1(n10159), .A2(n9439), .ZN(n5128) );
  INV_X1 U5571 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7394) );
  NOR2_X1 U5572 ( .A1(n10506), .A2(n7862), .ZN(n5123) );
  NAND2_X1 U5573 ( .A1(n10516), .A2(n7851), .ZN(n9634) );
  AND2_X1 U5574 ( .A1(n9630), .A2(n9634), .ZN(n10476) );
  INV_X1 U5575 ( .A(n7706), .ZN(n6162) );
  INV_X1 U5576 ( .A(n5211), .ZN(n5210) );
  INV_X1 U5577 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5412) );
  AND2_X1 U5578 ( .A1(n6877), .A2(n6868), .ZN(n6875) );
  AND2_X1 U5579 ( .A1(n6864), .A2(n6810), .ZN(n6862) );
  INV_X1 U5580 ( .A(SI_26_), .ZN(n7197) );
  INV_X1 U5581 ( .A(SI_27_), .ZN(n7194) );
  NOR2_X1 U5582 ( .A1(n6008), .A2(n5331), .ZN(n5330) );
  INV_X1 U5583 ( .A(n5983), .ZN(n5331) );
  INV_X1 U5584 ( .A(SI_23_), .ZN(n7105) );
  INV_X1 U5585 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5454) );
  INV_X1 U5586 ( .A(SI_21_), .ZN(n7118) );
  INV_X1 U5587 ( .A(n5140), .ZN(n5138) );
  INV_X1 U5588 ( .A(n5957), .ZN(n5137) );
  INV_X1 U5589 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U5590 ( .A1(n5402), .A2(n5141), .ZN(n5140) );
  AND2_X1 U5591 ( .A1(n5932), .A2(n5933), .ZN(n5939) );
  AOI21_X1 U5592 ( .B1(n4980), .B2(n5141), .A(n5935), .ZN(n4978) );
  INV_X1 U5593 ( .A(n4978), .ZN(n4975) );
  INV_X1 U5594 ( .A(n4980), .ZN(n4979) );
  INV_X1 U5595 ( .A(n5936), .ZN(n4976) );
  INV_X1 U5596 ( .A(SI_17_), .ZN(n7113) );
  INV_X1 U5597 ( .A(SI_18_), .ZN(n7107) );
  AOI21_X1 U5598 ( .B1(n4885), .B2(n4943), .A(n5307), .ZN(n5306) );
  INV_X1 U5599 ( .A(n5819), .ZN(n5307) );
  INV_X1 U5600 ( .A(SI_5_), .ZN(n7226) );
  NAND2_X1 U5601 ( .A1(n8017), .A2(n6489), .ZN(n8099) );
  NAND2_X1 U5602 ( .A1(n8099), .A2(n8100), .ZN(n8098) );
  NAND2_X1 U5603 ( .A1(n6760), .A2(n6717), .ZN(n5378) );
  INV_X1 U5604 ( .A(n6703), .ZN(n5002) );
  AOI21_X1 U5605 ( .B1(n8758), .B2(n5370), .A(n5369), .ZN(n5368) );
  INV_X1 U5606 ( .A(n6686), .ZN(n5369) );
  INV_X1 U5607 ( .A(n6670), .ZN(n5370) );
  AND2_X1 U5608 ( .A1(n6385), .A2(n6370), .ZN(n5389) );
  NAND2_X1 U5609 ( .A1(n6815), .A2(n6302), .ZN(n6286) );
  INV_X1 U5610 ( .A(n5385), .ZN(n5007) );
  INV_X1 U5611 ( .A(n6572), .ZN(n5005) );
  OR2_X1 U5612 ( .A1(n6464), .A2(n7988), .ZN(n6478) );
  INV_X1 U5613 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U5614 ( .A1(n8772), .A2(n8773), .ZN(n8771) );
  NOR2_X1 U5615 ( .A1(n6751), .A2(n6756), .ZN(n5319) );
  MUX2_X1 U5616 ( .A(n7051), .B(n7052), .S(n7028), .Z(n7033) );
  NOR2_X1 U5617 ( .A1(n5318), .A2(n5392), .ZN(n5317) );
  XNOR2_X1 U5618 ( .A(n7053), .B(n8993), .ZN(n5318) );
  NOR2_X1 U5619 ( .A1(n5332), .A2(n7049), .ZN(n7050) );
  OR2_X1 U5620 ( .A1(n6309), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6314) );
  INV_X1 U5621 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8186) );
  AND2_X1 U5622 ( .A1(n6704), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8942) );
  INV_X1 U5623 ( .A(n7049), .ZN(n7019) );
  OAI22_X1 U5624 ( .A1(n5238), .A2(n8952), .B1(n9176), .B2(n8392), .ZN(n5236)
         );
  NAND2_X1 U5625 ( .A1(n8990), .A2(n5216), .ZN(n8961) );
  OR2_X1 U5626 ( .A1(n6658), .A2(n8700), .ZN(n6674) );
  AND2_X1 U5627 ( .A1(n6634), .A2(n6633), .ZN(n9014) );
  NAND2_X1 U5628 ( .A1(n9071), .A2(n6832), .ZN(n9054) );
  AOI21_X1 U5629 ( .B1(n4883), .B2(n8443), .A(n4923), .ZN(n5252) );
  INV_X1 U5630 ( .A(n5230), .ZN(n8447) );
  INV_X1 U5631 ( .A(n8299), .ZN(n8303) );
  AOI22_X1 U5632 ( .A1(n7962), .A2(n7961), .B1(n5212), .B2(n8326), .ZN(n8120)
         );
  AND2_X1 U5633 ( .A1(n6959), .A2(n6960), .ZN(n8122) );
  NAND2_X1 U5634 ( .A1(n5213), .A2(n5212), .ZN(n8127) );
  AOI21_X1 U5635 ( .B1(n6822), .B2(n5071), .A(n5070), .ZN(n5069) );
  INV_X1 U5636 ( .A(n6945), .ZN(n5071) );
  INV_X1 U5637 ( .A(n6953), .ZN(n5070) );
  NAND2_X1 U5638 ( .A1(n7683), .A2(n6945), .ZN(n7886) );
  NOR2_X1 U5639 ( .A1(n5225), .A2(n7695), .ZN(n5223) );
  INV_X1 U5640 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8199) );
  NOR2_X1 U5641 ( .A1(n10445), .A2(n5225), .ZN(n7692) );
  NAND2_X1 U5642 ( .A1(n4887), .A2(n5086), .ZN(n5083) );
  OR2_X1 U5643 ( .A1(n10445), .A2(n8570), .ZN(n7635) );
  OR2_X1 U5644 ( .A1(n9156), .A2(n10374), .ZN(n9154) );
  OR2_X1 U5645 ( .A1(n7564), .A2(n7563), .ZN(n7566) );
  NAND2_X1 U5646 ( .A1(n6812), .A2(n6811), .ZN(n8941) );
  OR2_X1 U5647 ( .A1(n5251), .A2(n9272), .ZN(n6811) );
  NAND2_X1 U5648 ( .A1(n6688), .A2(n6687), .ZN(n9181) );
  OR2_X1 U5649 ( .A1(n5251), .A2(n9278), .ZN(n6687) );
  INV_X1 U5650 ( .A(n10613), .ZN(n10404) );
  OR2_X1 U5651 ( .A1(n6288), .A2(n7301), .ZN(n6292) );
  OR2_X1 U5652 ( .A1(n7564), .A2(n6852), .ZN(n6857) );
  NAND2_X1 U5653 ( .A1(n6735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U5654 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  INV_X1 U5655 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6733) );
  OR2_X1 U5656 ( .A1(n6235), .A2(n6214), .ZN(n6543) );
  AND2_X1 U5657 ( .A1(n6341), .A2(n6371), .ZN(n8160) );
  OR2_X1 U5658 ( .A1(n6095), .A2(n6094), .ZN(n5400) );
  NAND2_X1 U5659 ( .A1(n9378), .A2(n6004), .ZN(n5048) );
  NAND2_X1 U5660 ( .A1(n9312), .A2(n4916), .ZN(n5037) );
  INV_X1 U5661 ( .A(n5393), .ZN(n5039) );
  NAND2_X1 U5662 ( .A1(n5289), .A2(n8541), .ZN(n9339) );
  AND2_X1 U5663 ( .A1(n8542), .A2(n9340), .ZN(n5289) );
  OR2_X1 U5664 ( .A1(n5048), .A2(n6025), .ZN(n9301) );
  INV_X1 U5665 ( .A(n9378), .ZN(n5042) );
  AND2_X1 U5666 ( .A1(n5918), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5943) );
  AND2_X1 U5667 ( .A1(n5969), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5987) );
  OAI21_X1 U5668 ( .B1(n10364), .B2(n5639), .A(n5474), .ZN(n5479) );
  INV_X1 U5669 ( .A(n5858), .ZN(n5288) );
  AND2_X1 U5670 ( .A1(n5885), .A2(n9340), .ZN(n5287) );
  NAND2_X1 U5671 ( .A1(n5034), .A2(n5032), .ZN(n5840) );
  OR2_X1 U5672 ( .A1(n5817), .A2(n5033), .ZN(n5032) );
  NAND2_X1 U5673 ( .A1(n8410), .A2(n5030), .ZN(n5034) );
  INV_X1 U5674 ( .A(n9289), .ZN(n5033) );
  AND2_X1 U5675 ( .A1(n9782), .A2(n9669), .ZN(n9616) );
  NAND2_X1 U5676 ( .A1(n4958), .A2(n4957), .ZN(n9618) );
  AND2_X1 U5677 ( .A1(n9507), .A2(n9506), .ZN(n4957) );
  NAND2_X1 U5678 ( .A1(n9501), .A2(n4911), .ZN(n4958) );
  INV_X1 U5679 ( .A(n9616), .ZN(n9656) );
  OR2_X1 U5680 ( .A1(n7469), .A2(n7468), .ZN(n5017) );
  NAND2_X1 U5681 ( .A1(n7398), .A2(n4941), .ZN(n9702) );
  AND2_X1 U5682 ( .A1(n5025), .A2(n5024), .ZN(n10329) );
  NAND2_X1 U5683 ( .A1(n10312), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U5684 ( .A1(n8589), .A2(n10511), .ZN(n5156) );
  NAND2_X1 U5685 ( .A1(n5149), .A2(n5147), .ZN(n9792) );
  NAND2_X1 U5686 ( .A1(n5207), .A2(n5204), .ZN(n5149) );
  INV_X1 U5687 ( .A(n5148), .ZN(n5147) );
  AND2_X1 U5688 ( .A1(n9482), .A2(n9541), .ZN(n9791) );
  NAND2_X1 U5689 ( .A1(n9820), .A2(n9603), .ZN(n9797) );
  NAND2_X1 U5690 ( .A1(n4972), .A2(n9477), .ZN(n9820) );
  INV_X1 U5691 ( .A(n9816), .ZN(n4972) );
  AND2_X1 U5692 ( .A1(n6133), .A2(n6085), .ZN(n9832) );
  AOI21_X1 U5693 ( .B1(n4898), .B2(n5168), .A(n5164), .ZN(n5163) );
  NAND2_X1 U5694 ( .A1(n9861), .A2(n4898), .ZN(n5165) );
  INV_X1 U5695 ( .A(n9542), .ZN(n5168) );
  NAND2_X1 U5696 ( .A1(n9861), .A2(n9868), .ZN(n9862) );
  INV_X1 U5697 ( .A(n5194), .ZN(n5193) );
  OR2_X1 U5698 ( .A1(n10117), .A2(n9956), .ZN(n5197) );
  NAND2_X1 U5699 ( .A1(n9982), .A2(n9967), .ZN(n9964) );
  NAND2_X1 U5700 ( .A1(n10000), .A2(n8630), .ZN(n10001) );
  AND2_X1 U5701 ( .A1(n5904), .A2(n5903), .ZN(n9975) );
  NAND2_X1 U5702 ( .A1(n5169), .A2(n5171), .ZN(n9978) );
  AOI21_X1 U5703 ( .B1(n9994), .B2(n5173), .A(n5172), .ZN(n5171) );
  INV_X1 U5704 ( .A(n9575), .ZN(n5173) );
  AND2_X1 U5705 ( .A1(n9580), .A2(n9546), .ZN(n9977) );
  INV_X1 U5706 ( .A(n4872), .ZN(n5914) );
  AND2_X1 U5707 ( .A1(n5811), .A2(n5810), .ZN(n10017) );
  NAND2_X1 U5708 ( .A1(n8075), .A2(n5124), .ZN(n10024) );
  NOR2_X1 U5709 ( .A1(n5125), .A2(n10146), .ZN(n5124) );
  INV_X1 U5710 ( .A(n5126), .ZN(n5125) );
  NAND2_X1 U5711 ( .A1(n8374), .A2(n9566), .ZN(n8402) );
  NAND2_X1 U5712 ( .A1(n8075), .A2(n8081), .ZN(n8382) );
  NAND2_X1 U5713 ( .A1(n8075), .A2(n5128), .ZN(n8380) );
  NAND2_X1 U5714 ( .A1(n8071), .A2(n9434), .ZN(n8349) );
  OR2_X1 U5715 ( .A1(n5707), .A2(n8027), .ZN(n5736) );
  AND2_X1 U5716 ( .A1(n8045), .A2(n8044), .ZN(n8075) );
  NAND2_X1 U5717 ( .A1(n8042), .A2(n9518), .ZN(n8071) );
  AND2_X1 U5718 ( .A1(n10582), .A2(n10051), .ZN(n8045) );
  OR2_X1 U5719 ( .A1(n9431), .A2(n7916), .ZN(n9427) );
  NAND2_X1 U5720 ( .A1(n10037), .A2(n10033), .ZN(n8039) );
  NOR2_X1 U5721 ( .A1(n10049), .A2(n10560), .ZN(n10051) );
  AND2_X1 U5722 ( .A1(n7853), .A2(n7913), .ZN(n5191) );
  NAND2_X1 U5723 ( .A1(n5189), .A2(n4908), .ZN(n5188) );
  NAND2_X1 U5724 ( .A1(n5123), .A2(n5122), .ZN(n10049) );
  INV_X1 U5725 ( .A(n5123), .ZN(n10507) );
  AND2_X1 U5726 ( .A1(n9632), .A2(n7917), .ZN(n10509) );
  NAND2_X1 U5727 ( .A1(n7747), .A2(n7746), .ZN(n7749) );
  NAND2_X1 U5728 ( .A1(n5159), .A2(n5161), .ZN(n7747) );
  INV_X1 U5729 ( .A(n7720), .ZN(n5161) );
  INV_X1 U5730 ( .A(n10511), .ZN(n10479) );
  NAND2_X1 U5731 ( .A1(n7723), .A2(n8016), .ZN(n7715) );
  AND2_X1 U5732 ( .A1(n8016), .A2(n9900), .ZN(n7706) );
  NAND2_X1 U5733 ( .A1(n9497), .A2(n9496), .ZN(n10060) );
  AND3_X1 U5734 ( .A1(n5565), .A2(n5564), .A3(n5563), .ZN(n10434) );
  INV_X1 U5735 ( .A(n10562), .ZN(n10583) );
  AND2_X1 U5736 ( .A1(n5480), .A2(n9620), .ZN(n7728) );
  INV_X1 U5737 ( .A(n6149), .ZN(n7294) );
  INV_X1 U5738 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U5739 ( .A1(n5417), .A2(n5416), .ZN(n5464) );
  XNOR2_X1 U5740 ( .A(n6863), .B(n6862), .ZN(n9271) );
  NAND2_X1 U5741 ( .A1(n5435), .A2(n5434), .ZN(n5440) );
  NAND2_X1 U5742 ( .A1(n6057), .A2(n6056), .ZN(n6079) );
  NAND2_X1 U5743 ( .A1(n5455), .A2(n5454), .ZN(n5475) );
  NAND2_X1 U5744 ( .A1(n5842), .A2(n5841), .ZN(n5859) );
  AND2_X1 U5745 ( .A1(n5804), .A2(n5843), .ZN(n8003) );
  AOI21_X1 U5746 ( .B1(n5796), .B2(n5795), .A(n4885), .ZN(n5820) );
  INV_X1 U5747 ( .A(n5284), .ZN(n5282) );
  NAND2_X1 U5748 ( .A1(n5322), .A2(n5670), .ZN(n5697) );
  NAND2_X1 U5749 ( .A1(n5656), .A2(n5326), .ZN(n5322) );
  NAND2_X1 U5750 ( .A1(n5656), .A2(n5655), .ZN(n5672) );
  AND2_X1 U5751 ( .A1(n5655), .A2(n5631), .ZN(n5632) );
  AOI21_X1 U5752 ( .B1(n5591), .B2(n5294), .A(n5295), .ZN(n5292) );
  INV_X1 U5753 ( .A(n5605), .ZN(n5295) );
  AND2_X1 U5754 ( .A1(n5627), .A2(n5609), .ZN(n5610) );
  NAND2_X1 U5755 ( .A1(n5492), .A2(n5423), .ZN(n5428) );
  NOR2_X1 U5756 ( .A1(n10259), .A2(n8492), .ZN(n8493) );
  NAND2_X1 U5757 ( .A1(n8568), .A2(n6370), .ZN(n7653) );
  NAND2_X1 U5758 ( .A1(n8478), .A2(n6422), .ZN(n7075) );
  NAND2_X1 U5759 ( .A1(n5008), .A2(n5385), .ZN(n8674) );
  NOR2_X1 U5760 ( .A1(n6768), .A2(n6762), .ZN(n8766) );
  NAND2_X1 U5761 ( .A1(n7833), .A2(n6459), .ZN(n7995) );
  INV_X1 U5762 ( .A(n7612), .ZN(n6272) );
  INV_X1 U5763 ( .A(n10372), .ZN(n8782) );
  OAI21_X1 U5764 ( .B1(n6455), .B2(n4985), .A(n4984), .ZN(n8018) );
  INV_X1 U5765 ( .A(n4992), .ZN(n4985) );
  AOI21_X1 U5766 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n4984) );
  NAND2_X1 U5767 ( .A1(n6606), .A2(n6605), .ZN(n9210) );
  OR2_X1 U5768 ( .A1(n5251), .A2(n8480), .ZN(n6605) );
  INV_X1 U5769 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10383) );
  AND2_X1 U5770 ( .A1(n8766), .A2(n10448), .ZN(n10373) );
  AND2_X1 U5771 ( .A1(n8766), .A2(n10450), .ZN(n10372) );
  INV_X1 U5772 ( .A(n8740), .ZN(n8780) );
  NAND2_X1 U5773 ( .A1(n5367), .A2(n8758), .ZN(n8639) );
  INV_X1 U5774 ( .A(n10373), .ZN(n8778) );
  AND2_X1 U5775 ( .A1(n6583), .A2(n6582), .ZN(n9067) );
  AND4_X1 U5776 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n8709)
         );
  AND4_X1 U5777 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(n8338)
         );
  AND4_X1 U5778 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n6451), .ZN(n8322)
         );
  AND4_X1 U5779 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n8468)
         );
  AND4_X1 U5780 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n8328)
         );
  INV_X1 U5781 ( .A(n10449), .ZN(n8561) );
  NOR2_X1 U5782 ( .A1(n10625), .A2(n4904), .ZN(n8184) );
  NOR2_X1 U5783 ( .A1(n8184), .A2(n8185), .ZN(n8183) );
  AOI21_X1 U5784 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n8162), .A(n8267), .ZN(
        n8229) );
  AOI21_X1 U5785 ( .B1(n8201), .B2(P2_REG2_REG_6__SCAN_IN), .A(n8196), .ZN(
        n8197) );
  AOI21_X1 U5786 ( .B1(n8217), .B2(P2_REG2_REG_8__SCAN_IN), .A(n8255), .ZN(
        n8214) );
  AOI21_X1 U5787 ( .B1(n8789), .B2(P2_REG2_REG_10__SCAN_IN), .A(n8788), .ZN(
        n8790) );
  AND2_X1 U5788 ( .A1(n5094), .A2(n6338), .ZN(n6460) );
  XNOR2_X1 U5789 ( .A(n8873), .B(n8863), .ZN(n8852) );
  NAND2_X1 U5790 ( .A1(n8852), .A2(n8307), .ZN(n8875) );
  NAND2_X1 U5791 ( .A1(n8155), .A2(n8152), .ZN(n10636) );
  OR2_X1 U5792 ( .A1(n5251), .A2(n8528), .ZN(n6869) );
  XNOR2_X1 U5793 ( .A(n5242), .B(n7019), .ZN(n8950) );
  OAI21_X1 U5794 ( .B1(n8984), .B2(n5237), .A(n5235), .ZN(n5242) );
  OR2_X1 U5795 ( .A1(n5241), .A2(n8952), .ZN(n5237) );
  INV_X1 U5796 ( .A(n5236), .ZN(n5235) );
  NAND2_X1 U5797 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  XNOR2_X1 U5798 ( .A(n6861), .B(n7049), .ZN(n5089) );
  INV_X1 U5799 ( .A(n5234), .ZN(n8959) );
  OAI21_X1 U5800 ( .B1(n8984), .B2(n5241), .A(n5238), .ZN(n5234) );
  NAND2_X1 U5801 ( .A1(n8985), .A2(n7007), .ZN(n8974) );
  AND2_X1 U5802 ( .A1(n9000), .A2(n7004), .ZN(n8987) );
  OR2_X1 U5803 ( .A1(n5251), .A2(n9281), .ZN(n6671) );
  AND2_X1 U5804 ( .A1(n6642), .A2(n6641), .ZN(n9026) );
  OR2_X1 U5805 ( .A1(n5251), .A2(n8432), .ZN(n6641) );
  NAND2_X1 U5806 ( .A1(n5261), .A2(n5259), .ZN(n9019) );
  NAND2_X1 U5807 ( .A1(n5247), .A2(n4882), .ZN(n9073) );
  AND2_X1 U5808 ( .A1(n5247), .A2(n4934), .ZN(n9075) );
  NAND2_X1 U5809 ( .A1(n9086), .A2(n9091), .ZN(n9085) );
  NAND2_X1 U5810 ( .A1(n9108), .A2(n6894), .ZN(n9086) );
  NAND2_X1 U5811 ( .A1(n6557), .A2(n6556), .ZN(n6797) );
  NAND2_X1 U5812 ( .A1(n9123), .A2(n6974), .ZN(n9109) );
  AND2_X1 U5813 ( .A1(n9127), .A2(n9126), .ZN(n9234) );
  NAND2_X1 U5814 ( .A1(n5254), .A2(n4883), .ZN(n9136) );
  AND2_X1 U5815 ( .A1(n5254), .A2(n4895), .ZN(n9138) );
  NAND2_X1 U5816 ( .A1(n8085), .A2(n6901), .ZN(n8300) );
  NAND2_X1 U5817 ( .A1(n7882), .A2(n5397), .ZN(n7873) );
  NAND2_X1 U5818 ( .A1(n7671), .A2(n6940), .ZN(n7684) );
  NAND2_X1 U5819 ( .A1(n5262), .A2(n6791), .ZN(n7690) );
  NAND2_X1 U5820 ( .A1(n7570), .A2(n5087), .ZN(n5085) );
  NAND2_X1 U5821 ( .A1(n9164), .A2(n7578), .ZN(n10461) );
  NAND2_X1 U5822 ( .A1(n7569), .A2(n6922), .ZN(n10446) );
  OR2_X1 U5823 ( .A1(n10242), .A2(n6851), .ZN(n10470) );
  OAI211_X1 U5824 ( .C1(n6909), .C2(n9159), .A(n9158), .B(n10453), .ZN(n9163)
         );
  INV_X1 U5825 ( .A(n10461), .ZN(n9153) );
  NAND2_X1 U5826 ( .A1(n9164), .A2(n7596), .ZN(n10460) );
  OR3_X1 U5827 ( .A1(n9209), .A2(n9208), .A3(n9207), .ZN(n9257) );
  INV_X2 U5828 ( .A(n10621), .ZN(n10624) );
  XNOR2_X1 U5829 ( .A(n6737), .B(P2_IR_REG_24__SCAN_IN), .ZN(n10343) );
  NAND2_X1 U5830 ( .A1(n6736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U5831 ( .A1(n6748), .A2(n6747), .ZN(n6736) );
  NAND2_X1 U5832 ( .A1(n6218), .A2(n6215), .ZN(n6246) );
  AND2_X1 U5833 ( .A1(n6730), .A2(n6729), .ZN(n10342) );
  NOR2_X1 U5834 ( .A1(n6473), .A2(n6210), .ZN(n6731) );
  INV_X1 U5835 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U5836 ( .A1(n6241), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U5837 ( .A1(n6277), .A2(n6276), .ZN(n8167) );
  NOR2_X1 U5838 ( .A1(n7069), .A2(n8334), .ZN(n7313) );
  NAND2_X1 U5839 ( .A1(n5280), .A2(n5626), .ZN(n7908) );
  INV_X1 U5840 ( .A(n7642), .ZN(n5281) );
  AND2_X1 U5841 ( .A1(n5662), .A2(n5661), .ZN(n7919) );
  AND2_X1 U5842 ( .A1(n5782), .A2(n5781), .ZN(n9292) );
  NAND2_X1 U5843 ( .A1(n5036), .A2(n5817), .ZN(n9286) );
  OR2_X1 U5844 ( .A1(n5036), .A2(n5817), .ZN(n9287) );
  NAND2_X1 U5845 ( .A1(n5048), .A2(n6025), .ZN(n9305) );
  INV_X1 U5846 ( .A(n9299), .ZN(n6052) );
  INV_X1 U5847 ( .A(n5051), .ZN(n5050) );
  OAI21_X1 U5848 ( .B1(n4905), .B2(n5052), .A(n6195), .ZN(n5051) );
  NAND2_X1 U5849 ( .A1(n5037), .A2(n5038), .ZN(n9321) );
  AND2_X1 U5850 ( .A1(n5739), .A2(n5738), .ZN(n8379) );
  AND2_X1 U5851 ( .A1(n5584), .A2(n5583), .ZN(n10417) );
  NAND2_X1 U5852 ( .A1(n5942), .A2(n5941), .ZN(n10112) );
  NOR2_X1 U5853 ( .A1(n8059), .A2(n5060), .ZN(n5059) );
  NAND2_X1 U5854 ( .A1(n4893), .A2(n5267), .ZN(n8060) );
  NAND2_X1 U5855 ( .A1(n8024), .A2(n8025), .ZN(n5267) );
  NAND2_X1 U5856 ( .A1(n6178), .A2(n7449), .ZN(n9402) );
  INV_X1 U5857 ( .A(n9342), .ZN(n9401) );
  AND2_X1 U5858 ( .A1(n8541), .A2(n8542), .ZN(n8544) );
  NAND4_X1 U5859 ( .A1(n5685), .A2(n5684), .A3(n5683), .A4(n5682), .ZN(n10039)
         );
  NOR2_X1 U5860 ( .A1(n7364), .A2(n7457), .ZN(n7363) );
  INV_X1 U5861 ( .A(n5017), .ZN(n7467) );
  INV_X1 U5862 ( .A(n5015), .ZN(n7414) );
  NAND2_X1 U5863 ( .A1(n7326), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5014) );
  INV_X1 U5864 ( .A(n5027), .ZN(n7544) );
  INV_X1 U5865 ( .A(n5025), .ZN(n10306) );
  AND2_X1 U5866 ( .A1(n7542), .A2(n10330), .ZN(n10331) );
  NOR2_X1 U5867 ( .A1(n7800), .A2(n4954), .ZN(n7802) );
  NAND2_X1 U5868 ( .A1(n7802), .A2(n7803), .ZN(n8002) );
  NOR2_X1 U5869 ( .A1(n9771), .A2(n5023), .ZN(n5022) );
  AND2_X1 U5870 ( .A1(n9772), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5023) );
  INV_X1 U5871 ( .A(n10060), .ZN(n9787) );
  NAND2_X1 U5872 ( .A1(n6130), .A2(n6129), .ZN(n10066) );
  NAND2_X1 U5873 ( .A1(n9838), .A2(n8616), .ZN(n9810) );
  AND2_X1 U5874 ( .A1(n8614), .A2(n8613), .ZN(n9839) );
  NAND2_X1 U5875 ( .A1(n6011), .A2(n6010), .ZN(n10094) );
  NAND2_X1 U5876 ( .A1(n9896), .A2(n9641), .ZN(n9877) );
  NAND2_X1 U5877 ( .A1(n9942), .A2(n9586), .ZN(n9927) );
  NAND2_X1 U5878 ( .A1(n9953), .A2(n8603), .ZN(n9940) );
  AND2_X1 U5879 ( .A1(n9972), .A2(n8602), .ZN(n9955) );
  NAND2_X1 U5880 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  NAND2_X1 U5881 ( .A1(n8595), .A2(n8594), .ZN(n10013) );
  NAND2_X1 U5882 ( .A1(n8351), .A2(n8350), .ZN(n8371) );
  NAND2_X1 U5883 ( .A1(n10536), .A2(n10489), .ZN(n10530) );
  NAND2_X1 U5884 ( .A1(n10503), .A2(n7854), .ZN(n7914) );
  OR2_X1 U5885 ( .A1(n5536), .A2(n7302), .ZN(n5432) );
  NAND2_X1 U5886 ( .A1(n4872), .A2(n4888), .ZN(n5114) );
  NAND2_X1 U5887 ( .A1(n5700), .A2(n5451), .ZN(n5476) );
  INV_X1 U5888 ( .A(n7432), .ZN(n6171) );
  INV_X1 U5889 ( .A(n10530), .ZN(n10045) );
  INV_X1 U5890 ( .A(n10531), .ZN(n10491) );
  NAND2_X1 U5891 ( .A1(n10064), .A2(n10562), .ZN(n5133) );
  INV_X1 U5892 ( .A(n5131), .ZN(n5130) );
  NAND2_X1 U5893 ( .A1(n7069), .A2(n6169), .ZN(n10287) );
  AND2_X1 U5894 ( .A1(n10207), .A2(n8436), .ZN(n7296) );
  XNOR2_X1 U5895 ( .A(n6882), .B(n6881), .ZN(n10189) );
  INV_X1 U5896 ( .A(n7723), .ZN(n9620) );
  NAND2_X1 U5897 ( .A1(n5984), .A2(n5966), .ZN(n8056) );
  NAND2_X1 U5898 ( .A1(n4977), .A2(n4980), .ZN(n5913) );
  NAND2_X1 U5899 ( .A1(n5841), .A2(n5308), .ZN(n5822) );
  NAND2_X1 U5900 ( .A1(n5726), .A2(n5725), .ZN(n5729) );
  NAND2_X1 U5901 ( .A1(n5588), .A2(n5587), .ZN(n5592) );
  NAND2_X1 U5902 ( .A1(n5423), .A2(n5422), .ZN(n5490) );
  XNOR2_X1 U5903 ( .A(n5029), .B(n5487), .ZN(n7368) );
  NAND2_X1 U5904 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5029) );
  NOR2_X1 U5905 ( .A1(n8516), .A2(n8515), .ZN(n10276) );
  NOR2_X1 U5906 ( .A1(n10274), .A2(n10273), .ZN(n8515) );
  NAND2_X1 U5907 ( .A1(n4997), .A2(n4998), .ZN(n4996) );
  NAND2_X1 U5908 ( .A1(n5106), .A2(n7056), .ZN(n7062) );
  OR2_X1 U5909 ( .A1(n10620), .A2(n5220), .ZN(n5219) );
  INV_X1 U5910 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5220) );
  INV_X1 U5911 ( .A(n5221), .ZN(n9250) );
  NAND2_X1 U5912 ( .A1(n5271), .A2(n5273), .ZN(n5269) );
  OAI21_X1 U5913 ( .B1(n9663), .B2(n9662), .A(n9661), .ZN(n9668) );
  OAI21_X1 U5914 ( .B1(n5021), .B2(n10305), .A(n5018), .ZN(P1_U3260) );
  INV_X1 U5915 ( .A(n5019), .ZN(n5018) );
  XNOR2_X1 U5916 ( .A(n5022), .B(n9773), .ZN(n5021) );
  OAI21_X1 U5917 ( .B1(n9778), .B2(n10332), .A(n5020), .ZN(n5019) );
  INV_X1 U5918 ( .A(n5162), .ZN(n10364) );
  NOR2_X1 U5919 ( .A1(n7991), .A2(n4993), .ZN(n4992) );
  NAND2_X1 U5920 ( .A1(n10386), .A2(n8662), .ZN(n5233) );
  NAND2_X1 U5921 ( .A1(n8410), .A2(n8413), .ZN(n5036) );
  AND2_X1 U5922 ( .A1(n4900), .A2(n5400), .ZN(n4881) );
  AND2_X1 U5923 ( .A1(n9074), .A2(n4934), .ZN(n4882) );
  AND2_X1 U5924 ( .A1(n9137), .A2(n4895), .ZN(n4883) );
  INV_X1 U5925 ( .A(n6218), .ZN(n5264) );
  AND2_X1 U5926 ( .A1(n6920), .A2(n6919), .ZN(n4884) );
  NOR2_X1 U5927 ( .A1(n5794), .A2(n5793), .ZN(n4885) );
  AND2_X1 U5928 ( .A1(n6343), .A2(n6342), .ZN(n7662) );
  AND3_X1 U5929 ( .A1(n9798), .A2(n10511), .A3(n8620), .ZN(n4886) );
  AND2_X1 U5930 ( .A1(n6931), .A2(n5088), .ZN(n4887) );
  NAND4_X1 U5931 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n7711)
         );
  NAND2_X1 U5932 ( .A1(n6463), .A2(n6462), .ZN(n8000) );
  INV_X1 U5933 ( .A(n8000), .ZN(n5212) );
  AND2_X1 U5934 ( .A1(n6220), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5935 ( .A1(n5632), .A2(n5670), .ZN(n4889) );
  AND2_X1 U5936 ( .A1(n6051), .A2(n5044), .ZN(n4890) );
  AND2_X1 U5937 ( .A1(n4932), .A2(n5885), .ZN(n4891) );
  OR2_X1 U5938 ( .A1(n5459), .A2(n5749), .ZN(n5417) );
  AND2_X1 U5939 ( .A1(n6792), .A2(n6791), .ZN(n4892) );
  INV_X1 U5940 ( .A(n9176), .ZN(n6761) );
  OR2_X1 U5941 ( .A1(n5063), .A2(n5718), .ZN(n4893) );
  NAND2_X1 U5942 ( .A1(n5866), .A2(SI_17_), .ZN(n5887) );
  INV_X1 U5943 ( .A(n5887), .ZN(n5141) );
  NAND2_X1 U5944 ( .A1(n4947), .A2(n5144), .ZN(n5139) );
  INV_X1 U5945 ( .A(n9079), .ZN(n9164) );
  INV_X1 U5946 ( .A(n7831), .ZN(n4991) );
  OAI211_X1 U5947 ( .C1(n6819), .C2(n5086), .A(n5085), .B(n5088), .ZN(n7528)
         );
  INV_X1 U5948 ( .A(n5539), .ZN(n5639) );
  INV_X1 U5949 ( .A(n4873), .ZN(n5901) );
  OR2_X1 U5950 ( .A1(n5600), .A2(n5599), .ZN(n4894) );
  NAND2_X1 U5951 ( .A1(n5633), .A2(n5632), .ZN(n5656) );
  NAND2_X1 U5952 ( .A1(n9242), .A2(n6795), .ZN(n4895) );
  NAND2_X1 U5953 ( .A1(n5979), .A2(n5980), .ZN(n4896) );
  NAND2_X1 U5954 ( .A1(n10289), .A2(n7284), .ZN(n5536) );
  NAND2_X1 U5955 ( .A1(n9622), .A2(n7746), .ZN(n7721) );
  AND2_X1 U5956 ( .A1(n9622), .A2(n7746), .ZN(n5159) );
  AND2_X1 U5957 ( .A1(n6164), .A2(n5412), .ZN(n5437) );
  AND2_X1 U5958 ( .A1(n6794), .A2(n7887), .ZN(n4897) );
  NAND2_X1 U5959 ( .A1(n7615), .A2(n7614), .ZN(n7036) );
  AND2_X1 U5960 ( .A1(n6870), .A2(n6869), .ZN(n9175) );
  AND2_X1 U5961 ( .A1(n9855), .A2(n5166), .ZN(n4898) );
  OR2_X1 U5962 ( .A1(n9143), .A2(n9237), .ZN(n4899) );
  AND2_X1 U5963 ( .A1(n6190), .A2(n6118), .ZN(n4900) );
  AND2_X1 U5964 ( .A1(n7069), .A2(n5473), .ZN(n5686) );
  AND2_X1 U5965 ( .A1(n7004), .A2(n7003), .ZN(n9001) );
  INV_X1 U5966 ( .A(n9001), .ZN(n5081) );
  NAND2_X1 U5967 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4901) );
  NAND2_X1 U5968 ( .A1(n9846), .A2(n5116), .ZN(n4902) );
  AND2_X1 U5969 ( .A1(n8990), .A2(n5218), .ZN(n4903) );
  AND2_X1 U5970 ( .A1(n10629), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4904) );
  OR2_X2 U5971 ( .A1(n5468), .A2(n10192), .ZN(n5992) );
  NAND2_X1 U5972 ( .A1(n9862), .A2(n9542), .ZN(n9843) );
  AND2_X1 U5973 ( .A1(n4881), .A2(n6074), .ZN(n4905) );
  OR2_X1 U5974 ( .A1(n8604), .A2(n5195), .ZN(n4906) );
  AND2_X1 U5975 ( .A1(n9332), .A2(n9331), .ZN(n4907) );
  INV_X1 U5976 ( .A(n6934), .ZN(n5349) );
  AND2_X1 U5977 ( .A1(n5283), .A2(n5405), .ZN(n5700) );
  OR2_X1 U5978 ( .A1(n10548), .A2(n10513), .ZN(n4908) );
  AND4_X1 U5979 ( .A1(n5094), .A2(n5013), .A3(n6338), .A4(n5012), .ZN(n4909)
         );
  OR3_X1 U5980 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_IR_REG_1__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U5981 ( .A1(n4968), .A2(n9594), .ZN(n9861) );
  XNOR2_X1 U5982 ( .A(n9176), .B(n8392), .ZN(n8952) );
  NAND2_X1 U5983 ( .A1(n6657), .A2(n6656), .ZN(n9193) );
  NAND2_X1 U5984 ( .A1(n5592), .A2(n5591), .ZN(n5606) );
  OR2_X1 U5985 ( .A1(n9193), .A2(n9015), .ZN(n7004) );
  AND3_X1 U5986 ( .A1(n9500), .A2(n9608), .A3(n9654), .ZN(n4911) );
  AND4_X1 U5987 ( .A1(n6222), .A2(n6490), .A3(n6747), .A4(n6206), .ZN(n4912)
         );
  INV_X1 U5988 ( .A(n9586), .ZN(n5184) );
  AND2_X1 U5989 ( .A1(n5067), .A2(n4897), .ZN(n4913) );
  NAND2_X1 U5990 ( .A1(n5556), .A2(n5555), .ZN(n5588) );
  NAND2_X1 U5991 ( .A1(n5437), .A2(n5438), .ZN(n5433) );
  NAND2_X1 U5992 ( .A1(n5405), .A2(n5404), .ZN(n5635) );
  NAND2_X1 U5993 ( .A1(n6672), .A2(n6671), .ZN(n9187) );
  NAND2_X1 U5994 ( .A1(n5734), .A2(n5733), .ZN(n9439) );
  NAND2_X1 U5995 ( .A1(n8586), .A2(n9416), .ZN(n9895) );
  INV_X1 U5996 ( .A(n5387), .ZN(n5009) );
  NOR2_X1 U5997 ( .A1(n5388), .A2(n8532), .ZN(n5387) );
  NAND2_X1 U5998 ( .A1(n7662), .A2(n8561), .ZN(n4914) );
  INV_X1 U5999 ( .A(n9434), .ZN(n5177) );
  AND2_X1 U6000 ( .A1(n9603), .A2(n9539), .ZN(n9477) );
  OR2_X1 U6001 ( .A1(n5265), .A2(n5062), .ZN(n4915) );
  NAND2_X1 U6002 ( .A1(n5806), .A2(n5805), .ZN(n10146) );
  NAND2_X1 U6003 ( .A1(n8591), .A2(n8590), .ZN(n10063) );
  AND2_X1 U6004 ( .A1(n5039), .A2(n9311), .ZN(n4916) );
  AND2_X1 U6005 ( .A1(n9560), .A2(n9434), .ZN(n9518) );
  INV_X1 U6006 ( .A(n9518), .ZN(n8037) );
  AND2_X1 U6007 ( .A1(n9575), .A2(n9548), .ZN(n10019) );
  AND2_X1 U6008 ( .A1(n9564), .A2(n9566), .ZN(n9522) );
  AND2_X1 U6009 ( .A1(n8596), .A2(n8594), .ZN(n4917) );
  AND2_X1 U6010 ( .A1(n5015), .A2(n5014), .ZN(n4918) );
  OR2_X1 U6011 ( .A1(n4881), .A2(n5270), .ZN(n4919) );
  INV_X1 U6012 ( .A(n5204), .ZN(n5203) );
  NOR2_X1 U6013 ( .A1(n9477), .A2(n5205), .ZN(n5204) );
  NAND2_X1 U6014 ( .A1(n7877), .A2(n7987), .ZN(n4920) );
  NOR2_X1 U6015 ( .A1(n9175), .A2(n5360), .ZN(n5358) );
  INV_X1 U6016 ( .A(n9175), .ZN(n8937) );
  INV_X1 U6017 ( .A(n4999), .ZN(n4997) );
  NAND2_X1 U6018 ( .A1(n5000), .A2(n5379), .ZN(n4999) );
  AND2_X1 U6019 ( .A1(n5059), .A2(n4915), .ZN(n4921) );
  OR2_X1 U6020 ( .A1(n5156), .A2(n9532), .ZN(n4922) );
  NOR2_X1 U6021 ( .A1(n9237), .A2(n9124), .ZN(n4923) );
  NOR2_X1 U6022 ( .A1(n9197), .A2(n8724), .ZN(n4924) );
  NAND2_X1 U6023 ( .A1(n9305), .A2(n9303), .ZN(n9300) );
  OR2_X1 U6024 ( .A1(n8663), .A2(n10462), .ZN(n4925) );
  INV_X1 U6025 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5438) );
  AND2_X1 U6026 ( .A1(n6951), .A2(n6952), .ZN(n7872) );
  INV_X1 U6027 ( .A(n7872), .ZN(n5067) );
  AND2_X1 U6028 ( .A1(n5699), .A2(n7221), .ZN(n4926) );
  OR2_X1 U6029 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4927) );
  INV_X1 U6030 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6204) );
  OR2_X1 U6031 ( .A1(n7020), .A2(n5359), .ZN(n4928) );
  OR2_X1 U6032 ( .A1(n10084), .A2(n9863), .ZN(n4929) );
  OR2_X1 U6033 ( .A1(n9435), .A2(n5177), .ZN(n5176) );
  OR2_X1 U6034 ( .A1(n5046), .A2(n5043), .ZN(n4930) );
  AND2_X1 U6035 ( .A1(n5431), .A2(n5114), .ZN(n4931) );
  INV_X1 U6036 ( .A(n6336), .ZN(n5373) );
  OR2_X1 U6037 ( .A1(n5886), .A2(n5288), .ZN(n4932) );
  NAND2_X1 U6038 ( .A1(n9483), .A2(n9649), .ZN(n9532) );
  INV_X1 U6039 ( .A(n9532), .ZN(n8620) );
  NAND2_X1 U6040 ( .A1(n5165), .A2(n5163), .ZN(n9825) );
  OR2_X1 U6041 ( .A1(n8093), .A2(n8781), .ZN(n6901) );
  INV_X1 U6042 ( .A(n6901), .ZN(n5345) );
  NAND2_X1 U6043 ( .A1(n9222), .A2(n8678), .ZN(n4934) );
  AND2_X1 U6044 ( .A1(n6980), .A2(n6981), .ZN(n9091) );
  INV_X1 U6045 ( .A(n9091), .ZN(n5339) );
  AND2_X1 U6046 ( .A1(n5747), .A2(n5150), .ZN(n4935) );
  INV_X1 U6047 ( .A(n5670), .ZN(n5325) );
  AND2_X1 U6048 ( .A1(n5038), .A2(n4896), .ZN(n4936) );
  AND2_X1 U6049 ( .A1(n6336), .A2(n8666), .ZN(n4937) );
  AND2_X1 U6050 ( .A1(n6212), .A2(n5263), .ZN(n4938) );
  AND2_X1 U6051 ( .A1(n5271), .A2(n4919), .ZN(n4939) );
  INV_X1 U6052 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5012) );
  AND2_X1 U6053 ( .A1(n5405), .A2(n5282), .ZN(n4940) );
  INV_X1 U6054 ( .A(n6309), .ZN(n6550) );
  INV_X1 U6055 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6205) );
  INV_X1 U6056 ( .A(n5956), .ZN(n5143) );
  OR2_X1 U6057 ( .A1(n7399), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4941) );
  INV_X1 U6058 ( .A(n9641), .ZN(n5183) );
  AND2_X1 U6059 ( .A1(n7345), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6060 ( .A1(n9339), .A2(n5858), .ZN(n9347) );
  AND2_X1 U6061 ( .A1(n5819), .A2(n5799), .ZN(n4943) );
  NAND2_X1 U6062 ( .A1(n6104), .A2(n6103), .ZN(n10074) );
  INV_X1 U6063 ( .A(n10074), .ZN(n5120) );
  NAND2_X1 U6064 ( .A1(n9972), .A2(n5196), .ZN(n9953) );
  AND2_X1 U6065 ( .A1(n4978), .A2(n4976), .ZN(n4944) );
  INV_X1 U6066 ( .A(n5402), .ZN(n5144) );
  INV_X1 U6067 ( .A(n5115), .ZN(n9948) );
  NOR2_X1 U6068 ( .A1(n9964), .A2(n10117), .ZN(n5115) );
  AND2_X1 U6069 ( .A1(n4979), .A2(n4976), .ZN(n4945) );
  NAND2_X1 U6070 ( .A1(n5008), .A2(n5006), .ZN(n8675) );
  OR2_X1 U6071 ( .A1(n4979), .A2(n4976), .ZN(n4946) );
  NAND2_X1 U6072 ( .A1(n5939), .A2(n5142), .ZN(n4947) );
  NAND2_X1 U6073 ( .A1(n6081), .A2(n6080), .ZN(n10079) );
  OR2_X1 U6074 ( .A1(n8972), .A2(n8743), .ZN(n4948) );
  AND2_X1 U6075 ( .A1(n7067), .A2(n7068), .ZN(n4949) );
  AND2_X1 U6076 ( .A1(n7816), .A2(n6794), .ZN(n4950) );
  AND2_X1 U6077 ( .A1(n9958), .A2(n9583), .ZN(n4951) );
  AND2_X1 U6078 ( .A1(n5366), .A2(n8640), .ZN(n4952) );
  XNOR2_X1 U6079 ( .A(n5441), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U6080 ( .A(n6237), .B(n6236), .ZN(n8057) );
  INV_X1 U6081 ( .A(n8057), .ZN(n5392) );
  AND2_X1 U6082 ( .A1(n6259), .A2(n8057), .ZN(n6751) );
  AND2_X1 U6083 ( .A1(n7510), .A2(n6333), .ZN(n4953) );
  OR2_X1 U6084 ( .A1(n10445), .A2(n5226), .ZN(n5228) );
  NOR2_X1 U6085 ( .A1(n5703), .A2(n5210), .ZN(n6164) );
  AND2_X1 U6086 ( .A1(n7801), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4954) );
  NOR2_X2 U6087 ( .A1(n6768), .A2(n6753), .ZN(n10375) );
  NAND2_X1 U6088 ( .A1(n7722), .A2(n7723), .ZN(n6163) );
  NAND2_X1 U6089 ( .A1(n5256), .A2(n6784), .ZN(n7526) );
  NAND2_X1 U6090 ( .A1(n5601), .A2(n4894), .ZN(n7641) );
  AND2_X1 U6091 ( .A1(n9569), .A2(n9567), .ZN(n9523) );
  INV_X1 U6092 ( .A(n9523), .ZN(n8353) );
  INV_X1 U6093 ( .A(n8413), .ZN(n5031) );
  NAND2_X1 U6094 ( .A1(n6226), .A2(n6225), .ZN(n9242) );
  INV_X1 U6095 ( .A(n9242), .ZN(n5229) );
  OAI21_X1 U6096 ( .B1(n5266), .B2(n5062), .A(n4921), .ZN(n8061) );
  INV_X1 U6097 ( .A(n7994), .ZN(n4990) );
  AND2_X1 U6098 ( .A1(n7781), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U6099 ( .A1(n5200), .A2(n5201), .ZN(n8036) );
  NAND2_X1 U6100 ( .A1(n6455), .A2(n7831), .ZN(n7833) );
  INV_X1 U6101 ( .A(n6213), .ZN(n6727) );
  NAND2_X1 U6102 ( .A1(n6821), .A2(n6934), .ZN(n7670) );
  NAND2_X1 U6103 ( .A1(n8075), .A2(n5126), .ZN(n5129) );
  NAND2_X1 U6104 ( .A1(n7897), .A2(n7952), .ZN(n7963) );
  INV_X1 U6105 ( .A(n7963), .ZN(n5213) );
  INV_X1 U6106 ( .A(n5395), .ZN(n5265) );
  AND2_X1 U6107 ( .A1(n6007), .A2(n6006), .ZN(n4956) );
  NAND2_X1 U6108 ( .A1(n8663), .A2(n10462), .ZN(n5088) );
  NAND2_X1 U6109 ( .A1(n5335), .A2(n5334), .ZN(n6820) );
  INV_X1 U6110 ( .A(n6820), .ZN(n7570) );
  INV_X1 U6111 ( .A(n5315), .ZN(n5314) );
  NOR2_X1 U6112 ( .A1(n6078), .A2(n5316), .ZN(n5315) );
  XNOR2_X1 U6113 ( .A(n5417), .B(n5415), .ZN(n7315) );
  INV_X1 U6114 ( .A(n7634), .ZN(n5227) );
  NAND4_X1 U6115 ( .A1(n6270), .A2(n6269), .A3(n6268), .A4(n6267), .ZN(n7424)
         );
  NAND2_X1 U6116 ( .A1(n6321), .A2(n8666), .ZN(n7510) );
  NAND2_X1 U6117 ( .A1(n10377), .A2(n10376), .ZN(n8665) );
  INV_X1 U6118 ( .A(n10548), .ZN(n5122) );
  NAND2_X1 U6119 ( .A1(n6316), .A2(n6315), .ZN(n10451) );
  INV_X1 U6120 ( .A(n10451), .ZN(n6780) );
  INV_X1 U6121 ( .A(n5480), .ZN(n7722) );
  NAND2_X1 U6122 ( .A1(n10319), .A2(n7718), .ZN(n10305) );
  INV_X1 U6123 ( .A(n7662), .ZN(n8570) );
  INV_X1 U6124 ( .A(n8993), .ZN(n9106) );
  NAND2_X1 U6125 ( .A1(n6241), .A2(n6240), .ZN(n8993) );
  INV_X1 U6126 ( .A(n6750), .ZN(n6756) );
  INV_X1 U6127 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4965) );
  INV_X1 U6128 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5300) );
  INV_X1 U6129 ( .A(n5324), .ZN(n5323) );
  INV_X1 U6130 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U6131 ( .A1(n8695), .A2(n6670), .ZN(n5367) );
  NAND2_X1 U6132 ( .A1(n8704), .A2(n6528), .ZN(n8716) );
  NAND2_X1 U6133 ( .A1(n8725), .A2(n6655), .ZN(n8696) );
  NAND2_X1 U6134 ( .A1(n4959), .A2(n10019), .ZN(n9453) );
  NAND3_X1 U6135 ( .A1(n9449), .A2(n9448), .A3(n4960), .ZN(n4959) );
  OR2_X1 U6136 ( .A1(n9451), .A2(n9450), .ZN(n4960) );
  NAND2_X1 U6137 ( .A1(n9473), .A2(n9837), .ZN(n4962) );
  OAI21_X1 U6138 ( .B1(n5196), .B2(n4906), .A(n5197), .ZN(n5194) );
  NAND2_X1 U6139 ( .A1(n4933), .A2(n4983), .ZN(n10165) );
  INV_X1 U6140 ( .A(n5655), .ZN(n5327) );
  OAI21_X1 U6141 ( .B1(n5326), .B2(n5325), .A(n5696), .ZN(n5324) );
  OAI21_X1 U6142 ( .B1(n8614), .B2(n5203), .A(n8617), .ZN(n5148) );
  OAI21_X2 U6143 ( .B1(n9936), .B2(n8606), .A(n8605), .ZN(n9911) );
  NOR2_X2 U6144 ( .A1(n9792), .A2(n9791), .ZN(n9794) );
  NAND2_X1 U6145 ( .A1(n4969), .A2(n5181), .ZN(n4968) );
  NAND2_X1 U6146 ( .A1(n8586), .A2(n5179), .ZN(n4969) );
  NAND2_X2 U6147 ( .A1(n4971), .A2(n5821), .ZN(n5841) );
  NAND2_X1 U6148 ( .A1(n5889), .A2(n5887), .ZN(n4977) );
  OAI21_X1 U6149 ( .B1(n5889), .B2(n5888), .A(n5887), .ZN(n5940) );
  NAND3_X1 U6150 ( .A1(n8650), .A2(n8649), .A3(n4948), .ZN(P2_U3216) );
  NAND2_X1 U6151 ( .A1(n8652), .A2(n8651), .ZN(n6639) );
  NAND2_X1 U6152 ( .A1(n8687), .A2(n5394), .ZN(n8744) );
  NAND2_X1 U6153 ( .A1(n4989), .A2(n6455), .ZN(n4988) );
  NAND2_X1 U6154 ( .A1(n8643), .A2(n4995), .ZN(n4994) );
  OAI211_X1 U6155 ( .C1(n8643), .C2(n4996), .A(n6775), .B(n4994), .ZN(P2_U3222) );
  NAND2_X1 U6156 ( .A1(n8535), .A2(n5006), .ZN(n5003) );
  INV_X1 U6157 ( .A(n8535), .ZN(n5010) );
  NAND2_X1 U6158 ( .A1(n5003), .A2(n5004), .ZN(n6588) );
  NAND3_X1 U6159 ( .A1(n5094), .A2(n5013), .A3(n6338), .ZN(n6227) );
  NAND3_X1 U6160 ( .A1(n5094), .A2(n6338), .A3(n6204), .ZN(n6473) );
  NAND2_X1 U6161 ( .A1(n5037), .A2(n4936), .ZN(n9319) );
  NAND2_X1 U6162 ( .A1(n9312), .A2(n9311), .ZN(n9367) );
  OR2_X1 U6163 ( .A1(n5954), .A2(n5393), .ZN(n5038) );
  OAI21_X2 U6164 ( .B1(n5042), .B2(n4930), .A(n4890), .ZN(n9357) );
  INV_X1 U6165 ( .A(n6025), .ZN(n5047) );
  NAND2_X1 U6166 ( .A1(n5049), .A2(n5054), .ZN(n7063) );
  NAND2_X1 U6167 ( .A1(n9330), .A2(n4905), .ZN(n5049) );
  OAI21_X1 U6168 ( .B1(n9330), .B2(n5052), .A(n5050), .ZN(n6196) );
  INV_X1 U6169 ( .A(n5054), .ZN(n5052) );
  NAND2_X1 U6170 ( .A1(n9330), .A2(n6074), .ZN(n5053) );
  OAI21_X1 U6171 ( .B1(n9330), .B2(n4907), .A(n6074), .ZN(n9399) );
  NAND2_X1 U6172 ( .A1(n5064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5457) );
  NAND4_X1 U6173 ( .A1(n5451), .A2(n5283), .A3(n5065), .A4(n5405), .ZN(n5064)
         );
  NAND2_X1 U6174 ( .A1(n5068), .A2(n5066), .ZN(n6826) );
  NAND2_X1 U6175 ( .A1(n7683), .A2(n5069), .ZN(n5068) );
  OAI21_X1 U6176 ( .B1(n7683), .B2(n6947), .A(n5069), .ZN(n7869) );
  NAND2_X1 U6177 ( .A1(n5073), .A2(n5074), .ZN(n5072) );
  AND2_X1 U6178 ( .A1(n5075), .A2(n9091), .ZN(n5073) );
  AND2_X2 U6179 ( .A1(n6213), .A2(n4938), .ZN(n6218) );
  AND2_X2 U6180 ( .A1(n5361), .A2(n5362), .ZN(n6213) );
  NAND3_X1 U6181 ( .A1(n5084), .A2(n6930), .A3(n5083), .ZN(n7628) );
  NAND3_X1 U6182 ( .A1(n6819), .A2(n6820), .A3(n4887), .ZN(n5084) );
  NAND2_X1 U6183 ( .A1(n6819), .A2(n6820), .ZN(n7569) );
  NAND3_X1 U6184 ( .A1(n4880), .A2(n6283), .A3(n7613), .ZN(n6817) );
  AND2_X1 U6185 ( .A1(n6816), .A2(n6817), .ZN(n7615) );
  NOR2_X2 U6186 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6275) );
  NAND3_X1 U6187 ( .A1(n6978), .A2(n9091), .A3(n6979), .ZN(n5092) );
  NAND3_X1 U6188 ( .A1(n5094), .A2(n5093), .A3(n6338), .ZN(n5363) );
  AND4_X2 U6189 ( .A1(n6202), .A2(n6199), .A3(n6200), .A4(n6201), .ZN(n5094)
         );
  NAND2_X1 U6190 ( .A1(n8663), .A2(n7515), .ZN(n5099) );
  NAND3_X1 U6191 ( .A1(n5108), .A2(n7054), .A3(n5107), .ZN(n5106) );
  NAND3_X1 U6192 ( .A1(n5113), .A2(n6946), .A3(n7884), .ZN(n5112) );
  NAND3_X1 U6193 ( .A1(n6943), .A2(n6942), .A3(n7691), .ZN(n5113) );
  NOR2_X2 U6194 ( .A1(n7769), .A2(n7773), .ZN(n10423) );
  NAND3_X1 U6195 ( .A1(n10364), .A2(n7736), .A3(n7742), .ZN(n7769) );
  NAND2_X2 U6196 ( .A1(n4931), .A2(n5432), .ZN(n5162) );
  NAND2_X2 U6197 ( .A1(n4872), .A2(n6220), .ZN(n5548) );
  NOR2_X2 U6198 ( .A1(n10112), .A2(n9948), .ZN(n9930) );
  NOR2_X2 U6199 ( .A1(n10001), .A2(n10128), .ZN(n9982) );
  NAND2_X1 U6200 ( .A1(n9846), .A2(n9831), .ZN(n9828) );
  OR2_X2 U6201 ( .A1(n9828), .A2(n10074), .ZN(n9811) );
  INV_X1 U6202 ( .A(n5129), .ZN(n8398) );
  INV_X1 U6203 ( .A(n5888), .ZN(n5145) );
  NAND2_X1 U6204 ( .A1(n5748), .A2(n5747), .ZN(n5772) );
  NAND2_X1 U6205 ( .A1(n5748), .A2(n4935), .ZN(n5791) );
  NAND2_X1 U6206 ( .A1(n5155), .A2(n7226), .ZN(n5590) );
  MUX2_X1 U6207 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6220), .Z(n5589) );
  NAND3_X1 U6208 ( .A1(n9541), .A2(n9532), .A3(n10511), .ZN(n5157) );
  INV_X1 U6209 ( .A(n7748), .ZN(n9511) );
  XNOR2_X2 U6210 ( .A(n9679), .B(n5162), .ZN(n7748) );
  NAND2_X1 U6211 ( .A1(n10020), .A2(n5170), .ZN(n5169) );
  INV_X1 U6212 ( .A(n8376), .ZN(n5178) );
  NAND2_X1 U6213 ( .A1(n10037), .A2(n5187), .ZN(n8041) );
  NAND2_X1 U6214 ( .A1(n9559), .A2(n9554), .ZN(n10037) );
  AND2_X1 U6215 ( .A1(n8040), .A2(n10033), .ZN(n5187) );
  NAND2_X1 U6216 ( .A1(n7858), .A2(n9629), .ZN(n10478) );
  AOI21_X1 U6217 ( .B1(n8402), .B2(n9523), .A(n9444), .ZN(n8403) );
  NAND2_X1 U6218 ( .A1(n9926), .A2(n9413), .ZN(n9916) );
  NAND2_X1 U6219 ( .A1(n7764), .A2(n9510), .ZN(n7856) );
  NAND2_X1 U6220 ( .A1(n8403), .A2(n8404), .ZN(n8584) );
  NAND2_X1 U6221 ( .A1(n10510), .A2(n9632), .ZN(n7918) );
  NAND2_X1 U6222 ( .A1(n7856), .A2(n9624), .ZN(n10415) );
  NAND2_X1 U6223 ( .A1(n5211), .A2(n5290), .ZN(n5209) );
  INV_X2 U6224 ( .A(n5613), .ZN(n5405) );
  NAND2_X1 U6225 ( .A1(n7913), .A2(n5190), .ZN(n5189) );
  INV_X1 U6226 ( .A(n10505), .ZN(n5192) );
  NOR2_X2 U6227 ( .A1(n5703), .A2(n5209), .ZN(n5459) );
  NAND3_X1 U6228 ( .A1(n5405), .A2(n5283), .A3(n5444), .ZN(n5703) );
  NOR2_X2 U6229 ( .A1(n7895), .A2(n7900), .ZN(n7897) );
  OAI21_X1 U6230 ( .B1(n5221), .B2(n10619), .A(n5219), .ZN(P2_U3551) );
  INV_X1 U6231 ( .A(n10445), .ZN(n5224) );
  NAND2_X1 U6232 ( .A1(n5224), .A2(n5223), .ZN(n7822) );
  NOR2_X2 U6233 ( .A1(n4899), .A2(n9231), .ZN(n9118) );
  NAND2_X1 U6234 ( .A1(n6916), .A2(n5233), .ZN(n5334) );
  NAND3_X1 U6235 ( .A1(n7036), .A2(n6911), .A3(n5233), .ZN(n5335) );
  NAND2_X1 U6236 ( .A1(n9090), .A2(n4882), .ZN(n5246) );
  INV_X1 U6237 ( .A(n5247), .ZN(n9089) );
  AOI21_X2 U6238 ( .B1(n7816), .B2(n4913), .A(n5248), .ZN(n7962) );
  CLKBUF_X1 U6239 ( .A(n6288), .Z(n5251) );
  NAND2_X1 U6240 ( .A1(n8442), .A2(n4883), .ZN(n5253) );
  INV_X1 U6241 ( .A(n5254), .ZN(n8441) );
  NAND2_X1 U6242 ( .A1(n10442), .A2(n10447), .ZN(n5256) );
  NAND2_X1 U6243 ( .A1(n5256), .A2(n5255), .ZN(n6786) );
  AND2_X1 U6244 ( .A1(n4914), .A2(n6784), .ZN(n5255) );
  OAI21_X2 U6245 ( .B1(n9042), .B2(n5258), .A(n5257), .ZN(n8999) );
  NOR2_X1 U6246 ( .A1(n9202), .A2(n6800), .ZN(n9021) );
  NAND2_X1 U6247 ( .A1(n5262), .A2(n4892), .ZN(n7688) );
  NAND3_X1 U6248 ( .A1(n7937), .A2(n5691), .A3(n7978), .ZN(n5266) );
  NAND2_X1 U6249 ( .A1(n6096), .A2(n4939), .ZN(n5268) );
  OAI211_X1 U6250 ( .C1(n6096), .C2(n5269), .A(n5268), .B(n4949), .ZN(P1_U3212) );
  NAND2_X1 U6251 ( .A1(n5274), .A2(n5276), .ZN(n5693) );
  NAND3_X1 U6252 ( .A1(n5601), .A2(n4894), .A3(n5275), .ZN(n5274) );
  NAND3_X1 U6253 ( .A1(n5601), .A2(n4894), .A3(n5281), .ZN(n5280) );
  NOR2_X2 U6254 ( .A1(n5284), .A2(n4927), .ZN(n5283) );
  NAND2_X1 U6255 ( .A1(n5293), .A2(n5292), .ZN(n5611) );
  NAND3_X1 U6256 ( .A1(n5556), .A2(n5555), .A3(n5591), .ZN(n5293) );
  INV_X1 U6257 ( .A(n5587), .ZN(n5294) );
  NAND3_X1 U6258 ( .A1(n5423), .A2(n5422), .A3(n5488), .ZN(n5492) );
  NAND2_X2 U6259 ( .A1(n5298), .A2(n5296), .ZN(n5532) );
  NAND3_X1 U6260 ( .A1(n5297), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5296) );
  INV_X2 U6261 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5297) );
  NAND3_X1 U6262 ( .A1(n5301), .A2(n5300), .A3(n5299), .ZN(n5298) );
  NAND2_X1 U6263 ( .A1(n5842), .A2(n5310), .ZN(n5865) );
  NAND2_X1 U6264 ( .A1(n6035), .A2(n5315), .ZN(n5311) );
  NAND2_X1 U6265 ( .A1(n5963), .A2(n5962), .ZN(n5984) );
  NAND2_X1 U6266 ( .A1(n6027), .A2(n6026), .ZN(n6031) );
  NAND2_X1 U6267 ( .A1(n7036), .A2(n6911), .ZN(n6909) );
  NAND2_X1 U6268 ( .A1(n9063), .A2(n7044), .ZN(n9071) );
  NAND3_X1 U6269 ( .A1(n5342), .A2(n6964), .A3(n5340), .ZN(n8437) );
  NAND3_X1 U6270 ( .A1(n6965), .A2(n8087), .A3(n5343), .ZN(n5342) );
  NAND2_X1 U6271 ( .A1(n5347), .A2(n5350), .ZN(n7683) );
  NAND2_X1 U6272 ( .A1(n6821), .A2(n5348), .ZN(n5347) );
  NAND2_X1 U6273 ( .A1(n6861), .A2(n5354), .ZN(n5353) );
  NAND2_X1 U6274 ( .A1(n5353), .A2(n5356), .ZN(n6888) );
  INV_X1 U6275 ( .A(n6210), .ZN(n5361) );
  INV_X1 U6276 ( .A(n5363), .ZN(n5362) );
  NAND2_X2 U6277 ( .A1(n6252), .A2(n6251), .ZN(n6297) );
  AND2_X2 U6278 ( .A1(n6287), .A2(n7422), .ZN(n10377) );
  NAND2_X1 U6279 ( .A1(n7423), .A2(n7421), .ZN(n7422) );
  XNOR2_X1 U6280 ( .A(n6284), .B(n6286), .ZN(n7421) );
  NAND2_X1 U6281 ( .A1(n8695), .A2(n5368), .ZN(n5365) );
  NAND2_X1 U6282 ( .A1(n5365), .A2(n4952), .ZN(n8643) );
  NAND2_X1 U6283 ( .A1(n6321), .A2(n4937), .ZN(n5372) );
  NAND3_X1 U6284 ( .A1(n5372), .A2(n8576), .A3(n5371), .ZN(n8563) );
  OR2_X1 U6285 ( .A1(n6333), .A2(n5373), .ZN(n5371) );
  INV_X1 U6286 ( .A(n6717), .ZN(n5380) );
  NAND2_X1 U6287 ( .A1(n4909), .A2(n5383), .ZN(n5382) );
  INV_X1 U6288 ( .A(n6231), .ZN(n6239) );
  INV_X1 U6289 ( .A(n8533), .ZN(n5388) );
  NAND2_X1 U6290 ( .A1(n8568), .A2(n5389), .ZN(n7583) );
  NAND2_X1 U6291 ( .A1(n7583), .A2(n6386), .ZN(n6404) );
  NAND2_X1 U6292 ( .A1(n7073), .A2(n6444), .ZN(n6455) );
  NAND2_X1 U6293 ( .A1(n8478), .A2(n5390), .ZN(n7073) );
  NAND2_X1 U6294 ( .A1(n6750), .A2(n5392), .ZN(n5391) );
  INV_X1 U6295 ( .A(n9187), .ZN(n6848) );
  NOR2_X2 U6296 ( .A1(n9204), .A2(n9048), .ZN(n9034) );
  NAND2_X1 U6297 ( .A1(n9047), .A2(n9052), .ZN(n9048) );
  NAND2_X1 U6298 ( .A1(n7736), .A2(n7713), .ZN(n7737) );
  INV_X1 U6299 ( .A(n10192), .ZN(n5467) );
  NAND2_X1 U6300 ( .A1(n8373), .A2(n8352), .ZN(n8355) );
  INV_X1 U6301 ( .A(n6831), .ZN(n9116) );
  NAND2_X1 U6302 ( .A1(n5419), .A2(SI_1_), .ZN(n5423) );
  OR2_X1 U6303 ( .A1(n4868), .A2(n7613), .ZN(n6777) );
  INV_X4 U6304 ( .A(n5992), .ZN(n6182) );
  BUF_X2 U6305 ( .A(n6221), .Z(n6289) );
  AND2_X1 U6306 ( .A1(n6221), .A2(n6220), .ZN(n6279) );
  XNOR2_X1 U6307 ( .A(n5772), .B(n5771), .ZN(n5770) );
  NOR2_X2 U6308 ( .A1(n9092), .A2(n9216), .ZN(n9047) );
  OAI211_X1 U6309 ( .C1(n5532), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n5418), .B(
        SI_0_), .ZN(n5421) );
  NAND2_X1 U6310 ( .A1(n5532), .A2(n8319), .ZN(n5418) );
  OAI21_X1 U6311 ( .B1(n8950), .B2(n9245), .A(n6850), .ZN(n6858) );
  INV_X4 U6312 ( .A(n6325), .ZN(n6280) );
  OAI211_X2 U6313 ( .C1(n4872), .C2(n7413), .A(n5538), .B(n5537), .ZN(n7773)
         );
  OR2_X1 U6314 ( .A1(n5536), .A2(n7287), .ZN(n5537) );
  NOR2_X2 U6315 ( .A1(n9794), .A2(n8619), .ZN(n8621) );
  CLKBUF_X1 U6316 ( .A(n6763), .Z(n9275) );
  NAND2_X1 U6317 ( .A1(n6763), .A2(n6841), .ZN(n6221) );
  AND2_X1 U6318 ( .A1(n9369), .A2(n5953), .ZN(n5393) );
  NOR2_X1 U6319 ( .A1(n8751), .A2(n6618), .ZN(n5394) );
  INV_X1 U6320 ( .A(n9887), .ZN(n9894) );
  AND2_X1 U6321 ( .A1(n5695), .A2(n5694), .ZN(n5395) );
  NOR2_X1 U6322 ( .A1(n7938), .A2(n7939), .ZN(n5396) );
  INV_X1 U6323 ( .A(n8330), .ZN(n7056) );
  INV_X1 U6324 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6215) );
  OR2_X1 U6325 ( .A1(n6309), .A2(n7621), .ZN(n5398) );
  AND2_X1 U6326 ( .A1(n9121), .A2(n8718), .ZN(n5399) );
  INV_X1 U6327 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U6328 ( .A1(n6220), .A2(P1_U3084), .ZN(n10204) );
  INV_X1 U6329 ( .A(SI_15_), .ZN(n7202) );
  INV_X1 U6330 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5749) );
  AND2_X1 U6331 ( .A1(n5535), .A2(n5550), .ZN(n5401) );
  INV_X4 U6332 ( .A(n6220), .ZN(n7285) );
  INV_X2 U6333 ( .A(n5532), .ZN(n6220) );
  XOR2_X1 U6334 ( .A(n7283), .B(n7282), .Z(n8313) );
  OR2_X1 U6335 ( .A1(n7294), .A2(n10287), .ZN(n10210) );
  INV_X1 U6336 ( .A(n10019), .ZN(n8596) );
  NAND2_X2 U6337 ( .A1(n7864), .A2(n10531), .ZN(n10536) );
  OR2_X1 U6338 ( .A1(n7448), .A2(n6170), .ZN(n9410) );
  INV_X1 U6339 ( .A(n9410), .ZN(n9381) );
  NOR2_X1 U6340 ( .A1(n5938), .A2(n5937), .ZN(n5402) );
  NAND2_X1 U6341 ( .A1(n6545), .A2(n6544), .ZN(n6796) );
  INV_X1 U6342 ( .A(n9941), .ZN(n8585) );
  INV_X1 U6343 ( .A(n9837), .ZN(n8615) );
  INV_X1 U6344 ( .A(n10135), .ZN(n8630) );
  INV_X1 U6345 ( .A(n9047), .ZN(n9076) );
  INV_X1 U6346 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7179) );
  INV_X1 U6347 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7270) );
  INV_X1 U6348 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U6349 ( .A1(n9170), .A2(n8932), .ZN(n6887) );
  INV_X1 U6350 ( .A(n6617), .ZN(n6618) );
  OR4_X1 U6351 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6723) );
  INV_X1 U6352 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5413) );
  INV_X1 U6353 ( .A(SI_19_), .ZN(n7205) );
  INV_X1 U6354 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6243) );
  INV_X1 U6355 ( .A(n7076), .ZN(n6443) );
  INV_X1 U6356 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6532) );
  INV_X1 U6357 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7988) );
  INV_X1 U6358 ( .A(n9041), .ZN(n6833) );
  AND2_X1 U6359 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6327) );
  INV_X1 U6360 ( .A(n9359), .ZN(n6051) );
  INV_X1 U6361 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5640) );
  AND2_X1 U6362 ( .A1(n10066), .A2(n8618), .ZN(n8619) );
  OR2_X1 U6363 ( .A1(n5877), .A2(n9351), .ZN(n5898) );
  INV_X1 U6364 ( .A(SI_29_), .ZN(n7187) );
  INV_X1 U6365 ( .A(SI_16_), .ZN(n7108) );
  INV_X1 U6366 ( .A(SI_4_), .ZN(n7231) );
  NAND2_X1 U6367 ( .A1(n6626), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6643) );
  OR2_X1 U6368 ( .A1(n6517), .A2(n6243), .ZN(n6533) );
  NAND2_X1 U6369 ( .A1(n6639), .A2(n6638), .ZN(n6654) );
  OR2_X1 U6370 ( .A1(n6643), .A2(n7179), .ZN(n6658) );
  INV_X1 U6371 ( .A(n6311), .ZN(n6535) );
  OR2_X1 U6372 ( .A1(n6478), .A2(n7177), .ZN(n6496) );
  INV_X1 U6373 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7514) );
  NAND2_X2 U6374 ( .A1(n6289), .A2(n7285), .ZN(n6288) );
  AND2_X1 U6375 ( .A1(n9204), .A2(n9057), .ZN(n6800) );
  NAND2_X1 U6376 ( .A1(n6558), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6576) );
  INV_X1 U6377 ( .A(n8990), .ZN(n9005) );
  NAND2_X1 U6378 ( .A1(n6246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6247) );
  INV_X1 U6379 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6229) );
  INV_X1 U6380 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5807) );
  INV_X1 U6381 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5778) );
  INV_X1 U6382 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5735) );
  AND2_X1 U6383 ( .A1(n5827), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5847) );
  AND2_X1 U6384 ( .A1(n5943), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5969) );
  INV_X1 U6385 ( .A(n8627), .ZN(n8628) );
  OAI21_X1 U6386 ( .B1(n10475), .B2(n10476), .A(n7852), .ZN(n10505) );
  AOI21_X1 U6387 ( .B1(n5480), .B2(n7715), .A(n10494), .ZN(n5478) );
  INV_X1 U6388 ( .A(SI_20_), .ZN(n7111) );
  OR2_X1 U6389 ( .A1(n5843), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5844) );
  INV_X1 U6390 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8646) );
  INV_X1 U6391 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8655) );
  INV_X1 U6392 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8700) );
  XNOR2_X1 U6393 ( .A(n6654), .B(n6652), .ZN(n8723) );
  INV_X1 U6394 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8792) );
  OR2_X1 U6395 ( .A1(n7564), .A2(n6745), .ZN(n6768) );
  AND2_X1 U6396 ( .A1(n6627), .A2(n6610), .ZN(n9050) );
  INV_X1 U6397 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8102) );
  OR2_X1 U6398 ( .A1(n8175), .A2(n8174), .ZN(n10651) );
  NOR2_X1 U6399 ( .A1(n9193), .A2(n6801), .ZN(n6802) );
  AND2_X1 U6400 ( .A1(n8947), .A2(n6849), .ZN(n6850) );
  INV_X1 U6401 ( .A(n10611), .ZN(n10403) );
  INV_X1 U6402 ( .A(n7515), .ZN(n10462) );
  NOR2_X1 U6403 ( .A1(n6740), .A2(n10243), .ZN(n7564) );
  NOR2_X1 U6404 ( .A1(n5808), .A2(n5807), .ZN(n5827) );
  OR2_X1 U6405 ( .A1(n5779), .A2(n5778), .ZN(n5808) );
  INV_X1 U6406 ( .A(n9675), .ZN(n8064) );
  OR2_X1 U6407 ( .A1(n9349), .A2(n9348), .ZN(n5885) );
  NAND2_X1 U6408 ( .A1(n6186), .A2(n7718), .ZN(n9405) );
  INV_X1 U6409 ( .A(n5839), .ZN(n5835) );
  AND2_X1 U6410 ( .A1(n6136), .A2(n6135), .ZN(n9817) );
  INV_X1 U6411 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8027) );
  INV_X1 U6412 ( .A(n6181), .ZN(n7718) );
  INV_X1 U6413 ( .A(n9977), .ZN(n9973) );
  AND2_X1 U6414 ( .A1(n9592), .A2(n9641), .ZN(n9901) );
  NAND2_X1 U6415 ( .A1(n7718), .A2(n7717), .ZN(n10482) );
  AND2_X1 U6416 ( .A1(n5934), .A2(n5892), .ZN(n5932) );
  XNOR2_X1 U6417 ( .A(n7515), .B(n6325), .ZN(n8575) );
  AND2_X1 U6418 ( .A1(n7420), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8740) );
  OR2_X1 U6419 ( .A1(n8969), .A2(n4870), .ZN(n6697) );
  OR2_X1 U6420 ( .A1(n6258), .A2(n6257), .ZN(n6795) );
  INV_X1 U6421 ( .A(n10651), .ZN(n10653) );
  INV_X1 U6422 ( .A(n10636), .ZN(n10654) );
  NAND2_X1 U6423 ( .A1(n8313), .A2(n8175), .ZN(n8155) );
  INV_X1 U6424 ( .A(n7046), .ZN(n9055) );
  INV_X1 U6425 ( .A(n8345), .ZN(n9124) );
  AND2_X1 U6426 ( .A1(n8150), .A2(n9275), .ZN(n10448) );
  INV_X1 U6427 ( .A(n9164), .ZN(n10466) );
  NAND2_X1 U6428 ( .A1(n6742), .A2(n6741), .ZN(n7560) );
  NAND2_X1 U6429 ( .A1(n6769), .A2(n6751), .ZN(n10611) );
  AND2_X1 U6430 ( .A1(n9059), .A2(n9058), .ZN(n9213) );
  INV_X1 U6431 ( .A(n10596), .ZN(n10391) );
  INV_X1 U6432 ( .A(n9245), .ZN(n10617) );
  XNOR2_X1 U6433 ( .A(n6732), .B(P2_IR_REG_25__SCAN_IN), .ZN(n10241) );
  AND2_X1 U6434 ( .A1(n6445), .A2(n6428), .ZN(n8789) );
  AND2_X1 U6435 ( .A1(n6087), .A2(n6086), .ZN(n9818) );
  AND2_X1 U6436 ( .A1(n5850), .A2(n5849), .ZN(n10016) );
  INV_X1 U6437 ( .A(n9776), .ZN(n10324) );
  AND2_X1 U6438 ( .A1(n10319), .A2(n6181), .ZN(n10311) );
  INV_X1 U6439 ( .A(n9477), .ZN(n9815) );
  INV_X1 U6440 ( .A(n10482), .ZN(n10515) );
  AND2_X1 U6441 ( .A1(n10015), .A2(n10014), .ZN(n10138) );
  NAND2_X1 U6442 ( .A1(n7431), .A2(n6171), .ZN(n10531) );
  AND2_X1 U6443 ( .A1(n10536), .A2(n7707), .ZN(n10526) );
  AOI21_X1 U6444 ( .B1(n7294), .B2(n6150), .A(n7296), .ZN(n7436) );
  OR2_X1 U6445 ( .A1(n9485), .A2(n9659), .ZN(n10550) );
  AND2_X1 U6446 ( .A1(n10519), .A2(n10550), .ZN(n10162) );
  AND2_X1 U6447 ( .A1(n10285), .A2(n7434), .ZN(n7437) );
  INV_X1 U6448 ( .A(n10287), .ZN(n7431) );
  AND2_X1 U6449 ( .A1(n5893), .A2(n5874), .ZN(n9751) );
  AND2_X1 U6450 ( .A1(n5774), .A2(n5752), .ZN(n7781) );
  INV_X1 U6451 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8483) );
  NOR2_X1 U6452 ( .A1(n10270), .A2(n10269), .ZN(n8510) );
  AND2_X1 U6453 ( .A1(n8158), .A2(n8157), .ZN(n10655) );
  AND2_X1 U6454 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  INV_X1 U6455 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7494) );
  INV_X1 U6456 ( .A(n6759), .ZN(n8743) );
  INV_X1 U6457 ( .A(n10375), .ZN(n8759) );
  AND4_X1 U6458 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n8326)
         );
  NAND2_X1 U6459 ( .A1(n8155), .A2(n9275), .ZN(n10650) );
  AND2_X1 U6460 ( .A1(n8957), .A2(n8956), .ZN(n9179) );
  AND2_X1 U6461 ( .A1(n9088), .A2(n9087), .ZN(n9225) );
  AND2_X1 U6462 ( .A1(n7566), .A2(n10470), .ZN(n9079) );
  INV_X1 U6463 ( .A(n10620), .ZN(n10619) );
  OR2_X1 U6464 ( .A1(n6857), .A2(n6856), .ZN(n10621) );
  NAND2_X1 U6465 ( .A1(n10244), .A2(n10243), .ZN(n10344) );
  AND2_X1 U6466 ( .A1(n7055), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10347) );
  INV_X1 U6467 ( .A(n9402), .ZN(n9395) );
  INV_X1 U6468 ( .A(n9408), .ZN(n9388) );
  INV_X1 U6469 ( .A(n9818), .ZN(n9844) );
  INV_X1 U6470 ( .A(n10417), .ZN(n10516) );
  OR2_X1 U6471 ( .A1(P1_U3083), .A2(n7313), .ZN(n9776) );
  INV_X1 U6472 ( .A(n10315), .ZN(n10332) );
  NAND2_X1 U6473 ( .A1(n10536), .A2(n10499), .ZN(n10012) );
  AND2_X2 U6474 ( .A1(n7437), .A2(n7436), .ZN(n10591) );
  INV_X1 U6475 ( .A(n10591), .ZN(n10589) );
  OR2_X1 U6476 ( .A1(n10156), .A2(n10155), .ZN(n10183) );
  AND3_X1 U6477 ( .A1(n10569), .A2(n10568), .A3(n10567), .ZN(n10572) );
  AND2_X2 U6478 ( .A1(n7437), .A2(n7704), .ZN(n10595) );
  INV_X1 U6479 ( .A(n5468), .ZN(n8582) );
  NOR2_X1 U6480 ( .A1(n8511), .A2(n8510), .ZN(n10272) );
  NAND3_X1 U6481 ( .A1(n5430), .A2(n5558), .A3(n5403), .ZN(n5613) );
  NOR2_X1 U6482 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5409) );
  NOR2_X1 U6483 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5408) );
  NAND4_X1 U6484 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n5411)
         );
  NAND3_X1 U6485 ( .A1(n5445), .A2(n5869), .A3(n5872), .ZN(n5410) );
  NAND2_X1 U6486 ( .A1(n5434), .A2(n5413), .ZN(n5414) );
  NAND2_X1 U6487 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5416) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8314) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8319) );
  INV_X1 U6490 ( .A(n5421), .ZN(n5419) );
  INV_X1 U6491 ( .A(SI_1_), .ZN(n5420) );
  NAND2_X1 U6492 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  MUX2_X1 U6493 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5532), .Z(n5488) );
  INV_X1 U6494 ( .A(n5428), .ZN(n5425) );
  MUX2_X1 U6495 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5532), .Z(n5424) );
  NAND2_X1 U6496 ( .A1(n5424), .A2(SI_2_), .ZN(n5530) );
  OAI21_X1 U6497 ( .B1(n5424), .B2(SI_2_), .A(n5530), .ZN(n5426) );
  NAND2_X1 U6498 ( .A1(n5425), .A2(n5426), .ZN(n5429) );
  INV_X1 U6499 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U6500 ( .A1(n5429), .A2(n5531), .ZN(n7302) );
  OR2_X1 U6501 ( .A1(n5430), .A2(n5749), .ZN(n5560) );
  INV_X1 U6502 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5526) );
  XNOR2_X1 U6503 ( .A(n5560), .B(n5526), .ZN(n7466) );
  OR2_X1 U6504 ( .A1(n4872), .A2(n7466), .ZN(n5431) );
  NAND2_X1 U6505 ( .A1(n5433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5435) );
  OR2_X1 U6506 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  INV_X1 U6507 ( .A(n5437), .ZN(n6167) );
  NAND2_X1 U6508 ( .A1(n6167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5439) );
  INV_X1 U6509 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5443) );
  NAND4_X1 U6510 ( .A1(n5445), .A2(n5444), .A3(n5872), .A4(n5443), .ZN(n5450)
         );
  INV_X1 U6511 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5448) );
  INV_X1 U6512 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5447) );
  INV_X1 U6513 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5446) );
  NAND4_X1 U6514 ( .A1(n5869), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n5449)
         );
  NOR2_X1 U6515 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6516 ( .A1(n5457), .A2(n5452), .ZN(n5453) );
  AND2_X2 U6517 ( .A1(n7069), .A2(n7715), .ZN(n5539) );
  NOR3_X1 U6518 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6519 ( .A1(n5459), .A2(n5458), .ZN(n5465) );
  XNOR2_X2 U6520 ( .A(n5460), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6521 ( .A1(n4867), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5472) );
  NAND2_X2 U6522 ( .A1(n5467), .A2(n5468), .ZN(n5973) );
  NAND2_X1 U6523 ( .A1(n4869), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6524 ( .A1(n4875), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6525 ( .A1(n4874), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5469) );
  NAND4_X2 U6526 ( .A1(n5472), .A2(n5471), .A3(n5470), .A4(n5469), .ZN(n9679)
         );
  INV_X1 U6527 ( .A(n7715), .ZN(n5473) );
  INV_X2 U6528 ( .A(n5686), .ZN(n5907) );
  NAND2_X1 U6529 ( .A1(n9679), .A2(n5713), .ZN(n5474) );
  NAND2_X1 U6530 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X2 U6531 ( .A(n5477), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10494) );
  AND2_X2 U6532 ( .A1(n10519), .A2(n7715), .ZN(n5508) );
  XNOR2_X1 U6533 ( .A(n5479), .B(n5508), .ZN(n5520) );
  NAND2_X1 U6534 ( .A1(n5480), .A2(n7706), .ZN(n5481) );
  NAND2_X1 U6535 ( .A1(n9679), .A2(n6112), .ZN(n5482) );
  OAI21_X1 U6536 ( .B1(n10364), .B2(n5907), .A(n5482), .ZN(n5518) );
  XNOR2_X1 U6537 ( .A(n5520), .B(n5518), .ZN(n7476) );
  NAND2_X1 U6538 ( .A1(n5566), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6539 ( .A1(n4867), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6540 ( .A1(n4876), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6541 ( .A1(n5568), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6542 ( .A1(n7711), .A2(n6000), .ZN(n5497) );
  INV_X1 U6543 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5487) );
  INV_X1 U6544 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U6545 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U6546 ( .A1(n5492), .A2(n5491), .ZN(n7298) );
  INV_X1 U6547 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5493) );
  OR2_X1 U6548 ( .A1(n4878), .A2(n5493), .ZN(n5494) );
  NAND2_X1 U6549 ( .A1(n4879), .A2(n5539), .ZN(n5496) );
  NAND2_X1 U6550 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  XNOR2_X1 U6551 ( .A(n5498), .B(n5618), .ZN(n5514) );
  NAND2_X1 U6552 ( .A1(n9680), .A2(n6112), .ZN(n5500) );
  NAND2_X1 U6553 ( .A1(n4879), .A2(n5713), .ZN(n5499) );
  NAND2_X1 U6554 ( .A1(n5500), .A2(n5499), .ZN(n5515) );
  NAND2_X1 U6555 ( .A1(n5514), .A2(n5515), .ZN(n5513) );
  INV_X1 U6556 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U6557 ( .A1(n4867), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U6558 ( .A1(n4869), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6559 ( .A1(n4875), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U6560 ( .A1(n4873), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5501) );
  NAND4_X1 U6561 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n7714)
         );
  NAND2_X1 U6562 ( .A1(n7714), .A2(n5713), .ZN(n5507) );
  NAND2_X1 U6563 ( .A1(n7284), .A2(SI_0_), .ZN(n5505) );
  XNOR2_X1 U6564 ( .A(n5505), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10208) );
  MUX2_X1 U6565 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10208), .S(n4872), .Z(n7741)
         );
  NAND2_X1 U6566 ( .A1(n7741), .A2(n5539), .ZN(n5506) );
  OAI211_X1 U6567 ( .C1(n10293), .C2(n7069), .A(n5507), .B(n5506), .ZN(n7455)
         );
  OR2_X1 U6568 ( .A1(n7455), .A2(n5508), .ZN(n5512) );
  NAND2_X1 U6569 ( .A1(n7714), .A2(n6112), .ZN(n5511) );
  NAND2_X1 U6570 ( .A1(n7741), .A2(n5713), .ZN(n5510) );
  INV_X1 U6571 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10294) );
  OR2_X1 U6572 ( .A1(n7069), .A2(n10294), .ZN(n5509) );
  AND3_X1 U6573 ( .A1(n5511), .A2(n5510), .A3(n5509), .ZN(n7456) );
  NAND2_X1 U6574 ( .A1(n7456), .A2(n7455), .ZN(n7454) );
  NAND2_X1 U6575 ( .A1(n5512), .A2(n7454), .ZN(n7444) );
  NAND2_X1 U6576 ( .A1(n5513), .A2(n7444), .ZN(n5517) );
  INV_X1 U6577 ( .A(n5514), .ZN(n7446) );
  INV_X1 U6578 ( .A(n5515), .ZN(n7443) );
  NAND2_X1 U6579 ( .A1(n7446), .A2(n7443), .ZN(n5516) );
  NAND2_X1 U6580 ( .A1(n5517), .A2(n5516), .ZN(n7475) );
  NAND2_X1 U6581 ( .A1(n7476), .A2(n7475), .ZN(n5522) );
  INV_X1 U6582 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U6583 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  NAND2_X1 U6584 ( .A1(n5522), .A2(n5521), .ZN(n7484) );
  AOI22_X1 U6585 ( .A1(n6182), .A2(P1_REG1_REG_3__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_3__SCAN_IN), .ZN(n5525) );
  INV_X1 U6586 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5523) );
  AOI22_X1 U6587 ( .A1(n4869), .A2(n5523), .B1(n4874), .B2(
        P1_REG0_REG_3__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6588 ( .A1(n5560), .A2(n5526), .ZN(n5527) );
  NAND2_X1 U6589 ( .A1(n5527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5529) );
  INV_X1 U6590 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5528) );
  XNOR2_X1 U6591 ( .A(n5529), .B(n5528), .ZN(n7413) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7288) );
  OR2_X1 U6593 ( .A1(n5548), .A2(n7288), .ZN(n5538) );
  NAND2_X1 U6594 ( .A1(n5531), .A2(n5530), .ZN(n5549) );
  MUX2_X1 U6595 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5532), .Z(n5534) );
  INV_X1 U6596 ( .A(n5534), .ZN(n5533) );
  INV_X1 U6597 ( .A(SI_3_), .ZN(n7234) );
  NAND2_X1 U6598 ( .A1(n5533), .A2(n7234), .ZN(n5535) );
  NAND2_X1 U6599 ( .A1(n5534), .A2(SI_3_), .ZN(n5550) );
  XNOR2_X1 U6600 ( .A(n5549), .B(n5401), .ZN(n7287) );
  OAI22_X1 U6601 ( .A1(n10418), .A2(n5907), .B1(n7846), .B2(n5639), .ZN(n5540)
         );
  XNOR2_X1 U6602 ( .A(n5540), .B(n5508), .ZN(n5545) );
  OR2_X1 U6603 ( .A1(n10418), .A2(n6141), .ZN(n5542) );
  NAND2_X1 U6604 ( .A1(n7773), .A2(n5713), .ZN(n5541) );
  NAND2_X1 U6605 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  XNOR2_X1 U6606 ( .A(n5545), .B(n5543), .ZN(n7483) );
  NAND2_X1 U6607 ( .A1(n7484), .A2(n7483), .ZN(n5547) );
  INV_X1 U6608 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U6609 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  NAND2_X1 U6610 ( .A1(n5547), .A2(n5546), .ZN(n7504) );
  INV_X1 U6611 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8321) );
  OR2_X1 U6612 ( .A1(n5548), .A2(n8321), .ZN(n5565) );
  NAND2_X1 U6613 ( .A1(n5549), .A2(n5401), .ZN(n5551) );
  NAND2_X1 U6614 ( .A1(n5551), .A2(n5550), .ZN(n5556) );
  NAND2_X1 U6615 ( .A1(n5552), .A2(SI_4_), .ZN(n5587) );
  INV_X1 U6616 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U6617 ( .A1(n5553), .A2(n7231), .ZN(n5554) );
  OR2_X1 U6618 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  NAND2_X1 U6619 ( .A1(n5588), .A2(n5557), .ZN(n7293) );
  OR2_X1 U6620 ( .A1(n5536), .A2(n7293), .ZN(n5564) );
  OR2_X1 U6621 ( .A1(n5558), .A2(n5749), .ZN(n5559) );
  AND2_X1 U6622 ( .A1(n5560), .A2(n5559), .ZN(n5562) );
  INV_X1 U6623 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6624 ( .A1(n5562), .A2(n5561), .ZN(n5585) );
  OAI21_X1 U6625 ( .B1(n5562), .B2(n5561), .A(n5585), .ZN(n7329) );
  OR2_X1 U6626 ( .A1(n4872), .A2(n7329), .ZN(n5563) );
  INV_X1 U6627 ( .A(n10434), .ZN(n7857) );
  NAND2_X1 U6628 ( .A1(n7857), .A2(n5539), .ZN(n5574) );
  NAND2_X1 U6629 ( .A1(n6182), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5572) );
  INV_X1 U6630 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U6631 ( .A(n5567), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U6632 ( .A1(n5566), .A2(n7503), .ZN(n5571) );
  NAND2_X1 U6633 ( .A1(n4875), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6634 ( .A1(n4873), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5569) );
  NAND4_X1 U6635 ( .A1(n5572), .A2(n5571), .A3(n5570), .A4(n5569), .ZN(n9678)
         );
  NAND2_X1 U6636 ( .A1(n9678), .A2(n5713), .ZN(n5573) );
  NAND2_X1 U6637 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  XNOR2_X1 U6638 ( .A(n5575), .B(n5508), .ZN(n5579) );
  NAND2_X1 U6639 ( .A1(n9678), .A2(n6112), .ZN(n5576) );
  OAI21_X1 U6640 ( .B1(n10434), .B2(n5907), .A(n5576), .ZN(n5577) );
  XNOR2_X1 U6641 ( .A(n5579), .B(n5577), .ZN(n7505) );
  NAND2_X1 U6642 ( .A1(n7504), .A2(n7505), .ZN(n5581) );
  INV_X1 U6643 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U6644 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND2_X1 U6645 ( .A1(n5581), .A2(n5580), .ZN(n5600) );
  AOI22_X1 U6646 ( .A1(n6182), .A2(P1_REG1_REG_5__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n5584) );
  AOI21_X1 U6647 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5582) );
  NOR2_X1 U6648 ( .A1(n5582), .A2(n5602), .ZN(n10492) );
  AOI22_X1 U6649 ( .A1(n4869), .A2(n10492), .B1(n4873), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U6650 ( .A1(n5585), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5586) );
  XNOR2_X1 U6651 ( .A(n5586), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7374) );
  INV_X1 U6652 ( .A(n7374), .ZN(n7286) );
  NAND2_X1 U6653 ( .A1(n5589), .A2(SI_5_), .ZN(n5605) );
  AND2_X1 U6654 ( .A1(n5605), .A2(n5590), .ZN(n5591) );
  OR2_X1 U6655 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  NAND2_X1 U6656 ( .A1(n5606), .A2(n5593), .ZN(n7305) );
  INV_X1 U6657 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8325) );
  OR2_X1 U6658 ( .A1(n5548), .A2(n8325), .ZN(n5594) );
  OAI22_X1 U6659 ( .A1(n10417), .A2(n5907), .B1(n7851), .B2(n5639), .ZN(n5596)
         );
  XNOR2_X1 U6660 ( .A(n5596), .B(n5508), .ZN(n5599) );
  NAND2_X1 U6661 ( .A1(n5600), .A2(n5599), .ZN(n7604) );
  OR2_X1 U6662 ( .A1(n10417), .A2(n6141), .ZN(n5598) );
  NAND2_X1 U6663 ( .A1(n10490), .A2(n5713), .ZN(n5597) );
  NAND2_X1 U6664 ( .A1(n5598), .A2(n5597), .ZN(n7606) );
  NAND2_X1 U6665 ( .A1(n7604), .A2(n7606), .ZN(n5601) );
  AOI22_X1 U6666 ( .A1(n6182), .A2(P1_REG1_REG_6__SCAN_IN), .B1(n4876), .B2(
        P1_REG2_REG_6__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6667 ( .A1(n5602), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5641) );
  OAI21_X1 U6668 ( .B1(n5602), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5641), .ZN(
        n10532) );
  INV_X1 U6669 ( .A(n10532), .ZN(n7644) );
  AOI22_X1 U6670 ( .A1(n4869), .A2(n7644), .B1(n4874), .B2(
        P1_REG0_REG_6__SCAN_IN), .ZN(n5603) );
  MUX2_X1 U6671 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7284), .Z(n5607) );
  NAND2_X1 U6672 ( .A1(n5607), .A2(SI_6_), .ZN(n5627) );
  INV_X1 U6673 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U6674 ( .A1(n5608), .A2(n7227), .ZN(n5609) );
  NAND2_X1 U6675 ( .A1(n5611), .A2(n5610), .ZN(n5628) );
  OR2_X1 U6676 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U6677 ( .A1(n5628), .A2(n5612), .ZN(n7290) );
  OR2_X1 U6678 ( .A1(n7290), .A2(n5536), .ZN(n5616) );
  NAND2_X1 U6679 ( .A1(n5613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5614) );
  XNOR2_X1 U6680 ( .A(n5614), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7345) );
  AOI22_X1 U6681 ( .A1(n5915), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5914), .B2(
        n7345), .ZN(n5615) );
  NAND2_X1 U6682 ( .A1(n5616), .A2(n5615), .ZN(n7862) );
  NAND2_X1 U6683 ( .A1(n7862), .A2(n5539), .ZN(n5617) );
  OAI21_X1 U6684 ( .B1(n10483), .B2(n5907), .A(n5617), .ZN(n5619) );
  XNOR2_X1 U6685 ( .A(n5619), .B(n6090), .ZN(n5622) );
  OR2_X1 U6686 ( .A1(n10483), .A2(n6141), .ZN(n5621) );
  NAND2_X1 U6687 ( .A1(n7862), .A2(n5713), .ZN(n5620) );
  NAND2_X1 U6688 ( .A1(n5621), .A2(n5620), .ZN(n5623) );
  XNOR2_X1 U6689 ( .A(n5622), .B(n5623), .ZN(n7642) );
  INV_X1 U6690 ( .A(n5622), .ZN(n5625) );
  INV_X1 U6691 ( .A(n5623), .ZN(n5624) );
  NAND2_X1 U6692 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  MUX2_X1 U6693 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7284), .Z(n5629) );
  NAND2_X1 U6694 ( .A1(n5629), .A2(SI_7_), .ZN(n5655) );
  INV_X1 U6695 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U6696 ( .A1(n5630), .A2(n7220), .ZN(n5631) );
  OR2_X1 U6697 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  NAND2_X1 U6698 ( .A1(n5656), .A2(n5634), .ZN(n7300) );
  OR2_X1 U6699 ( .A1(n7300), .A2(n5536), .ZN(n5638) );
  NAND2_X1 U6700 ( .A1(n5635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5636) );
  XNOR2_X1 U6701 ( .A(n5636), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7399) );
  AOI22_X1 U6702 ( .A1(n5915), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5914), .B2(
        n7399), .ZN(n5637) );
  NAND2_X1 U6703 ( .A1(n5638), .A2(n5637), .ZN(n10548) );
  NAND2_X1 U6704 ( .A1(n10548), .A2(n5539), .ZN(n5648) );
  NOR2_X1 U6705 ( .A1(n5641), .A2(n5640), .ZN(n5659) );
  AND2_X1 U6706 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NOR2_X1 U6707 ( .A1(n5659), .A2(n5642), .ZN(n7904) );
  NAND2_X1 U6708 ( .A1(n4869), .A2(n7904), .ZN(n5646) );
  NAND2_X1 U6709 ( .A1(n6182), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6710 ( .A1(n4877), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U6711 ( .A1(n4874), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5643) );
  NAND4_X1 U6712 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(n10513)
         );
  NAND2_X1 U6713 ( .A1(n10513), .A2(n6000), .ZN(n5647) );
  NAND2_X1 U6714 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  XNOR2_X1 U6715 ( .A(n5649), .B(n6090), .ZN(n5651) );
  AND2_X1 U6716 ( .A1(n10513), .A2(n6112), .ZN(n5650) );
  AOI21_X1 U6717 ( .B1(n10548), .B2(n6000), .A(n5650), .ZN(n5652) );
  XNOR2_X1 U6718 ( .A(n5651), .B(n5652), .ZN(n7907) );
  INV_X1 U6719 ( .A(n5651), .ZN(n5653) );
  NAND2_X1 U6720 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  MUX2_X1 U6721 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7285), .Z(n5667) );
  XNOR2_X1 U6722 ( .A(n5667), .B(SI_8_), .ZN(n5671) );
  XNOR2_X1 U6723 ( .A(n5671), .B(n5672), .ZN(n7306) );
  NAND2_X1 U6724 ( .A1(n7306), .A2(n9493), .ZN(n5658) );
  OR2_X1 U6725 ( .A1(n4940), .A2(n5749), .ZN(n5674) );
  XNOR2_X1 U6726 ( .A(n5674), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U6727 ( .A1(n5915), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5914), .B2(
        n7400), .ZN(n5657) );
  AOI22_X1 U6728 ( .A1(n6182), .A2(P1_REG1_REG_8__SCAN_IN), .B1(n4876), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U6729 ( .A1(n5659), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5679) );
  OR2_X1 U6730 ( .A1(n5659), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5660) );
  AND2_X1 U6731 ( .A1(n5679), .A2(n5660), .ZN(n10042) );
  AOI22_X1 U6732 ( .A1(n5566), .A2(n10042), .B1(n4873), .B2(
        P1_REG0_REG_8__SCAN_IN), .ZN(n5661) );
  NOR2_X1 U6733 ( .A1(n7919), .A2(n6141), .ZN(n5663) );
  AOI21_X1 U6734 ( .B1(n10560), .B2(n6000), .A(n5663), .ZN(n5692) );
  NAND2_X1 U6735 ( .A1(n5693), .A2(n5692), .ZN(n7977) );
  NAND2_X1 U6736 ( .A1(n10560), .A2(n5539), .ZN(n5665) );
  OR2_X1 U6737 ( .A1(n7919), .A2(n5907), .ZN(n5664) );
  NAND2_X1 U6738 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X1 U6739 ( .A(n5666), .B(n6090), .ZN(n7980) );
  INV_X1 U6740 ( .A(n5667), .ZN(n5669) );
  INV_X1 U6741 ( .A(SI_8_), .ZN(n5668) );
  NAND2_X1 U6742 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  MUX2_X1 U6743 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7284), .Z(n5698) );
  XNOR2_X1 U6744 ( .A(n5698), .B(n7221), .ZN(n5696) );
  XNOR2_X1 U6745 ( .A(n5697), .B(n5696), .ZN(n7309) );
  NAND2_X1 U6746 ( .A1(n7309), .A2(n9493), .ZN(n5678) );
  INV_X1 U6747 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6748 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  NAND2_X1 U6749 ( .A1(n5675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U6750 ( .A(n5676), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7545) );
  AOI22_X1 U6751 ( .A1(n5915), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5914), .B2(
        n7545), .ZN(n5677) );
  NAND2_X1 U6752 ( .A1(n5678), .A2(n5677), .ZN(n8034) );
  NAND2_X1 U6753 ( .A1(n8034), .A2(n5539), .ZN(n5688) );
  NAND2_X1 U6754 ( .A1(n5679), .A2(n7394), .ZN(n5680) );
  AND2_X1 U6755 ( .A1(n5707), .A2(n5680), .ZN(n7941) );
  NAND2_X1 U6756 ( .A1(n5566), .A2(n7941), .ZN(n5685) );
  NAND2_X1 U6757 ( .A1(n6182), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U6758 ( .A1(n4875), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6759 ( .A1(n4873), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6760 ( .A1(n10039), .A2(n6000), .ZN(n5687) );
  NAND2_X1 U6761 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  XNOR2_X1 U6762 ( .A(n5689), .B(n5508), .ZN(n5695) );
  AND2_X1 U6763 ( .A1(n10039), .A2(n6112), .ZN(n5690) );
  AOI21_X1 U6764 ( .B1(n8034), .B2(n6000), .A(n5690), .ZN(n5694) );
  XNOR2_X1 U6765 ( .A(n5695), .B(n5694), .ZN(n7939) );
  INV_X1 U6766 ( .A(n7939), .ZN(n5691) );
  INV_X1 U6767 ( .A(n5698), .ZN(n5699) );
  MUX2_X1 U6768 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7284), .Z(n5722) );
  XNOR2_X1 U6769 ( .A(n5722), .B(n5723), .ZN(n5720) );
  XNOR2_X1 U6770 ( .A(n5721), .B(n5720), .ZN(n7354) );
  NAND2_X1 U6771 ( .A1(n7354), .A2(n9493), .ZN(n5706) );
  NOR2_X1 U6772 ( .A1(n5700), .A2(n5749), .ZN(n5701) );
  MUX2_X1 U6773 ( .A(n5749), .B(n5701), .S(P1_IR_REG_10__SCAN_IN), .Z(n5702)
         );
  INV_X1 U6774 ( .A(n5702), .ZN(n5704) );
  AND2_X1 U6775 ( .A1(n5704), .A2(n5703), .ZN(n10312) );
  AOI22_X1 U6776 ( .A1(n5915), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5914), .B2(
        n10312), .ZN(n5705) );
  NAND2_X1 U6777 ( .A1(n8109), .A2(n5539), .ZN(n5715) );
  NAND2_X1 U6778 ( .A1(n5707), .A2(n8027), .ZN(n5708) );
  AND2_X1 U6779 ( .A1(n5736), .A2(n5708), .ZN(n8047) );
  NAND2_X1 U6780 ( .A1(n4869), .A2(n8047), .ZN(n5712) );
  NAND2_X1 U6781 ( .A1(n6182), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6782 ( .A1(n4877), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6783 ( .A1(n4874), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5709) );
  NAND4_X1 U6784 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n9675)
         );
  NAND2_X1 U6785 ( .A1(n9675), .A2(n5713), .ZN(n5714) );
  NAND2_X1 U6786 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  XNOR2_X1 U6787 ( .A(n5716), .B(n6090), .ZN(n5718) );
  AND2_X1 U6788 ( .A1(n9675), .A2(n6112), .ZN(n5717) );
  AOI21_X1 U6789 ( .B1(n8109), .B2(n6000), .A(n5717), .ZN(n8025) );
  INV_X1 U6790 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U6791 ( .A1(n5721), .A2(n5720), .ZN(n5726) );
  INV_X1 U6792 ( .A(n5722), .ZN(n5724) );
  NAND2_X1 U6793 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  MUX2_X1 U6794 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7284), .Z(n5727) );
  NAND2_X1 U6795 ( .A1(n5727), .A2(SI_11_), .ZN(n5747) );
  OAI21_X1 U6796 ( .B1(n5727), .B2(SI_11_), .A(n5747), .ZN(n5730) );
  NAND2_X1 U6797 ( .A1(n5729), .A2(n5730), .ZN(n5731) );
  NAND2_X1 U6798 ( .A1(n5748), .A2(n5731), .ZN(n7383) );
  OR2_X1 U6799 ( .A1(n7383), .A2(n5536), .ZN(n5734) );
  NAND2_X1 U6800 ( .A1(n5703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5732) );
  XNOR2_X1 U6801 ( .A(n5732), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U6802 ( .A1(n5915), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5914), .B2(
        n10325), .ZN(n5733) );
  NAND2_X1 U6803 ( .A1(n9439), .A2(n5539), .ZN(n5741) );
  AOI22_X1 U6804 ( .A1(n6182), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n4876), .B2(
        P1_REG2_REG_11__SCAN_IN), .ZN(n5739) );
  AND2_X1 U6805 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  NOR2_X1 U6806 ( .A1(n5755), .A2(n5737), .ZN(n8078) );
  AOI22_X1 U6807 ( .A1(n4869), .A2(n8078), .B1(n4873), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n5738) );
  OR2_X1 U6808 ( .A1(n8379), .A2(n5907), .ZN(n5740) );
  NAND2_X1 U6809 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  XNOR2_X1 U6810 ( .A(n5742), .B(n5508), .ZN(n5745) );
  NOR2_X1 U6811 ( .A1(n8379), .A2(n6141), .ZN(n5743) );
  AOI21_X1 U6812 ( .B1(n9439), .B2(n6000), .A(n5743), .ZN(n5744) );
  XNOR2_X1 U6813 ( .A(n5745), .B(n5744), .ZN(n8059) );
  OR2_X1 U6814 ( .A1(n5745), .A2(n5744), .ZN(n5746) );
  NAND2_X1 U6815 ( .A1(n8061), .A2(n5746), .ZN(n8282) );
  MUX2_X1 U6816 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7284), .Z(n5771) );
  XNOR2_X1 U6817 ( .A(n5770), .B(SI_12_), .ZN(n7441) );
  NAND2_X1 U6818 ( .A1(n7441), .A2(n9493), .ZN(n5754) );
  NOR2_X1 U6819 ( .A1(n5703), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5801) );
  OR2_X1 U6820 ( .A1(n5801), .A2(n5749), .ZN(n5751) );
  INV_X1 U6821 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U6822 ( .A1(n5751), .A2(n5750), .ZN(n5774) );
  OR2_X1 U6823 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  AOI22_X1 U6824 ( .A1(n5915), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5914), .B2(
        n7781), .ZN(n5753) );
  NAND2_X1 U6825 ( .A1(n10159), .A2(n5539), .ZN(n5762) );
  OR2_X1 U6826 ( .A1(n5755), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6827 ( .A1(n5755), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5779) );
  AND2_X1 U6828 ( .A1(n5756), .A2(n5779), .ZN(n8383) );
  NAND2_X1 U6829 ( .A1(n5566), .A2(n8383), .ZN(n5760) );
  NAND2_X1 U6830 ( .A1(n6182), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U6831 ( .A1(n4875), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U6832 ( .A1(n4873), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5757) );
  NAND4_X1 U6833 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8357)
         );
  NAND2_X1 U6834 ( .A1(n8357), .A2(n6000), .ZN(n5761) );
  NAND2_X1 U6835 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  XNOR2_X1 U6836 ( .A(n5763), .B(n6090), .ZN(n8280) );
  INV_X1 U6837 ( .A(n8280), .ZN(n5766) );
  NAND2_X1 U6838 ( .A1(n10159), .A2(n6000), .ZN(n5765) );
  NAND2_X1 U6839 ( .A1(n8357), .A2(n6112), .ZN(n5764) );
  NAND2_X1 U6840 ( .A1(n5765), .A2(n5764), .ZN(n5767) );
  INV_X1 U6841 ( .A(n5767), .ZN(n8279) );
  NAND2_X1 U6842 ( .A1(n5766), .A2(n8279), .ZN(n5769) );
  AND2_X1 U6843 ( .A1(n8280), .A2(n5767), .ZN(n5768) );
  AOI21_X1 U6844 ( .B1(n8282), .B2(n5769), .A(n5768), .ZN(n8411) );
  NAND2_X1 U6845 ( .A1(n5796), .A2(n5791), .ZN(n5773) );
  MUX2_X1 U6846 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7284), .Z(n5789) );
  XNOR2_X1 U6847 ( .A(n5789), .B(n7215), .ZN(n5793) );
  XNOR2_X1 U6848 ( .A(n5773), .B(n5793), .ZN(n7480) );
  NAND2_X1 U6849 ( .A1(n7480), .A2(n9493), .ZN(n5777) );
  NAND2_X1 U6850 ( .A1(n5774), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  XNOR2_X1 U6851 ( .A(n5775), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7801) );
  AOI22_X1 U6852 ( .A1(n5915), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5914), .B2(
        n7801), .ZN(n5776) );
  NAND2_X1 U6853 ( .A1(n8409), .A2(n5539), .ZN(n5784) );
  AOI22_X1 U6854 ( .A1(n6182), .A2(P1_REG1_REG_13__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_13__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U6855 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  AND2_X1 U6856 ( .A1(n5808), .A2(n5780), .ZN(n8420) );
  AOI22_X1 U6857 ( .A1(n4869), .A2(n8420), .B1(n4874), .B2(
        P1_REG0_REG_13__SCAN_IN), .ZN(n5781) );
  OR2_X1 U6858 ( .A1(n9292), .A2(n5907), .ZN(n5783) );
  NAND2_X1 U6859 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  XNOR2_X1 U6860 ( .A(n5785), .B(n5508), .ZN(n5788) );
  NOR2_X1 U6861 ( .A1(n9292), .A2(n6141), .ZN(n5786) );
  AOI21_X1 U6862 ( .B1(n8409), .B2(n6000), .A(n5786), .ZN(n5787) );
  OR2_X1 U6863 ( .A1(n5788), .A2(n5787), .ZN(n8412) );
  NAND2_X1 U6864 ( .A1(n8411), .A2(n8412), .ZN(n8410) );
  NAND2_X1 U6865 ( .A1(n5788), .A2(n5787), .ZN(n8413) );
  INV_X1 U6866 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U6867 ( .A1(n5790), .A2(n7215), .ZN(n5792) );
  INV_X1 U6868 ( .A(n5792), .ZN(n5794) );
  MUX2_X1 U6869 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7285), .Z(n5797) );
  INV_X1 U6870 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U6871 ( .A1(n5798), .A2(n7114), .ZN(n5799) );
  XNOR2_X1 U6872 ( .A(n5820), .B(n4943), .ZN(n7523) );
  NAND2_X1 U6873 ( .A1(n7523), .A2(n9493), .ZN(n5806) );
  NOR2_X1 U6874 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5800) );
  NAND2_X1 U6875 ( .A1(n5801), .A2(n5800), .ZN(n5803) );
  NAND2_X1 U6876 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  MUX2_X1 U6877 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5802), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5804) );
  AOI22_X1 U6878 ( .A1(n5915), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5914), .B2(
        n8003), .ZN(n5805) );
  NAND2_X1 U6879 ( .A1(n10146), .A2(n5539), .ZN(n5813) );
  AOI22_X1 U6880 ( .A1(n6182), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n5811) );
  AND2_X1 U6881 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  NOR2_X1 U6882 ( .A1(n5827), .A2(n5809), .ZN(n9296) );
  AOI22_X1 U6883 ( .A1(n4869), .A2(n9296), .B1(n4874), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n5810) );
  OR2_X1 U6884 ( .A1(n10017), .A2(n5907), .ZN(n5812) );
  NAND2_X1 U6885 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  XNOR2_X1 U6886 ( .A(n5814), .B(n5508), .ZN(n5817) );
  NAND2_X1 U6887 ( .A1(n10146), .A2(n6000), .ZN(n5816) );
  OR2_X1 U6888 ( .A1(n10017), .A2(n6141), .ZN(n5815) );
  NAND2_X1 U6889 ( .A1(n5816), .A2(n5815), .ZN(n9289) );
  INV_X1 U6890 ( .A(n5817), .ZN(n5818) );
  INV_X1 U6891 ( .A(n5840), .ZN(n5836) );
  MUX2_X1 U6892 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7285), .Z(n5821) );
  NAND2_X1 U6893 ( .A1(n5822), .A2(n7202), .ZN(n5823) );
  NAND2_X1 U6894 ( .A1(n5842), .A2(n5823), .ZN(n7592) );
  OR2_X1 U6895 ( .A1(n7592), .A2(n5536), .ZN(n5826) );
  NAND2_X1 U6896 ( .A1(n5843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5824) );
  XNOR2_X1 U6897 ( .A(n5824), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U6898 ( .A1(n5915), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5914), .B2(
        n9716), .ZN(n5825) );
  NAND2_X2 U6899 ( .A1(n5826), .A2(n5825), .ZN(n10139) );
  NAND2_X1 U6900 ( .A1(n10139), .A2(n5539), .ZN(n5833) );
  AOI22_X1 U6901 ( .A1(n6182), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n5831) );
  NOR2_X1 U6902 ( .A1(n5827), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5828) );
  OR2_X1 U6903 ( .A1(n5847), .A2(n5828), .ZN(n10027) );
  INV_X1 U6904 ( .A(n10027), .ZN(n5829) );
  AOI22_X1 U6905 ( .A1(n5566), .A2(n5829), .B1(n4874), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n5830) );
  OR2_X1 U6906 ( .A1(n9996), .A2(n5907), .ZN(n5832) );
  NAND2_X1 U6907 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  XNOR2_X1 U6908 ( .A(n5834), .B(n6090), .ZN(n5839) );
  NAND2_X1 U6909 ( .A1(n5836), .A2(n5835), .ZN(n8545) );
  NAND2_X1 U6910 ( .A1(n10139), .A2(n6000), .ZN(n5838) );
  OR2_X1 U6911 ( .A1(n9996), .A2(n6141), .ZN(n5837) );
  NAND2_X1 U6912 ( .A1(n5838), .A2(n5837), .ZN(n8547) );
  NAND2_X1 U6913 ( .A1(n5840), .A2(n5839), .ZN(n8542) );
  MUX2_X1 U6914 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7284), .Z(n5862) );
  XNOR2_X1 U6915 ( .A(n5862), .B(SI_16_), .ZN(n5860) );
  XNOR2_X1 U6916 ( .A(n5859), .B(n5860), .ZN(n7681) );
  NAND2_X1 U6917 ( .A1(n7681), .A2(n9493), .ZN(n5846) );
  NAND2_X1 U6918 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U6919 ( .A(n5870), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9738) );
  AOI22_X1 U6920 ( .A1(n5915), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5914), .B2(
        n9738), .ZN(n5845) );
  NAND2_X2 U6921 ( .A1(n5846), .A2(n5845), .ZN(n10135) );
  NAND2_X1 U6922 ( .A1(n10135), .A2(n5539), .ZN(n5852) );
  AOI22_X1 U6923 ( .A1(n6182), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6924 ( .A1(n5847), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5877) );
  OR2_X1 U6925 ( .A1(n5847), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5848) );
  AND2_X1 U6926 ( .A1(n5877), .A2(n5848), .ZN(n10004) );
  AOI22_X1 U6927 ( .A1(n4869), .A2(n10004), .B1(n4874), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5849) );
  OR2_X1 U6928 ( .A1(n10016), .A2(n5907), .ZN(n5851) );
  NAND2_X1 U6929 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U6930 ( .A(n5853), .B(n6090), .ZN(n5855) );
  NOR2_X1 U6931 ( .A1(n10016), .A2(n6141), .ZN(n5854) );
  AOI21_X1 U6932 ( .B1(n10135), .B2(n6000), .A(n5854), .ZN(n5856) );
  XNOR2_X1 U6933 ( .A(n5855), .B(n5856), .ZN(n9340) );
  INV_X1 U6934 ( .A(n5855), .ZN(n5857) );
  NAND2_X1 U6935 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  INV_X1 U6936 ( .A(n5860), .ZN(n5861) );
  INV_X1 U6937 ( .A(n5862), .ZN(n5863) );
  NAND2_X1 U6938 ( .A1(n5863), .A2(n7108), .ZN(n5864) );
  MUX2_X1 U6939 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7285), .Z(n5866) );
  INV_X1 U6940 ( .A(n5866), .ZN(n5867) );
  NAND2_X1 U6941 ( .A1(n5867), .A2(n7113), .ZN(n5868) );
  NAND2_X1 U6942 ( .A1(n5887), .A2(n5868), .ZN(n5888) );
  XNOR2_X1 U6943 ( .A(n5889), .B(n5145), .ZN(n7829) );
  NAND2_X1 U6944 ( .A1(n7829), .A2(n9493), .ZN(n5876) );
  NAND2_X1 U6945 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U6946 ( .A1(n5871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6947 ( .A1(n5873), .A2(n5872), .ZN(n5893) );
  OR2_X1 U6948 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AOI22_X1 U6949 ( .A1(n5915), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5914), .B2(
        n9751), .ZN(n5875) );
  NAND2_X1 U6950 ( .A1(n10128), .A2(n5539), .ZN(n5882) );
  AOI22_X1 U6951 ( .A1(n6182), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n5880) );
  INV_X1 U6952 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U6953 ( .A1(n5877), .A2(n9351), .ZN(n5878) );
  AND2_X1 U6954 ( .A1(n5898), .A2(n5878), .ZN(n9983) );
  AOI22_X1 U6955 ( .A1(n5566), .A2(n9983), .B1(n4873), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5879) );
  OR2_X1 U6956 ( .A1(n9999), .A2(n5907), .ZN(n5881) );
  NAND2_X1 U6957 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  XNOR2_X1 U6958 ( .A(n5883), .B(n5508), .ZN(n9349) );
  NOR2_X1 U6959 ( .A1(n9999), .A2(n6141), .ZN(n5884) );
  AOI21_X1 U6960 ( .B1(n10128), .B2(n6000), .A(n5884), .ZN(n9348) );
  AND2_X1 U6961 ( .A1(n9349), .A2(n9348), .ZN(n5886) );
  MUX2_X1 U6962 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7285), .Z(n5890) );
  NAND2_X1 U6963 ( .A1(n5890), .A2(SI_18_), .ZN(n5934) );
  INV_X1 U6964 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U6965 ( .A1(n5891), .A2(n7107), .ZN(n5892) );
  OR2_X1 U6966 ( .A1(n8531), .A2(n5536), .ZN(n5896) );
  NAND2_X1 U6967 ( .A1(n5893), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5894) );
  XNOR2_X1 U6968 ( .A(n5894), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U6969 ( .A1(n5915), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9772), .B2(
        n5914), .ZN(n5895) );
  NAND2_X1 U6970 ( .A1(n10123), .A2(n6000), .ZN(n5906) );
  INV_X1 U6971 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5897) );
  AND2_X1 U6972 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  OR2_X1 U6973 ( .A1(n5899), .A2(n5918), .ZN(n9966) );
  INV_X1 U6974 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5900) );
  OAI22_X1 U6975 ( .A1(n9966), .A2(n5973), .B1(n5901), .B2(n5900), .ZN(n5902)
         );
  INV_X1 U6976 ( .A(n5902), .ZN(n5904) );
  AOI22_X1 U6977 ( .A1(n4867), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5903) );
  OR2_X1 U6978 ( .A1(n9975), .A2(n6141), .ZN(n5905) );
  NAND2_X1 U6979 ( .A1(n5906), .A2(n5905), .ZN(n9390) );
  NAND2_X1 U6980 ( .A1(n10123), .A2(n5539), .ZN(n5909) );
  OR2_X1 U6981 ( .A1(n9975), .A2(n5907), .ZN(n5908) );
  NAND2_X1 U6982 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  XNOR2_X1 U6983 ( .A(n5910), .B(n6090), .ZN(n9389) );
  OAI21_X1 U6984 ( .B1(n9392), .B2(n9390), .A(n9389), .ZN(n5912) );
  NAND2_X1 U6985 ( .A1(n9392), .A2(n9390), .ZN(n5911) );
  NAND2_X1 U6986 ( .A1(n5912), .A2(n5911), .ZN(n9312) );
  MUX2_X1 U6987 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7285), .Z(n5930) );
  XNOR2_X1 U6988 ( .A(n5930), .B(SI_19_), .ZN(n5936) );
  NAND2_X1 U6989 ( .A1(n7970), .A2(n9493), .ZN(n5917) );
  AOI22_X1 U6990 ( .A1(n5915), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10494), 
        .B2(n5914), .ZN(n5916) );
  NAND2_X1 U6991 ( .A1(n10117), .A2(n5539), .ZN(n5923) );
  NOR2_X1 U6992 ( .A1(n5918), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5919) );
  OR2_X1 U6993 ( .A1(n5943), .A2(n5919), .ZN(n9946) );
  AOI22_X1 U6994 ( .A1(n6182), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n4876), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U6995 ( .A1(n4874), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5920) );
  OAI211_X1 U6996 ( .C1(n9946), .C2(n5973), .A(n5921), .B(n5920), .ZN(n9956)
         );
  NAND2_X1 U6997 ( .A1(n9956), .A2(n6000), .ZN(n5922) );
  NAND2_X1 U6998 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  XNOR2_X1 U6999 ( .A(n5924), .B(n5508), .ZN(n5926) );
  AND2_X1 U7000 ( .A1(n9956), .A2(n6112), .ZN(n5925) );
  AOI21_X1 U7001 ( .B1(n10117), .B2(n6000), .A(n5925), .ZN(n5927) );
  NAND2_X1 U7002 ( .A1(n5926), .A2(n5927), .ZN(n9311) );
  INV_X1 U7003 ( .A(n5926), .ZN(n5929) );
  INV_X1 U7004 ( .A(n5927), .ZN(n5928) );
  NAND2_X1 U7005 ( .A1(n5929), .A2(n5928), .ZN(n9366) );
  INV_X1 U7006 ( .A(n5930), .ZN(n5931) );
  NAND2_X1 U7007 ( .A1(n5931), .A2(n7205), .ZN(n5933) );
  INV_X1 U7008 ( .A(n5933), .ZN(n5938) );
  INV_X1 U7009 ( .A(n5934), .ZN(n5935) );
  NOR2_X1 U7010 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  MUX2_X1 U7011 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7285), .Z(n5955) );
  XNOR2_X1 U7012 ( .A(n5955), .B(n7111), .ZN(n5957) );
  XNOR2_X1 U7013 ( .A(n5958), .B(n5957), .ZN(n8015) );
  NAND2_X1 U7014 ( .A1(n8015), .A2(n9493), .ZN(n5942) );
  INV_X1 U7015 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8348) );
  OR2_X1 U7016 ( .A1(n5548), .A2(n8348), .ZN(n5941) );
  NAND2_X1 U7017 ( .A1(n10112), .A2(n5539), .ZN(n5948) );
  NOR2_X1 U7018 ( .A1(n5943), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7019 ( .A1(n5969), .A2(n5944), .ZN(n9931) );
  AOI22_X1 U7020 ( .A1(n6182), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7021 ( .A1(n4874), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5945) );
  OAI211_X1 U7022 ( .C1(n9931), .C2(n5973), .A(n5946), .B(n5945), .ZN(n9944)
         );
  NAND2_X1 U7023 ( .A1(n9944), .A2(n6000), .ZN(n5947) );
  NAND2_X1 U7024 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  XNOR2_X1 U7025 ( .A(n5949), .B(n5508), .ZN(n9369) );
  INV_X1 U7026 ( .A(n9369), .ZN(n5951) );
  AND2_X1 U7027 ( .A1(n9944), .A2(n6112), .ZN(n5950) );
  AOI21_X1 U7028 ( .B1(n10112), .B2(n6000), .A(n5950), .ZN(n5953) );
  INV_X1 U7029 ( .A(n5953), .ZN(n9368) );
  NAND2_X1 U7030 ( .A1(n5951), .A2(n9368), .ZN(n5952) );
  AND2_X1 U7031 ( .A1(n9366), .A2(n5952), .ZN(n5954) );
  NOR2_X1 U7032 ( .A1(n5955), .A2(SI_20_), .ZN(n5956) );
  MUX2_X1 U7033 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7284), .Z(n5959) );
  NAND2_X1 U7034 ( .A1(n5959), .A2(SI_21_), .ZN(n5983) );
  INV_X1 U7035 ( .A(n5959), .ZN(n5960) );
  NAND2_X1 U7036 ( .A1(n5960), .A2(n7118), .ZN(n5961) );
  NAND2_X1 U7037 ( .A1(n5983), .A2(n5961), .ZN(n5964) );
  INV_X1 U7038 ( .A(n5964), .ZN(n5962) );
  INV_X1 U7039 ( .A(n5963), .ZN(n5965) );
  NAND2_X1 U7040 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  INV_X1 U7041 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8344) );
  OR2_X1 U7042 ( .A1(n5548), .A2(n8344), .ZN(n5967) );
  NAND2_X1 U7043 ( .A1(n10108), .A2(n5539), .ZN(n5975) );
  NOR2_X1 U7044 ( .A1(n5969), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7045 ( .A1(n5987), .A2(n5970), .ZN(n9918) );
  AOI22_X1 U7046 ( .A1(n6182), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7047 ( .A1(n4873), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5971) );
  OAI211_X1 U7048 ( .C1(n9918), .C2(n5973), .A(n5972), .B(n5971), .ZN(n9928)
         );
  NAND2_X1 U7049 ( .A1(n9928), .A2(n6000), .ZN(n5974) );
  NAND2_X1 U7050 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  XNOR2_X1 U7051 ( .A(n5976), .B(n6090), .ZN(n5979) );
  NAND2_X1 U7052 ( .A1(n10108), .A2(n6000), .ZN(n5978) );
  NAND2_X1 U7053 ( .A1(n9928), .A2(n6112), .ZN(n5977) );
  NAND2_X1 U7054 ( .A1(n5978), .A2(n5977), .ZN(n5980) );
  INV_X1 U7055 ( .A(n5979), .ZN(n5982) );
  INV_X1 U7056 ( .A(n5980), .ZN(n5981) );
  NAND2_X1 U7057 ( .A1(n5982), .A2(n5981), .ZN(n9322) );
  NAND2_X1 U7058 ( .A1(n9319), .A2(n9322), .ZN(n9379) );
  MUX2_X1 U7059 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7285), .Z(n6005) );
  XNOR2_X1 U7060 ( .A(n6005), .B(SI_22_), .ZN(n6008) );
  XNOR2_X1 U7061 ( .A(n6009), .B(n6008), .ZN(n8479) );
  NAND2_X1 U7062 ( .A1(n8479), .A2(n9493), .ZN(n5986) );
  INV_X1 U7063 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8481) );
  OR2_X1 U7064 ( .A1(n5548), .A2(n8481), .ZN(n5985) );
  NAND2_X1 U7065 ( .A1(n10102), .A2(n5539), .ZN(n5997) );
  OR2_X1 U7066 ( .A1(n5987), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7067 ( .A1(n5987), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6013) );
  AND2_X1 U7068 ( .A1(n5988), .A2(n6013), .ZN(n9903) );
  NAND2_X1 U7069 ( .A1(n9903), .A2(n4869), .ZN(n5995) );
  INV_X1 U7070 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7071 ( .A1(n4875), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7072 ( .A1(n4874), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7073 ( .C1(n5992), .C2(n5991), .A(n5990), .B(n5989), .ZN(n5993)
         );
  INV_X1 U7074 ( .A(n5993), .ZN(n5994) );
  NAND2_X1 U7075 ( .A1(n5995), .A2(n5994), .ZN(n9879) );
  NAND2_X1 U7076 ( .A1(n9879), .A2(n6000), .ZN(n5996) );
  NAND2_X1 U7077 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7078 ( .A(n5998), .B(n6090), .ZN(n6001) );
  AND2_X1 U7079 ( .A1(n9879), .A2(n6112), .ZN(n5999) );
  AOI21_X1 U7080 ( .B1(n10102), .B2(n6000), .A(n5999), .ZN(n6002) );
  XNOR2_X1 U7081 ( .A(n6001), .B(n6002), .ZN(n9380) );
  NAND2_X1 U7082 ( .A1(n9379), .A2(n9380), .ZN(n9378) );
  INV_X1 U7083 ( .A(n6001), .ZN(n6003) );
  NAND2_X1 U7084 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  INV_X1 U7085 ( .A(n6005), .ZN(n6007) );
  INV_X1 U7086 ( .A(SI_22_), .ZN(n6006) );
  MUX2_X1 U7087 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7285), .Z(n6028) );
  XNOR2_X1 U7088 ( .A(n6028), .B(n7105), .ZN(n6026) );
  XNOR2_X1 U7089 ( .A(n6027), .B(n6026), .ZN(n8333) );
  NAND2_X1 U7090 ( .A1(n8333), .A2(n9493), .ZN(n6011) );
  INV_X1 U7091 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8336) );
  OR2_X1 U7092 ( .A1(n5548), .A2(n8336), .ZN(n6010) );
  NAND2_X1 U7093 ( .A1(n10094), .A2(n5539), .ZN(n6021) );
  INV_X1 U7094 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U7095 ( .A1(n6012), .A2(n6013), .ZN(n6015) );
  INV_X1 U7096 ( .A(n6013), .ZN(n6014) );
  NAND2_X1 U7097 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6014), .ZN(n6041) );
  AND2_X1 U7098 ( .A1(n6015), .A2(n6041), .ZN(n9883) );
  NAND2_X1 U7099 ( .A1(n5566), .A2(n9883), .ZN(n6019) );
  NAND2_X1 U7100 ( .A1(n6182), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7101 ( .A1(n4875), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7102 ( .A1(n4873), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6016) );
  NAND4_X1 U7103 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n9897)
         );
  NAND2_X1 U7104 ( .A1(n9897), .A2(n6000), .ZN(n6020) );
  NAND2_X1 U7105 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  XNOR2_X1 U7106 ( .A(n6022), .B(n5508), .ZN(n6025) );
  NAND2_X1 U7107 ( .A1(n10094), .A2(n6000), .ZN(n6024) );
  NAND2_X1 U7108 ( .A1(n9897), .A2(n6112), .ZN(n6023) );
  NAND2_X1 U7109 ( .A1(n6024), .A2(n6023), .ZN(n9303) );
  INV_X1 U7110 ( .A(n6028), .ZN(n6029) );
  NAND2_X1 U7111 ( .A1(n6029), .A2(n7105), .ZN(n6030) );
  NAND2_X1 U7112 ( .A1(n6031), .A2(n6030), .ZN(n6035) );
  MUX2_X1 U7113 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7284), .Z(n6032) );
  NAND2_X1 U7114 ( .A1(n6032), .A2(SI_24_), .ZN(n6056) );
  OAI21_X1 U7115 ( .B1(n6032), .B2(SI_24_), .A(n6056), .ZN(n6034) );
  INV_X1 U7116 ( .A(n6034), .ZN(n6033) );
  NAND2_X1 U7117 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7118 ( .A1(n6057), .A2(n6036), .ZN(n8435) );
  OR2_X1 U7119 ( .A1(n8435), .A2(n5536), .ZN(n6038) );
  INV_X1 U7120 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8434) );
  OR2_X1 U7121 ( .A1(n5548), .A2(n8434), .ZN(n6037) );
  NAND2_X1 U7122 ( .A1(n10090), .A2(n5539), .ZN(n6048) );
  NAND2_X1 U7123 ( .A1(n4867), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6046) );
  INV_X1 U7124 ( .A(n6041), .ZN(n6039) );
  NAND2_X1 U7125 ( .A1(n6039), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6062) );
  INV_X1 U7126 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7127 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  AND2_X1 U7128 ( .A1(n6062), .A2(n6042), .ZN(n9869) );
  NAND2_X1 U7129 ( .A1(n4869), .A2(n9869), .ZN(n6045) );
  NAND2_X1 U7130 ( .A1(n4876), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7131 ( .A1(n4874), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6043) );
  NAND4_X1 U7132 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n9878)
         );
  NAND2_X1 U7133 ( .A1(n9878), .A2(n6000), .ZN(n6047) );
  NAND2_X1 U7134 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  XNOR2_X1 U7135 ( .A(n6049), .B(n5508), .ZN(n6054) );
  AND2_X1 U7136 ( .A1(n9878), .A2(n6112), .ZN(n6050) );
  AOI21_X1 U7137 ( .B1(n10090), .B2(n6000), .A(n6050), .ZN(n6053) );
  XNOR2_X1 U7138 ( .A(n6054), .B(n6053), .ZN(n9359) );
  NAND2_X1 U7139 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  NAND2_X1 U7140 ( .A1(n9357), .A2(n6055), .ZN(n9330) );
  MUX2_X1 U7141 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7285), .Z(n6075) );
  XNOR2_X1 U7142 ( .A(n6075), .B(SI_25_), .ZN(n6078) );
  XNOR2_X1 U7143 ( .A(n6079), .B(n6078), .ZN(n8453) );
  NAND2_X1 U7144 ( .A1(n8453), .A2(n9493), .ZN(n6059) );
  INV_X1 U7145 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8456) );
  OR2_X1 U7146 ( .A1(n5548), .A2(n8456), .ZN(n6058) );
  NAND2_X1 U7147 ( .A1(n10084), .A2(n5539), .ZN(n6069) );
  INV_X1 U7148 ( .A(n6062), .ZN(n6060) );
  NAND2_X1 U7149 ( .A1(n6060), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6084) );
  INV_X1 U7150 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7151 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  AND2_X1 U7152 ( .A1(n6084), .A2(n6063), .ZN(n9847) );
  NAND2_X1 U7153 ( .A1(n5566), .A2(n9847), .ZN(n6067) );
  NAND2_X1 U7154 ( .A1(n6182), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7155 ( .A1(n4877), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7156 ( .A1(n4873), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6064) );
  NAND4_X1 U7157 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n9863)
         );
  NAND2_X1 U7158 ( .A1(n9863), .A2(n6000), .ZN(n6068) );
  NAND2_X1 U7159 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  XNOR2_X1 U7160 ( .A(n6070), .B(n5508), .ZN(n9332) );
  AND2_X1 U7161 ( .A1(n9863), .A2(n6112), .ZN(n6071) );
  AOI21_X1 U7162 ( .B1(n10084), .B2(n6000), .A(n6071), .ZN(n9331) );
  INV_X1 U7163 ( .A(n9332), .ZN(n6073) );
  INV_X1 U7164 ( .A(n9331), .ZN(n6072) );
  NAND2_X1 U7165 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  INV_X1 U7166 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7167 ( .A1(n6076), .A2(n7092), .ZN(n6077) );
  MUX2_X1 U7168 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7285), .Z(n6099) );
  XNOR2_X1 U7169 ( .A(n6099), .B(n7197), .ZN(n6097) );
  XNOR2_X1 U7170 ( .A(n6098), .B(n6097), .ZN(n9279) );
  NAND2_X1 U7171 ( .A1(n9279), .A2(n9493), .ZN(n6081) );
  INV_X1 U7172 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10205) );
  OR2_X1 U7173 ( .A1(n5548), .A2(n10205), .ZN(n6080) );
  NAND2_X1 U7174 ( .A1(n10079), .A2(n5539), .ZN(n6089) );
  AOI22_X1 U7175 ( .A1(n6182), .A2(P1_REG1_REG_26__SCAN_IN), .B1(n4877), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n6087) );
  INV_X1 U7176 ( .A(n6084), .ZN(n6082) );
  NAND2_X1 U7177 ( .A1(n6082), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6133) );
  INV_X1 U7178 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7179 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  AOI22_X1 U7180 ( .A1(n5566), .A2(n9832), .B1(n4873), .B2(
        P1_REG0_REG_26__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7181 ( .A1(n9818), .A2(n5907), .ZN(n6088) );
  NAND2_X1 U7182 ( .A1(n6089), .A2(n6088), .ZN(n6091) );
  XNOR2_X1 U7183 ( .A(n6091), .B(n6090), .ZN(n6093) );
  NOR2_X1 U7184 ( .A1(n9818), .A2(n6141), .ZN(n6092) );
  AOI21_X1 U7185 ( .B1(n10079), .B2(n6000), .A(n6092), .ZN(n6094) );
  XNOR2_X1 U7186 ( .A(n6093), .B(n6094), .ZN(n9400) );
  INV_X1 U7187 ( .A(n6093), .ZN(n6095) );
  NAND2_X1 U7188 ( .A1(n6098), .A2(n6097), .ZN(n6102) );
  INV_X1 U7189 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7190 ( .A1(n6100), .A2(n7197), .ZN(n6101) );
  MUX2_X1 U7191 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7284), .Z(n6121) );
  XNOR2_X1 U7192 ( .A(n6121), .B(n7194), .ZN(n6119) );
  NAND2_X1 U7193 ( .A1(n10200), .A2(n9493), .ZN(n6104) );
  INV_X1 U7194 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10203) );
  OR2_X1 U7195 ( .A1(n5548), .A2(n10203), .ZN(n6103) );
  NAND2_X1 U7196 ( .A1(n10074), .A2(n5539), .ZN(n6110) );
  XNOR2_X1 U7197 ( .A(n6133), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U7198 ( .A1(n5566), .A2(n9813), .ZN(n6108) );
  NAND2_X1 U7199 ( .A1(n4867), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7200 ( .A1(n5681), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7201 ( .A1(n4874), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6105) );
  NAND4_X1 U7202 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n9826)
         );
  NAND2_X1 U7203 ( .A1(n9826), .A2(n6000), .ZN(n6109) );
  NAND2_X1 U7204 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  XNOR2_X1 U7205 ( .A(n6111), .B(n5508), .ZN(n6114) );
  AND2_X1 U7206 ( .A1(n9826), .A2(n6112), .ZN(n6113) );
  AOI21_X1 U7207 ( .B1(n10074), .B2(n6000), .A(n6113), .ZN(n6115) );
  NAND2_X1 U7208 ( .A1(n6114), .A2(n6115), .ZN(n6190) );
  INV_X1 U7209 ( .A(n6114), .ZN(n6117) );
  INV_X1 U7210 ( .A(n6115), .ZN(n6116) );
  NAND2_X1 U7211 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  NAND2_X1 U7212 ( .A1(n6120), .A2(n6119), .ZN(n6124) );
  INV_X1 U7213 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7214 ( .A1(n6122), .A2(n7194), .ZN(n6123) );
  NAND2_X1 U7215 ( .A1(n6124), .A2(n6123), .ZN(n6126) );
  MUX2_X1 U7216 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7285), .Z(n6804) );
  XNOR2_X1 U7217 ( .A(n6804), .B(n7191), .ZN(n6125) );
  NAND2_X1 U7218 ( .A1(n6126), .A2(n6125), .ZN(n6807) );
  OR2_X1 U7219 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7220 ( .A1(n6807), .A2(n6127), .ZN(n9274) );
  NAND2_X1 U7221 ( .A1(n9274), .A2(n9493), .ZN(n6130) );
  INV_X1 U7222 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n6128) );
  OR2_X1 U7223 ( .A1(n5548), .A2(n6128), .ZN(n6129) );
  NAND2_X1 U7224 ( .A1(n10066), .A2(n5539), .ZN(n6138) );
  AOI22_X1 U7225 ( .A1(n6182), .A2(P1_REG1_REG_28__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n6136) );
  INV_X1 U7226 ( .A(n6133), .ZN(n6132) );
  AND2_X1 U7227 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6131) );
  NAND2_X1 U7228 ( .A1(n6132), .A2(n6131), .ZN(n6183) );
  INV_X1 U7229 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7064) );
  INV_X1 U7230 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6187) );
  OAI21_X1 U7231 ( .B1(n6133), .B2(n7064), .A(n6187), .ZN(n6134) );
  AND2_X1 U7232 ( .A1(n6183), .A2(n6134), .ZN(n6179) );
  AOI22_X1 U7233 ( .A1(n4869), .A2(n6179), .B1(n4874), .B2(
        P1_REG0_REG_28__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7234 ( .A1(n9817), .A2(n5907), .ZN(n6137) );
  NAND2_X1 U7235 ( .A1(n6138), .A2(n6137), .ZN(n6139) );
  XNOR2_X1 U7236 ( .A(n6139), .B(n5508), .ZN(n6143) );
  NAND2_X1 U7237 ( .A1(n10066), .A2(n5713), .ZN(n6140) );
  OAI21_X1 U7238 ( .B1(n9817), .B2(n6141), .A(n6140), .ZN(n6142) );
  XNOR2_X1 U7239 ( .A(n6143), .B(n6142), .ZN(n6194) );
  INV_X1 U7240 ( .A(n6194), .ZN(n6191) );
  NAND2_X1 U7241 ( .A1(n8458), .A2(P1_B_REG_SCAN_IN), .ZN(n6145) );
  INV_X1 U7242 ( .A(n8436), .ZN(n6144) );
  MUX2_X1 U7243 ( .A(n6145), .B(P1_B_REG_SCAN_IN), .S(n6144), .Z(n6147) );
  NAND2_X1 U7244 ( .A1(n6147), .A2(n6146), .ZN(n6149) );
  INV_X1 U7245 ( .A(n8458), .ZN(n6148) );
  OAI22_X1 U7246 ( .A1(n6149), .A2(P1_D_REG_1__SCAN_IN), .B1(n6146), .B2(n6148), .ZN(n7700) );
  INV_X1 U7247 ( .A(n7700), .ZN(n6161) );
  INV_X1 U7248 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6150) );
  INV_X1 U7249 ( .A(n6146), .ZN(n10207) );
  NOR4_X1 U7250 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7251 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6153) );
  NOR4_X1 U7252 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6152) );
  NOR4_X1 U7253 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6151) );
  NAND4_X1 U7254 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n6160)
         );
  NOR2_X1 U7255 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6158) );
  NOR4_X1 U7256 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7257 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6156) );
  NOR4_X1 U7258 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6155) );
  NAND4_X1 U7259 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n6159)
         );
  OAI21_X1 U7260 ( .B1(n6160), .B2(n6159), .A(n7294), .ZN(n7702) );
  NAND3_X1 U7261 ( .A1(n6161), .A2(n7436), .A3(n7702), .ZN(n7448) );
  AND2_X2 U7262 ( .A1(n7728), .A2(n6162), .ZN(n10561) );
  INV_X1 U7263 ( .A(n6163), .ZN(n7717) );
  NOR2_X1 U7264 ( .A1(n10561), .A2(n7717), .ZN(n6173) );
  NAND2_X1 U7265 ( .A1(n6165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  MUX2_X1 U7266 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6166), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6168) );
  NAND2_X1 U7267 ( .A1(n6168), .A2(n6167), .ZN(n7070) );
  AND2_X1 U7268 ( .A1(n7070), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7269 ( .A1(n6173), .A2(n7431), .ZN(n6170) );
  NAND3_X1 U7270 ( .A1(n6191), .A2(n9381), .A3(n6190), .ZN(n6198) );
  NAND2_X1 U7271 ( .A1(n7728), .A2(n9659), .ZN(n7705) );
  OR2_X1 U7272 ( .A1(n10287), .A2(n7705), .ZN(n6176) );
  OR2_X1 U7273 ( .A1(n7448), .A2(n6176), .ZN(n6172) );
  NAND2_X1 U7274 ( .A1(n7448), .A2(n6173), .ZN(n6174) );
  OR2_X1 U7275 ( .A1(n6163), .A2(n7706), .ZN(n7433) );
  AND3_X1 U7276 ( .A1(n7069), .A2(n7070), .A3(n7433), .ZN(n7447) );
  NAND2_X1 U7277 ( .A1(n6174), .A2(n7447), .ZN(n6175) );
  NAND2_X1 U7278 ( .A1(n6175), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6178) );
  OR2_X1 U7279 ( .A1(n10287), .A2(n7428), .ZN(n9664) );
  NAND2_X1 U7280 ( .A1(n9664), .A2(n6176), .ZN(n6177) );
  NAND2_X1 U7281 ( .A1(n7448), .A2(n6177), .ZN(n7449) );
  INV_X1 U7282 ( .A(n6179), .ZN(n9802) );
  NOR2_X1 U7283 ( .A1(n7448), .A2(n9664), .ZN(n6186) );
  NAND2_X1 U7284 ( .A1(n6186), .A2(n6181), .ZN(n9342) );
  AOI22_X1 U7285 ( .A1(n4867), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n4875), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n6185) );
  INV_X1 U7286 ( .A(n6183), .ZN(n8633) );
  AOI22_X1 U7287 ( .A1(n5566), .A2(n8633), .B1(n4873), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n6184) );
  AND2_X1 U7288 ( .A1(n6185), .A2(n6184), .ZN(n8592) );
  INV_X1 U7289 ( .A(n8592), .ZN(n9795) );
  INV_X1 U7290 ( .A(n9826), .ZN(n8588) );
  OAI22_X1 U7291 ( .A1(n9405), .A2(n8588), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6187), .ZN(n6188) );
  AOI21_X1 U7292 ( .B1(n9401), .B2(n9795), .A(n6188), .ZN(n6189) );
  OAI21_X1 U7293 ( .B1(n9395), .B2(n9802), .A(n6189), .ZN(n6193) );
  NOR3_X1 U7294 ( .A1(n6191), .A2(n9410), .A3(n6190), .ZN(n6192) );
  AOI211_X1 U7295 ( .C1(n10066), .C2(n9408), .A(n6193), .B(n6192), .ZN(n6197)
         );
  AND2_X1 U7296 ( .A1(n6194), .A2(n9381), .ZN(n6195) );
  OAI211_X1 U7297 ( .C1(n7063), .C2(n6198), .A(n6197), .B(n6196), .ZN(P1_U3218) );
  NOR2_X1 U7298 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6202) );
  AND2_X2 U7299 ( .A1(n6275), .A2(n6203), .ZN(n6338) );
  NAND2_X1 U7300 ( .A1(n6230), .A2(n6205), .ZN(n6233) );
  INV_X1 U7301 ( .A(n6233), .ZN(n6209) );
  NOR2_X1 U7302 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6207) );
  NAND4_X1 U7303 ( .A1(n6209), .A2(n6208), .A3(n4912), .A4(n6207), .ZN(n6210)
         );
  INV_X1 U7304 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6214) );
  XNOR2_X1 U7305 ( .A(n6216), .B(n6215), .ZN(n6763) );
  NAND2_X1 U7306 ( .A1(n6729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7307 ( .A1(n7681), .A2(n6883), .ZN(n6226) );
  INV_X2 U7308 ( .A(n6288), .ZN(n6555) );
  INV_X2 U7309 ( .A(n6289), .ZN(n6554) );
  NAND3_X1 U7310 ( .A1(n6490), .A2(n6508), .A3(n6222), .ZN(n6223) );
  NAND2_X1 U7311 ( .A1(n6227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6224) );
  XNOR2_X1 U7312 ( .A(n6224), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8884) );
  AOI22_X1 U7313 ( .A1(n6555), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6554), .B2(
        n8884), .ZN(n6225) );
  NAND2_X1 U7314 ( .A1(n6231), .A2(n6230), .ZN(n6241) );
  NOR2_X1 U7315 ( .A1(n6233), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7316 ( .A1(n6235), .A2(n6234), .ZN(n6238) );
  NAND2_X1 U7317 ( .A1(n6238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7318 ( .A1(n6239), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7319 ( .A1(n7058), .A2(n8993), .ZN(n6242) );
  XNOR2_X1 U7320 ( .A(n9242), .B(n6280), .ZN(n6260) );
  NAND2_X1 U7321 ( .A1(n6327), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6360) );
  INV_X1 U7322 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U7323 ( .A1(n6360), .A2(n6359), .ZN(n6358) );
  NAND2_X1 U7324 ( .A1(n6358), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7325 ( .A1(n6495), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U7326 ( .A1(n6517), .A2(n6243), .ZN(n6244) );
  NAND2_X1 U7327 ( .A1(n6533), .A2(n6244), .ZN(n8708) );
  INV_X1 U7328 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7329 ( .A1(n6297), .A2(n8866), .ZN(n6250) );
  OAI21_X1 U7330 ( .B1(n8708), .B2(n6309), .A(n6250), .ZN(n6258) );
  INV_X1 U7331 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n6256) );
  NAND2_X2 U7332 ( .A1(n6253), .A2(n9273), .ZN(n6311) );
  INV_X1 U7333 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6254) );
  OR2_X1 U7334 ( .A1(n6311), .A2(n6254), .ZN(n6255) );
  OAI21_X1 U7335 ( .B1(n6295), .B2(n6256), .A(n6255), .ZN(n6257) );
  NAND2_X1 U7336 ( .A1(n6795), .A2(n6302), .ZN(n6261) );
  NAND2_X1 U7337 ( .A1(n6260), .A2(n6261), .ZN(n6528) );
  INV_X1 U7338 ( .A(n6260), .ZN(n6263) );
  INV_X1 U7339 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7340 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  AND2_X1 U7341 ( .A1(n6528), .A2(n6264), .ZN(n8706) );
  INV_X1 U7342 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7343 ( .A1(n6295), .A2(n6265), .ZN(n6268) );
  INV_X1 U7344 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7345 ( .A1(n6311), .A2(n6266), .ZN(n6267) );
  INV_X1 U7346 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10657) );
  NOR2_X1 U7347 ( .A1(n7285), .A2(n7233), .ZN(n6271) );
  XNOR2_X1 U7348 ( .A(n6271), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9284) );
  MUX2_X1 U7349 ( .A(n10657), .B(n9284), .S(n6289), .Z(n7622) );
  INV_X1 U7350 ( .A(n7622), .ZN(n7600) );
  NAND2_X1 U7351 ( .A1(n7424), .A2(n7600), .ZN(n7612) );
  NAND2_X1 U7352 ( .A1(n6272), .A2(n6302), .ZN(n7490) );
  NAND2_X1 U7353 ( .A1(n6280), .A2(n7622), .ZN(n6273) );
  NAND2_X1 U7354 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6274) );
  INV_X1 U7355 ( .A(n6275), .ZN(n6276) );
  OR2_X1 U7356 ( .A1(n6289), .A2(n8167), .ZN(n6278) );
  INV_X1 U7357 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U7358 ( .A1(n6561), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6283) );
  INV_X1 U7359 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7621) );
  INV_X1 U7360 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8168) );
  OR2_X1 U7361 ( .A1(n6297), .A2(n8168), .ZN(n6282) );
  INV_X1 U7362 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7627) );
  INV_X1 U7363 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U7364 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  OR2_X1 U7365 ( .A1(n6640), .A2(n7302), .ZN(n6293) );
  INV_X1 U7366 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7301) );
  OR2_X1 U7367 ( .A1(n6275), .A2(n6214), .ZN(n6290) );
  XNOR2_X1 U7368 ( .A(n6290), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10629) );
  INV_X1 U7369 ( .A(n10629), .ZN(n7303) );
  OR2_X1 U7370 ( .A1(n6289), .A2(n7303), .ZN(n6291) );
  AND3_X2 U7371 ( .A1(n6293), .A2(n6292), .A3(n6291), .ZN(n10386) );
  XNOR2_X1 U7372 ( .A(n10386), .B(n6325), .ZN(n8664) );
  INV_X1 U7373 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6294) );
  INV_X1 U7374 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6296) );
  INV_X1 U7375 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U7376 ( .A1(n8662), .A2(n6302), .ZN(n6303) );
  OR2_X1 U7377 ( .A1(n8664), .A2(n6303), .ZN(n6305) );
  NAND2_X1 U7378 ( .A1(n6303), .A2(n8664), .ZN(n6304) );
  AND2_X1 U7379 ( .A1(n6305), .A2(n6304), .ZN(n10376) );
  NAND2_X1 U7380 ( .A1(n8665), .A2(n6305), .ZN(n6321) );
  NAND2_X1 U7381 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4910), .ZN(n6306) );
  XNOR2_X1 U7382 ( .A(n6306), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8164) );
  AOI22_X1 U7383 ( .A1(n6555), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6554), .B2(
        n8164), .ZN(n6308) );
  OR2_X1 U7384 ( .A1(n7287), .A2(n6640), .ZN(n6307) );
  XNOR2_X1 U7385 ( .A(n6781), .B(n6280), .ZN(n6317) );
  INV_X1 U7386 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8165) );
  OR2_X1 U7387 ( .A1(n6297), .A2(n8165), .ZN(n6316) );
  INV_X1 U7388 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6310) );
  OR2_X1 U7389 ( .A1(n6311), .A2(n6310), .ZN(n6313) );
  NAND2_X1 U7390 ( .A1(n6561), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6312) );
  AND2_X1 U7391 ( .A1(n10451), .A2(n6302), .ZN(n6318) );
  NAND2_X1 U7392 ( .A1(n6317), .A2(n6318), .ZN(n6332) );
  INV_X1 U7393 ( .A(n6317), .ZN(n7511) );
  INV_X1 U7394 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7395 ( .A1(n7511), .A2(n6319), .ZN(n6320) );
  AND2_X1 U7396 ( .A1(n6332), .A2(n6320), .ZN(n8666) );
  OR2_X1 U7397 ( .A1(n7293), .A2(n6640), .ZN(n6324) );
  OR2_X1 U7398 ( .A1(n6338), .A2(n6214), .ZN(n6322) );
  XNOR2_X1 U7399 ( .A(n6322), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8162) );
  AOI22_X1 U7400 ( .A1(n6555), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6554), .B2(
        n8162), .ZN(n6323) );
  NAND2_X1 U7401 ( .A1(n6561), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6331) );
  INV_X1 U7402 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8163) );
  OR2_X1 U7403 ( .A1(n6297), .A2(n8163), .ZN(n6330) );
  INV_X1 U7404 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6326) );
  OR2_X1 U7405 ( .A1(n6311), .A2(n6326), .ZN(n6329) );
  INV_X1 U7406 ( .A(n6327), .ZN(n6345) );
  OAI21_X1 U7407 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n6345), .ZN(n10469) );
  OR2_X1 U7408 ( .A1(n4870), .A2(n10469), .ZN(n6328) );
  NAND2_X1 U7409 ( .A1(n8663), .A2(n6302), .ZN(n6334) );
  XNOR2_X1 U7410 ( .A(n8575), .B(n6334), .ZN(n7521) );
  AND2_X1 U7411 ( .A1(n7521), .A2(n6332), .ZN(n6333) );
  INV_X1 U7412 ( .A(n8575), .ZN(n6335) );
  NAND2_X1 U7413 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  OR2_X1 U7414 ( .A1(n7305), .A2(n6640), .ZN(n6343) );
  INV_X1 U7415 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7416 ( .A1(n6338), .A2(n6337), .ZN(n6340) );
  NAND2_X1 U7417 ( .A1(n6340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  MUX2_X1 U7418 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6339), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6341) );
  AOI22_X1 U7419 ( .A1(n6555), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6554), .B2(
        n8160), .ZN(n6342) );
  XNOR2_X1 U7420 ( .A(n7662), .B(n6280), .ZN(n6351) );
  NAND2_X1 U7421 ( .A1(n6561), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6350) );
  INV_X1 U7422 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8161) );
  OR2_X1 U7423 ( .A1(n6297), .A2(n8161), .ZN(n6349) );
  INV_X1 U7424 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6344) );
  OR2_X1 U7425 ( .A1(n6311), .A2(n6344), .ZN(n6348) );
  INV_X1 U7426 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U7427 ( .A1(n6345), .A2(n8574), .ZN(n6346) );
  NAND2_X1 U7428 ( .A1(n6360), .A2(n6346), .ZN(n7660) );
  OR2_X1 U7429 ( .A1(n4870), .A2(n7660), .ZN(n6347) );
  NAND4_X1 U7430 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n10449)
         );
  NAND2_X1 U7431 ( .A1(n10449), .A2(n6302), .ZN(n6352) );
  XNOR2_X1 U7432 ( .A(n6351), .B(n6352), .ZN(n8576) );
  INV_X1 U7433 ( .A(n6351), .ZN(n8560) );
  NAND2_X1 U7434 ( .A1(n8560), .A2(n6352), .ZN(n6353) );
  NAND2_X1 U7435 ( .A1(n8563), .A2(n6353), .ZN(n6366) );
  OR2_X1 U7436 ( .A1(n7290), .A2(n6640), .ZN(n6356) );
  NAND2_X1 U7437 ( .A1(n6371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6354) );
  XNOR2_X1 U7438 ( .A(n6354), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8201) );
  AOI22_X1 U7439 ( .A1(n6555), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6554), .B2(
        n8201), .ZN(n6355) );
  NAND2_X1 U7440 ( .A1(n6356), .A2(n6355), .ZN(n7634) );
  XNOR2_X1 U7441 ( .A(n7634), .B(n6280), .ZN(n6369) );
  NAND2_X1 U7442 ( .A1(n6561), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6365) );
  INV_X1 U7443 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8173) );
  OR2_X1 U7444 ( .A1(n6297), .A2(n8173), .ZN(n6364) );
  INV_X1 U7445 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6357) );
  OR2_X1 U7446 ( .A1(n6311), .A2(n6357), .ZN(n6363) );
  INV_X1 U7447 ( .A(n6358), .ZN(n6375) );
  NAND2_X1 U7448 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  NAND2_X1 U7449 ( .A1(n6375), .A2(n6361), .ZN(n8554) );
  OR2_X1 U7450 ( .A1(n6309), .A2(n8554), .ZN(n6362) );
  NOR2_X1 U7451 ( .A1(n8328), .A2(n6715), .ZN(n6367) );
  XNOR2_X1 U7452 ( .A(n6369), .B(n6367), .ZN(n8562) );
  NAND2_X1 U7453 ( .A1(n6366), .A2(n8562), .ZN(n8568) );
  INV_X1 U7454 ( .A(n6367), .ZN(n6368) );
  NAND2_X1 U7455 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  OR2_X1 U7456 ( .A1(n7300), .A2(n6640), .ZN(n6374) );
  NOR2_X1 U7457 ( .A1(n6371), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7458 ( .A1(n6388), .A2(n6214), .ZN(n6372) );
  XNOR2_X1 U7459 ( .A(n6372), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8213) );
  AOI22_X1 U7460 ( .A1(n6555), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6554), .B2(
        n8213), .ZN(n6373) );
  NAND2_X1 U7461 ( .A1(n6374), .A2(n6373), .ZN(n7792) );
  XNOR2_X1 U7462 ( .A(n7792), .B(n6325), .ZN(n6381) );
  NAND2_X1 U7463 ( .A1(n6561), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6380) );
  INV_X1 U7464 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8204) );
  OR2_X1 U7465 ( .A1(n6297), .A2(n8204), .ZN(n6379) );
  INV_X1 U7466 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7675) );
  OR2_X1 U7467 ( .A1(n6311), .A2(n7675), .ZN(n6378) );
  NAND2_X1 U7468 ( .A1(n6375), .A2(n8199), .ZN(n6376) );
  NAND2_X1 U7469 ( .A1(n6394), .A2(n6376), .ZN(n7674) );
  OR2_X1 U7470 ( .A1(n4870), .A2(n7674), .ZN(n6377) );
  NOR2_X1 U7471 ( .A1(n8556), .A2(n6715), .ZN(n6382) );
  NAND2_X1 U7472 ( .A1(n6381), .A2(n6382), .ZN(n6386) );
  INV_X1 U7473 ( .A(n6381), .ZN(n7586) );
  INV_X1 U7474 ( .A(n6382), .ZN(n6383) );
  NAND2_X1 U7475 ( .A1(n7586), .A2(n6383), .ZN(n6384) );
  NAND2_X1 U7476 ( .A1(n6386), .A2(n6384), .ZN(n7654) );
  INV_X1 U7477 ( .A(n7654), .ZN(n6385) );
  NAND2_X1 U7478 ( .A1(n7306), .A2(n6883), .ZN(n6391) );
  INV_X1 U7479 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U7480 ( .A1(n6388), .A2(n6387), .ZN(n6405) );
  NAND2_X1 U7481 ( .A1(n6405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6389) );
  XNOR2_X1 U7482 ( .A(n6389), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8217) );
  AOI22_X1 U7483 ( .A1(n6555), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6554), .B2(
        n8217), .ZN(n6390) );
  NAND2_X1 U7484 ( .A1(n6391), .A2(n6390), .ZN(n7695) );
  XNOR2_X1 U7485 ( .A(n7695), .B(n6325), .ZN(n6400) );
  NAND2_X1 U7486 ( .A1(n6561), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6399) );
  INV_X1 U7487 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8218) );
  OR2_X1 U7488 ( .A1(n6297), .A2(n8218), .ZN(n6398) );
  INV_X1 U7489 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6392) );
  OR2_X1 U7490 ( .A1(n6311), .A2(n6392), .ZN(n6397) );
  NAND2_X1 U7491 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U7492 ( .A1(n6411), .A2(n6395), .ZN(n7693) );
  OR2_X1 U7493 ( .A1(n4870), .A2(n7693), .ZN(n6396) );
  NOR2_X1 U7494 ( .A1(n8468), .A2(n6715), .ZN(n6401) );
  NAND2_X1 U7495 ( .A1(n6400), .A2(n6401), .ZN(n6417) );
  INV_X1 U7496 ( .A(n6400), .ZN(n8469) );
  INV_X1 U7497 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U7498 ( .A1(n8469), .A2(n6402), .ZN(n6403) );
  AND2_X1 U7499 ( .A1(n6417), .A2(n6403), .ZN(n7584) );
  NAND2_X1 U7500 ( .A1(n6404), .A2(n7584), .ZN(n7587) );
  NAND2_X1 U7501 ( .A1(n7309), .A2(n6883), .ZN(n6408) );
  NAND2_X1 U7502 ( .A1(n6406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6424) );
  XNOR2_X1 U7503 ( .A(n6424), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8242) );
  AOI22_X1 U7504 ( .A1(n6555), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6554), .B2(
        n8242), .ZN(n6407) );
  NAND2_X1 U7505 ( .A1(n6408), .A2(n6407), .ZN(n8476) );
  XNOR2_X1 U7506 ( .A(n8476), .B(n6280), .ZN(n6421) );
  NAND2_X1 U7507 ( .A1(n6561), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6416) );
  INV_X1 U7508 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8221) );
  OR2_X1 U7509 ( .A1(n6297), .A2(n8221), .ZN(n6415) );
  INV_X1 U7510 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7821) );
  OR2_X1 U7511 ( .A1(n6311), .A2(n7821), .ZN(n6414) );
  INV_X1 U7512 ( .A(n6409), .ZN(n6433) );
  NAND2_X1 U7513 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  NAND2_X1 U7514 ( .A1(n6433), .A2(n6412), .ZN(n8462) );
  OR2_X1 U7515 ( .A1(n6309), .A2(n8462), .ZN(n6413) );
  NOR2_X1 U7516 ( .A1(n8315), .A2(n6715), .ZN(n6419) );
  XNOR2_X1 U7517 ( .A(n6421), .B(n6419), .ZN(n8472) );
  AND2_X1 U7518 ( .A1(n8472), .A2(n6417), .ZN(n6418) );
  NAND2_X1 U7519 ( .A1(n7587), .A2(n6418), .ZN(n8478) );
  INV_X1 U7520 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U7521 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  NAND2_X1 U7522 ( .A1(n7354), .A2(n6883), .ZN(n6430) );
  INV_X1 U7523 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U7524 ( .A1(n6424), .A2(n6423), .ZN(n6425) );
  NAND2_X1 U7525 ( .A1(n6425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6427) );
  INV_X1 U7526 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7527 ( .A1(n6427), .A2(n6426), .ZN(n6445) );
  OR2_X1 U7528 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  AOI22_X1 U7529 ( .A1(n6555), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6554), .B2(
        n8789), .ZN(n6429) );
  NAND2_X1 U7530 ( .A1(n6430), .A2(n6429), .ZN(n7900) );
  XNOR2_X1 U7531 ( .A(n7900), .B(n6325), .ZN(n6439) );
  NAND2_X1 U7532 ( .A1(n6561), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6438) );
  INV_X1 U7533 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8248) );
  OR2_X1 U7534 ( .A1(n6297), .A2(n8248), .ZN(n6437) );
  INV_X1 U7535 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7894) );
  OR2_X1 U7536 ( .A1(n6311), .A2(n7894), .ZN(n6436) );
  INV_X1 U7537 ( .A(n6431), .ZN(n6449) );
  INV_X1 U7538 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7539 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  NAND2_X1 U7540 ( .A1(n6449), .A2(n6434), .ZN(n7893) );
  OR2_X1 U7541 ( .A1(n4870), .A2(n7893), .ZN(n6435) );
  NOR2_X1 U7542 ( .A1(n8460), .A2(n6715), .ZN(n6440) );
  NAND2_X1 U7543 ( .A1(n6439), .A2(n6440), .ZN(n6444) );
  INV_X1 U7544 ( .A(n6439), .ZN(n7832) );
  INV_X1 U7545 ( .A(n6440), .ZN(n6441) );
  NAND2_X1 U7546 ( .A1(n7832), .A2(n6441), .ZN(n6442) );
  NAND2_X1 U7547 ( .A1(n6444), .A2(n6442), .ZN(n7076) );
  OR2_X1 U7548 ( .A1(n7383), .A2(n6640), .ZN(n6448) );
  NAND2_X1 U7549 ( .A1(n6445), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U7550 ( .A(n6446), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8813) );
  AOI22_X1 U7551 ( .A1(n6555), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8813), .B2(
        n6554), .ZN(n6447) );
  NAND2_X1 U7552 ( .A1(n6448), .A2(n6447), .ZN(n7877) );
  XNOR2_X1 U7553 ( .A(n7877), .B(n6280), .ZN(n6456) );
  NAND2_X1 U7554 ( .A1(n6561), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6454) );
  INV_X1 U7555 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7875) );
  OR2_X1 U7556 ( .A1(n6311), .A2(n7875), .ZN(n6453) );
  NAND2_X1 U7557 ( .A1(n6449), .A2(n8792), .ZN(n6450) );
  NAND2_X1 U7558 ( .A1(n6464), .A2(n6450), .ZN(n7874) );
  OR2_X1 U7559 ( .A1(n4870), .A2(n7874), .ZN(n6452) );
  INV_X1 U7560 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8796) );
  OR2_X1 U7561 ( .A1(n6297), .A2(n8796), .ZN(n6451) );
  NOR2_X1 U7562 ( .A1(n8322), .A2(n6715), .ZN(n6457) );
  XNOR2_X1 U7563 ( .A(n6456), .B(n6457), .ZN(n7831) );
  INV_X1 U7564 ( .A(n6456), .ZN(n6458) );
  NAND2_X1 U7565 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  NAND2_X1 U7566 ( .A1(n7441), .A2(n6883), .ZN(n6463) );
  OR2_X1 U7567 ( .A1(n6460), .A2(n6214), .ZN(n6461) );
  XNOR2_X1 U7568 ( .A(n6461), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8820) );
  AOI22_X1 U7569 ( .A1(n6555), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6554), .B2(
        n8820), .ZN(n6462) );
  XNOR2_X1 U7570 ( .A(n8000), .B(n6325), .ZN(n7992) );
  NAND2_X1 U7571 ( .A1(n6561), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6469) );
  INV_X1 U7572 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7964) );
  OR2_X1 U7573 ( .A1(n6311), .A2(n7964), .ZN(n6468) );
  NAND2_X1 U7574 ( .A1(n6464), .A2(n7988), .ZN(n6465) );
  NAND2_X1 U7575 ( .A1(n6478), .A2(n6465), .ZN(n7985) );
  OR2_X1 U7576 ( .A1(n6309), .A2(n7985), .ZN(n6467) );
  INV_X1 U7577 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8806) );
  OR2_X1 U7578 ( .A1(n6297), .A2(n8806), .ZN(n6466) );
  NOR2_X1 U7579 ( .A1(n8326), .A2(n6715), .ZN(n6470) );
  AND2_X1 U7580 ( .A1(n7992), .A2(n6470), .ZN(n7991) );
  INV_X1 U7581 ( .A(n7992), .ZN(n6472) );
  INV_X1 U7582 ( .A(n6470), .ZN(n6471) );
  NAND2_X1 U7583 ( .A1(n6472), .A2(n6471), .ZN(n7994) );
  NAND2_X1 U7584 ( .A1(n7480), .A2(n6883), .ZN(n6475) );
  NAND2_X1 U7585 ( .A1(n6473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6491) );
  XNOR2_X1 U7586 ( .A(n6491), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8839) );
  AOI22_X1 U7587 ( .A1(n6555), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6554), .B2(
        n8839), .ZN(n6474) );
  XNOR2_X1 U7588 ( .A(n8128), .B(n6280), .ZN(n6484) );
  NAND2_X1 U7589 ( .A1(n6561), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6483) );
  INV_X1 U7590 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6476) );
  OR2_X1 U7591 ( .A1(n6297), .A2(n6476), .ZN(n6482) );
  INV_X1 U7592 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6477) );
  OR2_X1 U7593 ( .A1(n6311), .A2(n6477), .ZN(n6481) );
  NAND2_X1 U7594 ( .A1(n6478), .A2(n7177), .ZN(n6479) );
  NAND2_X1 U7595 ( .A1(n6496), .A2(n6479), .ZN(n8132) );
  OR2_X1 U7596 ( .A1(n4870), .A2(n8132), .ZN(n6480) );
  OR2_X1 U7597 ( .A1(n8338), .A2(n6715), .ZN(n6485) );
  NAND2_X1 U7598 ( .A1(n6484), .A2(n6485), .ZN(n6489) );
  INV_X1 U7599 ( .A(n6484), .ZN(n6487) );
  INV_X1 U7600 ( .A(n6485), .ZN(n6486) );
  NAND2_X1 U7601 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  AND2_X1 U7602 ( .A1(n6489), .A2(n6488), .ZN(n8019) );
  NAND2_X1 U7603 ( .A1(n7523), .A2(n6883), .ZN(n6494) );
  NAND2_X1 U7604 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  NAND2_X1 U7605 ( .A1(n6492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6509) );
  XNOR2_X1 U7606 ( .A(n6509), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8851) );
  AOI22_X1 U7607 ( .A1(n6555), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6554), .B2(
        n8851), .ZN(n6493) );
  XNOR2_X1 U7608 ( .A(n8093), .B(n6280), .ZN(n6502) );
  NAND2_X1 U7609 ( .A1(n6561), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6501) );
  INV_X1 U7610 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8842) );
  OR2_X1 U7611 ( .A1(n6297), .A2(n8842), .ZN(n6500) );
  INV_X1 U7612 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8091) );
  OR2_X1 U7613 ( .A1(n6311), .A2(n8091), .ZN(n6499) );
  INV_X1 U7614 ( .A(n6495), .ZN(n6515) );
  NAND2_X1 U7615 ( .A1(n6496), .A2(n8102), .ZN(n6497) );
  NAND2_X1 U7616 ( .A1(n6515), .A2(n6497), .ZN(n8103) );
  OR2_X1 U7617 ( .A1(n4870), .A2(n8103), .ZN(n6498) );
  OR2_X1 U7618 ( .A1(n8781), .A2(n6715), .ZN(n6503) );
  NAND2_X1 U7619 ( .A1(n6502), .A2(n6503), .ZN(n6507) );
  INV_X1 U7620 ( .A(n6502), .ZN(n6505) );
  INV_X1 U7621 ( .A(n6503), .ZN(n6504) );
  NAND2_X1 U7622 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  AND2_X1 U7623 ( .A1(n6507), .A2(n6506), .ZN(n8100) );
  NAND2_X1 U7624 ( .A1(n8098), .A2(n6507), .ZN(n8772) );
  OR2_X1 U7625 ( .A1(n7592), .A2(n6640), .ZN(n6513) );
  NAND2_X1 U7626 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  NAND2_X1 U7627 ( .A1(n6510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6511) );
  XNOR2_X1 U7628 ( .A(n6511), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8863) );
  AOI22_X1 U7629 ( .A1(n6555), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6554), .B2(
        n8863), .ZN(n6512) );
  XNOR2_X1 U7630 ( .A(n8785), .B(n6280), .ZN(n6522) );
  NAND2_X1 U7631 ( .A1(n6561), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6521) );
  INV_X1 U7632 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6514) );
  OR2_X1 U7633 ( .A1(n6297), .A2(n6514), .ZN(n6520) );
  INV_X1 U7634 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8307) );
  OR2_X1 U7635 ( .A1(n6311), .A2(n8307), .ZN(n6519) );
  NAND2_X1 U7636 ( .A1(n6515), .A2(n8775), .ZN(n6516) );
  NAND2_X1 U7637 ( .A1(n6517), .A2(n6516), .ZN(n8779) );
  OR2_X1 U7638 ( .A1(n6309), .A2(n8779), .ZN(n6518) );
  OR2_X1 U7639 ( .A1(n8709), .A2(n6715), .ZN(n6523) );
  NAND2_X1 U7640 ( .A1(n6522), .A2(n6523), .ZN(n6527) );
  INV_X1 U7641 ( .A(n6522), .ZN(n6525) );
  INV_X1 U7642 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U7643 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  AND2_X1 U7644 ( .A1(n6527), .A2(n6526), .ZN(n8773) );
  NAND2_X1 U7645 ( .A1(n8771), .A2(n6527), .ZN(n8705) );
  NAND2_X1 U7646 ( .A1(n8706), .A2(n8705), .ZN(n8704) );
  NAND2_X1 U7647 ( .A1(n7829), .A2(n6883), .ZN(n6531) );
  OR2_X1 U7648 ( .A1(n4909), .A2(n6214), .ZN(n6529) );
  XNOR2_X1 U7649 ( .A(n6529), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8899) );
  AOI22_X1 U7650 ( .A1(n6555), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6554), .B2(
        n8899), .ZN(n6530) );
  XNOR2_X1 U7651 ( .A(n9237), .B(n6280), .ZN(n6539) );
  INV_X1 U7652 ( .A(n6546), .ZN(n6548) );
  NAND2_X1 U7653 ( .A1(n6533), .A2(n6532), .ZN(n6534) );
  NAND2_X1 U7654 ( .A1(n6548), .A2(n6534), .ZN(n9141) );
  OR2_X1 U7655 ( .A1(n9141), .A2(n6309), .ZN(n6538) );
  AOI22_X1 U7656 ( .A1(n6871), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n6535), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7657 ( .A1(n6561), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7658 ( .A1(n9124), .A2(n6302), .ZN(n6540) );
  AND2_X1 U7659 ( .A1(n6539), .A2(n6540), .ZN(n8713) );
  INV_X1 U7660 ( .A(n6539), .ZN(n6542) );
  INV_X1 U7661 ( .A(n6540), .ZN(n6541) );
  NAND2_X1 U7662 ( .A1(n6542), .A2(n6541), .ZN(n8714) );
  OAI21_X2 U7663 ( .B1(n8716), .B2(n8713), .A(n8714), .ZN(n8535) );
  XNOR2_X1 U7664 ( .A(n6543), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8917) );
  AOI22_X1 U7665 ( .A1(n6555), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6554), .B2(
        n8917), .ZN(n6544) );
  XNOR2_X1 U7666 ( .A(n9231), .B(n6325), .ZN(n8533) );
  INV_X1 U7667 ( .A(n6558), .ZN(n6559) );
  INV_X1 U7668 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U7669 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  AND2_X1 U7670 ( .A1(n6559), .A2(n6549), .ZN(n9119) );
  NAND2_X1 U7671 ( .A1(n9119), .A2(n6550), .ZN(n6553) );
  AOI22_X1 U7672 ( .A1(n6871), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n6535), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U7673 ( .A1(n6561), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6551) );
  OR2_X1 U7674 ( .A1(n8718), .A2(n6715), .ZN(n8532) );
  NAND2_X1 U7675 ( .A1(n7970), .A2(n6883), .ZN(n6557) );
  AOI22_X1 U7676 ( .A1(n6555), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9106), .B2(
        n6554), .ZN(n6556) );
  XNOR2_X1 U7677 ( .A(n6797), .B(n6325), .ZN(n6568) );
  INV_X1 U7678 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U7679 ( .A1(n6559), .A2(n7147), .ZN(n6560) );
  NAND2_X1 U7680 ( .A1(n6576), .A2(n6560), .ZN(n9105) );
  OR2_X1 U7681 ( .A1(n9105), .A2(n4870), .ZN(n6567) );
  INV_X1 U7682 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U7683 ( .A1(n6871), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U7684 ( .A1(n6561), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U7685 ( .C1(n6311), .C2(n6564), .A(n6563), .B(n6562), .ZN(n6565)
         );
  INV_X1 U7686 ( .A(n6565), .ZN(n6566) );
  NOR2_X1 U7687 ( .A1(n8736), .A2(n6715), .ZN(n6569) );
  NAND2_X1 U7688 ( .A1(n6568), .A2(n6569), .ZN(n6572) );
  INV_X1 U7689 ( .A(n6568), .ZN(n8733) );
  INV_X1 U7690 ( .A(n6569), .ZN(n6570) );
  NAND2_X1 U7691 ( .A1(n8733), .A2(n6570), .ZN(n6571) );
  NAND2_X1 U7692 ( .A1(n6572), .A2(n6571), .ZN(n8673) );
  NAND2_X1 U7693 ( .A1(n8015), .A2(n6883), .ZN(n6575) );
  INV_X1 U7694 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6573) );
  XNOR2_X1 U7695 ( .A(n9222), .B(n6325), .ZN(n6584) );
  NAND2_X1 U7696 ( .A1(n6576), .A2(n7270), .ZN(n6577) );
  AND2_X1 U7697 ( .A1(n6592), .A2(n6577), .ZN(n9095) );
  NAND2_X1 U7698 ( .A1(n9095), .A2(n6550), .ZN(n6583) );
  INV_X1 U7699 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U7700 ( .A1(n6871), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U7701 ( .A1(n6535), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6578) );
  OAI211_X1 U7702 ( .C1(n6580), .C2(n6295), .A(n6579), .B(n6578), .ZN(n6581)
         );
  INV_X1 U7703 ( .A(n6581), .ZN(n6582) );
  NOR2_X1 U7704 ( .A1(n9067), .A2(n6715), .ZN(n6585) );
  NAND2_X1 U7705 ( .A1(n6584), .A2(n6585), .ZN(n6589) );
  INV_X1 U7706 ( .A(n6584), .ZN(n8686) );
  INV_X1 U7707 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U7708 ( .A1(n8686), .A2(n6586), .ZN(n6587) );
  AND2_X1 U7709 ( .A1(n6589), .A2(n6587), .ZN(n8731) );
  NAND2_X1 U7710 ( .A1(n6588), .A2(n8731), .ZN(n8684) );
  NAND2_X1 U7711 ( .A1(n8684), .A2(n6589), .ZN(n6604) );
  INV_X1 U7712 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8058) );
  XNOR2_X1 U7713 ( .A(n9216), .B(n6325), .ZN(n8749) );
  INV_X1 U7714 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8690) );
  INV_X1 U7715 ( .A(n6607), .ZN(n6609) );
  NAND2_X1 U7716 ( .A1(n6592), .A2(n8690), .ZN(n6593) );
  NAND2_X1 U7717 ( .A1(n6609), .A2(n6593), .ZN(n9077) );
  OR2_X1 U7718 ( .A1(n9077), .A2(n6309), .ZN(n6599) );
  INV_X1 U7719 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7720 ( .A1(n6535), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7721 ( .A1(n6871), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6594) );
  OAI211_X1 U7722 ( .C1(n6596), .C2(n6295), .A(n6595), .B(n6594), .ZN(n6597)
         );
  INV_X1 U7723 ( .A(n6597), .ZN(n6598) );
  NAND2_X1 U7724 ( .A1(n6599), .A2(n6598), .ZN(n9056) );
  AND2_X1 U7725 ( .A1(n9056), .A2(n6302), .ZN(n6600) );
  NAND2_X1 U7726 ( .A1(n8749), .A2(n6600), .ZN(n6617) );
  INV_X1 U7727 ( .A(n8749), .ZN(n6602) );
  INV_X1 U7728 ( .A(n6600), .ZN(n6601) );
  NAND2_X1 U7729 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  AND2_X1 U7730 ( .A1(n6617), .A2(n6603), .ZN(n8683) );
  NAND2_X1 U7731 ( .A1(n6604), .A2(n8683), .ZN(n8687) );
  NAND2_X1 U7732 ( .A1(n8479), .A2(n6883), .ZN(n6606) );
  INV_X1 U7733 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8480) );
  XNOR2_X1 U7734 ( .A(n9210), .B(n6325), .ZN(n6619) );
  INV_X1 U7735 ( .A(n6626), .ZN(n6627) );
  INV_X1 U7736 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7737 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  NAND2_X1 U7738 ( .A1(n9050), .A2(n6550), .ZN(n6616) );
  INV_X1 U7739 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U7740 ( .A1(n6535), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7741 ( .A1(n6871), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6611) );
  OAI211_X1 U7742 ( .C1(n6613), .C2(n6295), .A(n6612), .B(n6611), .ZN(n6614)
         );
  INV_X1 U7743 ( .A(n6614), .ZN(n6615) );
  NOR2_X1 U7744 ( .A1(n9069), .A2(n6715), .ZN(n6620) );
  XNOR2_X1 U7745 ( .A(n6619), .B(n6620), .ZN(n8751) );
  INV_X1 U7746 ( .A(n6619), .ZN(n6622) );
  INV_X1 U7747 ( .A(n6620), .ZN(n6621) );
  NAND2_X1 U7748 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  NAND2_X1 U7749 ( .A1(n8333), .A2(n6883), .ZN(n6625) );
  INV_X1 U7750 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U7751 ( .A(n9204), .B(n6325), .ZN(n6635) );
  NAND2_X1 U7752 ( .A1(n6627), .A2(n8655), .ZN(n6628) );
  NAND2_X1 U7753 ( .A1(n6643), .A2(n6628), .ZN(n9037) );
  OR2_X1 U7754 ( .A1(n9037), .A2(n4870), .ZN(n6634) );
  INV_X1 U7755 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U7756 ( .A1(n6871), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U7757 ( .A1(n6535), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6629) );
  OAI211_X1 U7758 ( .C1(n6631), .C2(n6295), .A(n6630), .B(n6629), .ZN(n6632)
         );
  INV_X1 U7759 ( .A(n6632), .ZN(n6633) );
  NAND2_X1 U7760 ( .A1(n9057), .A2(n6302), .ZN(n8651) );
  INV_X1 U7761 ( .A(n6635), .ZN(n6636) );
  NAND2_X1 U7762 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  OR2_X1 U7763 ( .A1(n8435), .A2(n6640), .ZN(n6642) );
  INV_X1 U7764 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8432) );
  XNOR2_X1 U7765 ( .A(n9026), .B(n6280), .ZN(n6652) );
  NAND2_X1 U7766 ( .A1(n6643), .A2(n7179), .ZN(n6644) );
  NAND2_X1 U7767 ( .A1(n6658), .A2(n6644), .ZN(n9022) );
  OR2_X1 U7768 ( .A1(n9022), .A2(n6309), .ZN(n6650) );
  INV_X1 U7769 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7770 ( .A1(n6871), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U7771 ( .A1(n6535), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6645) );
  OAI211_X1 U7772 ( .C1(n6647), .C2(n6295), .A(n6646), .B(n6645), .ZN(n6648)
         );
  INV_X1 U7773 ( .A(n6648), .ZN(n6649) );
  NOR2_X1 U7774 ( .A1(n9033), .A2(n6715), .ZN(n6651) );
  NAND2_X1 U7775 ( .A1(n8723), .A2(n6651), .ZN(n8725) );
  INV_X1 U7776 ( .A(n6652), .ZN(n6653) );
  OR2_X1 U7777 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  NAND2_X1 U7778 ( .A1(n8453), .A2(n6883), .ZN(n6657) );
  INV_X1 U7779 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8455) );
  XNOR2_X1 U7780 ( .A(n9193), .B(n6325), .ZN(n6666) );
  NAND2_X1 U7781 ( .A1(n6658), .A2(n8700), .ZN(n6659) );
  AND2_X1 U7782 ( .A1(n6674), .A2(n6659), .ZN(n9007) );
  NAND2_X1 U7783 ( .A1(n9007), .A2(n6550), .ZN(n6665) );
  INV_X1 U7784 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U7785 ( .A1(n6535), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U7786 ( .A1(n6871), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6660) );
  OAI211_X1 U7787 ( .C1(n6295), .C2(n6662), .A(n6661), .B(n6660), .ZN(n6663)
         );
  INV_X1 U7788 ( .A(n6663), .ZN(n6664) );
  NOR2_X1 U7789 ( .A1(n9015), .A2(n6715), .ZN(n6667) );
  NAND2_X1 U7790 ( .A1(n6666), .A2(n6667), .ZN(n6670) );
  INV_X1 U7791 ( .A(n6666), .ZN(n8762) );
  INV_X1 U7792 ( .A(n6667), .ZN(n6668) );
  NAND2_X1 U7793 ( .A1(n8762), .A2(n6668), .ZN(n6669) );
  AND2_X1 U7794 ( .A1(n6670), .A2(n6669), .ZN(n8697) );
  NAND2_X1 U7795 ( .A1(n8696), .A2(n8697), .ZN(n8695) );
  NAND2_X1 U7796 ( .A1(n9279), .A2(n6883), .ZN(n6672) );
  INV_X1 U7797 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9281) );
  XNOR2_X1 U7798 ( .A(n9187), .B(n6325), .ZN(n6682) );
  INV_X1 U7799 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6673) );
  INV_X1 U7800 ( .A(n6689), .ZN(n6690) );
  NAND2_X1 U7801 ( .A1(n6674), .A2(n6673), .ZN(n6675) );
  NAND2_X1 U7802 ( .A1(n6690), .A2(n6675), .ZN(n8995) );
  OR2_X1 U7803 ( .A1(n8995), .A2(n4870), .ZN(n6681) );
  INV_X1 U7804 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6678) );
  NAND2_X1 U7805 ( .A1(n6871), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U7806 ( .A1(n6535), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6676) );
  OAI211_X1 U7807 ( .C1(n6678), .C2(n6295), .A(n6677), .B(n6676), .ZN(n6679)
         );
  INV_X1 U7808 ( .A(n6679), .ZN(n6680) );
  NOR2_X1 U7809 ( .A1(n8975), .A2(n6715), .ZN(n6683) );
  NAND2_X1 U7810 ( .A1(n6682), .A2(n6683), .ZN(n6686) );
  INV_X1 U7811 ( .A(n6682), .ZN(n8642) );
  INV_X1 U7812 ( .A(n6683), .ZN(n6684) );
  NAND2_X1 U7813 ( .A1(n8642), .A2(n6684), .ZN(n6685) );
  AND2_X1 U7814 ( .A1(n6686), .A2(n6685), .ZN(n8758) );
  NAND2_X1 U7815 ( .A1(n10200), .A2(n6883), .ZN(n6688) );
  INV_X1 U7816 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9278) );
  XNOR2_X1 U7817 ( .A(n9181), .B(n6325), .ZN(n6698) );
  INV_X1 U7818 ( .A(n6704), .ZN(n6706) );
  NAND2_X1 U7819 ( .A1(n6690), .A2(n8646), .ZN(n6691) );
  NAND2_X1 U7820 ( .A1(n6706), .A2(n6691), .ZN(n8969) );
  INV_X1 U7821 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U7822 ( .A1(n6535), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U7823 ( .A1(n6871), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6692) );
  OAI211_X1 U7824 ( .C1(n6295), .C2(n6694), .A(n6693), .B(n6692), .ZN(n6695)
         );
  INV_X1 U7825 ( .A(n6695), .ZN(n6696) );
  NOR2_X1 U7826 ( .A1(n8765), .A2(n6715), .ZN(n6699) );
  NAND2_X1 U7827 ( .A1(n6698), .A2(n6699), .ZN(n6703) );
  INV_X1 U7828 ( .A(n6698), .ZN(n6701) );
  INV_X1 U7829 ( .A(n6699), .ZN(n6700) );
  NAND2_X1 U7830 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  AND2_X1 U7831 ( .A1(n6703), .A2(n6702), .ZN(n8640) );
  INV_X1 U7832 ( .A(n8942), .ZN(n6708) );
  INV_X1 U7833 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U7834 ( .A1(n6706), .A2(n6705), .ZN(n6707) );
  NAND2_X1 U7835 ( .A1(n8962), .A2(n6550), .ZN(n6714) );
  INV_X1 U7836 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U7837 ( .A1(n6871), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U7838 ( .A1(n6535), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6709) );
  OAI211_X1 U7839 ( .C1(n6711), .C2(n6295), .A(n6710), .B(n6709), .ZN(n6712)
         );
  INV_X1 U7840 ( .A(n6712), .ZN(n6713) );
  OAI21_X1 U7841 ( .B1(n6715), .B2(n6325), .A(n8392), .ZN(n6716) );
  OAI21_X1 U7842 ( .B1(n6325), .B2(n8392), .A(n6716), .ZN(n6717) );
  NOR4_X1 U7843 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6726) );
  NOR4_X1 U7844 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6725) );
  NOR4_X1 U7845 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6721) );
  NOR4_X1 U7846 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6720) );
  NOR4_X1 U7847 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6719) );
  NOR4_X1 U7848 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6718) );
  NAND4_X1 U7849 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6722)
         );
  NOR4_X1 U7850 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6723), .A4(n6722), .ZN(n6724) );
  AND3_X1 U7851 ( .A1(n6726), .A2(n6725), .A3(n6724), .ZN(n6740) );
  NAND2_X1 U7852 ( .A1(n6727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U7853 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6728), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6730) );
  OR2_X1 U7854 ( .A1(n6731), .A2(n6214), .ZN(n6732) );
  INV_X1 U7855 ( .A(n10343), .ZN(n8433) );
  INV_X1 U7856 ( .A(P2_B_REG_SCAN_IN), .ZN(n6842) );
  AOI22_X1 U7857 ( .A1(P2_B_REG_SCAN_IN), .A2(n8433), .B1(n10343), .B2(n6842), 
        .ZN(n6738) );
  OR2_X1 U7858 ( .A1(n10343), .A2(n10342), .ZN(n6742) );
  OR2_X1 U7859 ( .A1(n10243), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6741) );
  OR2_X1 U7860 ( .A1(n10243), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6744) );
  OR2_X1 U7861 ( .A1(n10342), .A2(n10241), .ZN(n6743) );
  NAND2_X1 U7862 ( .A1(n6744), .A2(n6743), .ZN(n7558) );
  OR2_X1 U7863 ( .A1(n7560), .A2(n7558), .ZN(n6745) );
  XNOR2_X1 U7864 ( .A(n6748), .B(n6747), .ZN(n7055) );
  INV_X1 U7865 ( .A(n10347), .ZN(n6749) );
  NAND2_X1 U7866 ( .A1(n6750), .A2(n8993), .ZN(n6769) );
  INV_X1 U7867 ( .A(n8150), .ZN(n8156) );
  NAND2_X1 U7868 ( .A1(n10611), .A2(n8156), .ZN(n6752) );
  OR2_X1 U7869 ( .A1(n10242), .A2(n6752), .ZN(n6753) );
  NAND2_X1 U7870 ( .A1(n9274), .A2(n6883), .ZN(n6755) );
  INV_X1 U7871 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U7872 ( .A1(n6756), .A2(n6751), .ZN(n7577) );
  OR2_X1 U7873 ( .A1(n10242), .A2(n7577), .ZN(n6758) );
  NAND2_X1 U7874 ( .A1(n9106), .A2(n6259), .ZN(n6757) );
  NAND2_X1 U7875 ( .A1(n10391), .A2(n8057), .ZN(n6851) );
  INV_X1 U7876 ( .A(n8765), .ZN(n8954) );
  OR2_X1 U7877 ( .A1(n10242), .A2(n6769), .ZN(n6762) );
  AOI22_X1 U7878 ( .A1(n8954), .A2(n10372), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6774) );
  INV_X1 U7879 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U7880 ( .A1(n6871), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U7881 ( .A1(n6535), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6764) );
  OAI211_X1 U7882 ( .C1(n6766), .C2(n6295), .A(n6765), .B(n6764), .ZN(n6767)
         );
  AOI21_X1 U7883 ( .B1(n8942), .B2(n6550), .A(n6767), .ZN(n8368) );
  INV_X1 U7884 ( .A(n8368), .ZN(n8955) );
  NAND2_X1 U7885 ( .A1(n6768), .A2(n6851), .ZN(n6772) );
  NAND2_X1 U7886 ( .A1(n6769), .A2(n8150), .ZN(n6770) );
  NAND2_X1 U7887 ( .A1(n6770), .A2(n7055), .ZN(n7057) );
  NOR2_X1 U7888 ( .A1(n8148), .A2(n7057), .ZN(n6771) );
  NAND2_X1 U7889 ( .A1(n6772), .A2(n6771), .ZN(n7420) );
  AOI22_X1 U7890 ( .A1(n8955), .A2(n10373), .B1(n8962), .B2(n8740), .ZN(n6773)
         );
  INV_X1 U7891 ( .A(n8709), .ZN(n8439) );
  INV_X1 U7892 ( .A(n8128), .ZN(n8135) );
  NAND2_X1 U7893 ( .A1(n4868), .A2(n7613), .ZN(n6776) );
  NAND2_X1 U7894 ( .A1(n7612), .A2(n6776), .ZN(n6778) );
  NAND2_X1 U7895 ( .A1(n6779), .A2(n10374), .ZN(n6915) );
  INV_X1 U7896 ( .A(n10386), .ZN(n10374) );
  OAI22_X2 U7897 ( .A1(n9151), .A2(n9159), .B1(n10374), .B2(n8662), .ZN(n7557)
         );
  NAND2_X1 U7898 ( .A1(n10451), .A2(n6781), .ZN(n6921) );
  NAND2_X1 U7899 ( .A1(n7557), .A2(n6818), .ZN(n6783) );
  OR2_X1 U7900 ( .A1(n10451), .A2(n10402), .ZN(n6782) );
  NAND2_X1 U7901 ( .A1(n6783), .A2(n6782), .ZN(n10442) );
  XNOR2_X1 U7902 ( .A(n8663), .B(n10462), .ZN(n10447) );
  NOR2_X1 U7903 ( .A1(n8663), .A2(n7515), .ZN(n6927) );
  INV_X1 U7904 ( .A(n6927), .ZN(n6784) );
  NAND2_X1 U7905 ( .A1(n7662), .A2(n10449), .ZN(n6931) );
  NAND2_X1 U7906 ( .A1(n8570), .A2(n8561), .ZN(n6930) );
  NAND2_X1 U7907 ( .A1(n7527), .A2(n10449), .ZN(n6785) );
  NAND2_X1 U7908 ( .A1(n6786), .A2(n6785), .ZN(n7633) );
  INV_X1 U7909 ( .A(n8328), .ZN(n7672) );
  OR2_X1 U7910 ( .A1(n7634), .A2(n7672), .ZN(n6787) );
  NAND2_X1 U7911 ( .A1(n7633), .A2(n6787), .ZN(n6789) );
  NAND2_X1 U7912 ( .A1(n7634), .A2(n7672), .ZN(n6788) );
  NAND2_X1 U7913 ( .A1(n6789), .A2(n6788), .ZN(n7669) );
  OR2_X1 U7914 ( .A1(n7792), .A2(n8556), .ZN(n6941) );
  NAND2_X1 U7915 ( .A1(n7792), .A2(n8556), .ZN(n6940) );
  NAND2_X1 U7916 ( .A1(n6941), .A2(n6940), .ZN(n7668) );
  INV_X1 U7917 ( .A(n7668), .ZN(n6790) );
  INV_X1 U7918 ( .A(n8556), .ZN(n7685) );
  OR2_X1 U7919 ( .A1(n7792), .A2(n7685), .ZN(n6791) );
  OR2_X1 U7920 ( .A1(n7695), .A2(n8468), .ZN(n6944) );
  NAND2_X1 U7921 ( .A1(n7695), .A2(n8468), .ZN(n6945) );
  INV_X1 U7922 ( .A(n7691), .ZN(n6792) );
  INV_X1 U7923 ( .A(n8468), .ZN(n8459) );
  NAND2_X1 U7924 ( .A1(n7695), .A2(n8459), .ZN(n6793) );
  OR2_X1 U7925 ( .A1(n8476), .A2(n8315), .ZN(n7884) );
  NAND2_X1 U7926 ( .A1(n8476), .A2(n8315), .ZN(n6823) );
  NAND2_X1 U7927 ( .A1(n7884), .A2(n6823), .ZN(n7885) );
  NAND2_X1 U7928 ( .A1(n7817), .A2(n7885), .ZN(n7816) );
  INV_X1 U7929 ( .A(n8315), .ZN(n7686) );
  OR2_X1 U7930 ( .A1(n8476), .A2(n7686), .ZN(n6794) );
  OR2_X1 U7931 ( .A1(n7900), .A2(n8460), .ZN(n6950) );
  NAND2_X1 U7932 ( .A1(n7900), .A2(n8460), .ZN(n6824) );
  NAND2_X1 U7933 ( .A1(n6950), .A2(n6824), .ZN(n7887) );
  INV_X1 U7934 ( .A(n7900), .ZN(n10598) );
  OR2_X1 U7935 ( .A1(n7877), .A2(n8322), .ZN(n6951) );
  NAND2_X1 U7936 ( .A1(n7877), .A2(n8322), .ZN(n6952) );
  INV_X1 U7937 ( .A(n8322), .ZN(n7987) );
  OR2_X1 U7938 ( .A1(n8000), .A2(n8326), .ZN(n6904) );
  NAND2_X1 U7939 ( .A1(n8000), .A2(n8326), .ZN(n6905) );
  NAND2_X1 U7940 ( .A1(n6904), .A2(n6905), .ZN(n7961) );
  OR2_X1 U7941 ( .A1(n8128), .A2(n8338), .ZN(n6959) );
  NAND2_X1 U7942 ( .A1(n8128), .A2(n8338), .ZN(n6960) );
  INV_X1 U7943 ( .A(n8122), .ZN(n8119) );
  OAI21_X1 U7944 ( .B1(n8135), .B2(n8338), .A(n8118), .ZN(n8084) );
  NAND2_X1 U7945 ( .A1(n8093), .A2(n8781), .ZN(n6900) );
  INV_X1 U7946 ( .A(n8781), .ZN(n8124) );
  OAI22_X1 U7947 ( .A1(n8084), .A2(n8086), .B1(n8093), .B2(n8124), .ZN(n8304)
         );
  OR2_X1 U7948 ( .A1(n8785), .A2(n8709), .ZN(n6964) );
  NAND2_X1 U7949 ( .A1(n8785), .A2(n8709), .ZN(n6965) );
  NAND2_X1 U7950 ( .A1(n8304), .A2(n8303), .ZN(n8302) );
  OAI21_X1 U7951 ( .B1(n8439), .B2(n8785), .A(n8302), .ZN(n8442) );
  OR2_X1 U7952 ( .A1(n9242), .A2(n8777), .ZN(n6898) );
  NAND2_X1 U7953 ( .A1(n9242), .A2(n8777), .ZN(n6899) );
  NAND2_X1 U7954 ( .A1(n9237), .A2(n8345), .ZN(n6897) );
  NAND2_X1 U7955 ( .A1(n6796), .A2(n8718), .ZN(n6973) );
  INV_X1 U7956 ( .A(n9231), .ZN(n9121) );
  NAND2_X1 U7957 ( .A1(n6797), .A2(n8736), .ZN(n6895) );
  INV_X1 U7958 ( .A(n8736), .ZN(n9125) );
  OAI22_X1 U7959 ( .A1(n9102), .A2(n9110), .B1(n6797), .B2(n9125), .ZN(n9090)
         );
  NAND2_X1 U7960 ( .A1(n9222), .A2(n9067), .ZN(n6981) );
  INV_X1 U7961 ( .A(n9067), .ZN(n8678) );
  NAND2_X1 U7962 ( .A1(n9216), .A2(n9056), .ZN(n6798) );
  NAND2_X1 U7963 ( .A1(n6799), .A2(n6798), .ZN(n7044) );
  NAND2_X1 U7964 ( .A1(n9210), .A2(n9069), .ZN(n6994) );
  NAND2_X1 U7965 ( .A1(n6988), .A2(n6994), .ZN(n7046) );
  INV_X1 U7966 ( .A(n9210), .ZN(n9052) );
  OR2_X1 U7967 ( .A1(n9204), .A2(n9014), .ZN(n6996) );
  NAND2_X1 U7968 ( .A1(n9204), .A2(n9014), .ZN(n6990) );
  NAND2_X1 U7969 ( .A1(n6996), .A2(n6990), .ZN(n9041) );
  NAND2_X1 U7970 ( .A1(n9197), .A2(n9033), .ZN(n6999) );
  INV_X1 U7971 ( .A(n9033), .ZN(n8724) );
  NAND2_X1 U7972 ( .A1(n9193), .A2(n9015), .ZN(n7003) );
  INV_X1 U7973 ( .A(n9193), .ZN(n9010) );
  INV_X1 U7974 ( .A(n9015), .ZN(n6801) );
  OR2_X1 U7975 ( .A1(n9187), .A2(n8975), .ZN(n7008) );
  NAND2_X1 U7976 ( .A1(n9187), .A2(n8975), .ZN(n7007) );
  NAND2_X1 U7977 ( .A1(n7008), .A2(n7007), .ZN(n8983) );
  INV_X1 U7978 ( .A(n8983), .ZN(n8986) );
  INV_X1 U7979 ( .A(n8975), .ZN(n8699) );
  NAND2_X1 U7980 ( .A1(n9181), .A2(n8765), .ZN(n7014) );
  INV_X1 U7981 ( .A(n9181), .ZN(n8972) );
  INV_X1 U7982 ( .A(n6804), .ZN(n6805) );
  NAND2_X1 U7983 ( .A1(n6805), .A2(n7191), .ZN(n6806) );
  NAND2_X1 U7984 ( .A1(n6807), .A2(n6806), .ZN(n6863) );
  INV_X1 U7985 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9272) );
  INV_X1 U7986 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U7987 ( .A(n9272), .B(n10191), .S(n7285), .Z(n6808) );
  NAND2_X1 U7988 ( .A1(n6808), .A2(n7187), .ZN(n6864) );
  INV_X1 U7989 ( .A(n6808), .ZN(n6809) );
  NAND2_X1 U7990 ( .A1(n6809), .A2(SI_29_), .ZN(n6810) );
  NAND2_X1 U7991 ( .A1(n9271), .A2(n6883), .ZN(n6812) );
  NAND2_X1 U7992 ( .A1(n8941), .A2(n8368), .ZN(n7023) );
  MUX2_X1 U7993 ( .A(n8156), .B(n7058), .S(n6756), .Z(n6814) );
  NOR2_X1 U7994 ( .A1(n6751), .A2(n9106), .ZN(n6813) );
  NAND2_X1 U7995 ( .A1(n6814), .A2(n6813), .ZN(n7892) );
  NAND2_X1 U7996 ( .A1(n4868), .A2(n6847), .ZN(n6816) );
  OR2_X1 U7997 ( .A1(n7424), .A2(n7622), .ZN(n7614) );
  NAND2_X1 U7998 ( .A1(n7424), .A2(n7622), .ZN(n7500) );
  NAND2_X1 U7999 ( .A1(n7500), .A2(n6816), .ZN(n6910) );
  NAND2_X1 U8000 ( .A1(n6910), .A2(n6817), .ZN(n6911) );
  INV_X1 U8001 ( .A(n6818), .ZN(n6819) );
  INV_X1 U8002 ( .A(n8663), .ZN(n8320) );
  OR2_X1 U8003 ( .A1(n7634), .A2(n8328), .ZN(n6935) );
  NAND2_X1 U8004 ( .A1(n7628), .A2(n6935), .ZN(n6821) );
  NAND2_X1 U8005 ( .A1(n7634), .A2(n8328), .ZN(n6934) );
  NAND2_X1 U8006 ( .A1(n6950), .A2(n7884), .ZN(n6947) );
  INV_X1 U8007 ( .A(n6947), .ZN(n6822) );
  AND2_X1 U8008 ( .A1(n6824), .A2(n6823), .ZN(n6949) );
  INV_X1 U8009 ( .A(n6949), .ZN(n6825) );
  NAND2_X1 U8010 ( .A1(n6825), .A2(n6950), .ZN(n6953) );
  NAND2_X1 U8011 ( .A1(n6826), .A2(n6952), .ZN(n7959) );
  INV_X1 U8012 ( .A(n7961), .ZN(n7041) );
  NAND2_X1 U8013 ( .A1(n7959), .A2(n7041), .ZN(n6827) );
  NAND2_X1 U8014 ( .A1(n6827), .A2(n6905), .ZN(n8121) );
  INV_X1 U8015 ( .A(n6960), .ZN(n6828) );
  NAND2_X1 U8016 ( .A1(n8437), .A2(n6899), .ZN(n6829) );
  NAND2_X1 U8017 ( .A1(n6829), .A2(n6898), .ZN(n9131) );
  NAND2_X1 U8018 ( .A1(n9131), .A2(n9133), .ZN(n6830) );
  NAND2_X1 U8019 ( .A1(n6830), .A2(n6896), .ZN(n9122) );
  INV_X1 U8020 ( .A(n9056), .ZN(n8752) );
  OR2_X1 U8021 ( .A1(n9216), .A2(n8752), .ZN(n6832) );
  INV_X1 U8022 ( .A(n9013), .ZN(n6835) );
  NAND2_X1 U8023 ( .A1(n6835), .A2(n6834), .ZN(n9017) );
  NAND2_X1 U8024 ( .A1(n8978), .A2(n7013), .ZN(n8953) );
  NAND2_X1 U8025 ( .A1(n8953), .A2(n8952), .ZN(n8951) );
  INV_X1 U8026 ( .A(n8392), .ZN(n8976) );
  OR2_X1 U8027 ( .A1(n9176), .A2(n8976), .ZN(n6837) );
  NAND2_X1 U8028 ( .A1(n6756), .A2(n5392), .ZN(n6890) );
  NAND2_X1 U8029 ( .A1(n9106), .A2(n7058), .ZN(n7034) );
  NAND2_X1 U8030 ( .A1(n8392), .A2(n10450), .ZN(n6845) );
  INV_X1 U8031 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8032 ( .A1(n6535), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U8033 ( .A1(n6871), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6838) );
  OAI211_X1 U8034 ( .C1(n6295), .C2(n6840), .A(n6839), .B(n6838), .ZN(n6886)
         );
  OR2_X1 U8035 ( .A1(n6841), .A2(n6842), .ZN(n6843) );
  AND2_X1 U8036 ( .A1(n10448), .A2(n6843), .ZN(n8931) );
  NAND2_X1 U8037 ( .A1(n6886), .A2(n8931), .ZN(n6844) );
  INV_X1 U8038 ( .A(n6797), .ZN(n9103) );
  INV_X1 U8039 ( .A(n7877), .ZN(n7952) );
  INV_X1 U8040 ( .A(n7695), .ZN(n10574) );
  NAND2_X1 U8041 ( .A1(n6847), .A2(n7622), .ZN(n9156) );
  NAND2_X1 U8042 ( .A1(n10443), .A2(n10462), .ZN(n10445) );
  INV_X1 U8043 ( .A(n7792), .ZN(n7676) );
  OR2_X2 U8044 ( .A1(n8093), .A2(n8090), .ZN(n8305) );
  NAND2_X1 U8045 ( .A1(n9103), .A2(n9118), .ZN(n9094) );
  OR2_X2 U8046 ( .A1(n9094), .A2(n9222), .ZN(n9092) );
  NAND2_X1 U8047 ( .A1(n9034), .A2(n9026), .ZN(n9006) );
  NOR2_X2 U8048 ( .A1(n9006), .A2(n9193), .ZN(n8990) );
  AOI21_X1 U8049 ( .B1(n8941), .B2(n8961), .A(n8935), .ZN(n8946) );
  AOI22_X1 U8050 ( .A1(n8946), .A2(n10404), .B1(n10403), .B2(n8941), .ZN(n6849) );
  NOR2_X1 U8051 ( .A1(n7057), .A2(P2_U3152), .ZN(n7562) );
  INV_X1 U8052 ( .A(n8148), .ZN(n7559) );
  NAND4_X1 U8053 ( .A1(n7562), .A2(n7558), .A3(n7559), .A4(n6851), .ZN(n6852)
         );
  NOR2_X4 U8054 ( .A1(n6857), .A2(n7560), .ZN(n10620) );
  NAND2_X1 U8055 ( .A1(n6858), .A2(n10620), .ZN(n6855) );
  INV_X1 U8056 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6853) );
  OR2_X1 U8057 ( .A1(n10620), .A2(n6853), .ZN(n6854) );
  NAND2_X1 U8058 ( .A1(n6855), .A2(n6854), .ZN(P2_U3549) );
  INV_X1 U8059 ( .A(n7560), .ZN(n6856) );
  NAND2_X1 U8060 ( .A1(n6858), .A2(n10624), .ZN(n6860) );
  OR2_X1 U8061 ( .A1(n10624), .A2(n6766), .ZN(n6859) );
  NAND2_X1 U8062 ( .A1(n6860), .A2(n6859), .ZN(P2_U3517) );
  NAND2_X1 U8063 ( .A1(n6863), .A2(n6862), .ZN(n6865) );
  NAND2_X1 U8064 ( .A1(n6865), .A2(n6864), .ZN(n6876) );
  INV_X1 U8065 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8528) );
  INV_X1 U8066 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9495) );
  MUX2_X1 U8067 ( .A(n8528), .B(n9495), .S(n7284), .Z(n6866) );
  NAND2_X1 U8068 ( .A1(n6866), .A2(n7186), .ZN(n6877) );
  INV_X1 U8069 ( .A(n6866), .ZN(n6867) );
  NAND2_X1 U8070 ( .A1(n6867), .A2(SI_30_), .ZN(n6868) );
  XNOR2_X1 U8071 ( .A(n6876), .B(n6875), .ZN(n9494) );
  NAND2_X1 U8072 ( .A1(n9494), .A2(n6883), .ZN(n6870) );
  AND2_X1 U8073 ( .A1(n9175), .A2(n6886), .ZN(n7020) );
  INV_X1 U8074 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8075 ( .A1(n6535), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8076 ( .A1(n6871), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6872) );
  OAI211_X1 U8077 ( .C1(n6295), .C2(n6874), .A(n6873), .B(n6872), .ZN(n8932)
         );
  NAND2_X1 U8078 ( .A1(n6876), .A2(n6875), .ZN(n6878) );
  NAND2_X1 U8079 ( .A1(n6878), .A2(n6877), .ZN(n6882) );
  MUX2_X1 U8080 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7285), .Z(n6880) );
  INV_X1 U8081 ( .A(SI_31_), .ZN(n6879) );
  XNOR2_X1 U8082 ( .A(n6880), .B(n6879), .ZN(n6881) );
  NAND2_X1 U8083 ( .A1(n10189), .A2(n6883), .ZN(n6885) );
  INV_X1 U8084 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9270) );
  INV_X1 U8085 ( .A(n6886), .ZN(n8342) );
  NAND2_X1 U8086 ( .A1(n8937), .A2(n8342), .ZN(n7025) );
  NOR2_X1 U8087 ( .A1(n9170), .A2(n8932), .ZN(n6893) );
  AOI21_X1 U8088 ( .B1(n6888), .B2(n7051), .A(n6893), .ZN(n6889) );
  XNOR2_X1 U8089 ( .A(n6889), .B(n8993), .ZN(n6892) );
  NAND2_X1 U8090 ( .A1(n6302), .A2(n6890), .ZN(n6891) );
  NAND2_X1 U8091 ( .A1(n6892), .A2(n6891), .ZN(n7054) );
  NOR2_X1 U8092 ( .A1(n6893), .A2(n7020), .ZN(n7052) );
  NOR2_X1 U8093 ( .A1(n8993), .A2(n8057), .ZN(n7565) );
  NAND2_X1 U8094 ( .A1(n7565), .A2(n6259), .ZN(n7028) );
  INV_X1 U8095 ( .A(n7028), .ZN(n7021) );
  MUX2_X1 U8096 ( .A(n6895), .B(n6894), .S(n7021), .Z(n6979) );
  MUX2_X1 U8097 ( .A(n6897), .B(n6896), .S(n7028), .Z(n6972) );
  MUX2_X1 U8098 ( .A(n6899), .B(n6898), .S(n7021), .Z(n6970) );
  INV_X1 U8099 ( .A(n6900), .ZN(n6902) );
  MUX2_X1 U8100 ( .A(n6902), .B(n5345), .S(n7021), .Z(n6968) );
  NAND2_X1 U8101 ( .A1(n6905), .A2(n6952), .ZN(n6903) );
  NAND2_X1 U8102 ( .A1(n6903), .A2(n6904), .ZN(n6908) );
  NAND2_X1 U8103 ( .A1(n6904), .A2(n6951), .ZN(n6906) );
  NAND2_X1 U8104 ( .A1(n6906), .A2(n6905), .ZN(n6907) );
  MUX2_X1 U8105 ( .A(n6908), .B(n6907), .S(n7021), .Z(n6958) );
  INV_X1 U8106 ( .A(n6911), .ZN(n6912) );
  MUX2_X1 U8107 ( .A(n6913), .B(n6912), .S(n7021), .Z(n6914) );
  NAND2_X1 U8108 ( .A1(n6914), .A2(n9159), .ZN(n6920) );
  INV_X1 U8109 ( .A(n6915), .ZN(n6916) );
  MUX2_X1 U8110 ( .A(n6917), .B(n6916), .S(n7028), .Z(n6918) );
  NOR2_X1 U8111 ( .A1(n6918), .A2(n6818), .ZN(n6919) );
  INV_X1 U8112 ( .A(n6921), .ZN(n6924) );
  INV_X1 U8113 ( .A(n6922), .ZN(n6923) );
  MUX2_X1 U8114 ( .A(n6924), .B(n6923), .S(n7021), .Z(n6925) );
  INV_X1 U8115 ( .A(n6925), .ZN(n6926) );
  MUX2_X1 U8116 ( .A(n7515), .B(n8663), .S(n7028), .Z(n6928) );
  NAND2_X1 U8117 ( .A1(n6929), .A2(n7527), .ZN(n6933) );
  AND2_X1 U8118 ( .A1(n6935), .A2(n6934), .ZN(n7632) );
  MUX2_X1 U8119 ( .A(n6931), .B(n6930), .S(n7028), .Z(n6932) );
  NAND3_X1 U8120 ( .A1(n6933), .A2(n7632), .A3(n6932), .ZN(n6939) );
  INV_X1 U8121 ( .A(n6935), .ZN(n6936) );
  MUX2_X1 U8122 ( .A(n5349), .B(n6936), .S(n7028), .Z(n6937) );
  NOR2_X1 U8123 ( .A1(n7668), .A2(n6937), .ZN(n6938) );
  NAND2_X1 U8124 ( .A1(n6939), .A2(n6938), .ZN(n6943) );
  MUX2_X1 U8125 ( .A(n6941), .B(n6940), .S(n7028), .Z(n6942) );
  MUX2_X1 U8126 ( .A(n6945), .B(n6944), .S(n7028), .Z(n6946) );
  NAND2_X1 U8127 ( .A1(n6947), .A2(n7021), .ZN(n6948) );
  NAND2_X1 U8128 ( .A1(n6951), .A2(n6950), .ZN(n6955) );
  NAND2_X1 U8129 ( .A1(n6953), .A2(n6952), .ZN(n6954) );
  MUX2_X1 U8130 ( .A(n6955), .B(n6954), .S(n7021), .Z(n6956) );
  NAND3_X1 U8131 ( .A1(n8122), .A2(n6958), .A3(n6957), .ZN(n6962) );
  MUX2_X1 U8132 ( .A(n6960), .B(n6959), .S(n7028), .Z(n6961) );
  NAND3_X1 U8133 ( .A1(n8086), .A2(n6962), .A3(n6961), .ZN(n6963) );
  NAND2_X1 U8134 ( .A1(n8299), .A2(n6963), .ZN(n6967) );
  MUX2_X1 U8135 ( .A(n6965), .B(n6964), .S(n7028), .Z(n6966) );
  OAI211_X1 U8136 ( .C1(n6968), .C2(n6967), .A(n8443), .B(n6966), .ZN(n6969)
         );
  NAND3_X1 U8137 ( .A1(n9133), .A2(n6970), .A3(n6969), .ZN(n6971) );
  NAND3_X1 U8138 ( .A1(n6831), .A2(n6972), .A3(n6971), .ZN(n6976) );
  MUX2_X1 U8139 ( .A(n6974), .B(n6973), .S(n7028), .Z(n6975) );
  NAND2_X1 U8140 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  NAND2_X1 U8141 ( .A1(n9110), .A2(n6977), .ZN(n6978) );
  MUX2_X1 U8142 ( .A(n6981), .B(n6980), .S(n7028), .Z(n6982) );
  NAND2_X1 U8143 ( .A1(n9216), .A2(n7021), .ZN(n6984) );
  OR2_X1 U8144 ( .A1(n9216), .A2(n7021), .ZN(n6983) );
  MUX2_X1 U8145 ( .A(n6984), .B(n6983), .S(n9056), .Z(n6985) );
  NOR2_X1 U8146 ( .A1(n6986), .A2(n7046), .ZN(n6987) );
  INV_X1 U8147 ( .A(n6988), .ZN(n6989) );
  NAND2_X1 U8148 ( .A1(n6991), .A2(n9026), .ZN(n6992) );
  OAI21_X1 U8149 ( .B1(n9033), .B2(n6993), .A(n6992), .ZN(n7002) );
  INV_X1 U8150 ( .A(n6994), .ZN(n6997) );
  OAI211_X1 U8151 ( .C1(n6998), .C2(n6997), .A(n6996), .B(n6995), .ZN(n7000)
         );
  NAND2_X1 U8152 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  AND2_X1 U8153 ( .A1(n7007), .A2(n7003), .ZN(n7006) );
  AND2_X1 U8154 ( .A1(n7008), .A2(n7004), .ZN(n7005) );
  MUX2_X1 U8155 ( .A(n7006), .B(n7005), .S(n7028), .Z(n7012) );
  INV_X1 U8156 ( .A(n7007), .ZN(n7010) );
  INV_X1 U8157 ( .A(n7008), .ZN(n7009) );
  MUX2_X1 U8158 ( .A(n7010), .B(n7009), .S(n7021), .Z(n7011) );
  MUX2_X1 U8159 ( .A(n7014), .B(n7013), .S(n7021), .Z(n7015) );
  OR3_X1 U8160 ( .A1(n9176), .A2(n8976), .A3(n7021), .ZN(n7017) );
  NAND3_X1 U8161 ( .A1(n9176), .A2(n8976), .A3(n7021), .ZN(n7016) );
  NAND4_X1 U8162 ( .A1(n7019), .A2(n7018), .A3(n7017), .A4(n7016), .ZN(n7027)
         );
  INV_X1 U8163 ( .A(n7020), .ZN(n7026) );
  MUX2_X1 U8164 ( .A(n7023), .B(n7022), .S(n7021), .Z(n7024) );
  NAND4_X1 U8165 ( .A1(n7027), .A2(n7026), .A3(n7025), .A4(n7024), .ZN(n7032)
         );
  INV_X1 U8166 ( .A(n9170), .ZN(n7029) );
  NAND2_X1 U8167 ( .A1(n7029), .A2(n8932), .ZN(n7031) );
  MUX2_X1 U8168 ( .A(n7029), .B(n8932), .S(n7028), .Z(n7030) );
  INV_X1 U8169 ( .A(n8952), .ZN(n8958) );
  INV_X1 U8170 ( .A(n8443), .ZN(n8438) );
  INV_X1 U8171 ( .A(n7527), .ZN(n7529) );
  INV_X1 U8172 ( .A(n7036), .ZN(n7616) );
  NAND4_X1 U8173 ( .A1(n7616), .A2(n9159), .A3(n6756), .A4(n7500), .ZN(n7037)
         );
  NOR4_X1 U8174 ( .A1(n10447), .A2(n7529), .A3(n7037), .A4(n6818), .ZN(n7038)
         );
  NAND4_X1 U8175 ( .A1(n6790), .A2(n7632), .A3(n7691), .A4(n7038), .ZN(n7039)
         );
  NOR4_X1 U8176 ( .A1(n5067), .A2(n7887), .A3(n7885), .A4(n7039), .ZN(n7040)
         );
  NAND4_X1 U8177 ( .A1(n8086), .A2(n8122), .A3(n7041), .A4(n7040), .ZN(n7042)
         );
  NOR4_X1 U8178 ( .A1(n9116), .A2(n8438), .A3(n8303), .A4(n7042), .ZN(n7043)
         );
  NAND4_X1 U8179 ( .A1(n7044), .A2(n9110), .A3(n9133), .A4(n7043), .ZN(n7045)
         );
  NOR4_X1 U8180 ( .A1(n9020), .A2(n7046), .A3(n5339), .A4(n7045), .ZN(n7047)
         );
  NAND4_X1 U8181 ( .A1(n8986), .A2(n9001), .A3(n6833), .A4(n7047), .ZN(n7048)
         );
  NAND3_X1 U8182 ( .A1(n7052), .A2(n7051), .A3(n7050), .ZN(n7053) );
  OR2_X1 U8183 ( .A1(n7055), .A2(P2_U3152), .ZN(n8330) );
  NOR4_X1 U8184 ( .A1(n10242), .A2(n7057), .A3(n6841), .A4(n9066), .ZN(n7060)
         );
  OAI21_X1 U8185 ( .B1(n8330), .B2(n7058), .A(P2_B_REG_SCAN_IN), .ZN(n7059) );
  OR2_X1 U8186 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  NAND2_X1 U8187 ( .A1(n7062), .A2(n7061), .ZN(P2_U3244) );
  NOR2_X1 U8188 ( .A1(n9342), .A2(n9817), .ZN(n7066) );
  OAI22_X1 U8189 ( .A1(n9405), .A2(n9818), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7064), .ZN(n7065) );
  AOI211_X1 U8190 ( .C1(n9813), .C2(n9402), .A(n7066), .B(n7065), .ZN(n7068)
         );
  NAND2_X1 U8191 ( .A1(n10074), .A2(n9408), .ZN(n7067) );
  INV_X1 U8192 ( .A(n7070), .ZN(n8334) );
  NAND2_X1 U8193 ( .A1(n7069), .A2(n6163), .ZN(n7071) );
  NAND2_X1 U8194 ( .A1(n7071), .A2(n7070), .ZN(n10288) );
  NAND2_X1 U8195 ( .A1(n10288), .A2(n4872), .ZN(n7072) );
  NAND2_X1 U8196 ( .A1(n7072), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U8197 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U8198 ( .A(n7073), .ZN(n7074) );
  AOI211_X1 U8199 ( .C1(n7076), .C2(n7075), .A(n8759), .B(n7074), .ZN(n7080)
         );
  NOR2_X1 U8200 ( .A1(n10598), .A2(n8743), .ZN(n7079) );
  OAI22_X1 U8201 ( .A1(n8778), .A2(n8322), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6432), .ZN(n7078) );
  OAI22_X1 U8202 ( .A1(n8782), .A2(n8315), .B1(n8780), .B2(n7893), .ZN(n7077)
         );
  OR4_X1 U8203 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(P2_U3219)
         );
  NAND2_X1 U8204 ( .A1(n8148), .A2(n10347), .ZN(n7283) );
  XNOR2_X1 U8205 ( .A(n10383), .B(keyinput_59), .ZN(n7175) );
  OAI22_X1 U8206 ( .A1(n6608), .A2(keyinput_57), .B1(keyinput_56), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n7081) );
  AOI221_X1 U8207 ( .B1(n6608), .B2(keyinput_57), .C1(P2_REG3_REG_13__SCAN_IN), 
        .C2(keyinput_56), .A(n7081), .ZN(n7168) );
  INV_X1 U8208 ( .A(keyinput_55), .ZN(n7166) );
  INV_X1 U8209 ( .A(keyinput_54), .ZN(n7164) );
  OAI22_X1 U8210 ( .A1(n8700), .A2(keyinput_47), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(keyinput_48), .ZN(n7082) );
  AOI221_X1 U8211 ( .B1(n8700), .B2(keyinput_47), .C1(keyinput_48), .C2(
        P2_REG3_REG_16__SCAN_IN), .A(n7082), .ZN(n7158) );
  INV_X1 U8212 ( .A(keyinput_46), .ZN(n7154) );
  OAI22_X1 U8213 ( .A1(n8655), .A2(keyinput_38), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(keyinput_39), .ZN(n7083) );
  AOI221_X1 U8214 ( .B1(n8655), .B2(keyinput_38), .C1(keyinput_39), .C2(
        P2_REG3_REG_10__SCAN_IN), .A(n7083), .ZN(n7144) );
  OAI22_X1 U8215 ( .A1(n8646), .A2(keyinput_36), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(keyinput_35), .ZN(n7084) );
  AOI221_X1 U8216 ( .B1(n8646), .B2(keyinput_36), .C1(keyinput_35), .C2(
        P2_REG3_REG_7__SCAN_IN), .A(n7084), .ZN(n7141) );
  INV_X1 U8217 ( .A(SI_0_), .ZN(n7233) );
  OAI22_X1 U8218 ( .A1(n5297), .A2(keyinput_33), .B1(n7233), .B2(keyinput_32), 
        .ZN(n7085) );
  AOI221_X1 U8219 ( .B1(n5297), .B2(keyinput_33), .C1(keyinput_32), .C2(n7233), 
        .A(n7085), .ZN(n7089) );
  XNOR2_X1 U8220 ( .A(SI_1_), .B(keyinput_31), .ZN(n7088) );
  XNOR2_X1 U8221 ( .A(SI_2_), .B(keyinput_30), .ZN(n7087) );
  OR2_X1 U8222 ( .A1(SI_3_), .A2(keyinput_29), .ZN(n7086) );
  NAND4_X1 U8223 ( .A1(n7089), .A2(n7088), .A3(n7087), .A4(n7086), .ZN(n7090)
         );
  AOI21_X1 U8224 ( .B1(SI_3_), .B2(keyinput_29), .A(n7090), .ZN(n7138) );
  INV_X1 U8225 ( .A(keyinput_19), .ZN(n7124) );
  INV_X1 U8226 ( .A(SI_24_), .ZN(n7183) );
  AOI22_X1 U8227 ( .A1(n7183), .A2(keyinput_8), .B1(n7092), .B2(keyinput_7), 
        .ZN(n7091) );
  OAI221_X1 U8228 ( .B1(n7183), .B2(keyinput_8), .C1(n7092), .C2(keyinput_7), 
        .A(n7091), .ZN(n7103) );
  INV_X1 U8229 ( .A(keyinput_6), .ZN(n7101) );
  INV_X1 U8230 ( .A(keyinput_5), .ZN(n7099) );
  AOI22_X1 U8231 ( .A1(keyinput_0), .A2(P2_WR_REG_SCAN_IN), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n7093) );
  OAI221_X1 U8232 ( .B1(keyinput_0), .B2(P2_WR_REG_SCAN_IN), .C1(SI_31_), .C2(
        keyinput_1), .A(n7093), .ZN(n7096) );
  INV_X1 U8233 ( .A(SI_30_), .ZN(n7186) );
  AOI22_X1 U8234 ( .A1(n7187), .A2(keyinput_3), .B1(n7186), .B2(keyinput_2), 
        .ZN(n7094) );
  OAI221_X1 U8235 ( .B1(n7187), .B2(keyinput_3), .C1(n7186), .C2(keyinput_2), 
        .A(n7094), .ZN(n7095) );
  OAI22_X1 U8236 ( .A1(keyinput_4), .A2(n7191), .B1(n7096), .B2(n7095), .ZN(
        n7097) );
  AOI21_X1 U8237 ( .B1(keyinput_4), .B2(n7191), .A(n7097), .ZN(n7098) );
  AOI221_X1 U8238 ( .B1(SI_27_), .B2(keyinput_5), .C1(n7194), .C2(n7099), .A(
        n7098), .ZN(n7100) );
  AOI221_X1 U8239 ( .B1(SI_26_), .B2(n7101), .C1(n7197), .C2(keyinput_6), .A(
        n7100), .ZN(n7102) );
  OAI22_X1 U8240 ( .A1(keyinput_9), .A2(n7105), .B1(n7103), .B2(n7102), .ZN(
        n7104) );
  AOI21_X1 U8241 ( .B1(keyinput_9), .B2(n7105), .A(n7104), .ZN(n7122) );
  AOI22_X1 U8242 ( .A1(n7108), .A2(keyinput_16), .B1(n7107), .B2(keyinput_14), 
        .ZN(n7106) );
  OAI221_X1 U8243 ( .B1(n7108), .B2(keyinput_16), .C1(n7107), .C2(keyinput_14), 
        .A(n7106), .ZN(n7121) );
  AOI22_X1 U8244 ( .A1(SI_19_), .A2(keyinput_13), .B1(SI_22_), .B2(keyinput_10), .ZN(n7109) );
  OAI221_X1 U8245 ( .B1(SI_19_), .B2(keyinput_13), .C1(SI_22_), .C2(
        keyinput_10), .A(n7109), .ZN(n7120) );
  OAI22_X1 U8246 ( .A1(n7111), .A2(keyinput_12), .B1(keyinput_17), .B2(SI_15_), 
        .ZN(n7110) );
  AOI221_X1 U8247 ( .B1(n7111), .B2(keyinput_12), .C1(SI_15_), .C2(keyinput_17), .A(n7110), .ZN(n7117) );
  AOI22_X1 U8248 ( .A1(n7114), .A2(keyinput_18), .B1(n7113), .B2(keyinput_15), 
        .ZN(n7112) );
  OAI221_X1 U8249 ( .B1(n7114), .B2(keyinput_18), .C1(n7113), .C2(keyinput_15), 
        .A(n7112), .ZN(n7115) );
  AOI21_X1 U8250 ( .B1(keyinput_11), .B2(n7118), .A(n7115), .ZN(n7116) );
  OAI211_X1 U8251 ( .C1(keyinput_11), .C2(n7118), .A(n7117), .B(n7116), .ZN(
        n7119) );
  NOR4_X1 U8252 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7123)
         );
  AOI221_X1 U8253 ( .B1(SI_13_), .B2(n7124), .C1(n7215), .C2(keyinput_19), .A(
        n7123), .ZN(n7131) );
  AOI22_X1 U8254 ( .A1(SI_8_), .A2(keyinput_24), .B1(SI_10_), .B2(keyinput_22), 
        .ZN(n7125) );
  OAI221_X1 U8255 ( .B1(SI_8_), .B2(keyinput_24), .C1(SI_10_), .C2(keyinput_22), .A(n7125), .ZN(n7130) );
  AOI22_X1 U8256 ( .A1(SI_12_), .A2(keyinput_20), .B1(SI_11_), .B2(keyinput_21), .ZN(n7126) );
  OAI221_X1 U8257 ( .B1(SI_12_), .B2(keyinput_20), .C1(SI_11_), .C2(
        keyinput_21), .A(n7126), .ZN(n7129) );
  AOI22_X1 U8258 ( .A1(n7220), .A2(keyinput_25), .B1(n7221), .B2(keyinput_23), 
        .ZN(n7127) );
  OAI221_X1 U8259 ( .B1(n7220), .B2(keyinput_25), .C1(n7221), .C2(keyinput_23), 
        .A(n7127), .ZN(n7128) );
  NOR4_X1 U8260 ( .A1(n7131), .A2(n7130), .A3(n7129), .A4(n7128), .ZN(n7134)
         );
  XNOR2_X1 U8261 ( .A(n7226), .B(keyinput_27), .ZN(n7133) );
  XNOR2_X1 U8262 ( .A(SI_6_), .B(keyinput_26), .ZN(n7132) );
  OR3_X1 U8263 ( .A1(n7134), .A2(n7133), .A3(n7132), .ZN(n7136) );
  NAND2_X1 U8264 ( .A1(SI_4_), .A2(keyinput_28), .ZN(n7135) );
  OAI211_X1 U8265 ( .C1(SI_4_), .C2(keyinput_28), .A(n7136), .B(n7135), .ZN(
        n7137) );
  AOI22_X1 U8266 ( .A1(keyinput_34), .A2(P2_U3152), .B1(n7138), .B2(n7137), 
        .ZN(n7139) );
  OAI21_X1 U8267 ( .B1(P2_U3152), .B2(keyinput_34), .A(n7139), .ZN(n7140) );
  AOI22_X1 U8268 ( .A1(keyinput_37), .A2(n8102), .B1(n7141), .B2(n7140), .ZN(
        n7142) );
  OAI21_X1 U8269 ( .B1(n8102), .B2(keyinput_37), .A(n7142), .ZN(n7143) );
  OAI211_X1 U8270 ( .C1(n8186), .C2(keyinput_40), .A(n7144), .B(n7143), .ZN(
        n7145) );
  AOI21_X1 U8271 ( .B1(n8186), .B2(keyinput_40), .A(n7145), .ZN(n7152) );
  AOI22_X1 U8272 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_42), .B1(n7147), 
        .B2(keyinput_41), .ZN(n7146) );
  OAI221_X1 U8273 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .C1(n7147), 
        .C2(keyinput_41), .A(n7146), .ZN(n7151) );
  OAI22_X1 U8274 ( .A1(n6393), .A2(keyinput_43), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(keyinput_45), .ZN(n7148) );
  AOI221_X1 U8275 ( .B1(n6393), .B2(keyinput_43), .C1(keyinput_45), .C2(
        P2_REG3_REG_21__SCAN_IN), .A(n7148), .ZN(n7150) );
  XOR2_X1 U8276 ( .A(n7621), .B(keyinput_44), .Z(n7149) );
  OAI211_X1 U8277 ( .C1(n7152), .C2(n7151), .A(n7150), .B(n7149), .ZN(n7153)
         );
  OAI221_X1 U8278 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .C1(n7988), 
        .C2(n7154), .A(n7153), .ZN(n7157) );
  AOI22_X1 U8279 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_50), .ZN(n7155) );
  OAI221_X1 U8280 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_50), .A(n7155), .ZN(n7156) );
  AOI21_X1 U8281 ( .B1(n7158), .B2(n7157), .A(n7156), .ZN(n7161) );
  AOI22_X1 U8282 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(n7514), 
        .B2(keyinput_52), .ZN(n7159) );
  OAI221_X1 U8283 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n7514), 
        .C2(keyinput_52), .A(n7159), .ZN(n7160) );
  AOI211_X1 U8284 ( .C1(n7179), .C2(keyinput_51), .A(n7161), .B(n7160), .ZN(
        n7162) );
  OAI21_X1 U8285 ( .B1(n7179), .B2(keyinput_51), .A(n7162), .ZN(n7163) );
  OAI221_X1 U8286 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n7494), 
        .C2(n7164), .A(n7163), .ZN(n7165) );
  OAI221_X1 U8287 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(n7166), .C1(n7270), .C2(
        keyinput_55), .A(n7165), .ZN(n7167) );
  AOI22_X1 U8288 ( .A1(n7168), .A2(n7167), .B1(keyinput_58), .B2(
        P2_REG3_REG_11__SCAN_IN), .ZN(n7169) );
  OAI21_X1 U8289 ( .B1(keyinput_58), .B2(P2_REG3_REG_11__SCAN_IN), .A(n7169), 
        .ZN(n7174) );
  AOI22_X1 U8290 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_61), .B1(n8775), 
        .B2(keyinput_63), .ZN(n7170) );
  OAI221_X1 U8291 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .C1(n8775), 
        .C2(keyinput_63), .A(n7170), .ZN(n7173) );
  AOI22_X1 U8292 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .ZN(n7171) );
  OAI221_X1 U8293 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_62), .A(n7171), .ZN(n7172) );
  INV_X1 U8294 ( .A(keyinput_123), .ZN(n7275) );
  AOI22_X1 U8295 ( .A1(n6608), .A2(keyinput_121), .B1(keyinput_120), .B2(n7177), .ZN(n7176) );
  OAI221_X1 U8296 ( .B1(n6608), .B2(keyinput_121), .C1(n7177), .C2(
        keyinput_120), .A(n7176), .ZN(n7272) );
  INV_X1 U8297 ( .A(keyinput_119), .ZN(n7269) );
  INV_X1 U8298 ( .A(keyinput_118), .ZN(n7267) );
  OAI22_X1 U8299 ( .A1(n7179), .A2(keyinput_115), .B1(n7514), .B2(keyinput_116), .ZN(n7178) );
  AOI221_X1 U8300 ( .B1(n7179), .B2(keyinput_115), .C1(keyinput_116), .C2(
        n7514), .A(n7178), .ZN(n7264) );
  INV_X1 U8301 ( .A(keyinput_110), .ZN(n7257) );
  OAI22_X1 U8302 ( .A1(n6705), .A2(keyinput_106), .B1(keyinput_105), .B2(
        P2_REG3_REG_19__SCAN_IN), .ZN(n7180) );
  AOI221_X1 U8303 ( .B1(n6705), .B2(keyinput_106), .C1(P2_REG3_REG_19__SCAN_IN), .C2(keyinput_105), .A(n7180), .ZN(n7255) );
  AOI22_X1 U8304 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(n8199), 
        .B2(keyinput_99), .ZN(n7181) );
  OAI221_X1 U8305 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(n8199), .C2(keyinput_99), .A(n7181), .ZN(n7245) );
  INV_X1 U8306 ( .A(keyinput_83), .ZN(n7216) );
  AOI22_X1 U8307 ( .A1(SI_25_), .A2(keyinput_71), .B1(n7183), .B2(keyinput_72), 
        .ZN(n7182) );
  OAI221_X1 U8308 ( .B1(SI_25_), .B2(keyinput_71), .C1(n7183), .C2(keyinput_72), .A(n7182), .ZN(n7199) );
  INV_X1 U8309 ( .A(keyinput_70), .ZN(n7196) );
  INV_X1 U8310 ( .A(keyinput_69), .ZN(n7193) );
  AOI22_X1 U8311 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), .B2(
        keyinput_65), .ZN(n7184) );
  OAI221_X1 U8312 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n7184), .ZN(n7189) );
  AOI22_X1 U8313 ( .A1(n7187), .A2(keyinput_67), .B1(n7186), .B2(keyinput_66), 
        .ZN(n7185) );
  OAI221_X1 U8314 ( .B1(n7187), .B2(keyinput_67), .C1(n7186), .C2(keyinput_66), 
        .A(n7185), .ZN(n7188) );
  OAI22_X1 U8315 ( .A1(keyinput_68), .A2(n7191), .B1(n7189), .B2(n7188), .ZN(
        n7190) );
  AOI21_X1 U8316 ( .B1(keyinput_68), .B2(n7191), .A(n7190), .ZN(n7192) );
  AOI221_X1 U8317 ( .B1(SI_27_), .B2(keyinput_69), .C1(n7194), .C2(n7193), .A(
        n7192), .ZN(n7195) );
  AOI221_X1 U8318 ( .B1(SI_26_), .B2(keyinput_70), .C1(n7197), .C2(n7196), .A(
        n7195), .ZN(n7198) );
  OAI22_X1 U8319 ( .A1(n7199), .A2(n7198), .B1(keyinput_73), .B2(SI_23_), .ZN(
        n7200) );
  AOI21_X1 U8320 ( .B1(keyinput_73), .B2(SI_23_), .A(n7200), .ZN(n7213) );
  AOI22_X1 U8321 ( .A1(SI_18_), .A2(keyinput_78), .B1(n7202), .B2(keyinput_81), 
        .ZN(n7201) );
  OAI221_X1 U8322 ( .B1(SI_18_), .B2(keyinput_78), .C1(n7202), .C2(keyinput_81), .A(n7201), .ZN(n7212) );
  AOI22_X1 U8323 ( .A1(SI_20_), .A2(keyinput_76), .B1(SI_21_), .B2(keyinput_75), .ZN(n7203) );
  OAI221_X1 U8324 ( .B1(SI_20_), .B2(keyinput_76), .C1(SI_21_), .C2(
        keyinput_75), .A(n7203), .ZN(n7211) );
  AOI22_X1 U8325 ( .A1(SI_17_), .A2(keyinput_79), .B1(n7205), .B2(keyinput_77), 
        .ZN(n7204) );
  OAI221_X1 U8326 ( .B1(SI_17_), .B2(keyinput_79), .C1(n7205), .C2(keyinput_77), .A(n7204), .ZN(n7208) );
  AOI22_X1 U8327 ( .A1(SI_14_), .A2(keyinput_82), .B1(SI_16_), .B2(keyinput_80), .ZN(n7206) );
  OAI221_X1 U8328 ( .B1(SI_14_), .B2(keyinput_82), .C1(SI_16_), .C2(
        keyinput_80), .A(n7206), .ZN(n7207) );
  AOI211_X1 U8329 ( .C1(keyinput_74), .C2(SI_22_), .A(n7208), .B(n7207), .ZN(
        n7209) );
  OAI21_X1 U8330 ( .B1(keyinput_74), .B2(SI_22_), .A(n7209), .ZN(n7210) );
  NOR4_X1 U8331 ( .A1(n7213), .A2(n7212), .A3(n7211), .A4(n7210), .ZN(n7214)
         );
  AOI221_X1 U8332 ( .B1(SI_13_), .B2(n7216), .C1(n7215), .C2(keyinput_83), .A(
        n7214), .ZN(n7225) );
  AOI22_X1 U8333 ( .A1(SI_12_), .A2(keyinput_84), .B1(SI_10_), .B2(keyinput_86), .ZN(n7217) );
  OAI221_X1 U8334 ( .B1(SI_12_), .B2(keyinput_84), .C1(SI_10_), .C2(
        keyinput_86), .A(n7217), .ZN(n7224) );
  AOI22_X1 U8335 ( .A1(SI_8_), .A2(keyinput_88), .B1(SI_11_), .B2(keyinput_85), 
        .ZN(n7218) );
  OAI221_X1 U8336 ( .B1(SI_8_), .B2(keyinput_88), .C1(SI_11_), .C2(keyinput_85), .A(n7218), .ZN(n7223) );
  AOI22_X1 U8337 ( .A1(n7221), .A2(keyinput_87), .B1(keyinput_89), .B2(n7220), 
        .ZN(n7219) );
  OAI221_X1 U8338 ( .B1(n7221), .B2(keyinput_87), .C1(n7220), .C2(keyinput_89), 
        .A(n7219), .ZN(n7222) );
  NOR4_X1 U8339 ( .A1(n7225), .A2(n7224), .A3(n7223), .A4(n7222), .ZN(n7230)
         );
  XNOR2_X1 U8340 ( .A(n7226), .B(keyinput_91), .ZN(n7229) );
  XNOR2_X1 U8341 ( .A(n7227), .B(keyinput_90), .ZN(n7228) );
  NOR3_X1 U8342 ( .A1(n7230), .A2(n7229), .A3(n7228), .ZN(n7241) );
  XNOR2_X1 U8343 ( .A(n7231), .B(keyinput_92), .ZN(n7240) );
  AOI22_X1 U8344 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_97), .B1(n7233), .B2(
        keyinput_96), .ZN(n7232) );
  OAI221_X1 U8345 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_97), .C1(n7233), .C2(
        keyinput_96), .A(n7232), .ZN(n7238) );
  XNOR2_X1 U8346 ( .A(n7234), .B(keyinput_93), .ZN(n7237) );
  XNOR2_X1 U8347 ( .A(SI_1_), .B(keyinput_95), .ZN(n7236) );
  XNOR2_X1 U8348 ( .A(SI_2_), .B(keyinput_94), .ZN(n7235) );
  NOR4_X1 U8349 ( .A1(n7238), .A2(n7237), .A3(n7236), .A4(n7235), .ZN(n7239)
         );
  OAI21_X1 U8350 ( .B1(n7241), .B2(n7240), .A(n7239), .ZN(n7242) );
  OAI21_X1 U8351 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_98), .A(n7242), 
        .ZN(n7243) );
  AOI21_X1 U8352 ( .B1(keyinput_98), .B2(P2_STATE_REG_SCAN_IN), .A(n7243), 
        .ZN(n7244) );
  OAI22_X1 U8353 ( .A1(keyinput_101), .A2(n8102), .B1(n7245), .B2(n7244), .ZN(
        n7246) );
  AOI21_X1 U8354 ( .B1(keyinput_101), .B2(n8102), .A(n7246), .ZN(n7249) );
  AOI22_X1 U8355 ( .A1(n8655), .A2(keyinput_102), .B1(keyinput_104), .B2(n8186), .ZN(n7247) );
  OAI221_X1 U8356 ( .B1(n8655), .B2(keyinput_102), .C1(n8186), .C2(
        keyinput_104), .A(n7247), .ZN(n7248) );
  AOI211_X1 U8357 ( .C1(n6432), .C2(keyinput_103), .A(n7249), .B(n7248), .ZN(
        n7250) );
  OAI21_X1 U8358 ( .B1(n6432), .B2(keyinput_103), .A(n7250), .ZN(n7254) );
  XNOR2_X1 U8359 ( .A(n7621), .B(keyinput_108), .ZN(n7253) );
  AOI22_X1 U8360 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(n6393), 
        .B2(keyinput_107), .ZN(n7251) );
  OAI221_X1 U8361 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(n6393), .C2(keyinput_107), .A(n7251), .ZN(n7252) );
  AOI211_X1 U8362 ( .C1(n7255), .C2(n7254), .A(n7253), .B(n7252), .ZN(n7256)
         );
  AOI221_X1 U8363 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n7257), .C1(n7988), .C2(
        keyinput_110), .A(n7256), .ZN(n7262) );
  AOI22_X1 U8364 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_112), .B1(n8700), 
        .B2(keyinput_111), .ZN(n7258) );
  OAI221_X1 U8365 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_112), .C1(n8700), .C2(keyinput_111), .A(n7258), .ZN(n7261) );
  OAI22_X1 U8366 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_114), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .ZN(n7259) );
  AOI221_X1 U8367 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .C1(
        keyinput_113), .C2(P2_REG3_REG_5__SCAN_IN), .A(n7259), .ZN(n7260) );
  OAI21_X1 U8368 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n7263) );
  OAI211_X1 U8369 ( .C1(P2_REG3_REG_9__SCAN_IN), .C2(keyinput_117), .A(n7264), 
        .B(n7263), .ZN(n7265) );
  AOI21_X1 U8370 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .A(n7265), 
        .ZN(n7266) );
  AOI221_X1 U8371 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(n7494), 
        .C2(n7267), .A(n7266), .ZN(n7268) );
  AOI221_X1 U8372 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(n7270), .C2(n7269), .A(n7268), .ZN(n7271) );
  OAI22_X1 U8373 ( .A1(keyinput_122), .A2(n8792), .B1(n7272), .B2(n7271), .ZN(
        n7273) );
  AOI22_X1 U8374 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_125), .B1(n6673), 
        .B2(keyinput_126), .ZN(n7276) );
  OAI221_X1 U8375 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .C1(n6673), 
        .C2(keyinput_126), .A(n7276), .ZN(n7279) );
  AOI22_X1 U8376 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(n8775), 
        .B2(keyinput_127), .ZN(n7277) );
  OAI221_X1 U8377 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(n8775), .C2(keyinput_127), .A(n7277), .ZN(n7278) );
  AND2_X1 U8378 ( .A1(n7285), .A2(P1_U3084), .ZN(n10199) );
  INV_X2 U8379 ( .A(n10199), .ZN(n10197) );
  OAI222_X1 U8380 ( .A1(n10204), .A2(n8314), .B1(n10197), .B2(n7302), .C1(
        P1_U3084), .C2(n7466), .ZN(P1_U3351) );
  INV_X1 U8381 ( .A(n8164), .ZN(n8192) );
  NOR2_X1 U8382 ( .A1(n7285), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9265) );
  INV_X1 U8383 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7389) );
  OAI222_X1 U8384 ( .A1(P2_U3152), .A2(n8192), .B1(n8529), .B2(n7287), .C1(
        n9280), .C2(n7389), .ZN(P2_U3355) );
  OAI222_X1 U8385 ( .A1(P1_U3084), .A2(n7368), .B1(n10197), .B2(n7298), .C1(
        n5493), .C2(n10204), .ZN(P1_U3352) );
  OAI222_X1 U8386 ( .A1(P1_U3084), .A2(n7286), .B1(n10197), .B2(n7305), .C1(
        n8325), .C2(n10204), .ZN(P1_U3348) );
  OAI222_X1 U8387 ( .A1(n10204), .A2(n8321), .B1(n10197), .B2(n7293), .C1(
        P1_U3084), .C2(n7329), .ZN(P1_U3349) );
  OAI222_X1 U8388 ( .A1(n10204), .A2(n7288), .B1(n10197), .B2(n7287), .C1(
        n7413), .C2(P1_U3084), .ZN(P1_U3350) );
  INV_X1 U8389 ( .A(n10204), .ZN(n10195) );
  AOI22_X1 U8390 ( .A1(n10195), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7345), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7289) );
  OAI21_X1 U8391 ( .B1(n7290), .B2(n10197), .A(n7289), .ZN(P1_U3347) );
  INV_X1 U8392 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7291) );
  INV_X1 U8393 ( .A(n8201), .ZN(n8180) );
  OAI222_X1 U8394 ( .A1(n9280), .A2(n7291), .B1(n8529), .B2(n7290), .C1(n8180), 
        .C2(P2_U3152), .ZN(P2_U3352) );
  AOI22_X1 U8395 ( .A1(n7399), .A2(P1_STATE_REG_SCAN_IN), .B1(n10195), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n7292) );
  OAI21_X1 U8396 ( .B1(n7300), .B2(n10197), .A(n7292), .ZN(P1_U3346) );
  INV_X1 U8397 ( .A(n8162), .ZN(n8276) );
  OAI222_X1 U8398 ( .A1(n9280), .A2(n4965), .B1(n8529), .B2(n7293), .C1(n8276), 
        .C2(P2_U3152), .ZN(P2_U3354) );
  NAND2_X1 U8399 ( .A1(n10210), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7295) );
  OAI21_X1 U8400 ( .B1(n10210), .B2(n7296), .A(n7295), .ZN(P1_U3440) );
  OAI222_X1 U8401 ( .A1(P2_U3152), .A2(n8167), .B1(n8529), .B2(n7298), .C1(
        n7297), .C2(n9280), .ZN(P2_U3357) );
  INV_X1 U8402 ( .A(n8213), .ZN(n8220) );
  INV_X1 U8403 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7299) );
  OAI222_X1 U8404 ( .A1(P2_U3152), .A2(n8220), .B1(n8529), .B2(n7300), .C1(
        n7299), .C2(n9280), .ZN(P2_U3351) );
  OAI222_X1 U8405 ( .A1(P2_U3152), .A2(n7303), .B1(n8529), .B2(n7302), .C1(
        n7301), .C2(n9280), .ZN(P2_U3356) );
  INV_X1 U8406 ( .A(n8160), .ZN(n8237) );
  INV_X1 U8407 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7304) );
  OAI222_X1 U8408 ( .A1(P2_U3152), .A2(n8237), .B1(n8529), .B2(n7305), .C1(
        n7304), .C2(n9280), .ZN(P2_U3353) );
  INV_X1 U8409 ( .A(n7400), .ZN(n9694) );
  INV_X1 U8410 ( .A(n7306), .ZN(n7307) );
  INV_X1 U8411 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8367) );
  OAI222_X1 U8412 ( .A1(n9694), .A2(P1_U3084), .B1(n10197), .B2(n7307), .C1(
        n10204), .C2(n8367), .ZN(P1_U3345) );
  INV_X1 U8413 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7308) );
  INV_X1 U8414 ( .A(n8217), .ZN(n8264) );
  OAI222_X1 U8415 ( .A1(n9280), .A2(n7308), .B1(n8529), .B2(n7307), .C1(
        P2_U3152), .C2(n8264), .ZN(P2_U3350) );
  INV_X1 U8416 ( .A(n7309), .ZN(n7312) );
  AOI22_X1 U8417 ( .A1(n7545), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10195), .ZN(n7310) );
  OAI21_X1 U8418 ( .B1(n7312), .B2(n10197), .A(n7310), .ZN(P1_U3344) );
  INV_X1 U8419 ( .A(n8242), .ZN(n8247) );
  INV_X1 U8420 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7311) );
  OAI222_X1 U8421 ( .A1(P2_U3152), .A2(n8247), .B1(n8529), .B2(n7312), .C1(
        n7311), .C2(n9280), .ZN(P2_U3349) );
  XNOR2_X1 U8422 ( .A(n7345), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7318) );
  INV_X1 U8423 ( .A(n7329), .ZN(n9687) );
  INV_X1 U8424 ( .A(n7413), .ZN(n7326) );
  INV_X1 U8425 ( .A(n7466), .ZN(n7324) );
  INV_X1 U8426 ( .A(n7368), .ZN(n7322) );
  NAND2_X1 U8427 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7457) );
  AOI21_X1 U8428 ( .B1(n7322), .B2(P1_REG2_REG_1__SCAN_IN), .A(n7363), .ZN(
        n7469) );
  XOR2_X1 U8429 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7466), .Z(n7468) );
  INV_X1 U8430 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7768) );
  XNOR2_X1 U8431 ( .A(n7413), .B(n7768), .ZN(n7415) );
  XNOR2_X1 U8432 ( .A(n7329), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U8433 ( .A1(n4918), .A2(n9689), .ZN(n9688) );
  OAI21_X1 U8434 ( .B1(n9687), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9688), .ZN(
        n7376) );
  NOR2_X1 U8435 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7374), .ZN(n7314) );
  AOI21_X1 U8436 ( .B1(n7374), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7314), .ZN(
        n7377) );
  NAND2_X1 U8437 ( .A1(n7376), .A2(n7377), .ZN(n7375) );
  OAI21_X1 U8438 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7374), .A(n7375), .ZN(
        n7317) );
  CLKBUF_X1 U8439 ( .A(n7315), .Z(n10295) );
  OR2_X1 U8440 ( .A1(n10295), .A2(P1_U3084), .ZN(n10201) );
  INV_X1 U8441 ( .A(n10201), .ZN(n7316) );
  AND2_X1 U8442 ( .A1(n10288), .A2(n7316), .ZN(n10319) );
  NOR2_X1 U8443 ( .A1(n7317), .A2(n7318), .ZN(n7340) );
  AOI211_X1 U8444 ( .C1(n7318), .C2(n7317), .A(n10305), .B(n7340), .ZN(n7319)
         );
  AOI21_X1 U8445 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n10324), .A(n7319), .ZN(
        n7339) );
  INV_X1 U8446 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7320) );
  NOR2_X1 U8447 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7320), .ZN(n7643) );
  NOR2_X1 U8448 ( .A1(n6181), .A2(P1_U3084), .ZN(n10194) );
  AND3_X1 U8449 ( .A1(n10288), .A2(n10194), .A3(n10295), .ZN(n10315) );
  XNOR2_X1 U8450 ( .A(n7466), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7463) );
  XNOR2_X1 U8451 ( .A(n7368), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n7357) );
  AND2_X1 U8452 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7321) );
  NAND2_X1 U8453 ( .A1(n7357), .A2(n7321), .ZN(n7358) );
  NAND2_X1 U8454 ( .A1(n7322), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7323) );
  NAND2_X1 U8455 ( .A1(n7358), .A2(n7323), .ZN(n7462) );
  NAND2_X1 U8456 ( .A1(n7463), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U8457 ( .A1(n7324), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U8458 ( .A1(n7461), .A2(n7325), .ZN(n7409) );
  XNOR2_X1 U8459 ( .A(n7413), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U8460 ( .A1(n7409), .A2(n7410), .ZN(n7408) );
  NAND2_X1 U8461 ( .A1(n7326), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U8462 ( .A1(n7408), .A2(n7327), .ZN(n9682) );
  INV_X1 U8463 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7328) );
  XNOR2_X1 U8464 ( .A(n7329), .B(n7328), .ZN(n9683) );
  NOR2_X1 U8465 ( .A1(n9682), .A2(n9683), .ZN(n9681) );
  AND2_X1 U8466 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  OR2_X1 U8467 ( .A1(n9681), .A2(n7330), .ZN(n7372) );
  OR2_X1 U8468 ( .A1(n7374), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8469 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7374), .ZN(n7332) );
  NAND2_X1 U8470 ( .A1(n7331), .A2(n7332), .ZN(n7371) );
  OR2_X1 U8471 ( .A1(n7372), .A2(n7371), .ZN(n7369) );
  NAND2_X1 U8472 ( .A1(n7369), .A2(n7332), .ZN(n7335) );
  INV_X1 U8473 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7333) );
  XNOR2_X1 U8474 ( .A(n7345), .B(n7333), .ZN(n7334) );
  AND2_X1 U8475 ( .A1(n7335), .A2(n7334), .ZN(n7344) );
  NOR2_X1 U8476 ( .A1(n7335), .A2(n7334), .ZN(n7336) );
  NOR3_X1 U8477 ( .A1(n10332), .A2(n7344), .A3(n7336), .ZN(n7337) );
  AOI211_X1 U8478 ( .C1(n10311), .C2(n7345), .A(n7643), .B(n7337), .ZN(n7338)
         );
  NAND2_X1 U8479 ( .A1(n7339), .A2(n7338), .ZN(P1_U3247) );
  INV_X1 U8480 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7353) );
  NOR2_X1 U8481 ( .A1(n7399), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7341) );
  AOI21_X1 U8482 ( .B1(n7399), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7341), .ZN(
        n7342) );
  OAI21_X1 U8483 ( .B1(n7343), .B2(n7342), .A(n7398), .ZN(n7350) );
  INV_X1 U8484 ( .A(n10305), .ZN(n10336) );
  AOI21_X1 U8485 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n7345), .A(n7344), .ZN(
        n7348) );
  NOR2_X1 U8486 ( .A1(n7399), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7346) );
  AOI21_X1 U8487 ( .B1(n7399), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7346), .ZN(
        n7347) );
  NAND2_X1 U8488 ( .A1(n7348), .A2(n7347), .ZN(n7391) );
  OAI21_X1 U8489 ( .B1(n7348), .B2(n7347), .A(n7391), .ZN(n7349) );
  AOI22_X1 U8490 ( .A1(n7350), .A2(n10336), .B1(n10315), .B2(n7349), .ZN(n7352) );
  AND2_X1 U8491 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7903) );
  AOI21_X1 U8492 ( .B1(n10311), .B2(n7399), .A(n7903), .ZN(n7351) );
  OAI211_X1 U8493 ( .C1(n9776), .C2(n7353), .A(n7352), .B(n7351), .ZN(P1_U3248) );
  INV_X1 U8494 ( .A(n10312), .ZN(n7538) );
  INV_X1 U8495 ( .A(n7354), .ZN(n7356) );
  INV_X1 U8496 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8324) );
  OAI222_X1 U8497 ( .A1(P1_U3084), .A2(n7538), .B1(n10197), .B2(n7356), .C1(
        n8324), .C2(n10204), .ZN(P1_U3343) );
  INV_X1 U8498 ( .A(n8789), .ZN(n8795) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7355) );
  OAI222_X1 U8500 ( .A1(P2_U3152), .A2(n8795), .B1(n8529), .B2(n7356), .C1(
        n7355), .C2(n9280), .ZN(P2_U3348) );
  INV_X1 U8501 ( .A(n10311), .ZN(n10316) );
  NAND2_X1 U8502 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7361) );
  INV_X1 U8503 ( .A(n7357), .ZN(n7360) );
  INV_X1 U8504 ( .A(n7358), .ZN(n7359) );
  AOI211_X1 U8505 ( .C1(n7361), .C2(n7360), .A(n7359), .B(n10332), .ZN(n7362)
         );
  AOI21_X1 U8506 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n7362), .ZN(
        n7367) );
  AOI211_X1 U8507 ( .C1(n7457), .C2(n7364), .A(n7363), .B(n10305), .ZN(n7365)
         );
  AOI21_X1 U8508 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n10324), .A(n7365), .ZN(
        n7366) );
  OAI211_X1 U8509 ( .C1(n7368), .C2(n10316), .A(n7367), .B(n7366), .ZN(
        P1_U3242) );
  INV_X1 U8510 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7381) );
  AND2_X1 U8511 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7608) );
  INV_X1 U8512 ( .A(n7369), .ZN(n7370) );
  AOI211_X1 U8513 ( .C1(n7372), .C2(n7371), .A(n7370), .B(n10332), .ZN(n7373)
         );
  AOI211_X1 U8514 ( .C1(n10311), .C2(n7374), .A(n7608), .B(n7373), .ZN(n7380)
         );
  OAI21_X1 U8515 ( .B1(n7377), .B2(n7376), .A(n7375), .ZN(n7378) );
  NAND2_X1 U8516 ( .A1(n7378), .A2(n10336), .ZN(n7379) );
  OAI211_X1 U8517 ( .C1(n7381), .C2(n9776), .A(n7380), .B(n7379), .ZN(P1_U3246) );
  INV_X1 U8518 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7382) );
  INV_X1 U8519 ( .A(n8813), .ZN(n8805) );
  OAI222_X1 U8520 ( .A1(n9280), .A2(n7382), .B1(n8529), .B2(n7383), .C1(n8805), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8521 ( .A(n10325), .ZN(n10340) );
  INV_X1 U8522 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8323) );
  OAI222_X1 U8523 ( .A1(P1_U3084), .A2(n10340), .B1(n10197), .B2(n7383), .C1(
        n8323), .C2(n10204), .ZN(P1_U3342) );
  INV_X1 U8524 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7473) );
  NAND2_X1 U8525 ( .A1(n8357), .A2(P1_U4006), .ZN(n7384) );
  OAI21_X1 U8526 ( .B1(n7473), .B2(P1_U4006), .A(n7384), .ZN(P1_U3567) );
  INV_X1 U8527 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7842) );
  INV_X1 U8528 ( .A(n9999), .ZN(n9957) );
  NAND2_X1 U8529 ( .A1(n9957), .A2(P1_U4006), .ZN(n7385) );
  OAI21_X1 U8530 ( .B1(n7842), .B2(P1_U4006), .A(n7385), .ZN(P1_U3572) );
  NAND2_X1 U8531 ( .A1(n9944), .A2(P1_U4006), .ZN(n7386) );
  OAI21_X1 U8532 ( .B1(n6573), .B2(P1_U4006), .A(n7386), .ZN(P1_U3575) );
  INV_X1 U8533 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7525) );
  INV_X1 U8534 ( .A(n10017), .ZN(n8593) );
  NAND2_X1 U8535 ( .A1(n8593), .A2(P1_U4006), .ZN(n7387) );
  OAI21_X1 U8536 ( .B1(n7525), .B2(P1_U4006), .A(n7387), .ZN(P1_U3569) );
  NAND2_X1 U8537 ( .A1(n7760), .A2(P1_U4006), .ZN(n7388) );
  OAI21_X1 U8538 ( .B1(P1_U4006), .B2(n7389), .A(n7388), .ZN(P1_U3558) );
  NOR2_X1 U8539 ( .A1(n7545), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7390) );
  AOI21_X1 U8540 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7545), .A(n7390), .ZN(
        n7393) );
  INV_X1 U8541 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U8542 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7400), .B1(n9694), .B2(
        n10570), .ZN(n9699) );
  OAI21_X1 U8543 ( .B1(n7399), .B2(P1_REG1_REG_7__SCAN_IN), .A(n7391), .ZN(
        n9698) );
  NAND2_X1 U8544 ( .A1(n9699), .A2(n9698), .ZN(n9697) );
  OAI21_X1 U8545 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7400), .A(n9697), .ZN(
        n7392) );
  NAND2_X1 U8546 ( .A1(n7393), .A2(n7392), .ZN(n7539) );
  OAI21_X1 U8547 ( .B1(n7393), .B2(n7392), .A(n7539), .ZN(n7406) );
  INV_X1 U8548 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7396) );
  NOR2_X1 U8549 ( .A1(n7394), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7940) );
  AOI21_X1 U8550 ( .B1(n10311), .B2(n7545), .A(n7940), .ZN(n7395) );
  OAI21_X1 U8551 ( .B1(n9776), .B2(n7396), .A(n7395), .ZN(n7405) );
  INV_X1 U8552 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7397) );
  AOI22_X1 U8553 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7400), .B1(n9694), .B2(
        n7397), .ZN(n9703) );
  OAI21_X1 U8554 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7400), .A(n9701), .ZN(
        n7403) );
  NAND2_X1 U8555 ( .A1(n7545), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7401) );
  OAI21_X1 U8556 ( .B1(n7545), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7401), .ZN(
        n7402) );
  AOI211_X1 U8557 ( .C1(n7403), .C2(n7402), .A(n7544), .B(n10305), .ZN(n7404)
         );
  AOI211_X1 U8558 ( .C1(n7406), .C2(n10315), .A(n7405), .B(n7404), .ZN(n7407)
         );
  INV_X1 U8559 ( .A(n7407), .ZN(P1_U3250) );
  AND2_X1 U8560 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7487) );
  INV_X1 U8561 ( .A(n7487), .ZN(n7412) );
  OAI211_X1 U8562 ( .C1(n7410), .C2(n7409), .A(n10315), .B(n7408), .ZN(n7411)
         );
  OAI211_X1 U8563 ( .C1(n10316), .C2(n7413), .A(n7412), .B(n7411), .ZN(n7418)
         );
  AOI211_X1 U8564 ( .C1(n7416), .C2(n7415), .A(n7414), .B(n10305), .ZN(n7417)
         );
  AOI211_X1 U8565 ( .C1(n10324), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n7418), .B(
        n7417), .ZN(n7419) );
  INV_X1 U8566 ( .A(n7419), .ZN(P1_U3244) );
  NOR2_X1 U8567 ( .A1(n7420), .A2(P2_U3152), .ZN(n10384) );
  OAI21_X1 U8568 ( .B1(n7423), .B2(n7421), .A(n7422), .ZN(n7425) );
  INV_X1 U8569 ( .A(n7424), .ZN(n8318) );
  OAI22_X1 U8570 ( .A1(n8318), .A2(n9066), .B1(n6779), .B2(n9068), .ZN(n7619)
         );
  AOI22_X1 U8571 ( .A1(n10375), .A2(n7425), .B1(n8766), .B2(n7619), .ZN(n7427)
         );
  NAND2_X1 U8572 ( .A1(n6759), .A2(n7613), .ZN(n7426) );
  OAI211_X1 U8573 ( .C1(n10384), .C2(n7621), .A(n7427), .B(n7426), .ZN(
        P2_U3224) );
  INV_X1 U8574 ( .A(n7714), .ZN(n7727) );
  NAND2_X1 U8575 ( .A1(n7727), .A2(n7741), .ZN(n7720) );
  INV_X1 U8576 ( .A(n7741), .ZN(n7742) );
  NAND2_X1 U8577 ( .A1(n7714), .A2(n7742), .ZN(n9621) );
  AND2_X1 U8578 ( .A1(n7720), .A2(n9621), .ZN(n9509) );
  INV_X1 U8579 ( .A(n7728), .ZN(n7429) );
  NAND2_X1 U8580 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  INV_X1 U8581 ( .A(n10514), .ZN(n10484) );
  OAI22_X1 U8582 ( .A1(n9509), .A2(n7430), .B1(n7713), .B2(n10484), .ZN(n7699)
         );
  AOI21_X1 U8583 ( .B1(n7741), .B2(n7728), .A(n7699), .ZN(n7440) );
  AND2_X1 U8584 ( .A1(n7700), .A2(n7431), .ZN(n10285) );
  AND3_X1 U8585 ( .A1(n7702), .A2(n7433), .A3(n7432), .ZN(n7434) );
  NAND2_X1 U8586 ( .A1(n10589), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7435) );
  OAI21_X1 U8587 ( .B1(n7440), .B2(n10589), .A(n7435), .ZN(P1_U3523) );
  INV_X1 U8588 ( .A(n7436), .ZN(n7704) );
  INV_X1 U8589 ( .A(n10595), .ZN(n10592) );
  INV_X1 U8590 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7438) );
  OR2_X1 U8591 ( .A1(n10595), .A2(n7438), .ZN(n7439) );
  OAI21_X1 U8592 ( .B1(n7440), .B2(n10592), .A(n7439), .ZN(P1_U3454) );
  INV_X1 U8593 ( .A(n7441), .ZN(n7474) );
  AOI22_X1 U8594 ( .A1(n7781), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10195), .ZN(n7442) );
  OAI21_X1 U8595 ( .B1(n7474), .B2(n10197), .A(n7442), .ZN(P1_U3341) );
  XNOR2_X1 U8596 ( .A(n7444), .B(n7443), .ZN(n7445) );
  XNOR2_X1 U8597 ( .A(n7446), .B(n7445), .ZN(n7453) );
  INV_X1 U8598 ( .A(n9405), .ZN(n8028) );
  AOI22_X1 U8599 ( .A1(n8028), .A2(n7714), .B1(n4879), .B2(n9408), .ZN(n7452)
         );
  INV_X1 U8600 ( .A(n10561), .ZN(n10581) );
  INV_X1 U8601 ( .A(n7447), .ZN(n7701) );
  AOI211_X1 U8602 ( .C1(n7448), .C2(n10581), .A(P1_U3084), .B(n7701), .ZN(
        n7450) );
  NAND2_X1 U8603 ( .A1(n7450), .A2(n7449), .ZN(n7497) );
  AOI22_X1 U8604 ( .A1(n9401), .A2(n9679), .B1(n7497), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7451) );
  OAI211_X1 U8605 ( .C1(n7453), .C2(n9410), .A(n7452), .B(n7451), .ZN(P1_U3220) );
  OAI21_X1 U8606 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7495) );
  MUX2_X1 U8607 ( .A(n7457), .B(n7495), .S(n10295), .Z(n7460) );
  NOR2_X1 U8608 ( .A1(n10295), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7458) );
  OR2_X1 U8609 ( .A1(n6181), .A2(n7458), .ZN(n10290) );
  AND2_X1 U8610 ( .A1(n10290), .A2(n10294), .ZN(n10300) );
  INV_X1 U8611 ( .A(n10300), .ZN(n7459) );
  OAI211_X1 U8612 ( .C1(n7460), .C2(n6181), .A(P1_U4006), .B(n7459), .ZN(n9693) );
  NAND2_X1 U8613 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7465) );
  OAI211_X1 U8614 ( .C1(n7463), .C2(n7462), .A(n10315), .B(n7461), .ZN(n7464)
         );
  OAI211_X1 U8615 ( .C1(n10316), .C2(n7466), .A(n7465), .B(n7464), .ZN(n7471)
         );
  AOI211_X1 U8616 ( .C1(n7469), .C2(n7468), .A(n7467), .B(n10305), .ZN(n7470)
         );
  AOI211_X1 U8617 ( .C1(n10324), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n7471), .B(
        n7470), .ZN(n7472) );
  NAND2_X1 U8618 ( .A1(n9693), .A2(n7472), .ZN(P1_U3243) );
  INV_X1 U8619 ( .A(n8820), .ZN(n8826) );
  OAI222_X1 U8620 ( .A1(P2_U3152), .A2(n8826), .B1(n8529), .B2(n7474), .C1(
        n9280), .C2(n7473), .ZN(P2_U3346) );
  XOR2_X1 U8621 ( .A(n7476), .B(n7475), .Z(n7479) );
  AOI22_X1 U8622 ( .A1(n8028), .A2(n9680), .B1(n5162), .B2(n9408), .ZN(n7478)
         );
  AOI22_X1 U8623 ( .A1(n9401), .A2(n7760), .B1(n7497), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7477) );
  OAI211_X1 U8624 ( .C1(n7479), .C2(n9410), .A(n7478), .B(n7477), .ZN(P1_U3235) );
  INV_X1 U8625 ( .A(n7801), .ZN(n7807) );
  INV_X1 U8626 ( .A(n7480), .ZN(n7481) );
  INV_X1 U8627 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8339) );
  OAI222_X1 U8628 ( .A1(P1_U3084), .A2(n7807), .B1(n10197), .B2(n7481), .C1(
        n8339), .C2(n10204), .ZN(P1_U3340) );
  INV_X1 U8629 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7482) );
  INV_X1 U8630 ( .A(n8839), .ZN(n8834) );
  OAI222_X1 U8631 ( .A1(n9280), .A2(n7482), .B1(n8529), .B2(n7481), .C1(n8834), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XNOR2_X1 U8632 ( .A(n7483), .B(n7484), .ZN(n7485) );
  NAND2_X1 U8633 ( .A1(n7485), .A2(n9381), .ZN(n7489) );
  INV_X1 U8634 ( .A(n9678), .ZN(n10481) );
  INV_X1 U8635 ( .A(n9679), .ZN(n7761) );
  OAI22_X1 U8636 ( .A1(n10481), .A2(n9342), .B1(n9405), .B2(n7761), .ZN(n7486)
         );
  AOI211_X1 U8637 ( .C1(n7773), .C2(n9408), .A(n7487), .B(n7486), .ZN(n7488)
         );
  OAI211_X1 U8638 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9395), .A(n7489), .B(
        n7488), .ZN(P1_U3216) );
  NAND2_X1 U8639 ( .A1(n10375), .A2(n6302), .ZN(n8761) );
  OAI22_X1 U8640 ( .A1(n8318), .A2(n8761), .B1(n8759), .B2(n7622), .ZN(n7491)
         );
  NAND2_X1 U8641 ( .A1(n7491), .A2(n7490), .ZN(n7493) );
  AOI22_X1 U8642 ( .A1(n10373), .A2(n4868), .B1(n7600), .B2(n6759), .ZN(n7492)
         );
  OAI211_X1 U8643 ( .C1(n7494), .C2(n10384), .A(n7493), .B(n7492), .ZN(
        P2_U3234) );
  INV_X1 U8644 ( .A(n7495), .ZN(n7499) );
  OAI22_X1 U8645 ( .A1(n7713), .A2(n9342), .B1(n9388), .B2(n7742), .ZN(n7496)
         );
  AOI21_X1 U8646 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7497), .A(n7496), .ZN(
        n7498) );
  OAI21_X1 U8647 ( .B1(n7499), .B2(n9410), .A(n7498), .ZN(P1_U3230) );
  NAND2_X1 U8648 ( .A1(n7614), .A2(n7500), .ZN(n7594) );
  AOI22_X1 U8649 ( .A1(n7594), .A2(n10453), .B1(n10448), .B2(n4868), .ZN(n7597) );
  AOI22_X1 U8650 ( .A1(n10617), .A2(n7594), .B1(n6751), .B2(n7600), .ZN(n7501)
         );
  NAND2_X1 U8651 ( .A1(n7597), .A2(n7501), .ZN(n7650) );
  NAND2_X1 U8652 ( .A1(n10624), .A2(n7650), .ZN(n7502) );
  OAI21_X1 U8653 ( .B1(n10624), .B2(n6265), .A(n7502), .ZN(P2_U3451) );
  INV_X1 U8654 ( .A(n7503), .ZN(n10435) );
  XNOR2_X1 U8655 ( .A(n7505), .B(n7504), .ZN(n7506) );
  NAND2_X1 U8656 ( .A1(n7506), .A2(n9381), .ZN(n7509) );
  AND2_X1 U8657 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9686) );
  OAI22_X1 U8658 ( .A1(n10418), .A2(n9405), .B1(n9342), .B2(n10417), .ZN(n7507) );
  AOI211_X1 U8659 ( .C1(n7857), .C2(n9408), .A(n9686), .B(n7507), .ZN(n7508)
         );
  OAI211_X1 U8660 ( .C1(n9395), .C2(n10435), .A(n7509), .B(n7508), .ZN(
        P1_U3228) );
  INV_X1 U8661 ( .A(n7510), .ZN(n7513) );
  NOR3_X1 U8662 ( .A1(n8761), .A2(n7511), .A3(n6780), .ZN(n7512) );
  AOI21_X1 U8663 ( .B1(n10375), .B2(n7513), .A(n7512), .ZN(n7522) );
  NOR2_X1 U8664 ( .A1(n7514), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8270) );
  INV_X1 U8665 ( .A(n8270), .ZN(n7517) );
  NAND2_X1 U8666 ( .A1(n6759), .A2(n7515), .ZN(n7516) );
  OAI211_X1 U8667 ( .C1(n8780), .C2(n10469), .A(n7517), .B(n7516), .ZN(n7519)
         );
  OAI22_X1 U8668 ( .A1(n8561), .A2(n8778), .B1(n8782), .B2(n6780), .ZN(n7518)
         );
  AOI211_X1 U8669 ( .C1(n4953), .C2(n10375), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI21_X1 U8670 ( .B1(n7522), .B2(n7521), .A(n7520), .ZN(P2_U3232) );
  INV_X1 U8671 ( .A(n8003), .ZN(n8008) );
  INV_X1 U8672 ( .A(n7523), .ZN(n7524) );
  INV_X1 U8673 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8341) );
  OAI222_X1 U8674 ( .A1(P1_U3084), .A2(n8008), .B1(n10197), .B2(n7524), .C1(
        n8341), .C2(n10204), .ZN(P1_U3339) );
  INV_X1 U8675 ( .A(n8851), .ZN(n8855) );
  OAI222_X1 U8676 ( .A1(P2_U3152), .A2(n8855), .B1(n9280), .B2(n7525), .C1(
        n7524), .C2(n8529), .ZN(P2_U3344) );
  INV_X1 U8677 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7536) );
  XNOR2_X1 U8678 ( .A(n7526), .B(n7527), .ZN(n7659) );
  XNOR2_X1 U8679 ( .A(n7528), .B(n7529), .ZN(n7532) );
  OR2_X1 U8680 ( .A1(n8328), .A2(n9068), .ZN(n7531) );
  NAND2_X1 U8681 ( .A1(n8663), .A2(n10450), .ZN(n7530) );
  NAND2_X1 U8682 ( .A1(n7531), .A2(n7530), .ZN(n8571) );
  AOI21_X1 U8683 ( .B1(n7532), .B2(n10453), .A(n8571), .ZN(n7667) );
  INV_X1 U8684 ( .A(n7635), .ZN(n7533) );
  AOI211_X1 U8685 ( .C1(n8570), .C2(n10445), .A(n10613), .B(n7533), .ZN(n7665)
         );
  AOI21_X1 U8686 ( .B1(n10403), .B2(n8570), .A(n7665), .ZN(n7534) );
  OAI211_X1 U8687 ( .C1(n9245), .C2(n7659), .A(n7667), .B(n7534), .ZN(n9249)
         );
  NAND2_X1 U8688 ( .A1(n9249), .A2(n10624), .ZN(n7535) );
  OAI21_X1 U8689 ( .B1(n10624), .B2(n7536), .A(n7535), .ZN(P2_U3466) );
  INV_X1 U8690 ( .A(n9817), .ZN(n8618) );
  NAND2_X1 U8691 ( .A1(n8618), .A2(P1_U4006), .ZN(n7537) );
  OAI21_X1 U8692 ( .B1(P1_U4006), .B2(n9276), .A(n7537), .ZN(P1_U3583) );
  INV_X1 U8693 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8117) );
  AOI22_X1 U8694 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n10312), .B1(n7538), .B2(
        n8117), .ZN(n10303) );
  OAI21_X1 U8695 ( .B1(n7545), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7539), .ZN(
        n10302) );
  NAND2_X1 U8696 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OR2_X1 U8697 ( .A1(n10312), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U8698 ( .A1(n10301), .A2(n7540), .ZN(n10333) );
  NAND2_X1 U8699 ( .A1(n10325), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U8700 ( .A1(n10333), .A2(n7541), .ZN(n7542) );
  OR2_X1 U8701 ( .A1(n10325), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10330) );
  XNOR2_X1 U8702 ( .A(n7781), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7543) );
  NOR2_X1 U8703 ( .A1(n10331), .A2(n7543), .ZN(n7782) );
  AOI21_X1 U8704 ( .B1(n10331), .B2(n7543), .A(n7782), .ZN(n7556) );
  AND2_X1 U8705 ( .A1(n10325), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10327) );
  INV_X1 U8706 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7547) );
  NAND2_X1 U8707 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n10312), .ZN(n7546) );
  OAI21_X1 U8708 ( .B1(n10312), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7546), .ZN(
        n10307) );
  AOI21_X1 U8709 ( .B1(n10340), .B2(n7547), .A(n10329), .ZN(n10326) );
  NOR2_X1 U8710 ( .A1(n10327), .A2(n10326), .ZN(n7550) );
  NAND2_X1 U8711 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7781), .ZN(n7548) );
  OAI21_X1 U8712 ( .B1(n7781), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7548), .ZN(
        n7549) );
  NOR2_X1 U8713 ( .A1(n7550), .A2(n7549), .ZN(n7776) );
  AOI211_X1 U8714 ( .C1(n7550), .C2(n7549), .A(n7776), .B(n10305), .ZN(n7551)
         );
  INV_X1 U8715 ( .A(n7551), .ZN(n7555) );
  INV_X1 U8716 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7552) );
  NOR2_X1 U8717 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7552), .ZN(n8283) );
  INV_X1 U8718 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8509) );
  NOR2_X1 U8719 ( .A1(n9776), .A2(n8509), .ZN(n7553) );
  AOI211_X1 U8720 ( .C1(n7781), .C2(n10311), .A(n8283), .B(n7553), .ZN(n7554)
         );
  OAI211_X1 U8721 ( .C1(n7556), .C2(n10332), .A(n7555), .B(n7554), .ZN(
        P1_U3253) );
  XNOR2_X1 U8722 ( .A(n7557), .B(n6818), .ZN(n7574) );
  INV_X1 U8723 ( .A(n7574), .ZN(n10408) );
  INV_X1 U8724 ( .A(n7558), .ZN(n7561) );
  NAND4_X1 U8725 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n7563)
         );
  NAND2_X1 U8726 ( .A1(n6750), .A2(n7565), .ZN(n7595) );
  OR2_X1 U8727 ( .A1(n9079), .A2(n7595), .ZN(n9150) );
  NOR2_X2 U8728 ( .A1(n7566), .A2(n6302), .ZN(n10465) );
  AND2_X1 U8729 ( .A1(n9154), .A2(n10402), .ZN(n7567) );
  NOR2_X1 U8730 ( .A1(n10443), .A2(n7567), .ZN(n10405) );
  NAND2_X1 U8731 ( .A1(n10465), .A2(n10405), .ZN(n7568) );
  OAI21_X1 U8732 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10470), .A(n7568), .ZN(
        n7576) );
  INV_X1 U8733 ( .A(n7892), .ZN(n9160) );
  OAI22_X1 U8734 ( .A1(n8320), .A2(n9068), .B1(n6779), .B2(n9066), .ZN(n7573)
         );
  NAND2_X1 U8735 ( .A1(n7570), .A2(n6818), .ZN(n7571) );
  AOI21_X1 U8736 ( .B1(n7569), .B2(n7571), .A(n9064), .ZN(n7572) );
  AOI211_X1 U8737 ( .C1(n9160), .C2(n7574), .A(n7573), .B(n7572), .ZN(n10407)
         );
  NOR2_X1 U8738 ( .A1(n10407), .A2(n9079), .ZN(n7575) );
  AOI211_X1 U8739 ( .C1(n9079), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7576), .B(
        n7575), .ZN(n7580) );
  INV_X1 U8740 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U8741 ( .A1(n9153), .A2(n10402), .ZN(n7579) );
  OAI211_X1 U8742 ( .C1(n10408), .C2(n9150), .A(n7580), .B(n7579), .ZN(
        P2_U3293) );
  OAI22_X1 U8743 ( .A1(n8778), .A2(n8315), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6393), .ZN(n7582) );
  OAI22_X1 U8744 ( .A1(n8782), .A2(n8556), .B1(n8780), .B2(n7693), .ZN(n7581)
         );
  AOI211_X1 U8745 ( .C1(n7695), .C2(n6759), .A(n7582), .B(n7581), .ZN(n7591)
         );
  INV_X1 U8746 ( .A(n7584), .ZN(n7585) );
  AOI21_X1 U8747 ( .B1(n7583), .B2(n7585), .A(n8759), .ZN(n7589) );
  NOR3_X1 U8748 ( .A1(n8761), .A2(n7586), .A3(n8556), .ZN(n7588) );
  OAI21_X1 U8749 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7590) );
  NAND2_X1 U8750 ( .A1(n7591), .A2(n7590), .ZN(P2_U3223) );
  INV_X1 U8751 ( .A(n9716), .ZN(n9709) );
  INV_X1 U8752 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8337) );
  OAI222_X1 U8753 ( .A1(P1_U3084), .A2(n9709), .B1(n10197), .B2(n7592), .C1(
        n8337), .C2(n10204), .ZN(P1_U3338) );
  INV_X1 U8754 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7593) );
  INV_X1 U8755 ( .A(n8863), .ZN(n8874) );
  OAI222_X1 U8756 ( .A1(n9280), .A2(n7593), .B1(n8529), .B2(n7592), .C1(n8874), 
        .C2(P2_U3152), .ZN(P2_U3343) );
  INV_X1 U8757 ( .A(n7594), .ZN(n7603) );
  NAND2_X1 U8758 ( .A1(n7892), .A2(n7595), .ZN(n7596) );
  OAI21_X1 U8759 ( .B1(n7494), .B2(n10470), .A(n7597), .ZN(n7599) );
  NOR2_X1 U8760 ( .A1(n9164), .A2(n6266), .ZN(n7598) );
  AOI21_X1 U8761 ( .B1(n9164), .B2(n7599), .A(n7598), .ZN(n7602) );
  OAI21_X1 U8762 ( .B1(n9153), .B2(n10465), .A(n7600), .ZN(n7601) );
  OAI211_X1 U8763 ( .C1(n7603), .C2(n10460), .A(n7602), .B(n7601), .ZN(
        P2_U3296) );
  NAND2_X1 U8764 ( .A1(n4894), .A2(n7604), .ZN(n7605) );
  XOR2_X1 U8765 ( .A(n7606), .B(n7605), .Z(n7611) );
  OAI22_X1 U8766 ( .A1(n10481), .A2(n9405), .B1(n9342), .B2(n10483), .ZN(n7607) );
  AOI211_X1 U8767 ( .C1(n10490), .C2(n9408), .A(n7608), .B(n7607), .ZN(n7610)
         );
  NAND2_X1 U8768 ( .A1(n9402), .A2(n10492), .ZN(n7609) );
  OAI211_X1 U8769 ( .C1(n7611), .C2(n9410), .A(n7610), .B(n7609), .ZN(P1_U3225) );
  XOR2_X1 U8770 ( .A(n7612), .B(n7615), .Z(n10360) );
  AOI22_X1 U8771 ( .A1(n9100), .A2(n10360), .B1(n9153), .B2(n7613), .ZN(n7626)
         );
  INV_X1 U8772 ( .A(n7614), .ZN(n7618) );
  INV_X1 U8773 ( .A(n7615), .ZN(n7617) );
  AOI211_X1 U8774 ( .C1(n7618), .C2(n7617), .A(n9064), .B(n7616), .ZN(n7620)
         );
  NOR2_X1 U8775 ( .A1(n7620), .A2(n7619), .ZN(n10357) );
  OAI21_X1 U8776 ( .B1(n7621), .B2(n10470), .A(n10357), .ZN(n7624) );
  OAI21_X1 U8777 ( .B1(n6847), .B2(n7622), .A(n9156), .ZN(n10356) );
  INV_X1 U8778 ( .A(n10356), .ZN(n7623) );
  AOI22_X1 U8779 ( .A1(n7624), .A2(n9164), .B1(n7623), .B2(n10465), .ZN(n7625)
         );
  OAI211_X1 U8780 ( .C1(n7627), .C2(n9164), .A(n7626), .B(n7625), .ZN(P2_U3295) );
  XNOR2_X1 U8781 ( .A(n7628), .B(n7632), .ZN(n7631) );
  NAND2_X1 U8782 ( .A1(n10449), .A2(n10450), .ZN(n7629) );
  OAI21_X1 U8783 ( .B1(n8556), .B2(n9068), .A(n7629), .ZN(n7630) );
  AOI21_X1 U8784 ( .B1(n7631), .B2(n10453), .A(n7630), .ZN(n10544) );
  XNOR2_X1 U8785 ( .A(n7633), .B(n7632), .ZN(n10542) );
  INV_X1 U8786 ( .A(n10465), .ZN(n9040) );
  NAND2_X1 U8787 ( .A1(n7635), .A2(n7634), .ZN(n7636) );
  NAND2_X1 U8788 ( .A1(n5228), .A2(n7636), .ZN(n10540) );
  OAI22_X1 U8789 ( .A1(n9040), .A2(n10540), .B1(n8554), .B2(n10470), .ZN(n7637) );
  AOI21_X1 U8790 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10466), .A(n7637), .ZN(
        n7638) );
  OAI21_X1 U8791 ( .B1(n5227), .B2(n10461), .A(n7638), .ZN(n7639) );
  AOI21_X1 U8792 ( .B1(n9100), .B2(n10542), .A(n7639), .ZN(n7640) );
  OAI21_X1 U8793 ( .B1(n10466), .B2(n10544), .A(n7640), .ZN(P2_U3290) );
  XNOR2_X1 U8794 ( .A(n7641), .B(n7642), .ZN(n7648) );
  INV_X1 U8795 ( .A(n10513), .ZN(n7855) );
  AOI21_X1 U8796 ( .B1(n8028), .B2(n10516), .A(n7643), .ZN(n7646) );
  AOI22_X1 U8797 ( .A1(n9402), .A2(n7644), .B1(n7862), .B2(n9408), .ZN(n7645)
         );
  OAI211_X1 U8798 ( .C1(n7855), .C2(n9342), .A(n7646), .B(n7645), .ZN(n7647)
         );
  AOI21_X1 U8799 ( .B1(n7648), .B2(n9381), .A(n7647), .ZN(n7649) );
  INV_X1 U8800 ( .A(n7649), .ZN(P1_U3237) );
  INV_X1 U8801 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U8802 ( .A1(n10620), .A2(n7650), .ZN(n7651) );
  OAI21_X1 U8803 ( .B1(n10620), .B2(n10643), .A(n7651), .ZN(P2_U3520) );
  INV_X1 U8804 ( .A(n7583), .ZN(n7652) );
  AOI211_X1 U8805 ( .C1(n7654), .C2(n7653), .A(n8759), .B(n7652), .ZN(n7658)
         );
  AOI22_X1 U8806 ( .A1(n10372), .A2(n7672), .B1(n10373), .B2(n8459), .ZN(n7656) );
  AOI22_X1 U8807 ( .A1(n6759), .A2(n7792), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n7655) );
  OAI211_X1 U8808 ( .C1(n7674), .C2(n8780), .A(n7656), .B(n7655), .ZN(n7657)
         );
  OR2_X1 U8809 ( .A1(n7658), .A2(n7657), .ZN(P2_U3215) );
  NOR2_X1 U8810 ( .A1(n10466), .A2(n9106), .ZN(n9145) );
  NOR2_X1 U8811 ( .A1(n10460), .A2(n7659), .ZN(n7664) );
  INV_X1 U8812 ( .A(n7660), .ZN(n8580) );
  INV_X1 U8813 ( .A(n10470), .ZN(n9157) );
  AOI22_X1 U8814 ( .A1(n10466), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8580), .B2(
        n9157), .ZN(n7661) );
  OAI21_X1 U8815 ( .B1(n10461), .B2(n7662), .A(n7661), .ZN(n7663) );
  AOI211_X1 U8816 ( .C1(n7665), .C2(n9145), .A(n7664), .B(n7663), .ZN(n7666)
         );
  OAI21_X1 U8817 ( .B1(n9079), .B2(n7667), .A(n7666), .ZN(P2_U3291) );
  XNOR2_X1 U8818 ( .A(n7669), .B(n7668), .ZN(n7796) );
  OAI21_X1 U8819 ( .B1(n6790), .B2(n7670), .A(n7671), .ZN(n7673) );
  AOI222_X1 U8820 ( .A1(n10453), .A2(n7673), .B1(n8459), .B2(n10448), .C1(
        n7672), .C2(n10450), .ZN(n7795) );
  OR2_X1 U8821 ( .A1(n7795), .A2(n9079), .ZN(n7680) );
  AOI21_X1 U8822 ( .B1(n7792), .B2(n5228), .A(n7692), .ZN(n7793) );
  OAI22_X1 U8823 ( .A1(n9164), .A2(n7675), .B1(n7674), .B2(n10470), .ZN(n7678)
         );
  NOR2_X1 U8824 ( .A1(n10461), .A2(n7676), .ZN(n7677) );
  AOI211_X1 U8825 ( .C1(n7793), .C2(n10465), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI211_X1 U8826 ( .C1(n7796), .C2(n10460), .A(n7680), .B(n7679), .ZN(
        P2_U3289) );
  INV_X1 U8827 ( .A(n7681), .ZN(n7755) );
  AOI22_X1 U8828 ( .A1(n9738), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10195), .ZN(n7682) );
  OAI21_X1 U8829 ( .B1(n7755), .B2(n10197), .A(n7682), .ZN(P1_U3337) );
  OAI21_X1 U8830 ( .B1(n7691), .B2(n7684), .A(n7683), .ZN(n7687) );
  AOI222_X1 U8831 ( .A1(n10453), .A2(n7687), .B1(n7686), .B2(n10448), .C1(
        n7685), .C2(n10450), .ZN(n10575) );
  INV_X1 U8832 ( .A(n7688), .ZN(n7689) );
  AOI21_X1 U8833 ( .B1(n7691), .B2(n7690), .A(n7689), .ZN(n10578) );
  INV_X1 U8834 ( .A(n9145), .ZN(n7879) );
  OAI211_X1 U8835 ( .C1(n10574), .C2(n7692), .A(n10404), .B(n7822), .ZN(n10573) );
  OAI22_X1 U8836 ( .A1(n9164), .A2(n6392), .B1(n7693), .B2(n10470), .ZN(n7694)
         );
  AOI21_X1 U8837 ( .B1(n9153), .B2(n7695), .A(n7694), .ZN(n7696) );
  OAI21_X1 U8838 ( .B1(n7879), .B2(n10573), .A(n7696), .ZN(n7697) );
  AOI21_X1 U8839 ( .B1(n10578), .B2(n9100), .A(n7697), .ZN(n7698) );
  OAI21_X1 U8840 ( .B1(n10575), .B2(n9079), .A(n7698), .ZN(P2_U3288) );
  INV_X1 U8841 ( .A(n7699), .ZN(n7710) );
  NOR2_X1 U8842 ( .A1(n7701), .A2(n7700), .ZN(n7703) );
  NAND4_X1 U8843 ( .A1(n7704), .A2(P1_STATE_REG_SCAN_IN), .A3(n7703), .A4(
        n7702), .ZN(n7864) );
  AOI22_X1 U8844 ( .A1(n10502), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n10491), .ZN(n7709) );
  INV_X1 U8845 ( .A(n7705), .ZN(n10489) );
  AND2_X1 U8846 ( .A1(n7728), .A2(n7706), .ZN(n7707) );
  OAI21_X1 U8847 ( .B1(n10045), .B2(n10526), .A(n7741), .ZN(n7708) );
  OAI211_X1 U8848 ( .C1(n7710), .C2(n10502), .A(n7709), .B(n7708), .ZN(
        P1_U3291) );
  INV_X1 U8849 ( .A(n7711), .ZN(n7713) );
  NAND2_X1 U8850 ( .A1(n7714), .A2(n7741), .ZN(n7734) );
  XNOR2_X1 U8851 ( .A(n5159), .B(n7734), .ZN(n10348) );
  NOR2_X1 U8852 ( .A1(n7715), .A2(n9900), .ZN(n7716) );
  NAND2_X1 U8853 ( .A1(n10536), .A2(n7716), .ZN(n10431) );
  INV_X1 U8854 ( .A(n7747), .ZN(n7719) );
  AOI21_X1 U8855 ( .B1(n7721), .B2(n7720), .A(n7719), .ZN(n7726) );
  NAND2_X1 U8856 ( .A1(n7722), .A2(n10494), .ZN(n7725) );
  NAND2_X1 U8857 ( .A1(n7723), .A2(n9659), .ZN(n7724) );
  OAI222_X1 U8858 ( .A1(n10482), .A2(n7727), .B1(n10519), .B2(n10348), .C1(
        n7726), .C2(n10479), .ZN(n10350) );
  XNOR2_X1 U8859 ( .A(n7742), .B(n4879), .ZN(n7729) );
  AOI22_X1 U8860 ( .A1(n7729), .A2(n10562), .B1(n10514), .B2(n9679), .ZN(
        n10349) );
  INV_X1 U8861 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7730) );
  OAI22_X1 U8862 ( .A1(n10349), .A2(n10494), .B1(n10531), .B2(n7730), .ZN(
        n7731) );
  OAI21_X1 U8863 ( .B1(n10350), .B2(n7731), .A(n10536), .ZN(n7733) );
  INV_X2 U8864 ( .A(n10536), .ZN(n10502) );
  AOI22_X1 U8865 ( .A1(n10045), .A2(n4879), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n10502), .ZN(n7732) );
  OAI211_X1 U8866 ( .C1(n10348), .C2(n10431), .A(n7733), .B(n7732), .ZN(
        P1_U3290) );
  NAND2_X1 U8867 ( .A1(n9680), .A2(n4879), .ZN(n7735) );
  NAND2_X1 U8868 ( .A1(n7735), .A2(n7734), .ZN(n7738) );
  NAND2_X1 U8869 ( .A1(n7738), .A2(n7737), .ZN(n7757) );
  XNOR2_X1 U8870 ( .A(n7757), .B(n7748), .ZN(n10363) );
  INV_X1 U8871 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7740) );
  INV_X1 U8872 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7739) );
  OAI22_X1 U8873 ( .A1(n10536), .A2(n7740), .B1(n7739), .B2(n10531), .ZN(n7745) );
  INV_X1 U8874 ( .A(n10526), .ZN(n10430) );
  OAI21_X1 U8875 ( .B1(n7741), .B2(n4879), .A(n5162), .ZN(n7743) );
  NAND2_X1 U8876 ( .A1(n7743), .A2(n7769), .ZN(n10365) );
  NOR2_X1 U8877 ( .A1(n10430), .A2(n10365), .ZN(n7744) );
  AOI211_X1 U8878 ( .C1(n10045), .C2(n5162), .A(n7745), .B(n7744), .ZN(n7754)
         );
  OAI21_X1 U8879 ( .B1(n7749), .B2(n7748), .A(n7763), .ZN(n7750) );
  NAND2_X1 U8880 ( .A1(n7750), .A2(n10511), .ZN(n7752) );
  AOI22_X1 U8881 ( .A1(n7760), .A2(n10514), .B1(n10515), .B2(n9680), .ZN(n7751) );
  OAI211_X1 U8882 ( .C1(n10363), .C2(n10519), .A(n7752), .B(n7751), .ZN(n10366) );
  NAND2_X1 U8883 ( .A1(n10366), .A2(n10536), .ZN(n7753) );
  OAI211_X1 U8884 ( .C1(n10363), .C2(n10431), .A(n7754), .B(n7753), .ZN(
        P1_U3289) );
  INV_X1 U8885 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7756) );
  INV_X1 U8886 ( .A(n8884), .ZN(n8889) );
  OAI222_X1 U8887 ( .A1(n9280), .A2(n7756), .B1(n8529), .B2(n7755), .C1(
        P2_U3152), .C2(n8889), .ZN(P2_U3342) );
  NAND2_X1 U8888 ( .A1(n7757), .A2(n9511), .ZN(n7759) );
  NAND2_X1 U8889 ( .A1(n7761), .A2(n10364), .ZN(n7758) );
  NAND2_X1 U8890 ( .A1(n7759), .A2(n7758), .ZN(n7845) );
  NAND2_X1 U8891 ( .A1(n10418), .A2(n7773), .ZN(n9624) );
  NAND2_X1 U8892 ( .A1(n7760), .A2(n7846), .ZN(n9627) );
  NAND2_X1 U8893 ( .A1(n9624), .A2(n9627), .ZN(n7844) );
  INV_X1 U8894 ( .A(n7844), .ZN(n9510) );
  XNOR2_X1 U8895 ( .A(n7845), .B(n9510), .ZN(n10393) );
  NAND2_X1 U8896 ( .A1(n7761), .A2(n5162), .ZN(n7762) );
  NAND2_X1 U8897 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  OAI21_X1 U8898 ( .B1(n9510), .B2(n7764), .A(n7856), .ZN(n7765) );
  NAND2_X1 U8899 ( .A1(n7765), .A2(n10511), .ZN(n7767) );
  AOI22_X1 U8900 ( .A1(n10514), .A2(n9678), .B1(n9679), .B2(n10515), .ZN(n7766) );
  OAI211_X1 U8901 ( .C1(n10393), .C2(n10519), .A(n7767), .B(n7766), .ZN(n10398) );
  NAND2_X1 U8902 ( .A1(n10398), .A2(n10536), .ZN(n7775) );
  OAI22_X1 U8903 ( .A1(n10536), .A2(n7768), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10531), .ZN(n7772) );
  AND2_X1 U8904 ( .A1(n7769), .A2(n7773), .ZN(n7770) );
  OR2_X1 U8905 ( .A1(n7770), .A2(n10423), .ZN(n10395) );
  NOR2_X1 U8906 ( .A1(n10430), .A2(n10395), .ZN(n7771) );
  AOI211_X1 U8907 ( .C1(n10045), .C2(n7773), .A(n7772), .B(n7771), .ZN(n7774)
         );
  OAI211_X1 U8908 ( .C1(n10393), .C2(n10431), .A(n7775), .B(n7774), .ZN(
        P1_U3288) );
  INV_X1 U8909 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U8910 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7801), .ZN(n7777) );
  OAI21_X1 U8911 ( .B1(n7801), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7777), .ZN(
        n7778) );
  AOI211_X1 U8912 ( .C1(n7779), .C2(n7778), .A(n7800), .B(n10305), .ZN(n7780)
         );
  AOI21_X1 U8913 ( .B1(n10311), .B2(n7801), .A(n7780), .ZN(n7790) );
  XNOR2_X1 U8914 ( .A(n7801), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7786) );
  INV_X1 U8915 ( .A(n7781), .ZN(n7784) );
  INV_X1 U8916 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7783) );
  AOI21_X1 U8917 ( .B1(n7784), .B2(n7783), .A(n7782), .ZN(n7785) );
  NOR2_X1 U8918 ( .A1(n7785), .A2(n7786), .ZN(n7806) );
  AOI21_X1 U8919 ( .B1(n7786), .B2(n7785), .A(n7806), .ZN(n7787) );
  NOR2_X1 U8920 ( .A1(n10332), .A2(n7787), .ZN(n7788) );
  AND2_X1 U8921 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8416) );
  NOR2_X1 U8922 ( .A1(n7788), .A2(n8416), .ZN(n7789) );
  OAI211_X1 U8923 ( .C1(n7791), .C2(n9776), .A(n7790), .B(n7789), .ZN(P1_U3254) );
  INV_X1 U8924 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7798) );
  AOI22_X1 U8925 ( .A1(n7793), .A2(n10404), .B1(n10403), .B2(n7792), .ZN(n7794) );
  OAI211_X1 U8926 ( .C1(n9245), .C2(n7796), .A(n7795), .B(n7794), .ZN(n9248)
         );
  NAND2_X1 U8927 ( .A1(n9248), .A2(n10624), .ZN(n7797) );
  OAI21_X1 U8928 ( .B1(n10624), .B2(n7798), .A(n7797), .ZN(P2_U3472) );
  NOR2_X1 U8929 ( .A1(n8003), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7799) );
  AOI21_X1 U8930 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8003), .A(n7799), .ZN(
        n7803) );
  OAI21_X1 U8931 ( .B1(n7803), .B2(n7802), .A(n8002), .ZN(n7814) );
  INV_X1 U8932 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U8933 ( .A1(n10311), .A2(n8003), .ZN(n7804) );
  NAND2_X1 U8934 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9290) );
  OAI211_X1 U8935 ( .C1(n9776), .C2(n7805), .A(n7804), .B(n9290), .ZN(n7813)
         );
  INV_X1 U8936 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7808) );
  AOI21_X1 U8937 ( .B1(n7808), .B2(n7807), .A(n7806), .ZN(n7810) );
  INV_X1 U8938 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8007) );
  AOI22_X1 U8939 ( .A1(n8003), .A2(n8007), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8008), .ZN(n7809) );
  NOR2_X1 U8940 ( .A1(n7810), .A2(n7809), .ZN(n8006) );
  AOI21_X1 U8941 ( .B1(n7810), .B2(n7809), .A(n8006), .ZN(n7811) );
  NOR2_X1 U8942 ( .A1(n7811), .A2(n10332), .ZN(n7812) );
  AOI211_X1 U8943 ( .C1(n7814), .C2(n10336), .A(n7813), .B(n7812), .ZN(n7815)
         );
  INV_X1 U8944 ( .A(n7815), .ZN(P1_U3255) );
  OAI21_X1 U8945 ( .B1(n7817), .B2(n7885), .A(n7816), .ZN(n7934) );
  INV_X1 U8946 ( .A(n7934), .ZN(n7828) );
  XNOR2_X1 U8947 ( .A(n7886), .B(n7885), .ZN(n7820) );
  OAI22_X1 U8948 ( .A1(n8468), .A2(n9066), .B1(n8460), .B2(n9068), .ZN(n7818)
         );
  AOI21_X1 U8949 ( .B1(n7934), .B2(n9160), .A(n7818), .ZN(n7819) );
  OAI21_X1 U8950 ( .B1(n7820), .B2(n9064), .A(n7819), .ZN(n7932) );
  NAND2_X1 U8951 ( .A1(n7932), .A2(n9164), .ZN(n7827) );
  OAI22_X1 U8952 ( .A1(n9164), .A2(n7821), .B1(n8462), .B2(n10470), .ZN(n7825)
         );
  INV_X1 U8953 ( .A(n7822), .ZN(n7823) );
  INV_X1 U8954 ( .A(n8476), .ZN(n7930) );
  OAI21_X1 U8955 ( .B1(n7823), .B2(n7930), .A(n7895), .ZN(n7931) );
  NOR2_X1 U8956 ( .A1(n7931), .A2(n9040), .ZN(n7824) );
  AOI211_X1 U8957 ( .C1(n9153), .C2(n8476), .A(n7825), .B(n7824), .ZN(n7826)
         );
  OAI211_X1 U8958 ( .C1(n7828), .C2(n9150), .A(n7827), .B(n7826), .ZN(P2_U3287) );
  INV_X1 U8959 ( .A(n7829), .ZN(n7841) );
  AOI22_X1 U8960 ( .A1(n9751), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10195), .ZN(n7830) );
  OAI21_X1 U8961 ( .B1(n7841), .B2(n10197), .A(n7830), .ZN(P1_U3336) );
  AOI21_X1 U8962 ( .B1(n7073), .B2(n4991), .A(n8759), .ZN(n7835) );
  NOR3_X1 U8963 ( .A1(n7832), .A2(n8460), .A3(n8761), .ZN(n7834) );
  OAI21_X1 U8964 ( .B1(n7835), .B2(n7834), .A(n7833), .ZN(n7840) );
  INV_X1 U8965 ( .A(n7874), .ZN(n7838) );
  INV_X1 U8966 ( .A(n8766), .ZN(n8738) );
  OAI22_X1 U8967 ( .A1(n8460), .A2(n9066), .B1(n8326), .B2(n9068), .ZN(n7870)
         );
  INV_X1 U8968 ( .A(n7870), .ZN(n7836) );
  OAI22_X1 U8969 ( .A1(n8738), .A2(n7836), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8792), .ZN(n7837) );
  AOI21_X1 U8970 ( .B1(n7838), .B2(n8740), .A(n7837), .ZN(n7839) );
  OAI211_X1 U8971 ( .C1(n7952), .C2(n8743), .A(n7840), .B(n7839), .ZN(P2_U3238) );
  INV_X1 U8972 ( .A(n8899), .ZN(n8905) );
  OAI222_X1 U8973 ( .A1(P2_U3152), .A2(n8905), .B1(n9280), .B2(n7842), .C1(
        n7841), .C2(n8529), .ZN(P2_U3341) );
  AND2_X1 U8974 ( .A1(n10519), .A2(n9900), .ZN(n7843) );
  NOR2_X1 U8975 ( .A1(n5508), .A2(n7843), .ZN(n10499) );
  NAND2_X1 U8976 ( .A1(n7845), .A2(n7844), .ZN(n7848) );
  NAND2_X1 U8977 ( .A1(n10418), .A2(n7846), .ZN(n7847) );
  NAND2_X1 U8978 ( .A1(n7848), .A2(n7847), .ZN(n10412) );
  NAND2_X1 U8979 ( .A1(n10412), .A2(n10413), .ZN(n7850) );
  NAND2_X1 U8980 ( .A1(n10481), .A2(n10434), .ZN(n7849) );
  NAND2_X1 U8981 ( .A1(n7850), .A2(n7849), .ZN(n10475) );
  NAND2_X1 U8982 ( .A1(n10417), .A2(n10490), .ZN(n9630) );
  NAND2_X1 U8983 ( .A1(n10516), .A2(n10490), .ZN(n7852) );
  NAND2_X1 U8984 ( .A1(n10483), .A2(n7862), .ZN(n9632) );
  INV_X1 U8985 ( .A(n10483), .ZN(n9677) );
  NAND2_X1 U8986 ( .A1(n10529), .A2(n9677), .ZN(n7917) );
  NAND2_X1 U8987 ( .A1(n10483), .A2(n10529), .ZN(n7854) );
  OR2_X1 U8988 ( .A1(n10548), .A2(n7855), .ZN(n9423) );
  NAND2_X1 U8989 ( .A1(n10548), .A2(n7855), .ZN(n9422) );
  NAND2_X1 U8990 ( .A1(n9423), .A2(n9422), .ZN(n7913) );
  INV_X1 U8991 ( .A(n7913), .ZN(n9513) );
  XNOR2_X1 U8992 ( .A(n7914), .B(n9513), .ZN(n10551) );
  NAND2_X1 U8993 ( .A1(n9678), .A2(n10434), .ZN(n9626) );
  NAND2_X1 U8994 ( .A1(n10415), .A2(n9626), .ZN(n7858) );
  NAND2_X1 U8995 ( .A1(n10481), .A2(n7857), .ZN(n9629) );
  INV_X1 U8996 ( .A(n10476), .ZN(n7859) );
  OAI21_X2 U8997 ( .B1(n10478), .B2(n7859), .A(n9634), .ZN(n10510) );
  NAND2_X1 U8998 ( .A1(n7918), .A2(n7917), .ZN(n7860) );
  XNOR2_X1 U8999 ( .A(n7860), .B(n9513), .ZN(n7861) );
  OAI222_X1 U9000 ( .A1(n10484), .A2(n7919), .B1(n10482), .B2(n10483), .C1(
        n10479), .C2(n7861), .ZN(n10552) );
  NAND2_X1 U9001 ( .A1(n10552), .A2(n10536), .ZN(n7868) );
  AND2_X1 U9002 ( .A1(n10423), .A2(n10434), .ZN(n10477) );
  NAND2_X1 U9003 ( .A1(n10477), .A2(n7851), .ZN(n10506) );
  INV_X1 U9004 ( .A(n10049), .ZN(n7863) );
  AOI211_X1 U9005 ( .C1(n10548), .C2(n10507), .A(n10583), .B(n7863), .ZN(
        n10547) );
  OR2_X1 U9006 ( .A1(n7864), .A2(n10494), .ZN(n8052) );
  INV_X1 U9007 ( .A(n8052), .ZN(n10003) );
  AOI22_X1 U9008 ( .A1(n10502), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7904), .B2(
        n10491), .ZN(n7865) );
  OAI21_X1 U9009 ( .B1(n5122), .B2(n10530), .A(n7865), .ZN(n7866) );
  AOI21_X1 U9010 ( .B1(n10547), .B2(n10003), .A(n7866), .ZN(n7867) );
  OAI211_X1 U9011 ( .C1(n10012), .C2(n10551), .A(n7868), .B(n7867), .ZN(
        P1_U3284) );
  XNOR2_X1 U9012 ( .A(n7869), .B(n7872), .ZN(n7871) );
  AOI21_X1 U9013 ( .B1(n7871), .B2(n10453), .A(n7870), .ZN(n7951) );
  XNOR2_X1 U9014 ( .A(n7873), .B(n7872), .ZN(n7954) );
  OAI211_X1 U9015 ( .C1(n7952), .C2(n7897), .A(n10404), .B(n7963), .ZN(n7950)
         );
  OAI22_X1 U9016 ( .A1(n9164), .A2(n7875), .B1(n7874), .B2(n10470), .ZN(n7876)
         );
  AOI21_X1 U9017 ( .B1(n7877), .B2(n9153), .A(n7876), .ZN(n7878) );
  OAI21_X1 U9018 ( .B1(n7950), .B2(n7879), .A(n7878), .ZN(n7880) );
  AOI21_X1 U9019 ( .B1(n7954), .B2(n9100), .A(n7880), .ZN(n7881) );
  OAI21_X1 U9020 ( .B1(n9079), .B2(n7951), .A(n7881), .ZN(P2_U3285) );
  OAI21_X1 U9021 ( .B1(n4950), .B2(n7887), .A(n7882), .ZN(n10597) );
  OAI22_X1 U9022 ( .A1(n8322), .A2(n9068), .B1(n8315), .B2(n9066), .ZN(n7883)
         );
  INV_X1 U9023 ( .A(n7883), .ZN(n7891) );
  OAI21_X1 U9024 ( .B1(n7886), .B2(n7885), .A(n7884), .ZN(n7888) );
  XNOR2_X1 U9025 ( .A(n7888), .B(n7887), .ZN(n7889) );
  NAND2_X1 U9026 ( .A1(n7889), .A2(n10453), .ZN(n7890) );
  OAI211_X1 U9027 ( .C1(n10597), .C2(n7892), .A(n7891), .B(n7890), .ZN(n10602)
         );
  NAND2_X1 U9028 ( .A1(n10602), .A2(n9164), .ZN(n7902) );
  OAI22_X1 U9029 ( .A1(n9164), .A2(n7894), .B1(n7893), .B2(n10470), .ZN(n7899)
         );
  AND2_X1 U9030 ( .A1(n7900), .A2(n7895), .ZN(n7896) );
  OR2_X1 U9031 ( .A1(n7897), .A2(n7896), .ZN(n10599) );
  NOR2_X1 U9032 ( .A1(n10599), .A2(n9040), .ZN(n7898) );
  AOI211_X1 U9033 ( .C1(n9153), .C2(n7900), .A(n7899), .B(n7898), .ZN(n7901)
         );
  OAI211_X1 U9034 ( .C1(n10597), .C2(n9150), .A(n7902), .B(n7901), .ZN(
        P2_U3286) );
  AOI21_X1 U9035 ( .B1(n8028), .B2(n9677), .A(n7903), .ZN(n7906) );
  NAND2_X1 U9036 ( .A1(n9402), .A2(n7904), .ZN(n7905) );
  OAI211_X1 U9037 ( .C1(n7919), .C2(n9342), .A(n7906), .B(n7905), .ZN(n7911)
         );
  XOR2_X1 U9038 ( .A(n7908), .B(n7907), .Z(n7909) );
  NOR2_X1 U9039 ( .A1(n7909), .A2(n9410), .ZN(n7910) );
  AOI211_X1 U9040 ( .C1(n10548), .C2(n9408), .A(n7911), .B(n7910), .ZN(n7912)
         );
  INV_X1 U9041 ( .A(n7912), .ZN(P1_U3211) );
  NAND2_X1 U9042 ( .A1(n10560), .A2(n7919), .ZN(n9428) );
  NAND2_X1 U9043 ( .A1(n10033), .A2(n9428), .ZN(n10046) );
  NAND2_X1 U9044 ( .A1(n10047), .A2(n10046), .ZN(n10565) );
  INV_X1 U9045 ( .A(n7919), .ZN(n9676) );
  NAND2_X1 U9046 ( .A1(n10560), .A2(n9676), .ZN(n7915) );
  INV_X1 U9047 ( .A(n8034), .ZN(n10582) );
  AND2_X1 U9048 ( .A1(n10582), .A2(n10039), .ZN(n9431) );
  INV_X1 U9049 ( .A(n10039), .ZN(n7976) );
  NAND2_X1 U9050 ( .A1(n8034), .A2(n7976), .ZN(n9550) );
  INV_X1 U9051 ( .A(n9550), .ZN(n7916) );
  XNOR2_X1 U9052 ( .A(n8035), .B(n9427), .ZN(n7923) );
  AND2_X1 U9053 ( .A1(n9423), .A2(n7917), .ZN(n9636) );
  NAND2_X1 U9054 ( .A1(n7918), .A2(n9636), .ZN(n9559) );
  AND2_X1 U9055 ( .A1(n9428), .A2(n9422), .ZN(n9554) );
  XNOR2_X1 U9056 ( .A(n8039), .B(n9427), .ZN(n7921) );
  OAI22_X1 U9057 ( .A1(n8064), .A2(n10484), .B1(n7919), .B2(n10482), .ZN(n7920) );
  AOI21_X1 U9058 ( .B1(n7921), .B2(n10511), .A(n7920), .ZN(n7922) );
  OAI21_X1 U9059 ( .B1(n10519), .B2(n7923), .A(n7922), .ZN(n10585) );
  INV_X1 U9060 ( .A(n10585), .ZN(n7929) );
  INV_X1 U9061 ( .A(n7923), .ZN(n10587) );
  INV_X1 U9062 ( .A(n10431), .ZN(n10527) );
  NOR2_X1 U9063 ( .A1(n10051), .A2(n10582), .ZN(n7924) );
  OR2_X1 U9064 ( .A1(n8045), .A2(n7924), .ZN(n10584) );
  AOI22_X1 U9065 ( .A1(n10502), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7941), .B2(
        n10491), .ZN(n7926) );
  NAND2_X1 U9066 ( .A1(n8034), .A2(n10045), .ZN(n7925) );
  OAI211_X1 U9067 ( .C1(n10584), .C2(n10430), .A(n7926), .B(n7925), .ZN(n7927)
         );
  AOI21_X1 U9068 ( .B1(n10587), .B2(n10527), .A(n7927), .ZN(n7928) );
  OAI21_X1 U9069 ( .B1(n7929), .B2(n10502), .A(n7928), .ZN(P1_U3282) );
  OAI22_X1 U9070 ( .A1(n7931), .A2(n10613), .B1(n7930), .B2(n10611), .ZN(n7933) );
  AOI211_X1 U9071 ( .C1(n10391), .C2(n7934), .A(n7933), .B(n7932), .ZN(n7947)
         );
  NAND2_X1 U9072 ( .A1(n10619), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7935) );
  OAI21_X1 U9073 ( .B1(n7947), .B2(n10619), .A(n7935), .ZN(P2_U3529) );
  INV_X1 U9074 ( .A(n8917), .ZN(n8915) );
  INV_X1 U9075 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7936) );
  OAI222_X1 U9076 ( .A1(P2_U3152), .A2(n8915), .B1(n8529), .B2(n8531), .C1(
        n7936), .C2(n9280), .ZN(P2_U3340) );
  NAND2_X1 U9077 ( .A1(n7937), .A2(n7978), .ZN(n7938) );
  AOI21_X1 U9078 ( .B1(n7939), .B2(n7938), .A(n5396), .ZN(n7946) );
  AOI21_X1 U9079 ( .B1(n8028), .B2(n9676), .A(n7940), .ZN(n7943) );
  NAND2_X1 U9080 ( .A1(n9402), .A2(n7941), .ZN(n7942) );
  OAI211_X1 U9081 ( .C1(n8064), .C2(n9342), .A(n7943), .B(n7942), .ZN(n7944)
         );
  AOI21_X1 U9082 ( .B1(n8034), .B2(n9408), .A(n7944), .ZN(n7945) );
  OAI21_X1 U9083 ( .B1(n7946), .B2(n9410), .A(n7945), .ZN(P1_U3229) );
  INV_X1 U9084 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7949) );
  OR2_X1 U9085 ( .A1(n7947), .A2(n10621), .ZN(n7948) );
  OAI21_X1 U9086 ( .B1(n10624), .B2(n7949), .A(n7948), .ZN(P2_U3478) );
  OAI211_X1 U9087 ( .C1(n7952), .C2(n10611), .A(n7951), .B(n7950), .ZN(n7953)
         );
  AOI21_X1 U9088 ( .B1(n7954), .B2(n10617), .A(n7953), .ZN(n7958) );
  NAND2_X1 U9089 ( .A1(n10619), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7955) );
  OAI21_X1 U9090 ( .B1(n7958), .B2(n10619), .A(n7955), .ZN(P2_U3531) );
  INV_X1 U9091 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7956) );
  OR2_X1 U9092 ( .A1(n10624), .A2(n7956), .ZN(n7957) );
  OAI21_X1 U9093 ( .B1(n7958), .B2(n10621), .A(n7957), .ZN(P2_U3484) );
  XNOR2_X1 U9094 ( .A(n7959), .B(n7961), .ZN(n7960) );
  OAI222_X1 U9095 ( .A1(n9068), .A2(n8338), .B1(n9066), .B2(n8322), .C1(n7960), 
        .C2(n9064), .ZN(n10606) );
  INV_X1 U9096 ( .A(n10606), .ZN(n7969) );
  XNOR2_X1 U9097 ( .A(n7962), .B(n7961), .ZN(n10608) );
  OAI21_X1 U9098 ( .B1(n5212), .B2(n5213), .A(n8127), .ZN(n10605) );
  OAI22_X1 U9099 ( .A1(n9164), .A2(n7964), .B1(n7985), .B2(n10470), .ZN(n7965)
         );
  AOI21_X1 U9100 ( .B1(n8000), .B2(n9153), .A(n7965), .ZN(n7966) );
  OAI21_X1 U9101 ( .B1(n10605), .B2(n9040), .A(n7966), .ZN(n7967) );
  AOI21_X1 U9102 ( .B1(n10608), .B2(n9100), .A(n7967), .ZN(n7968) );
  OAI21_X1 U9103 ( .B1(n7969), .B2(n9079), .A(n7968), .ZN(P2_U3284) );
  INV_X1 U9104 ( .A(n7970), .ZN(n7971) );
  INV_X1 U9105 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8369) );
  OAI222_X1 U9106 ( .A1(n9900), .A2(P1_U3084), .B1(n10197), .B2(n7971), .C1(
        n10204), .C2(n8369), .ZN(P1_U3334) );
  INV_X1 U9107 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7972) );
  OAI222_X1 U9108 ( .A1(n9280), .A2(n7972), .B1(n8529), .B2(n7971), .C1(n8993), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U9109 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7973) );
  NOR2_X1 U9110 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7973), .ZN(n9696) );
  AOI21_X1 U9111 ( .B1(n8028), .B2(n10513), .A(n9696), .ZN(n7975) );
  NAND2_X1 U9112 ( .A1(n9402), .A2(n10042), .ZN(n7974) );
  OAI211_X1 U9113 ( .C1(n7976), .C2(n9342), .A(n7975), .B(n7974), .ZN(n7983)
         );
  NAND2_X1 U9114 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  XOR2_X1 U9115 ( .A(n7980), .B(n7979), .Z(n7981) );
  NOR2_X1 U9116 ( .A1(n7981), .A2(n9410), .ZN(n7982) );
  AOI211_X1 U9117 ( .C1(n10560), .C2(n9408), .A(n7983), .B(n7982), .ZN(n7984)
         );
  INV_X1 U9118 ( .A(n7984), .ZN(P1_U3219) );
  INV_X1 U9119 ( .A(n7985), .ZN(n7986) );
  AOI22_X1 U9120 ( .A1(n10372), .A2(n7987), .B1(n8740), .B2(n7986), .ZN(n7990)
         );
  NOR2_X1 U9121 ( .A1(n7988), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8809) );
  INV_X1 U9122 ( .A(n8809), .ZN(n7989) );
  OAI211_X1 U9123 ( .C1(n8338), .C2(n8778), .A(n7990), .B(n7989), .ZN(n7999)
         );
  NOR3_X1 U9124 ( .A1(n4990), .A2(n7991), .A3(n8759), .ZN(n7997) );
  INV_X1 U9125 ( .A(n8761), .ZN(n8750) );
  INV_X1 U9126 ( .A(n8326), .ZN(n8123) );
  NAND3_X1 U9127 ( .A1(n7992), .A2(n8750), .A3(n8123), .ZN(n7993) );
  OAI21_X1 U9128 ( .B1(n7994), .B2(n8759), .A(n7993), .ZN(n7996) );
  MUX2_X1 U9129 ( .A(n7997), .B(n7996), .S(n7995), .Z(n7998) );
  AOI211_X1 U9130 ( .C1(n8000), .C2(n6759), .A(n7999), .B(n7998), .ZN(n8001)
         );
  INV_X1 U9131 ( .A(n8001), .ZN(P2_U3226) );
  OAI21_X1 U9132 ( .B1(n8003), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8002), .ZN(
        n9708) );
  XNOR2_X1 U9133 ( .A(n9708), .B(n9709), .ZN(n8005) );
  INV_X1 U9134 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8004) );
  NOR2_X1 U9135 ( .A1(n8004), .A2(n8005), .ZN(n9710) );
  AOI211_X1 U9136 ( .C1(n8005), .C2(n8004), .A(n9710), .B(n10305), .ZN(n8014)
         );
  INV_X1 U9137 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8517) );
  AOI21_X1 U9138 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n9715) );
  XNOR2_X1 U9139 ( .A(n9715), .B(n9709), .ZN(n8009) );
  NAND2_X1 U9140 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n8009), .ZN(n9717) );
  OAI211_X1 U9141 ( .C1(n8009), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10315), .B(
        n9717), .ZN(n8012) );
  NAND2_X1 U9142 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8548) );
  INV_X1 U9143 ( .A(n8548), .ZN(n8010) );
  AOI21_X1 U9144 ( .B1(n10311), .B2(n9716), .A(n8010), .ZN(n8011) );
  OAI211_X1 U9145 ( .C1(n8517), .C2(n9776), .A(n8012), .B(n8011), .ZN(n8013)
         );
  OR2_X1 U9146 ( .A1(n8014), .A2(n8013), .ZN(P1_U3256) );
  INV_X1 U9147 ( .A(n8015), .ZN(n8569) );
  OAI222_X1 U9148 ( .A1(P1_U3084), .A2(n8016), .B1(n10197), .B2(n8569), .C1(
        n8348), .C2(n10204), .ZN(P1_U3333) );
  OAI21_X1 U9149 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8020) );
  NAND2_X1 U9150 ( .A1(n8020), .A2(n10375), .ZN(n8023) );
  AND2_X1 U9151 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8831) );
  OAI22_X1 U9152 ( .A1(n8782), .A2(n8326), .B1(n8780), .B2(n8132), .ZN(n8021)
         );
  AOI211_X1 U9153 ( .C1(n10373), .C2(n8124), .A(n8831), .B(n8021), .ZN(n8022)
         );
  OAI211_X1 U9154 ( .C1(n8135), .C2(n8743), .A(n8023), .B(n8022), .ZN(P2_U3236) );
  NAND2_X1 U9155 ( .A1(n8024), .A2(n4893), .ZN(n8026) );
  XNOR2_X1 U9156 ( .A(n8026), .B(n8025), .ZN(n8033) );
  NOR2_X1 U9157 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8027), .ZN(n10310) );
  AOI21_X1 U9158 ( .B1(n8028), .B2(n10039), .A(n10310), .ZN(n8030) );
  NAND2_X1 U9159 ( .A1(n9402), .A2(n8047), .ZN(n8029) );
  OAI211_X1 U9160 ( .C1(n8379), .C2(n9342), .A(n8030), .B(n8029), .ZN(n8031)
         );
  AOI21_X1 U9161 ( .B1(n8109), .B2(n9408), .A(n8031), .ZN(n8032) );
  OAI21_X1 U9162 ( .B1(n8033), .B2(n9410), .A(n8032), .ZN(P1_U3215) );
  OAI222_X1 U9163 ( .A1(P1_U3084), .A2(n9620), .B1(n10197), .B2(n8056), .C1(
        n8344), .C2(n10204), .ZN(P1_U3332) );
  OR2_X1 U9164 ( .A1(n8109), .A2(n8064), .ZN(n9560) );
  NAND2_X1 U9165 ( .A1(n8109), .A2(n8064), .ZN(n9434) );
  INV_X1 U9166 ( .A(n8069), .ZN(n8038) );
  AOI21_X1 U9167 ( .B1(n9518), .B2(n8036), .A(n8038), .ZN(n8112) );
  INV_X1 U9168 ( .A(n9431), .ZN(n8040) );
  NAND2_X1 U9169 ( .A1(n8041), .A2(n9550), .ZN(n8042) );
  OAI21_X1 U9170 ( .B1(n9518), .B2(n8042), .A(n8071), .ZN(n8043) );
  INV_X1 U9171 ( .A(n8379), .ZN(n9674) );
  AOI222_X1 U9172 ( .A1(n10511), .A2(n8043), .B1(n10039), .B2(n10515), .C1(
        n9674), .C2(n10514), .ZN(n8111) );
  INV_X1 U9173 ( .A(n8111), .ZN(n8054) );
  INV_X1 U9174 ( .A(n8109), .ZN(n8044) );
  OAI21_X1 U9175 ( .B1(n8045), .B2(n8044), .A(n10562), .ZN(n8046) );
  OR2_X1 U9176 ( .A1(n8075), .A2(n8046), .ZN(n8107) );
  INV_X1 U9177 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8049) );
  INV_X1 U9178 ( .A(n8047), .ZN(n8048) );
  OAI22_X1 U9179 ( .A1(n10536), .A2(n8049), .B1(n8048), .B2(n10531), .ZN(n8050) );
  AOI21_X1 U9180 ( .B1(n8109), .B2(n10045), .A(n8050), .ZN(n8051) );
  OAI21_X1 U9181 ( .B1(n8107), .B2(n8052), .A(n8051), .ZN(n8053) );
  AOI21_X1 U9182 ( .B1(n8054), .B2(n10536), .A(n8053), .ZN(n8055) );
  OAI21_X1 U9183 ( .B1(n10012), .B2(n8112), .A(n8055), .ZN(P1_U3281) );
  OAI222_X1 U9184 ( .A1(n9280), .A2(n8058), .B1(P2_U3152), .B2(n8057), .C1(
        n8529), .C2(n8056), .ZN(P2_U3337) );
  INV_X1 U9185 ( .A(n9439), .ZN(n8081) );
  AOI21_X1 U9186 ( .B1(n8060), .B2(n8059), .A(n9410), .ZN(n8062) );
  NAND2_X1 U9187 ( .A1(n8062), .A2(n8061), .ZN(n8067) );
  AND2_X1 U9188 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10323) );
  AOI21_X1 U9189 ( .B1(n9401), .B2(n8357), .A(n10323), .ZN(n8063) );
  OAI21_X1 U9190 ( .B1(n8064), .B2(n9405), .A(n8063), .ZN(n8065) );
  AOI21_X1 U9191 ( .B1(n8078), .B2(n9402), .A(n8065), .ZN(n8066) );
  OAI211_X1 U9192 ( .C1(n8081), .C2(n9388), .A(n8067), .B(n8066), .ZN(P1_U3234) );
  INV_X1 U9193 ( .A(n10519), .ZN(n10555) );
  OR2_X1 U9194 ( .A1(n8109), .A2(n9675), .ZN(n8068) );
  NAND2_X1 U9195 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  XNOR2_X1 U9196 ( .A(n9439), .B(n8379), .ZN(n9520) );
  OAI21_X1 U9197 ( .B1(n8070), .B2(n9520), .A(n8351), .ZN(n8289) );
  XNOR2_X1 U9198 ( .A(n8349), .B(n9520), .ZN(n8073) );
  AOI22_X1 U9199 ( .A1(n10514), .A2(n8357), .B1(n9675), .B2(n10515), .ZN(n8072) );
  OAI21_X1 U9200 ( .B1(n8073), .B2(n10479), .A(n8072), .ZN(n8074) );
  AOI21_X1 U9201 ( .B1(n10555), .B2(n8289), .A(n8074), .ZN(n8292) );
  INV_X1 U9202 ( .A(n8075), .ZN(n8077) );
  INV_X1 U9203 ( .A(n8382), .ZN(n8076) );
  AOI21_X1 U9204 ( .B1(n9439), .B2(n8077), .A(n8076), .ZN(n8290) );
  NAND2_X1 U9205 ( .A1(n8290), .A2(n10526), .ZN(n8080) );
  AOI22_X1 U9206 ( .A1(n10502), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8078), .B2(
        n10491), .ZN(n8079) );
  OAI211_X1 U9207 ( .C1(n8081), .C2(n10530), .A(n8080), .B(n8079), .ZN(n8082)
         );
  AOI21_X1 U9208 ( .B1(n8289), .B2(n10527), .A(n8082), .ZN(n8083) );
  OAI21_X1 U9209 ( .B1(n8292), .B2(n10502), .A(n8083), .ZN(P1_U3280) );
  XNOR2_X1 U9210 ( .A(n8084), .B(n8086), .ZN(n10618) );
  INV_X1 U9211 ( .A(n10618), .ZN(n8097) );
  OAI211_X1 U9212 ( .C1(n8087), .C2(n8086), .A(n10453), .B(n8085), .ZN(n8089)
         );
  NAND2_X1 U9213 ( .A1(n8439), .A2(n10448), .ZN(n8088) );
  OAI211_X1 U9214 ( .C1(n8338), .C2(n9066), .A(n8089), .B(n8088), .ZN(n10616)
         );
  INV_X1 U9215 ( .A(n8093), .ZN(n10612) );
  INV_X1 U9216 ( .A(n8090), .ZN(n8126) );
  OAI21_X1 U9217 ( .B1(n10612), .B2(n8126), .A(n8305), .ZN(n10614) );
  OAI22_X1 U9218 ( .A1(n9164), .A2(n8091), .B1(n8103), .B2(n10470), .ZN(n8092)
         );
  AOI21_X1 U9219 ( .B1(n8093), .B2(n9153), .A(n8092), .ZN(n8094) );
  OAI21_X1 U9220 ( .B1(n10614), .B2(n9040), .A(n8094), .ZN(n8095) );
  AOI21_X1 U9221 ( .B1(n10616), .B2(n9164), .A(n8095), .ZN(n8096) );
  OAI21_X1 U9222 ( .B1(n8097), .B2(n10460), .A(n8096), .ZN(P2_U3282) );
  OAI21_X1 U9223 ( .B1(n8100), .B2(n8099), .A(n8098), .ZN(n8101) );
  NAND2_X1 U9224 ( .A1(n8101), .A2(n10375), .ZN(n8106) );
  NOR2_X1 U9225 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8102), .ZN(n8847) );
  OAI22_X1 U9226 ( .A1(n8782), .A2(n8338), .B1(n8780), .B2(n8103), .ZN(n8104)
         );
  AOI211_X1 U9227 ( .C1(n10373), .C2(n8439), .A(n8847), .B(n8104), .ZN(n8105)
         );
  OAI211_X1 U9228 ( .C1(n10612), .C2(n8743), .A(n8106), .B(n8105), .ZN(
        P2_U3217) );
  INV_X1 U9229 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8114) );
  INV_X1 U9230 ( .A(n8107), .ZN(n8108) );
  AOI21_X1 U9231 ( .B1(n10561), .B2(n8109), .A(n8108), .ZN(n8110) );
  OAI211_X1 U9232 ( .C1(n10162), .C2(n8112), .A(n8111), .B(n8110), .ZN(n8115)
         );
  NAND2_X1 U9233 ( .A1(n8115), .A2(n10595), .ZN(n8113) );
  OAI21_X1 U9234 ( .B1(n10595), .B2(n8114), .A(n8113), .ZN(P1_U3484) );
  NAND2_X1 U9235 ( .A1(n8115), .A2(n10591), .ZN(n8116) );
  OAI21_X1 U9236 ( .B1(n10591), .B2(n8117), .A(n8116), .ZN(P1_U3533) );
  INV_X1 U9237 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8131) );
  OAI21_X1 U9238 ( .B1(n8120), .B2(n8119), .A(n8118), .ZN(n8136) );
  XNOR2_X1 U9239 ( .A(n8121), .B(n8122), .ZN(n8125) );
  AOI222_X1 U9240 ( .A1(n10453), .A2(n8125), .B1(n8124), .B2(n10448), .C1(
        n8123), .C2(n10450), .ZN(n8141) );
  AOI21_X1 U9241 ( .B1(n8128), .B2(n8127), .A(n8126), .ZN(n8139) );
  AOI22_X1 U9242 ( .A1(n8139), .A2(n10404), .B1(n10403), .B2(n8128), .ZN(n8129) );
  OAI211_X1 U9243 ( .C1(n8136), .C2(n9245), .A(n8141), .B(n8129), .ZN(n9247)
         );
  NAND2_X1 U9244 ( .A1(n9247), .A2(n10624), .ZN(n8130) );
  OAI21_X1 U9245 ( .B1(n10624), .B2(n8131), .A(n8130), .ZN(P2_U3490) );
  INV_X1 U9246 ( .A(n8132), .ZN(n8133) );
  AOI22_X1 U9247 ( .A1(n10466), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8133), .B2(
        n9157), .ZN(n8134) );
  OAI21_X1 U9248 ( .B1(n8135), .B2(n10461), .A(n8134), .ZN(n8138) );
  NOR2_X1 U9249 ( .A1(n8136), .A2(n10460), .ZN(n8137) );
  AOI211_X1 U9250 ( .C1(n8139), .C2(n10465), .A(n8138), .B(n8137), .ZN(n8140)
         );
  OAI21_X1 U9251 ( .B1(n9079), .B2(n8141), .A(n8140), .ZN(P2_U3283) );
  NAND2_X1 U9252 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n8201), .ZN(n8142) );
  OAI21_X1 U9253 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n8201), .A(n8142), .ZN(
        n8154) );
  INV_X1 U9254 ( .A(n8167), .ZN(n10641) );
  NAND2_X1 U9255 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10638) );
  NAND2_X1 U9256 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n10641), .ZN(n8143) );
  OAI21_X1 U9257 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n10641), .A(n8143), .ZN(
        n10639) );
  NOR2_X1 U9258 ( .A1(n10638), .A2(n10639), .ZN(n10637) );
  NAND2_X1 U9259 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n10629), .ZN(n8144) );
  OAI21_X1 U9260 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10629), .A(n8144), .ZN(
        n10627) );
  NOR2_X1 U9261 ( .A1(n10626), .A2(n10627), .ZN(n10625) );
  AOI22_X1 U9262 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n8192), .B1(n8164), .B2(
        n6310), .ZN(n8185) );
  AOI21_X1 U9263 ( .B1(n8164), .B2(P2_REG2_REG_3__SCAN_IN), .A(n8183), .ZN(
        n8268) );
  NAND2_X1 U9264 ( .A1(n8162), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8145) );
  OAI21_X1 U9265 ( .B1(n8162), .B2(P2_REG2_REG_4__SCAN_IN), .A(n8145), .ZN(
        n8269) );
  NOR2_X1 U9266 ( .A1(n8268), .A2(n8269), .ZN(n8267) );
  NAND2_X1 U9267 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n8160), .ZN(n8146) );
  OAI21_X1 U9268 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n8160), .A(n8146), .ZN(
        n8230) );
  NOR2_X1 U9269 ( .A1(n8229), .A2(n8230), .ZN(n8228) );
  AOI21_X1 U9270 ( .B1(n8160), .B2(P2_REG2_REG_5__SCAN_IN), .A(n8228), .ZN(
        n8153) );
  NOR2_X1 U9271 ( .A1(n8153), .A2(n8154), .ZN(n8196) );
  NOR2_X1 U9272 ( .A1(n9275), .A2(P2_U3152), .ZN(n8147) );
  AOI21_X1 U9273 ( .B1(n8148), .B2(n8147), .A(n7056), .ZN(n8149) );
  OAI21_X1 U9274 ( .B1(n10242), .B2(n8150), .A(n8149), .ZN(n8151) );
  NAND2_X1 U9275 ( .A1(n8151), .A2(n6289), .ZN(n8175) );
  NOR2_X1 U9276 ( .A1(n9275), .A2(n6841), .ZN(n8152) );
  AOI211_X1 U9277 ( .C1(n8154), .C2(n8153), .A(n8196), .B(n10636), .ZN(n8182)
         );
  OAI21_X1 U9278 ( .B1(n10242), .B2(n8156), .A(n6289), .ZN(n8158) );
  NAND2_X1 U9279 ( .A1(n10242), .A2(n8330), .ZN(n8157) );
  NAND2_X1 U9280 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8555) );
  INV_X1 U9281 ( .A(n8555), .ZN(n8159) );
  AOI21_X1 U9282 ( .B1(n10655), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8159), .ZN(
        n8179) );
  NAND2_X1 U9283 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n8160), .ZN(n8172) );
  MUX2_X1 U9284 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n8161), .S(n8160), .Z(n8233)
         );
  NAND2_X1 U9285 ( .A1(n8162), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8171) );
  MUX2_X1 U9286 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n8163), .S(n8162), .Z(n8273)
         );
  MUX2_X1 U9287 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8165), .S(n8164), .Z(n8188)
         );
  NAND2_X1 U9288 ( .A1(P2_REG1_REG_2__SCAN_IN), .A2(n10629), .ZN(n8170) );
  MUX2_X1 U9289 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8166), .S(n10629), .Z(n10631) );
  NAND2_X1 U9290 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(n10641), .ZN(n8169) );
  MUX2_X1 U9291 ( .A(n8168), .B(P2_REG1_REG_1__SCAN_IN), .S(n8167), .Z(n10645)
         );
  NAND3_X1 U9292 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10645), .ZN(n10644) );
  NAND2_X1 U9293 ( .A1(n8169), .A2(n10644), .ZN(n10632) );
  NAND2_X1 U9294 ( .A1(n10631), .A2(n10632), .ZN(n10630) );
  NAND2_X1 U9295 ( .A1(n8170), .A2(n10630), .ZN(n8189) );
  NAND2_X1 U9296 ( .A1(n8188), .A2(n8189), .ZN(n8187) );
  OAI21_X1 U9297 ( .B1(n8192), .B2(n8165), .A(n8187), .ZN(n8272) );
  NAND2_X1 U9298 ( .A1(n8273), .A2(n8272), .ZN(n8271) );
  NAND2_X1 U9299 ( .A1(n8171), .A2(n8271), .ZN(n8234) );
  NAND2_X1 U9300 ( .A1(n8233), .A2(n8234), .ZN(n8232) );
  NAND2_X1 U9301 ( .A1(n8172), .A2(n8232), .ZN(n8177) );
  MUX2_X1 U9302 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8173), .S(n8201), .Z(n8176)
         );
  INV_X1 U9303 ( .A(n6841), .ZN(n8174) );
  NAND2_X1 U9304 ( .A1(n8176), .A2(n8177), .ZN(n8202) );
  OAI211_X1 U9305 ( .C1(n8177), .C2(n8176), .A(n10653), .B(n8202), .ZN(n8178)
         );
  OAI211_X1 U9306 ( .C1(n10650), .C2(n8180), .A(n8179), .B(n8178), .ZN(n8181)
         );
  OR2_X1 U9307 ( .A1(n8182), .A2(n8181), .ZN(P2_U3251) );
  AOI211_X1 U9308 ( .C1(n8185), .C2(n8184), .A(n8183), .B(n10636), .ZN(n8194)
         );
  NOR2_X1 U9309 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8186), .ZN(n8661) );
  AOI21_X1 U9310 ( .B1(n10655), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8661), .ZN(
        n8191) );
  OAI211_X1 U9311 ( .C1(n8189), .C2(n8188), .A(n10653), .B(n8187), .ZN(n8190)
         );
  OAI211_X1 U9312 ( .C1(n10650), .C2(n8192), .A(n8191), .B(n8190), .ZN(n8193)
         );
  OR2_X1 U9313 ( .A1(n8194), .A2(n8193), .ZN(P2_U3248) );
  NAND2_X1 U9314 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(n8213), .ZN(n8195) );
  OAI21_X1 U9315 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n8213), .A(n8195), .ZN(
        n8198) );
  NOR2_X1 U9316 ( .A1(n8197), .A2(n8198), .ZN(n8212) );
  AOI211_X1 U9317 ( .C1(n8198), .C2(n8197), .A(n8212), .B(n10636), .ZN(n8210)
         );
  NOR2_X1 U9318 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8199), .ZN(n8200) );
  AOI21_X1 U9319 ( .B1(n10655), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8200), .ZN(
        n8208) );
  NAND2_X1 U9320 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n8201), .ZN(n8203) );
  NAND2_X1 U9321 ( .A1(n8203), .A2(n8202), .ZN(n8206) );
  MUX2_X1 U9322 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8204), .S(n8213), .Z(n8205)
         );
  NAND2_X1 U9323 ( .A1(n8205), .A2(n8206), .ZN(n8219) );
  OAI211_X1 U9324 ( .C1(n8206), .C2(n8205), .A(n10653), .B(n8219), .ZN(n8207)
         );
  OAI211_X1 U9325 ( .C1(n10650), .C2(n8220), .A(n8208), .B(n8207), .ZN(n8209)
         );
  OR2_X1 U9326 ( .A1(n8210), .A2(n8209), .ZN(P2_U3252) );
  NAND2_X1 U9327 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n8242), .ZN(n8211) );
  OAI21_X1 U9328 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8242), .A(n8211), .ZN(
        n8215) );
  AOI21_X1 U9329 ( .B1(n8213), .B2(P2_REG2_REG_7__SCAN_IN), .A(n8212), .ZN(
        n8256) );
  AOI22_X1 U9330 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n8264), .B1(n8217), .B2(
        n6392), .ZN(n8257) );
  NOR2_X1 U9331 ( .A1(n8256), .A2(n8257), .ZN(n8255) );
  NOR2_X1 U9332 ( .A1(n8214), .A2(n8215), .ZN(n8241) );
  AOI211_X1 U9333 ( .C1(n8215), .C2(n8214), .A(n8241), .B(n10636), .ZN(n8227)
         );
  NAND2_X1 U9334 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8465) );
  INV_X1 U9335 ( .A(n8465), .ZN(n8216) );
  AOI21_X1 U9336 ( .B1(n10655), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8216), .ZN(
        n8225) );
  MUX2_X1 U9337 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8218), .S(n8217), .Z(n8260)
         );
  OAI21_X1 U9338 ( .B1(n8220), .B2(n8204), .A(n8219), .ZN(n8261) );
  NAND2_X1 U9339 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  OAI21_X1 U9340 ( .B1(n8264), .B2(n8218), .A(n8259), .ZN(n8223) );
  MUX2_X1 U9341 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8221), .S(n8242), .Z(n8222)
         );
  NAND2_X1 U9342 ( .A1(n8222), .A2(n8223), .ZN(n8246) );
  OAI211_X1 U9343 ( .C1(n8223), .C2(n8222), .A(n10653), .B(n8246), .ZN(n8224)
         );
  OAI211_X1 U9344 ( .C1(n10650), .C2(n8247), .A(n8225), .B(n8224), .ZN(n8226)
         );
  OR2_X1 U9345 ( .A1(n8227), .A2(n8226), .ZN(P2_U3254) );
  AOI211_X1 U9346 ( .C1(n8230), .C2(n8229), .A(n8228), .B(n10636), .ZN(n8239)
         );
  NOR2_X1 U9347 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8574), .ZN(n8231) );
  AOI21_X1 U9348 ( .B1(n10655), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8231), .ZN(
        n8236) );
  OAI211_X1 U9349 ( .C1(n8234), .C2(n8233), .A(n10653), .B(n8232), .ZN(n8235)
         );
  OAI211_X1 U9350 ( .C1(n10650), .C2(n8237), .A(n8236), .B(n8235), .ZN(n8238)
         );
  OR2_X1 U9351 ( .A1(n8239), .A2(n8238), .ZN(P2_U3250) );
  NAND2_X1 U9352 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8789), .ZN(n8240) );
  OAI21_X1 U9353 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8789), .A(n8240), .ZN(
        n8244) );
  AOI21_X1 U9354 ( .B1(n8242), .B2(P2_REG2_REG_9__SCAN_IN), .A(n8241), .ZN(
        n8243) );
  NOR2_X1 U9355 ( .A1(n8243), .A2(n8244), .ZN(n8788) );
  AOI211_X1 U9356 ( .C1(n8244), .C2(n8243), .A(n8788), .B(n10636), .ZN(n8254)
         );
  NOR2_X1 U9357 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6432), .ZN(n8245) );
  AOI21_X1 U9358 ( .B1(n10655), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8245), .ZN(
        n8252) );
  OAI21_X1 U9359 ( .B1(n8247), .B2(n8221), .A(n8246), .ZN(n8250) );
  MUX2_X1 U9360 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8248), .S(n8789), .Z(n8249)
         );
  NAND2_X1 U9361 ( .A1(n8249), .A2(n8250), .ZN(n8794) );
  OAI211_X1 U9362 ( .C1(n8250), .C2(n8249), .A(n10653), .B(n8794), .ZN(n8251)
         );
  OAI211_X1 U9363 ( .C1(n10650), .C2(n8795), .A(n8252), .B(n8251), .ZN(n8253)
         );
  OR2_X1 U9364 ( .A1(n8254), .A2(n8253), .ZN(P2_U3255) );
  AOI211_X1 U9365 ( .C1(n8257), .C2(n8256), .A(n8255), .B(n10636), .ZN(n8266)
         );
  NOR2_X1 U9366 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6393), .ZN(n8258) );
  AOI21_X1 U9367 ( .B1(n10655), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8258), .ZN(
        n8263) );
  OAI211_X1 U9368 ( .C1(n8261), .C2(n8260), .A(n10653), .B(n8259), .ZN(n8262)
         );
  OAI211_X1 U9369 ( .C1(n10650), .C2(n8264), .A(n8263), .B(n8262), .ZN(n8265)
         );
  OR2_X1 U9370 ( .A1(n8266), .A2(n8265), .ZN(P2_U3253) );
  AOI211_X1 U9371 ( .C1(n8269), .C2(n8268), .A(n8267), .B(n10636), .ZN(n8278)
         );
  AOI21_X1 U9372 ( .B1(n10655), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8270), .ZN(
        n8275) );
  OAI211_X1 U9373 ( .C1(n8273), .C2(n8272), .A(n10653), .B(n8271), .ZN(n8274)
         );
  OAI211_X1 U9374 ( .C1(n10650), .C2(n8276), .A(n8275), .B(n8274), .ZN(n8277)
         );
  OR2_X1 U9375 ( .A1(n8278), .A2(n8277), .ZN(P2_U3249) );
  XNOR2_X1 U9376 ( .A(n8280), .B(n8279), .ZN(n8281) );
  XNOR2_X1 U9377 ( .A(n8282), .B(n8281), .ZN(n8288) );
  INV_X1 U9378 ( .A(n9292), .ZN(n9673) );
  AOI21_X1 U9379 ( .B1(n9401), .B2(n9673), .A(n8283), .ZN(n8285) );
  NAND2_X1 U9380 ( .A1(n9402), .A2(n8383), .ZN(n8284) );
  OAI211_X1 U9381 ( .C1(n8379), .C2(n9405), .A(n8285), .B(n8284), .ZN(n8286)
         );
  AOI21_X1 U9382 ( .B1(n10159), .B2(n9408), .A(n8286), .ZN(n8287) );
  OAI21_X1 U9383 ( .B1(n8288), .B2(n9410), .A(n8287), .ZN(P1_U3222) );
  AOI22_X1 U9384 ( .A1(n8370), .A2(n10205), .B1(P2_U3966), .B2(n8975), .ZN(
        P2_U3578) );
  AOI22_X1 U9385 ( .A1(n8370), .A2(n8456), .B1(P2_U3966), .B2(n9015), .ZN(
        P2_U3577) );
  AOI22_X1 U9386 ( .A1(n8370), .A2(n10203), .B1(P2_U3966), .B2(n8765), .ZN(
        P2_U3579) );
  AOI22_X1 U9387 ( .A1(n8370), .A2(n8434), .B1(P2_U3966), .B2(n9033), .ZN(
        P2_U3576) );
  INV_X1 U9388 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8295) );
  INV_X1 U9389 ( .A(n8289), .ZN(n8293) );
  AOI22_X1 U9390 ( .A1(n8290), .A2(n10562), .B1(n10561), .B2(n9439), .ZN(n8291) );
  OAI211_X1 U9391 ( .C1(n8293), .C2(n10550), .A(n8292), .B(n8291), .ZN(n8296)
         );
  NAND2_X1 U9392 ( .A1(n8296), .A2(n10595), .ZN(n8294) );
  OAI21_X1 U9393 ( .B1(n10595), .B2(n8295), .A(n8294), .ZN(P1_U3487) );
  INV_X1 U9394 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U9395 ( .A1(n8296), .A2(n10591), .ZN(n8297) );
  OAI21_X1 U9396 ( .B1(n10591), .B2(n8298), .A(n8297), .ZN(P1_U3534) );
  XNOR2_X1 U9397 ( .A(n8300), .B(n8299), .ZN(n8301) );
  OAI222_X1 U9398 ( .A1(n9068), .A2(n8777), .B1(n9066), .B2(n8781), .C1(n9064), 
        .C2(n8301), .ZN(n8425) );
  INV_X1 U9399 ( .A(n8425), .ZN(n8312) );
  OAI21_X1 U9400 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8427) );
  INV_X1 U9401 ( .A(n8785), .ZN(n8423) );
  INV_X1 U9402 ( .A(n8305), .ZN(n8306) );
  OAI21_X1 U9403 ( .B1(n8423), .B2(n8306), .A(n8447), .ZN(n8424) );
  OAI22_X1 U9404 ( .A1(n9164), .A2(n8307), .B1(n8779), .B2(n10470), .ZN(n8308)
         );
  AOI21_X1 U9405 ( .B1(n8785), .B2(n9153), .A(n8308), .ZN(n8309) );
  OAI21_X1 U9406 ( .B1(n8424), .B2(n9040), .A(n8309), .ZN(n8310) );
  AOI21_X1 U9407 ( .B1(n8427), .B2(n9100), .A(n8310), .ZN(n8311) );
  OAI21_X1 U9408 ( .B1(n8312), .B2(n9079), .A(n8311), .ZN(P2_U3281) );
  NOR2_X1 U9409 ( .A1(n10655), .A2(P2_U3966), .ZN(P2_U3151) );
  CLKBUF_X3 U9410 ( .A(n8313), .Z(n8370) );
  AOI22_X1 U9411 ( .A1(n8370), .A2(n8314), .B1(P2_U3966), .B2(n6779), .ZN(
        P2_U3554) );
  INV_X1 U9412 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8316) );
  AOI22_X1 U9413 ( .A1(n8370), .A2(n8316), .B1(P2_U3966), .B2(n8315), .ZN(
        P2_U3561) );
  INV_X1 U9414 ( .A(n4868), .ZN(n8317) );
  AOI22_X1 U9415 ( .A1(n8370), .A2(n5493), .B1(P2_U3966), .B2(n8317), .ZN(
        P2_U3553) );
  AOI22_X1 U9416 ( .A1(n8370), .A2(n8319), .B1(P2_U3966), .B2(n8318), .ZN(
        P2_U3552) );
  AOI22_X1 U9417 ( .A1(n8370), .A2(n8321), .B1(P2_U3966), .B2(n8320), .ZN(
        P2_U3556) );
  AOI22_X1 U9418 ( .A1(n8370), .A2(n8323), .B1(P2_U3966), .B2(n8322), .ZN(
        P2_U3563) );
  AOI22_X1 U9419 ( .A1(n8370), .A2(n8324), .B1(P2_U3966), .B2(n8460), .ZN(
        P2_U3562) );
  AOI22_X1 U9420 ( .A1(n8370), .A2(n8325), .B1(P2_U3966), .B2(n8561), .ZN(
        P2_U3557) );
  INV_X1 U9421 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8327) );
  AOI22_X1 U9422 ( .A1(n8370), .A2(n8327), .B1(P2_U3966), .B2(n8326), .ZN(
        P2_U3564) );
  INV_X1 U9423 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8329) );
  AOI22_X1 U9424 ( .A1(n8370), .A2(n8329), .B1(P2_U3966), .B2(n8328), .ZN(
        P2_U3558) );
  NAND2_X1 U9425 ( .A1(n8333), .A2(n9265), .ZN(n8331) );
  OAI211_X1 U9426 ( .C1(n8332), .C2(n9280), .A(n8331), .B(n8330), .ZN(P2_U3335) );
  NAND2_X1 U9427 ( .A1(n8333), .A2(n10199), .ZN(n8335) );
  NAND2_X1 U9428 ( .A1(n8334), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9667) );
  OAI211_X1 U9429 ( .C1(n8336), .C2(n10204), .A(n8335), .B(n9667), .ZN(
        P1_U3330) );
  AOI22_X1 U9430 ( .A1(n8370), .A2(n8481), .B1(P2_U3966), .B2(n9069), .ZN(
        P2_U3574) );
  AOI22_X1 U9431 ( .A1(n8370), .A2(n8337), .B1(P2_U3966), .B2(n8709), .ZN(
        P2_U3567) );
  AOI22_X1 U9432 ( .A1(n8370), .A2(n8339), .B1(P2_U3966), .B2(n8338), .ZN(
        P2_U3565) );
  INV_X1 U9433 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8340) );
  AOI22_X1 U9434 ( .A1(n8370), .A2(n8340), .B1(P2_U3966), .B2(n8556), .ZN(
        P2_U3559) );
  AOI22_X1 U9435 ( .A1(n8370), .A2(n8341), .B1(P2_U3966), .B2(n8781), .ZN(
        P2_U3566) );
  AOI22_X1 U9436 ( .A1(n8370), .A2(n9495), .B1(P2_U3966), .B2(n8342), .ZN(
        P2_U3582) );
  INV_X1 U9437 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8343) );
  AOI22_X1 U9438 ( .A1(n8370), .A2(n8343), .B1(P2_U3966), .B2(n8718), .ZN(
        P2_U3570) );
  AOI22_X1 U9439 ( .A1(n8370), .A2(n8344), .B1(P2_U3966), .B2(n8752), .ZN(
        P2_U3573) );
  INV_X1 U9440 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8346) );
  AOI22_X1 U9441 ( .A1(n8370), .A2(n8346), .B1(P2_U3966), .B2(n8345), .ZN(
        P2_U3569) );
  INV_X1 U9442 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8347) );
  AOI22_X1 U9443 ( .A1(n8370), .A2(n8347), .B1(P2_U3966), .B2(n8777), .ZN(
        P2_U3568) );
  AOI22_X1 U9444 ( .A1(n8370), .A2(n8348), .B1(P2_U3966), .B2(n9067), .ZN(
        P2_U3572) );
  AND2_X1 U9445 ( .A1(n9439), .A2(n8379), .ZN(n9435) );
  OR2_X1 U9446 ( .A1(n9439), .A2(n8379), .ZN(n9563) );
  INV_X1 U9447 ( .A(n8357), .ZN(n8418) );
  OR2_X1 U9448 ( .A1(n10159), .A2(n8418), .ZN(n9564) );
  NAND2_X1 U9449 ( .A1(n10159), .A2(n8418), .ZN(n9566) );
  INV_X1 U9450 ( .A(n9522), .ZN(n8377) );
  NAND2_X1 U9451 ( .A1(n8409), .A2(n9292), .ZN(n9567) );
  XNOR2_X1 U9452 ( .A(n8402), .B(n8353), .ZN(n8360) );
  OR2_X1 U9453 ( .A1(n9439), .A2(n9674), .ZN(n8350) );
  NAND2_X1 U9454 ( .A1(n10159), .A2(n8357), .ZN(n8352) );
  INV_X1 U9455 ( .A(n8355), .ZN(n8354) );
  NAND2_X1 U9456 ( .A1(n8354), .A2(n8353), .ZN(n8395) );
  NAND2_X1 U9457 ( .A1(n8355), .A2(n9523), .ZN(n8356) );
  NAND2_X1 U9458 ( .A1(n8395), .A2(n8356), .ZN(n10149) );
  NAND2_X1 U9459 ( .A1(n10149), .A2(n10555), .ZN(n8359) );
  AOI22_X1 U9460 ( .A1(n8593), .A2(n10514), .B1(n10515), .B2(n8357), .ZN(n8358) );
  OAI211_X1 U9461 ( .C1(n10479), .C2(n8360), .A(n8359), .B(n8358), .ZN(n10156)
         );
  INV_X1 U9462 ( .A(n10156), .ZN(n8366) );
  AND2_X1 U9463 ( .A1(n8409), .A2(n8380), .ZN(n8361) );
  OR2_X1 U9464 ( .A1(n8361), .A2(n8398), .ZN(n10151) );
  AOI22_X1 U9465 ( .A1(n10502), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8420), .B2(
        n10491), .ZN(n8363) );
  NAND2_X1 U9466 ( .A1(n8409), .A2(n10045), .ZN(n8362) );
  OAI211_X1 U9467 ( .C1(n10151), .C2(n10430), .A(n8363), .B(n8362), .ZN(n8364)
         );
  AOI21_X1 U9468 ( .B1(n10149), .B2(n10527), .A(n8364), .ZN(n8365) );
  OAI21_X1 U9469 ( .B1(n8366), .B2(n10502), .A(n8365), .ZN(P1_U3278) );
  AOI22_X1 U9470 ( .A1(n8370), .A2(n8367), .B1(n8468), .B2(P2_U3966), .ZN(
        P2_U3560) );
  AOI22_X1 U9471 ( .A1(n8370), .A2(n10191), .B1(n8368), .B2(P2_U3966), .ZN(
        P2_U3581) );
  AOI22_X1 U9472 ( .A1(n8370), .A2(n8369), .B1(n8736), .B2(P2_U3966), .ZN(
        P2_U3571) );
  NAND2_X1 U9473 ( .A1(n8371), .A2(n9522), .ZN(n8372) );
  NAND2_X1 U9474 ( .A1(n8373), .A2(n8372), .ZN(n10161) );
  INV_X1 U9475 ( .A(n8374), .ZN(n8375) );
  AOI21_X1 U9476 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8378) );
  OAI222_X1 U9477 ( .A1(n10484), .A2(n9292), .B1(n10482), .B2(n8379), .C1(
        n10479), .C2(n8378), .ZN(n10157) );
  NAND2_X1 U9478 ( .A1(n10157), .A2(n10536), .ZN(n8388) );
  INV_X1 U9479 ( .A(n8380), .ZN(n8381) );
  AOI211_X1 U9480 ( .C1(n10159), .C2(n8382), .A(n10583), .B(n8381), .ZN(n10158) );
  INV_X1 U9481 ( .A(n10159), .ZN(n8385) );
  AOI22_X1 U9482 ( .A1(n10502), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8383), .B2(
        n10491), .ZN(n8384) );
  OAI21_X1 U9483 ( .B1(n8385), .B2(n10530), .A(n8384), .ZN(n8386) );
  AOI21_X1 U9484 ( .B1(n10158), .B2(n10003), .A(n8386), .ZN(n8387) );
  OAI211_X1 U9485 ( .C1(n10012), .C2(n10161), .A(n8388), .B(n8387), .ZN(
        P1_U3279) );
  OAI22_X1 U9486 ( .A1(n8370), .A2(n9057), .B1(P2_DATAO_REG_23__SCAN_IN), .B2(
        P2_U3966), .ZN(n8389) );
  INV_X1 U9487 ( .A(n8389), .ZN(P2_U3575) );
  OAI22_X1 U9488 ( .A1(n8370), .A2(n10451), .B1(P2_DATAO_REG_3__SCAN_IN), .B2(
        P2_U3966), .ZN(n8390) );
  INV_X1 U9489 ( .A(n8390), .ZN(P2_U3555) );
  OAI22_X1 U9490 ( .A1(n8370), .A2(n8932), .B1(P2_DATAO_REG_31__SCAN_IN), .B2(
        P2_U3966), .ZN(n8391) );
  INV_X1 U9491 ( .A(n8391), .ZN(P2_U3583) );
  OAI22_X1 U9492 ( .A1(n8370), .A2(n8392), .B1(P2_DATAO_REG_28__SCAN_IN), .B2(
        P2_U3966), .ZN(n8393) );
  INV_X1 U9493 ( .A(n8393), .ZN(P2_U3580) );
  OR2_X1 U9494 ( .A1(n8409), .A2(n9673), .ZN(n8394) );
  NAND2_X1 U9495 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  NAND2_X1 U9496 ( .A1(n10146), .A2(n10017), .ZN(n9547) );
  NAND2_X1 U9497 ( .A1(n9570), .A2(n9547), .ZN(n9525) );
  OAI21_X1 U9498 ( .B1(n8396), .B2(n9525), .A(n8595), .ZN(n8397) );
  INV_X1 U9499 ( .A(n8397), .ZN(n10148) );
  INV_X1 U9500 ( .A(n10146), .ZN(n9293) );
  INV_X1 U9501 ( .A(n10024), .ZN(n8399) );
  AOI211_X1 U9502 ( .C1(n10146), .C2(n5129), .A(n10583), .B(n8399), .ZN(n10145) );
  AOI22_X1 U9503 ( .A1(n10502), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9296), .B2(
        n10491), .ZN(n8400) );
  OAI21_X1 U9504 ( .B1(n9293), .B2(n10530), .A(n8400), .ZN(n8401) );
  AOI21_X1 U9505 ( .B1(n10145), .B2(n10003), .A(n8401), .ZN(n8408) );
  INV_X1 U9506 ( .A(n9567), .ZN(n9444) );
  INV_X1 U9507 ( .A(n9525), .ZN(n8404) );
  OAI211_X1 U9508 ( .C1(n8403), .C2(n8404), .A(n8584), .B(n10511), .ZN(n8406)
         );
  INV_X1 U9509 ( .A(n9996), .ZN(n9672) );
  AOI22_X1 U9510 ( .A1(n10515), .A2(n9673), .B1(n9672), .B2(n10514), .ZN(n8405) );
  NAND2_X1 U9511 ( .A1(n8406), .A2(n8405), .ZN(n10144) );
  NAND2_X1 U9512 ( .A1(n10144), .A2(n10536), .ZN(n8407) );
  OAI211_X1 U9513 ( .C1(n10148), .C2(n10012), .A(n8408), .B(n8407), .ZN(
        P1_U3277) );
  INV_X1 U9514 ( .A(n8409), .ZN(n10150) );
  NOR2_X1 U9515 ( .A1(n8410), .A2(n5031), .ZN(n8415) );
  AOI21_X1 U9516 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  OAI21_X1 U9517 ( .B1(n8415), .B2(n8414), .A(n9381), .ZN(n8422) );
  AOI21_X1 U9518 ( .B1(n9401), .B2(n8593), .A(n8416), .ZN(n8417) );
  OAI21_X1 U9519 ( .B1(n8418), .B2(n9405), .A(n8417), .ZN(n8419) );
  AOI21_X1 U9520 ( .B1(n8420), .B2(n9402), .A(n8419), .ZN(n8421) );
  OAI211_X1 U9521 ( .C1(n10150), .C2(n9388), .A(n8422), .B(n8421), .ZN(
        P1_U3232) );
  OAI22_X1 U9522 ( .A1(n8424), .A2(n10613), .B1(n8423), .B2(n10611), .ZN(n8426) );
  AOI211_X1 U9523 ( .C1(n10617), .C2(n8427), .A(n8426), .B(n8425), .ZN(n8429)
         );
  MUX2_X1 U9524 ( .A(n6514), .B(n8429), .S(n10620), .Z(n8428) );
  INV_X1 U9525 ( .A(n8428), .ZN(P2_U3535) );
  INV_X1 U9526 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8430) );
  MUX2_X1 U9527 ( .A(n8430), .B(n8429), .S(n10624), .Z(n8431) );
  INV_X1 U9528 ( .A(n8431), .ZN(P2_U3496) );
  OAI222_X1 U9529 ( .A1(P2_U3152), .A2(n8433), .B1(n8529), .B2(n8435), .C1(
        n8432), .C2(n9280), .ZN(P2_U3334) );
  OAI222_X1 U9530 ( .A1(n8436), .A2(P1_U3084), .B1(n10197), .B2(n8435), .C1(
        n8434), .C2(n10204), .ZN(P1_U3329) );
  XNOR2_X1 U9531 ( .A(n8437), .B(n8438), .ZN(n8440) );
  AOI222_X1 U9532 ( .A1(n10453), .A2(n8440), .B1(n9124), .B2(n10448), .C1(
        n8439), .C2(n10450), .ZN(n9244) );
  AOI21_X1 U9533 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8444) );
  INV_X1 U9534 ( .A(n8444), .ZN(n9246) );
  NAND2_X1 U9535 ( .A1(n10466), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8445) );
  OAI21_X1 U9536 ( .B1(n10470), .B2(n8708), .A(n8445), .ZN(n8446) );
  AOI21_X1 U9537 ( .B1(n9242), .B2(n9153), .A(n8446), .ZN(n8450) );
  AOI21_X1 U9538 ( .B1(n9242), .B2(n8447), .A(n10613), .ZN(n8448) );
  AND2_X1 U9539 ( .A1(n8448), .A2(n9143), .ZN(n9241) );
  NAND2_X1 U9540 ( .A1(n9241), .A2(n9145), .ZN(n8449) );
  OAI211_X1 U9541 ( .C1(n9246), .C2(n10460), .A(n8450), .B(n8449), .ZN(n8451)
         );
  INV_X1 U9542 ( .A(n8451), .ZN(n8452) );
  OAI21_X1 U9543 ( .B1(n9079), .B2(n9244), .A(n8452), .ZN(P2_U3280) );
  INV_X1 U9544 ( .A(n8453), .ZN(n8457) );
  INV_X1 U9545 ( .A(n10241), .ZN(n8454) );
  OAI222_X1 U9546 ( .A1(n9280), .A2(n8455), .B1(n8529), .B2(n8457), .C1(
        P2_U3152), .C2(n8454), .ZN(P2_U3333) );
  OAI222_X1 U9547 ( .A1(P1_U3084), .A2(n8458), .B1(n10197), .B2(n8457), .C1(
        n8456), .C2(n10204), .ZN(P1_U3328) );
  NAND2_X1 U9548 ( .A1(n10372), .A2(n8459), .ZN(n8467) );
  INV_X1 U9549 ( .A(n8460), .ZN(n8461) );
  NAND2_X1 U9550 ( .A1(n10373), .A2(n8461), .ZN(n8466) );
  INV_X1 U9551 ( .A(n8462), .ZN(n8463) );
  NAND2_X1 U9552 ( .A1(n8740), .A2(n8463), .ZN(n8464) );
  NAND4_X1 U9553 ( .A1(n8467), .A2(n8466), .A3(n8465), .A4(n8464), .ZN(n8475)
         );
  INV_X1 U9554 ( .A(n7587), .ZN(n8471) );
  NOR3_X1 U9555 ( .A1(n8761), .A2(n8469), .A3(n8468), .ZN(n8470) );
  AOI21_X1 U9556 ( .B1(n8471), .B2(n10375), .A(n8470), .ZN(n8473) );
  NOR2_X1 U9557 ( .A1(n8473), .A2(n8472), .ZN(n8474) );
  AOI211_X1 U9558 ( .C1(n8476), .C2(n6759), .A(n8475), .B(n8474), .ZN(n8477)
         );
  OAI21_X1 U9559 ( .B1(n8478), .B2(n8759), .A(n8477), .ZN(P2_U3233) );
  INV_X1 U9560 ( .A(n8479), .ZN(n8482) );
  OAI222_X1 U9561 ( .A1(n9280), .A2(n8480), .B1(n8529), .B2(n8482), .C1(n6259), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  OAI222_X1 U9562 ( .A1(n5480), .A2(P1_U3084), .B1(n10197), .B2(n8482), .C1(
        n8481), .C2(n10204), .ZN(P1_U3331) );
  NOR2_X1 U9563 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8523) );
  NOR2_X1 U9564 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8521) );
  NOR2_X1 U9565 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8519) );
  NOR2_X1 U9566 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8516) );
  NOR2_X1 U9567 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8514) );
  NOR2_X1 U9568 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8511) );
  NAND2_X1 U9569 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8508) );
  XOR2_X1 U9570 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10268) );
  NAND2_X1 U9571 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8506) );
  XOR2_X1 U9572 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10266) );
  NOR2_X1 U9573 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n8490) );
  XOR2_X1 U9574 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n8483), .Z(n10257) );
  NAND2_X1 U9575 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8488) );
  XOR2_X1 U9576 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10255) );
  NAND2_X1 U9577 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8486) );
  INV_X1 U9578 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8484) );
  XNOR2_X1 U9579 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n8484), .ZN(n10253) );
  AOI21_X1 U9580 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10247) );
  INV_X1 U9581 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10251) );
  NAND3_X1 U9582 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10249) );
  OAI21_X1 U9583 ( .B1(n10247), .B2(n10251), .A(n10249), .ZN(n10252) );
  NAND2_X1 U9584 ( .A1(n10253), .A2(n10252), .ZN(n8485) );
  NAND2_X1 U9585 ( .A1(n8486), .A2(n8485), .ZN(n10254) );
  NAND2_X1 U9586 ( .A1(n10255), .A2(n10254), .ZN(n8487) );
  NAND2_X1 U9587 ( .A1(n8488), .A2(n8487), .ZN(n10256) );
  NOR2_X1 U9588 ( .A1(n10257), .A2(n10256), .ZN(n8489) );
  NOR2_X1 U9589 ( .A1(n8490), .A2(n8489), .ZN(n8491) );
  NOR2_X1 U9590 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8491), .ZN(n10259) );
  AND2_X1 U9591 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8491), .ZN(n10258) );
  NOR2_X1 U9592 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10258), .ZN(n8492) );
  NAND2_X1 U9593 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8493), .ZN(n8495) );
  XOR2_X1 U9594 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8493), .Z(n10261) );
  NAND2_X1 U9595 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10261), .ZN(n8494) );
  NAND2_X1 U9596 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  NAND2_X1 U9597 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8496), .ZN(n8498) );
  XOR2_X1 U9598 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8496), .Z(n10262) );
  NAND2_X1 U9599 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10262), .ZN(n8497) );
  NAND2_X1 U9600 ( .A1(n8498), .A2(n8497), .ZN(n8499) );
  NAND2_X1 U9601 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8499), .ZN(n8501) );
  XOR2_X1 U9602 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8499), .Z(n10263) );
  NAND2_X1 U9603 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10263), .ZN(n8500) );
  NAND2_X1 U9604 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  NAND2_X1 U9605 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8502), .ZN(n8504) );
  XOR2_X1 U9606 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8502), .Z(n10264) );
  NAND2_X1 U9607 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10264), .ZN(n8503) );
  NAND2_X1 U9608 ( .A1(n8504), .A2(n8503), .ZN(n10265) );
  NAND2_X1 U9609 ( .A1(n10266), .A2(n10265), .ZN(n8505) );
  NAND2_X1 U9610 ( .A1(n8506), .A2(n8505), .ZN(n10267) );
  NAND2_X1 U9611 ( .A1(n10268), .A2(n10267), .ZN(n8507) );
  NAND2_X1 U9612 ( .A1(n8508), .A2(n8507), .ZN(n10270) );
  XOR2_X1 U9613 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n8509), .Z(n10269) );
  INV_X1 U9614 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8512) );
  XOR2_X1 U9615 ( .A(n8512), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10271) );
  XNOR2_X1 U9616 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10273) );
  XOR2_X1 U9617 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n8517), .Z(n10275) );
  NOR2_X1 U9618 ( .A1(n10276), .A2(n10275), .ZN(n8518) );
  NOR2_X1 U9619 ( .A1(n8519), .A2(n8518), .ZN(n10278) );
  INV_X1 U9620 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9725) );
  XOR2_X1 U9621 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n9725), .Z(n10277) );
  NOR2_X1 U9622 ( .A1(n10278), .A2(n10277), .ZN(n8520) );
  NOR2_X1 U9623 ( .A1(n8521), .A2(n8520), .ZN(n10280) );
  INV_X1 U9624 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9736) );
  XOR2_X1 U9625 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n9736), .Z(n10279) );
  NOR2_X1 U9626 ( .A1(n10280), .A2(n10279), .ZN(n8522) );
  NOR2_X1 U9627 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  AND2_X1 U9628 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8524), .ZN(n10281) );
  NOR2_X1 U9629 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10281), .ZN(n8525) );
  NOR2_X1 U9630 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8524), .ZN(n10282) );
  NOR2_X1 U9631 ( .A1(n8525), .A2(n10282), .ZN(n8527) );
  XNOR2_X1 U9632 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8526) );
  XNOR2_X1 U9633 ( .A(n8527), .B(n8526), .ZN(ADD_1071_U4) );
  INV_X1 U9634 ( .A(n9494), .ZN(n8583) );
  OAI222_X1 U9635 ( .A1(n8529), .A2(n8583), .B1(P2_U3152), .B2(n6252), .C1(
        n8528), .C2(n9280), .ZN(P2_U3328) );
  AOI22_X1 U9636 ( .A1(n9772), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10195), .ZN(n8530) );
  OAI21_X1 U9637 ( .B1(n8531), .B2(n10197), .A(n8530), .ZN(P1_U3335) );
  XNOR2_X1 U9638 ( .A(n8533), .B(n8532), .ZN(n8534) );
  XNOR2_X1 U9639 ( .A(n8535), .B(n8534), .ZN(n8540) );
  AND2_X1 U9640 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8912) );
  INV_X1 U9641 ( .A(n9119), .ZN(n8536) );
  OAI22_X1 U9642 ( .A1(n8778), .A2(n8736), .B1(n8780), .B2(n8536), .ZN(n8537)
         );
  AOI211_X1 U9643 ( .C1(n10372), .C2(n9124), .A(n8912), .B(n8537), .ZN(n8539)
         );
  NAND2_X1 U9644 ( .A1(n9231), .A2(n6759), .ZN(n8538) );
  OAI211_X1 U9645 ( .C1(n8540), .C2(n8759), .A(n8539), .B(n8538), .ZN(P2_U3240) );
  INV_X1 U9646 ( .A(n8541), .ZN(n8543) );
  NAND2_X1 U9647 ( .A1(n8543), .A2(n8542), .ZN(n8546) );
  AOI22_X1 U9648 ( .A1(n8547), .A2(n8546), .B1(n8544), .B2(n8545), .ZN(n8553)
         );
  INV_X1 U9649 ( .A(n10016), .ZN(n9671) );
  OAI21_X1 U9650 ( .B1(n9405), .B2(n10017), .A(n8548), .ZN(n8549) );
  AOI21_X1 U9651 ( .B1(n9401), .B2(n9671), .A(n8549), .ZN(n8550) );
  OAI21_X1 U9652 ( .B1(n9395), .B2(n10027), .A(n8550), .ZN(n8551) );
  AOI21_X1 U9653 ( .B1(n10139), .B2(n9408), .A(n8551), .ZN(n8552) );
  OAI21_X1 U9654 ( .B1(n8553), .B2(n9410), .A(n8552), .ZN(P1_U3239) );
  INV_X1 U9655 ( .A(n8554), .ZN(n8559) );
  OAI21_X1 U9656 ( .B1(n8743), .B2(n5227), .A(n8555), .ZN(n8558) );
  OAI22_X1 U9657 ( .A1(n8561), .A2(n8782), .B1(n8778), .B2(n8556), .ZN(n8557)
         );
  AOI211_X1 U9658 ( .C1(n8559), .C2(n8740), .A(n8558), .B(n8557), .ZN(n8567)
         );
  OAI22_X1 U9659 ( .A1(n8561), .A2(n8761), .B1(n8759), .B2(n8560), .ZN(n8565)
         );
  INV_X1 U9660 ( .A(n8562), .ZN(n8564) );
  NAND3_X1 U9661 ( .A1(n8565), .A2(n8564), .A3(n8563), .ZN(n8566) );
  OAI211_X1 U9662 ( .C1(n8759), .C2(n8568), .A(n8567), .B(n8566), .ZN(P2_U3241) );
  OAI222_X1 U9663 ( .A1(n8529), .A2(n8569), .B1(n9280), .B2(n6573), .C1(n6750), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U9664 ( .A1(n6759), .A2(n8570), .ZN(n8573) );
  NAND2_X1 U9665 ( .A1(n8766), .A2(n8571), .ZN(n8572) );
  OAI211_X1 U9666 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8579) );
  AOI22_X1 U9667 ( .A1(n8750), .A2(n8663), .B1(n10375), .B2(n8575), .ZN(n8577)
         );
  NOR3_X1 U9668 ( .A1(n8577), .A2(n4953), .A3(n8576), .ZN(n8578) );
  AOI211_X1 U9669 ( .C1(n8740), .C2(n8580), .A(n8579), .B(n8578), .ZN(n8581)
         );
  OAI21_X1 U9670 ( .B1(n8563), .B2(n8759), .A(n8581), .ZN(P2_U3229) );
  OAI222_X1 U9671 ( .A1(n10197), .A2(n8583), .B1(n8582), .B2(P1_U3084), .C1(
        n9495), .C2(n10204), .ZN(P1_U3323) );
  NAND2_X1 U9672 ( .A1(n8584), .A2(n9570), .ZN(n10020) );
  NAND2_X1 U9673 ( .A1(n10139), .A2(n9996), .ZN(n9548) );
  NAND2_X1 U9674 ( .A1(n10135), .A2(n10016), .ZN(n9545) );
  NAND2_X1 U9675 ( .A1(n9576), .A2(n9545), .ZN(n9991) );
  INV_X1 U9676 ( .A(n9991), .ZN(n9994) );
  NAND2_X1 U9677 ( .A1(n10128), .A2(n9999), .ZN(n9546) );
  NAND2_X1 U9678 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U9679 ( .A1(n9976), .A2(n9580), .ZN(n9960) );
  NAND2_X1 U9680 ( .A1(n10123), .A2(n9975), .ZN(n9582) );
  INV_X1 U9681 ( .A(n9954), .ZN(n9959) );
  NAND2_X1 U9682 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  INV_X1 U9683 ( .A(n9956), .ZN(n9373) );
  OR2_X1 U9684 ( .A1(n10117), .A2(n9373), .ZN(n9587) );
  NAND2_X1 U9685 ( .A1(n10117), .A2(n9373), .ZN(n9586) );
  NAND2_X1 U9686 ( .A1(n9587), .A2(n9586), .ZN(n9941) );
  INV_X1 U9687 ( .A(n9944), .ZN(n9325) );
  OR2_X1 U9688 ( .A1(n10112), .A2(n9325), .ZN(n9412) );
  NAND2_X1 U9689 ( .A1(n10112), .A2(n9325), .ZN(n9413) );
  INV_X1 U9690 ( .A(n9928), .ZN(n9384) );
  OR2_X1 U9691 ( .A1(n10108), .A2(n9384), .ZN(n9415) );
  NAND2_X1 U9692 ( .A1(n10108), .A2(n9384), .ZN(n9416) );
  NAND2_X1 U9693 ( .A1(n9415), .A2(n9416), .ZN(n9910) );
  INV_X1 U9694 ( .A(n9910), .ZN(n9915) );
  NAND2_X1 U9695 ( .A1(n9916), .A2(n9915), .ZN(n8586) );
  INV_X1 U9696 ( .A(n9879), .ZN(n9919) );
  OR2_X1 U9697 ( .A1(n10102), .A2(n9919), .ZN(n9592) );
  NAND2_X1 U9698 ( .A1(n10102), .A2(n9919), .ZN(n9641) );
  INV_X1 U9699 ( .A(n9897), .ZN(n9362) );
  OR2_X1 U9700 ( .A1(n10094), .A2(n9362), .ZN(n9470) );
  NAND2_X1 U9701 ( .A1(n10094), .A2(n9362), .ZN(n9594) );
  NAND2_X1 U9702 ( .A1(n9470), .A2(n9594), .ZN(n9881) );
  INV_X1 U9703 ( .A(n9881), .ZN(n9876) );
  XNOR2_X1 U9704 ( .A(n10090), .B(n9878), .ZN(n9868) );
  INV_X1 U9705 ( .A(n9878), .ZN(n9469) );
  NAND2_X1 U9706 ( .A1(n10090), .A2(n9469), .ZN(n9542) );
  INV_X1 U9707 ( .A(n9863), .ZN(n9406) );
  OR2_X1 U9708 ( .A1(n10084), .A2(n9406), .ZN(n9598) );
  NAND2_X1 U9709 ( .A1(n10084), .A2(n9406), .ZN(n9543) );
  OR2_X1 U9710 ( .A1(n10079), .A2(n9818), .ZN(n9599) );
  NAND2_X1 U9711 ( .A1(n10079), .A2(n9818), .ZN(n9537) );
  NAND2_X1 U9712 ( .A1(n9825), .A2(n9837), .ZN(n8587) );
  NAND2_X1 U9713 ( .A1(n8587), .A2(n9537), .ZN(n9816) );
  NAND2_X1 U9714 ( .A1(n10074), .A2(n8588), .ZN(n9539) );
  OR2_X1 U9715 ( .A1(n10066), .A2(n9817), .ZN(n9482) );
  NAND2_X1 U9716 ( .A1(n10066), .A2(n9817), .ZN(n9541) );
  INV_X1 U9717 ( .A(n9791), .ZN(n9796) );
  INV_X1 U9718 ( .A(n9541), .ZN(n8589) );
  NAND2_X1 U9719 ( .A1(n9271), .A2(n9493), .ZN(n8591) );
  OR2_X1 U9720 ( .A1(n5548), .A2(n10191), .ZN(n8590) );
  NAND2_X1 U9721 ( .A1(n10063), .A2(n8592), .ZN(n9649) );
  OR2_X1 U9722 ( .A1(n10146), .A2(n8593), .ZN(n8594) );
  NAND2_X1 U9723 ( .A1(n10139), .A2(n9672), .ZN(n9990) );
  NAND2_X1 U9724 ( .A1(n10135), .A2(n9671), .ZN(n8598) );
  AND2_X1 U9725 ( .A1(n9990), .A2(n8598), .ZN(n8597) );
  NAND2_X1 U9726 ( .A1(n10015), .A2(n8597), .ZN(n8601) );
  INV_X1 U9727 ( .A(n8598), .ZN(n8599) );
  OR2_X1 U9728 ( .A1(n8599), .A2(n9991), .ZN(n8600) );
  NAND2_X1 U9729 ( .A1(n8601), .A2(n8600), .ZN(n9974) );
  OR2_X1 U9730 ( .A1(n9957), .A2(n10128), .ZN(n8602) );
  INV_X1 U9731 ( .A(n9975), .ZN(n9943) );
  NAND2_X1 U9732 ( .A1(n10123), .A2(n9943), .ZN(n8603) );
  AND2_X1 U9733 ( .A1(n10117), .A2(n9956), .ZN(n8604) );
  NOR2_X1 U9734 ( .A1(n10112), .A2(n9944), .ZN(n8606) );
  NAND2_X1 U9735 ( .A1(n10112), .A2(n9944), .ZN(n8605) );
  AND2_X1 U9736 ( .A1(n10108), .A2(n9928), .ZN(n8607) );
  AOI21_X1 U9737 ( .B1(n9911), .B2(n9910), .A(n8607), .ZN(n9902) );
  NAND2_X1 U9738 ( .A1(n10102), .A2(n9879), .ZN(n8609) );
  NOR2_X1 U9739 ( .A1(n10102), .A2(n9879), .ZN(n8608) );
  AOI21_X1 U9740 ( .B1(n9902), .B2(n8609), .A(n8608), .ZN(n9882) );
  NAND2_X1 U9741 ( .A1(n9882), .A2(n9881), .ZN(n9850) );
  NAND2_X1 U9742 ( .A1(n10094), .A2(n9897), .ZN(n9866) );
  NAND2_X1 U9743 ( .A1(n10090), .A2(n9878), .ZN(n8610) );
  AND2_X1 U9744 ( .A1(n9866), .A2(n8610), .ZN(n9851) );
  INV_X1 U9745 ( .A(n9855), .ZN(n8611) );
  AND2_X1 U9746 ( .A1(n9851), .A2(n8611), .ZN(n8612) );
  NAND2_X1 U9747 ( .A1(n9850), .A2(n8612), .ZN(n8614) );
  OR2_X1 U9748 ( .A1(n10090), .A2(n9878), .ZN(n9852) );
  NAND2_X1 U9749 ( .A1(n10079), .A2(n9844), .ZN(n8616) );
  OR2_X1 U9750 ( .A1(n10074), .A2(n9826), .ZN(n8617) );
  XNOR2_X2 U9751 ( .A(n8621), .B(n8620), .ZN(n10065) );
  NAND2_X1 U9752 ( .A1(n6182), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U9753 ( .A1(n4876), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U9754 ( .A1(n4874), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8622) );
  AND3_X1 U9755 ( .A1(n8624), .A2(n8623), .A3(n8622), .ZN(n9508) );
  INV_X1 U9756 ( .A(n10295), .ZN(n8625) );
  NAND2_X1 U9757 ( .A1(n8625), .A2(P1_B_REG_SCAN_IN), .ZN(n8626) );
  NAND2_X1 U9758 ( .A1(n10514), .A2(n8626), .ZN(n9779) );
  OAI22_X1 U9759 ( .A1(n9817), .A2(n10482), .B1(n9508), .B2(n9779), .ZN(n8627)
         );
  OAI21_X1 U9760 ( .B1(n10065), .B2(n10519), .A(n8628), .ZN(n8629) );
  INV_X1 U9761 ( .A(n10079), .ZN(n9831) );
  INV_X1 U9762 ( .A(n10108), .ZN(n8631) );
  INV_X1 U9763 ( .A(n10123), .ZN(n9967) );
  NAND2_X1 U9764 ( .A1(n8631), .A2(n9930), .ZN(n9912) );
  NOR2_X2 U9765 ( .A1(n9912), .A2(n10102), .ZN(n9887) );
  OR2_X2 U9766 ( .A1(n10090), .A2(n9889), .ZN(n9859) );
  NOR2_X2 U9767 ( .A1(n10084), .A2(n9859), .ZN(n9846) );
  INV_X1 U9768 ( .A(n10063), .ZN(n8635) );
  AOI21_X1 U9769 ( .B1(n10063), .B2(n4902), .A(n9786), .ZN(n10064) );
  AOI22_X1 U9770 ( .A1(n10502), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8633), .B2(
        n10491), .ZN(n8634) );
  OAI21_X1 U9771 ( .B1(n8635), .B2(n10530), .A(n8634), .ZN(n8637) );
  NOR2_X1 U9772 ( .A1(n10065), .A2(n10431), .ZN(n8636) );
  AOI211_X1 U9773 ( .C1(n10064), .C2(n10526), .A(n8637), .B(n8636), .ZN(n8638)
         );
  OAI21_X1 U9774 ( .B1(n4933), .B2(n10502), .A(n8638), .ZN(P1_U3355) );
  INV_X1 U9775 ( .A(n8640), .ZN(n8641) );
  AOI21_X1 U9776 ( .B1(n8639), .B2(n8641), .A(n8759), .ZN(n8645) );
  NOR3_X1 U9777 ( .A1(n8642), .A2(n8975), .A3(n8761), .ZN(n8644) );
  OAI21_X1 U9778 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8650) );
  NOR2_X1 U9779 ( .A1(n8969), .A2(n8780), .ZN(n8648) );
  OAI22_X1 U9780 ( .A1(n8976), .A2(n8778), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8646), .ZN(n8647) );
  AOI211_X1 U9781 ( .C1(n10372), .C2(n8699), .A(n8648), .B(n8647), .ZN(n8649)
         );
  NAND2_X1 U9782 ( .A1(n8750), .A2(n9057), .ZN(n8654) );
  NAND2_X1 U9783 ( .A1(n8651), .A2(n10375), .ZN(n8653) );
  MUX2_X1 U9784 ( .A(n8654), .B(n8653), .S(n8652), .Z(n8659) );
  OAI22_X1 U9785 ( .A1(n8782), .A2(n9069), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8655), .ZN(n8657) );
  OAI22_X1 U9786 ( .A1(n8778), .A2(n9033), .B1(n8780), .B2(n9037), .ZN(n8656)
         );
  AOI211_X1 U9787 ( .C1(n9204), .C2(n6759), .A(n8657), .B(n8656), .ZN(n8658)
         );
  NAND2_X1 U9788 ( .A1(n8659), .A2(n8658), .ZN(P2_U3218) );
  NOR2_X1 U9789 ( .A1(n8780), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8660) );
  AOI211_X1 U9790 ( .C1(n10402), .C2(n6759), .A(n8661), .B(n8660), .ZN(n8672)
         );
  AOI22_X1 U9791 ( .A1(n10373), .A2(n8663), .B1(n10372), .B2(n8662), .ZN(n8671) );
  NOR3_X1 U9792 ( .A1(n8761), .A2(n8664), .A3(n6779), .ZN(n8669) );
  INV_X1 U9793 ( .A(n8666), .ZN(n8667) );
  AOI21_X1 U9794 ( .B1(n8665), .B2(n8667), .A(n8759), .ZN(n8668) );
  OAI21_X1 U9795 ( .B1(n8669), .B2(n8668), .A(n7510), .ZN(n8670) );
  NAND3_X1 U9796 ( .A1(n8672), .A2(n8671), .A3(n8670), .ZN(P2_U3220) );
  AOI21_X1 U9797 ( .B1(n8674), .B2(n8673), .A(n8759), .ZN(n8676) );
  NAND2_X1 U9798 ( .A1(n8676), .A2(n8675), .ZN(n8682) );
  INV_X1 U9799 ( .A(n9105), .ZN(n8680) );
  INV_X1 U9800 ( .A(n8718), .ZN(n8677) );
  AOI22_X1 U9801 ( .A1(n8678), .A2(n10448), .B1(n10450), .B2(n8677), .ZN(n9111) );
  NAND2_X1 U9802 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8926) );
  OAI21_X1 U9803 ( .B1(n8738), .B2(n9111), .A(n8926), .ZN(n8679) );
  AOI21_X1 U9804 ( .B1(n8680), .B2(n8740), .A(n8679), .ZN(n8681) );
  OAI211_X1 U9805 ( .C1(n9103), .C2(n8743), .A(n8682), .B(n8681), .ZN(P2_U3221) );
  INV_X1 U9806 ( .A(n8683), .ZN(n8685) );
  AOI21_X1 U9807 ( .B1(n8685), .B2(n8684), .A(n8759), .ZN(n8689) );
  NOR3_X1 U9808 ( .A1(n8686), .A2(n9067), .A3(n8761), .ZN(n8688) );
  OAI21_X1 U9809 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8694) );
  OAI22_X1 U9810 ( .A1(n8778), .A2(n9069), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8690), .ZN(n8692) );
  OAI22_X1 U9811 ( .A1(n8782), .A2(n9067), .B1(n8780), .B2(n9077), .ZN(n8691)
         );
  AOI211_X1 U9812 ( .C1(n9216), .C2(n6759), .A(n8692), .B(n8691), .ZN(n8693)
         );
  NAND2_X1 U9813 ( .A1(n8694), .A2(n8693), .ZN(P2_U3225) );
  OAI211_X1 U9814 ( .C1(n8697), .C2(n8696), .A(n8695), .B(n10375), .ZN(n8703)
         );
  NOR2_X1 U9815 ( .A1(n9033), .A2(n9066), .ZN(n8698) );
  AOI21_X1 U9816 ( .B1(n8699), .B2(n10448), .A(n8698), .ZN(n9003) );
  OAI22_X1 U9817 ( .A1(n9003), .A2(n8738), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8700), .ZN(n8701) );
  AOI21_X1 U9818 ( .B1(n9007), .B2(n8740), .A(n8701), .ZN(n8702) );
  OAI211_X1 U9819 ( .C1(n9010), .C2(n8743), .A(n8703), .B(n8702), .ZN(P2_U3227) );
  OAI21_X1 U9820 ( .B1(n8706), .B2(n8705), .A(n8704), .ZN(n8707) );
  NAND2_X1 U9821 ( .A1(n8707), .A2(n10375), .ZN(n8712) );
  AND2_X1 U9822 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8870) );
  OAI22_X1 U9823 ( .A1(n8782), .A2(n8709), .B1(n8780), .B2(n8708), .ZN(n8710)
         );
  AOI211_X1 U9824 ( .C1(n10373), .C2(n9124), .A(n8870), .B(n8710), .ZN(n8711)
         );
  OAI211_X1 U9825 ( .C1(n5229), .C2(n8743), .A(n8712), .B(n8711), .ZN(P2_U3228) );
  INV_X1 U9826 ( .A(n8713), .ZN(n8715) );
  NAND2_X1 U9827 ( .A1(n8715), .A2(n8714), .ZN(n8717) );
  XNOR2_X1 U9828 ( .A(n8717), .B(n8716), .ZN(n8722) );
  OAI22_X1 U9829 ( .A1(n8718), .A2(n9068), .B1(n8777), .B2(n9066), .ZN(n9134)
         );
  AOI22_X1 U9830 ( .A1(n8766), .A2(n9134), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8719) );
  OAI21_X1 U9831 ( .B1(n8780), .B2(n9141), .A(n8719), .ZN(n8720) );
  AOI21_X1 U9832 ( .B1(n9237), .B2(n6759), .A(n8720), .ZN(n8721) );
  OAI21_X1 U9833 ( .B1(n8722), .B2(n8759), .A(n8721), .ZN(P2_U3230) );
  AOI22_X1 U9834 ( .A1(n8723), .A2(n10375), .B1(n8750), .B2(n8724), .ZN(n8730)
         );
  INV_X1 U9835 ( .A(n8725), .ZN(n8729) );
  OAI22_X1 U9836 ( .A1(n9015), .A2(n8778), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7179), .ZN(n8727) );
  OAI22_X1 U9837 ( .A1(n8782), .A2(n9014), .B1(n8780), .B2(n9022), .ZN(n8726)
         );
  AOI211_X1 U9838 ( .C1(n9197), .C2(n6759), .A(n8727), .B(n8726), .ZN(n8728)
         );
  OAI21_X1 U9839 ( .B1(n8730), .B2(n8729), .A(n8728), .ZN(P2_U3231) );
  INV_X1 U9840 ( .A(n9222), .ZN(n9098) );
  INV_X1 U9841 ( .A(n8731), .ZN(n8732) );
  AOI21_X1 U9842 ( .B1(n8732), .B2(n8675), .A(n8759), .ZN(n8735) );
  NOR3_X1 U9843 ( .A1(n8733), .A2(n8736), .A3(n8761), .ZN(n8734) );
  OAI21_X1 U9844 ( .B1(n8735), .B2(n8734), .A(n8684), .ZN(n8742) );
  NOR2_X1 U9845 ( .A1(n8736), .A2(n9066), .ZN(n8737) );
  AOI21_X1 U9846 ( .B1(n9056), .B2(n10448), .A(n8737), .ZN(n9087) );
  OAI22_X1 U9847 ( .A1(n8738), .A2(n9087), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7270), .ZN(n8739) );
  AOI21_X1 U9848 ( .B1(n9095), .B2(n8740), .A(n8739), .ZN(n8741) );
  OAI211_X1 U9849 ( .C1(n9098), .C2(n8743), .A(n8742), .B(n8741), .ZN(P2_U3235) );
  INV_X1 U9850 ( .A(n8687), .ZN(n8746) );
  INV_X1 U9851 ( .A(n8744), .ZN(n8745) );
  AOI21_X1 U9852 ( .B1(n8746), .B2(n8751), .A(n8745), .ZN(n8757) );
  INV_X1 U9853 ( .A(n9050), .ZN(n8748) );
  AOI22_X1 U9854 ( .A1(n10373), .A2(n9057), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8747) );
  OAI21_X1 U9855 ( .B1(n8748), .B2(n8780), .A(n8747), .ZN(n8755) );
  NAND3_X1 U9856 ( .A1(n8751), .A2(n8750), .A3(n8749), .ZN(n8753) );
  AOI21_X1 U9857 ( .B1(n8753), .B2(n8782), .A(n8752), .ZN(n8754) );
  AOI211_X1 U9858 ( .C1(n9210), .C2(n6759), .A(n8755), .B(n8754), .ZN(n8756)
         );
  OAI21_X1 U9859 ( .B1(n8757), .B2(n8759), .A(n8756), .ZN(P2_U3237) );
  INV_X1 U9860 ( .A(n8758), .ZN(n8760) );
  AOI21_X1 U9861 ( .B1(n8695), .B2(n8760), .A(n8759), .ZN(n8764) );
  NOR3_X1 U9862 ( .A1(n8762), .A2(n9015), .A3(n8761), .ZN(n8763) );
  OAI21_X1 U9863 ( .B1(n8764), .B2(n8763), .A(n8639), .ZN(n8770) );
  OAI22_X1 U9864 ( .A1(n8765), .A2(n9068), .B1(n9015), .B2(n9066), .ZN(n8988)
         );
  AOI22_X1 U9865 ( .A1(n8988), .A2(n8766), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8767) );
  OAI21_X1 U9866 ( .B1(n8995), .B2(n8780), .A(n8767), .ZN(n8768) );
  AOI21_X1 U9867 ( .B1(n9187), .B2(n6759), .A(n8768), .ZN(n8769) );
  NAND2_X1 U9868 ( .A1(n8770), .A2(n8769), .ZN(P2_U3242) );
  OAI21_X1 U9869 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(n8774) );
  NAND2_X1 U9870 ( .A1(n8774), .A2(n10375), .ZN(n8787) );
  NOR2_X1 U9871 ( .A1(n8775), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8853) );
  INV_X1 U9872 ( .A(n8853), .ZN(n8776) );
  OAI21_X1 U9873 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8784) );
  OAI22_X1 U9874 ( .A1(n8782), .A2(n8781), .B1(n8780), .B2(n8779), .ZN(n8783)
         );
  AOI211_X1 U9875 ( .C1(n8785), .C2(n6759), .A(n8784), .B(n8783), .ZN(n8786)
         );
  NAND2_X1 U9876 ( .A1(n8787), .A2(n8786), .ZN(P2_U3243) );
  AOI22_X1 U9877 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n8813), .B1(n8805), .B2(
        n7875), .ZN(n8791) );
  NAND2_X1 U9878 ( .A1(n8790), .A2(n8791), .ZN(n8812) );
  OAI21_X1 U9879 ( .B1(n8791), .B2(n8790), .A(n8812), .ZN(n8802) );
  NOR2_X1 U9880 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8792), .ZN(n8793) );
  AOI21_X1 U9881 ( .B1(n10655), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8793), .ZN(
        n8800) );
  OAI21_X1 U9882 ( .B1(n8795), .B2(n8248), .A(n8794), .ZN(n8798) );
  MUX2_X1 U9883 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8796), .S(n8813), .Z(n8797)
         );
  NAND2_X1 U9884 ( .A1(n8797), .A2(n8798), .ZN(n8804) );
  OAI211_X1 U9885 ( .C1(n8798), .C2(n8797), .A(n10653), .B(n8804), .ZN(n8799)
         );
  OAI211_X1 U9886 ( .C1(n10650), .C2(n8805), .A(n8800), .B(n8799), .ZN(n8801)
         );
  AOI21_X1 U9887 ( .B1(n10654), .B2(n8802), .A(n8801), .ZN(n8803) );
  INV_X1 U9888 ( .A(n8803), .ZN(P2_U3256) );
  INV_X1 U9889 ( .A(n10650), .ZN(n10642) );
  OAI21_X1 U9890 ( .B1(n8805), .B2(n8796), .A(n8804), .ZN(n8808) );
  MUX2_X1 U9891 ( .A(n8806), .B(P2_REG1_REG_12__SCAN_IN), .S(n8820), .Z(n8807)
         );
  NOR2_X1 U9892 ( .A1(n8808), .A2(n8807), .ZN(n8825) );
  AOI21_X1 U9893 ( .B1(n8808), .B2(n8807), .A(n8825), .ZN(n8811) );
  AOI21_X1 U9894 ( .B1(n10655), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8809), .ZN(
        n8810) );
  OAI21_X1 U9895 ( .B1(n10651), .B2(n8811), .A(n8810), .ZN(n8817) );
  AOI22_X1 U9896 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8826), .B1(n8820), .B2(
        n7964), .ZN(n8815) );
  OAI21_X1 U9897 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8813), .A(n8812), .ZN(
        n8814) );
  NOR2_X1 U9898 ( .A1(n8814), .A2(n8815), .ZN(n8819) );
  AOI211_X1 U9899 ( .C1(n8815), .C2(n8814), .A(n8819), .B(n10636), .ZN(n8816)
         );
  AOI211_X1 U9900 ( .C1(n10642), .C2(n8820), .A(n8817), .B(n8816), .ZN(n8818)
         );
  INV_X1 U9901 ( .A(n8818), .ZN(P2_U3257) );
  NOR2_X1 U9902 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n8839), .ZN(n8821) );
  AOI21_X1 U9903 ( .B1(n8839), .B2(P2_REG2_REG_13__SCAN_IN), .A(n8821), .ZN(
        n8822) );
  NAND2_X1 U9904 ( .A1(n8823), .A2(n8822), .ZN(n8835) );
  OAI21_X1 U9905 ( .B1(n8823), .B2(n8822), .A(n8835), .ZN(n8824) );
  NAND2_X1 U9906 ( .A1(n10654), .A2(n8824), .ZN(n8833) );
  AOI21_X1 U9907 ( .B1(n8806), .B2(n8826), .A(n8825), .ZN(n8828) );
  AOI22_X1 U9908 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n8834), .B1(n8839), .B2(
        n6476), .ZN(n8827) );
  NOR2_X1 U9909 ( .A1(n8828), .A2(n8827), .ZN(n8841) );
  AOI21_X1 U9910 ( .B1(n8828), .B2(n8827), .A(n8841), .ZN(n8829) );
  NOR2_X1 U9911 ( .A1(n8829), .A2(n10651), .ZN(n8830) );
  AOI211_X1 U9912 ( .C1(n10655), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n8831), .B(
        n8830), .ZN(n8832) );
  OAI211_X1 U9913 ( .C1(n8834), .C2(n10650), .A(n8833), .B(n8832), .ZN(
        P2_U3258) );
  AOI22_X1 U9914 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8851), .B1(n8855), .B2(
        n8091), .ZN(n8836) );
  NAND2_X1 U9915 ( .A1(n8836), .A2(n8837), .ZN(n8850) );
  OAI21_X1 U9916 ( .B1(n8837), .B2(n8836), .A(n8850), .ZN(n8838) );
  NAND2_X1 U9917 ( .A1(n10654), .A2(n8838), .ZN(n8849) );
  NOR2_X1 U9918 ( .A1(n8839), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8840) );
  NOR2_X1 U9919 ( .A1(n8841), .A2(n8840), .ZN(n8844) );
  MUX2_X1 U9920 ( .A(n8842), .B(P2_REG1_REG_14__SCAN_IN), .S(n8851), .Z(n8843)
         );
  NOR2_X1 U9921 ( .A1(n8844), .A2(n8843), .ZN(n8854) );
  AOI21_X1 U9922 ( .B1(n8844), .B2(n8843), .A(n8854), .ZN(n8845) );
  NOR2_X1 U9923 ( .A1(n8845), .A2(n10651), .ZN(n8846) );
  AOI211_X1 U9924 ( .C1(n10655), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8847), .B(
        n8846), .ZN(n8848) );
  OAI211_X1 U9925 ( .C1(n10650), .C2(n8855), .A(n8849), .B(n8848), .ZN(
        P2_U3259) );
  OAI21_X1 U9926 ( .B1(n8852), .B2(n8307), .A(n8875), .ZN(n8860) );
  AOI21_X1 U9927 ( .B1(n10655), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8853), .ZN(
        n8858) );
  AOI21_X1 U9928 ( .B1(n8842), .B2(n8855), .A(n8854), .ZN(n8862) );
  XNOR2_X1 U9929 ( .A(n8874), .B(n8862), .ZN(n8856) );
  NAND2_X1 U9930 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8856), .ZN(n8864) );
  OAI211_X1 U9931 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n8856), .A(n10653), .B(
        n8864), .ZN(n8857) );
  OAI211_X1 U9932 ( .C1(n10650), .C2(n8874), .A(n8858), .B(n8857), .ZN(n8859)
         );
  AOI21_X1 U9933 ( .B1(n10654), .B2(n8860), .A(n8859), .ZN(n8861) );
  INV_X1 U9934 ( .A(n8861), .ZN(P2_U3260) );
  NAND2_X1 U9935 ( .A1(n8863), .A2(n8862), .ZN(n8865) );
  NAND2_X1 U9936 ( .A1(n8865), .A2(n8864), .ZN(n8869) );
  NOR2_X1 U9937 ( .A1(n8884), .A2(n8866), .ZN(n8867) );
  AOI21_X1 U9938 ( .B1(n8884), .B2(n8866), .A(n8867), .ZN(n8868) );
  NOR2_X1 U9939 ( .A1(n8869), .A2(n8868), .ZN(n8888) );
  AOI21_X1 U9940 ( .B1(n8869), .B2(n8868), .A(n8888), .ZN(n8872) );
  AOI21_X1 U9941 ( .B1(n10655), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8870), .ZN(
        n8871) );
  OAI21_X1 U9942 ( .B1(n8872), .B2(n10651), .A(n8871), .ZN(n8880) );
  AOI22_X1 U9943 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8889), .B1(n8884), .B2(
        n6254), .ZN(n8878) );
  NAND2_X1 U9944 ( .A1(n8874), .A2(n8873), .ZN(n8876) );
  NAND2_X1 U9945 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  NOR2_X1 U9946 ( .A1(n8877), .A2(n8878), .ZN(n8883) );
  AOI211_X1 U9947 ( .C1(n8878), .C2(n8877), .A(n8883), .B(n10636), .ZN(n8879)
         );
  AOI211_X1 U9948 ( .C1(n10642), .C2(n8884), .A(n8880), .B(n8879), .ZN(n8881)
         );
  INV_X1 U9949 ( .A(n8881), .ZN(P2_U3261) );
  INV_X1 U9950 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8882) );
  AOI22_X1 U9951 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8905), .B1(n8899), .B2(
        n8882), .ZN(n8886) );
  NOR2_X1 U9952 ( .A1(n8885), .A2(n8886), .ZN(n8898) );
  AOI211_X1 U9953 ( .C1(n8886), .C2(n8885), .A(n8898), .B(n10636), .ZN(n8895)
         );
  AND2_X1 U9954 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8887) );
  AOI21_X1 U9955 ( .B1(n10655), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8887), .ZN(
        n8893) );
  XNOR2_X1 U9956 ( .A(n8905), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8891) );
  AOI21_X1 U9957 ( .B1(n8889), .B2(n8866), .A(n8888), .ZN(n8890) );
  NAND2_X1 U9958 ( .A1(n8891), .A2(n8890), .ZN(n8903) );
  OAI211_X1 U9959 ( .C1(n8891), .C2(n8890), .A(n10653), .B(n8903), .ZN(n8892)
         );
  OAI211_X1 U9960 ( .C1(n10650), .C2(n8905), .A(n8893), .B(n8892), .ZN(n8894)
         );
  OR2_X1 U9961 ( .A1(n8895), .A2(n8894), .ZN(P2_U3262) );
  INV_X1 U9962 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8896) );
  NOR2_X1 U9963 ( .A1(n8915), .A2(n8896), .ZN(n8897) );
  AOI21_X1 U9964 ( .B1(n8896), .B2(n8915), .A(n8897), .ZN(n8901) );
  AOI21_X1 U9965 ( .B1(n8899), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8898), .ZN(
        n8900) );
  NAND2_X1 U9966 ( .A1(n8901), .A2(n8900), .ZN(n8916) );
  OAI21_X1 U9967 ( .B1(n8901), .B2(n8900), .A(n8916), .ZN(n8902) );
  NAND2_X1 U9968 ( .A1(n10654), .A2(n8902), .ZN(n8914) );
  INV_X1 U9969 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8904) );
  OAI21_X1 U9970 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8909) );
  INV_X1 U9971 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U9972 ( .A1(n8915), .A2(n8906), .ZN(n8920) );
  NAND2_X1 U9973 ( .A1(n8917), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U9974 ( .A1(n8920), .A2(n8907), .ZN(n8908) );
  NOR2_X1 U9975 ( .A1(n8908), .A2(n8909), .ZN(n8922) );
  AOI21_X1 U9976 ( .B1(n8909), .B2(n8908), .A(n8922), .ZN(n8910) );
  NOR2_X1 U9977 ( .A1(n10651), .A2(n8910), .ZN(n8911) );
  AOI211_X1 U9978 ( .C1(n10655), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8912), .B(
        n8911), .ZN(n8913) );
  OAI211_X1 U9979 ( .C1(n10650), .C2(n8915), .A(n8914), .B(n8913), .ZN(
        P2_U3263) );
  MUX2_X1 U9980 ( .A(n6564), .B(P2_REG2_REG_19__SCAN_IN), .S(n8993), .Z(n8919)
         );
  OAI21_X1 U9981 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8917), .A(n8916), .ZN(
        n8918) );
  XOR2_X1 U9982 ( .A(n8919), .B(n8918), .Z(n8930) );
  INV_X1 U9983 ( .A(n8920), .ZN(n8921) );
  NOR2_X1 U9984 ( .A1(n8922), .A2(n8921), .ZN(n8924) );
  XNOR2_X1 U9985 ( .A(n8993), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8923) );
  XNOR2_X1 U9986 ( .A(n8924), .B(n8923), .ZN(n8927) );
  NAND2_X1 U9987 ( .A1(n10655), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8925) );
  OAI211_X1 U9988 ( .C1(n10651), .C2(n8927), .A(n8926), .B(n8925), .ZN(n8928)
         );
  AOI21_X1 U9989 ( .B1(n10642), .B2(n9106), .A(n8928), .ZN(n8929) );
  OAI21_X1 U9990 ( .B1(n10636), .B2(n8930), .A(n8929), .ZN(P2_U3264) );
  NAND2_X1 U9991 ( .A1(n9175), .A2(n8935), .ZN(n9171) );
  NAND2_X1 U9992 ( .A1(n9169), .A2(n10465), .ZN(n8934) );
  NAND2_X1 U9993 ( .A1(n8932), .A2(n8931), .ZN(n9173) );
  NOR2_X1 U9994 ( .A1(n9079), .A2(n9173), .ZN(n8938) );
  AOI21_X1 U9995 ( .B1(n9079), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8938), .ZN(
        n8933) );
  OAI211_X1 U9996 ( .C1(n9170), .C2(n10461), .A(n8934), .B(n8933), .ZN(
        P2_U3265) );
  INV_X1 U9997 ( .A(n8935), .ZN(n8936) );
  NAND2_X1 U9998 ( .A1(n8937), .A2(n8936), .ZN(n9172) );
  NAND3_X1 U9999 ( .A1(n9172), .A2(n10465), .A3(n9171), .ZN(n8940) );
  AOI21_X1 U10000 ( .B1(n9079), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8938), .ZN(
        n8939) );
  OAI211_X1 U10001 ( .C1(n9175), .C2(n10461), .A(n8940), .B(n8939), .ZN(
        P2_U3266) );
  INV_X1 U10002 ( .A(n8941), .ZN(n8944) );
  AOI22_X1 U10003 ( .A1(n8942), .A2(n9157), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10466), .ZN(n8943) );
  OAI21_X1 U10004 ( .B1(n8944), .B2(n10461), .A(n8943), .ZN(n8945) );
  AOI21_X1 U10005 ( .B1(n8946), .B2(n10465), .A(n8945), .ZN(n8949) );
  OR2_X1 U10006 ( .A1(n8947), .A2(n10466), .ZN(n8948) );
  OAI211_X1 U10007 ( .C1(n8950), .C2(n10460), .A(n8949), .B(n8948), .ZN(
        P2_U3267) );
  OAI211_X1 U10008 ( .C1(n8953), .C2(n8952), .A(n8951), .B(n10453), .ZN(n8957)
         );
  AOI22_X1 U10009 ( .A1(n8955), .A2(n10448), .B1(n8954), .B2(n10450), .ZN(
        n8956) );
  XNOR2_X1 U10010 ( .A(n8959), .B(n8958), .ZN(n9180) );
  INV_X1 U10011 ( .A(n9180), .ZN(n8966) );
  OR2_X1 U10012 ( .A1(n6761), .A2(n4903), .ZN(n8960) );
  AND2_X1 U10013 ( .A1(n8961), .A2(n8960), .ZN(n9177) );
  NAND2_X1 U10014 ( .A1(n9177), .A2(n10465), .ZN(n8964) );
  AOI22_X1 U10015 ( .A1(n8962), .A2(n9157), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10466), .ZN(n8963) );
  OAI211_X1 U10016 ( .C1(n6761), .C2(n10461), .A(n8964), .B(n8963), .ZN(n8965)
         );
  AOI21_X1 U10017 ( .B1(n8966), .B2(n9100), .A(n8965), .ZN(n8967) );
  OAI21_X1 U10018 ( .B1(n9179), .B2(n9079), .A(n8967), .ZN(P2_U3268) );
  XOR2_X1 U10019 ( .A(n8973), .B(n8968), .Z(n9185) );
  AOI21_X1 U10020 ( .B1(n9181), .B2(n8991), .A(n4903), .ZN(n9182) );
  INV_X1 U10021 ( .A(n8969), .ZN(n8970) );
  AOI22_X1 U10022 ( .A1(n8970), .A2(n9157), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10466), .ZN(n8971) );
  OAI21_X1 U10023 ( .B1(n8972), .B2(n10461), .A(n8971), .ZN(n8981) );
  AOI21_X1 U10024 ( .B1(n8974), .B2(n8973), .A(n9064), .ZN(n8979) );
  OAI22_X1 U10025 ( .A1(n8976), .A2(n9068), .B1(n8975), .B2(n9066), .ZN(n8977)
         );
  AOI21_X1 U10026 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n9184) );
  NOR2_X1 U10027 ( .A1(n9184), .A2(n9079), .ZN(n8980) );
  AOI211_X1 U10028 ( .C1(n9182), .C2(n10465), .A(n8981), .B(n8980), .ZN(n8982)
         );
  OAI21_X1 U10029 ( .B1(n9185), .B2(n10460), .A(n8982), .ZN(P2_U3269) );
  XNOR2_X1 U10030 ( .A(n8984), .B(n8983), .ZN(n9190) );
  AOI22_X1 U10031 ( .A1(n9187), .A2(n9153), .B1(n10466), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8998) );
  OAI21_X1 U10032 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(n8989) );
  AOI21_X1 U10033 ( .B1(n8989), .B2(n10453), .A(n8988), .ZN(n9189) );
  INV_X1 U10034 ( .A(n8991), .ZN(n8992) );
  AOI211_X1 U10035 ( .C1(n9187), .C2(n9005), .A(n10613), .B(n8992), .ZN(n9186)
         );
  NAND2_X1 U10036 ( .A1(n9186), .A2(n8993), .ZN(n8994) );
  OAI211_X1 U10037 ( .C1(n10470), .C2(n8995), .A(n9189), .B(n8994), .ZN(n8996)
         );
  NAND2_X1 U10038 ( .A1(n8996), .A2(n9164), .ZN(n8997) );
  OAI211_X1 U10039 ( .C1(n9190), .C2(n10460), .A(n8998), .B(n8997), .ZN(
        P2_U3270) );
  XNOR2_X1 U10040 ( .A(n8999), .B(n9001), .ZN(n9195) );
  OAI211_X1 U10041 ( .C1(n9002), .C2(n9001), .A(n9000), .B(n10453), .ZN(n9004)
         );
  NAND2_X1 U10042 ( .A1(n9004), .A2(n9003), .ZN(n9192) );
  AOI211_X1 U10043 ( .C1(n9193), .C2(n9006), .A(n10613), .B(n8990), .ZN(n9191)
         );
  NAND2_X1 U10044 ( .A1(n9191), .A2(n9145), .ZN(n9009) );
  AOI22_X1 U10045 ( .A1(n9007), .A2(n9157), .B1(n10466), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9008) );
  OAI211_X1 U10046 ( .C1(n9010), .C2(n10461), .A(n9009), .B(n9008), .ZN(n9011)
         );
  AOI21_X1 U10047 ( .B1(n9164), .B2(n9192), .A(n9011), .ZN(n9012) );
  OAI21_X1 U10048 ( .B1(n9195), .B2(n10460), .A(n9012), .ZN(P2_U3271) );
  AOI21_X1 U10049 ( .B1(n9013), .B2(n9020), .A(n9064), .ZN(n9018) );
  OAI22_X1 U10050 ( .A1(n9015), .A2(n9068), .B1(n9014), .B2(n9066), .ZN(n9016)
         );
  AOI21_X1 U10051 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9200) );
  OAI21_X1 U10052 ( .B1(n9021), .B2(n9020), .A(n9019), .ZN(n9196) );
  XNOR2_X1 U10053 ( .A(n9197), .B(n9034), .ZN(n9198) );
  NAND2_X1 U10054 ( .A1(n9198), .A2(n10465), .ZN(n9025) );
  INV_X1 U10055 ( .A(n9022), .ZN(n9023) );
  AOI22_X1 U10056 ( .A1(n9023), .A2(n9157), .B1(n10466), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n9024) );
  OAI211_X1 U10057 ( .C1(n9026), .C2(n10461), .A(n9025), .B(n9024), .ZN(n9027)
         );
  AOI21_X1 U10058 ( .B1(n9196), .B2(n9100), .A(n9027), .ZN(n9028) );
  OAI21_X1 U10059 ( .B1(n9079), .B2(n9200), .A(n9028), .ZN(P2_U3272) );
  INV_X1 U10060 ( .A(n9029), .ZN(n9030) );
  AOI21_X1 U10061 ( .B1(n9041), .B2(n9031), .A(n9030), .ZN(n9032) );
  OAI222_X1 U10062 ( .A1(n9066), .A2(n9069), .B1(n9068), .B2(n9033), .C1(n9064), .C2(n9032), .ZN(n9208) );
  AND2_X1 U10063 ( .A1(n9204), .A2(n9048), .ZN(n9035) );
  OR2_X1 U10064 ( .A1(n9035), .A2(n9034), .ZN(n9206) );
  NAND2_X1 U10065 ( .A1(n10466), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9036) );
  OAI21_X1 U10066 ( .B1(n10470), .B2(n9037), .A(n9036), .ZN(n9038) );
  AOI21_X1 U10067 ( .B1(n9204), .B2(n9153), .A(n9038), .ZN(n9039) );
  OAI21_X1 U10068 ( .B1(n9206), .B2(n9040), .A(n9039), .ZN(n9044) );
  NOR2_X1 U10069 ( .A1(n9042), .A2(n9041), .ZN(n9203) );
  NOR3_X1 U10070 ( .A1(n9203), .A2(n9202), .A3(n10460), .ZN(n9043) );
  AOI211_X1 U10071 ( .C1(n9164), .C2(n9208), .A(n9044), .B(n9043), .ZN(n9045)
         );
  INV_X1 U10072 ( .A(n9045), .ZN(P2_U3273) );
  XNOR2_X1 U10073 ( .A(n9046), .B(n9055), .ZN(n9214) );
  INV_X1 U10074 ( .A(n9048), .ZN(n9049) );
  AOI21_X1 U10075 ( .B1(n9210), .B2(n9076), .A(n9049), .ZN(n9211) );
  AOI22_X1 U10076 ( .A1(n10466), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9050), 
        .B2(n9157), .ZN(n9051) );
  OAI21_X1 U10077 ( .B1(n9052), .B2(n10461), .A(n9051), .ZN(n9061) );
  OAI211_X1 U10078 ( .C1(n9055), .C2(n9054), .A(n10453), .B(n9053), .ZN(n9059)
         );
  AOI22_X1 U10079 ( .A1(n9057), .A2(n10448), .B1(n10450), .B2(n9056), .ZN(
        n9058) );
  NOR2_X1 U10080 ( .A1(n9213), .A2(n9079), .ZN(n9060) );
  AOI211_X1 U10081 ( .C1(n9211), .C2(n10465), .A(n9061), .B(n9060), .ZN(n9062)
         );
  OAI21_X1 U10082 ( .B1(n9214), .B2(n10460), .A(n9062), .ZN(P2_U3274) );
  INV_X1 U10083 ( .A(n9063), .ZN(n9065) );
  AOI21_X1 U10084 ( .B1(n9065), .B2(n9074), .A(n9064), .ZN(n9072) );
  OAI22_X1 U10085 ( .A1(n9069), .A2(n9068), .B1(n9067), .B2(n9066), .ZN(n9070)
         );
  AOI21_X1 U10086 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n9219) );
  OAI21_X1 U10087 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9215) );
  INV_X1 U10088 ( .A(n9216), .ZN(n9082) );
  AOI21_X1 U10089 ( .B1(n9216), .B2(n9092), .A(n9047), .ZN(n9217) );
  NAND2_X1 U10090 ( .A1(n9217), .A2(n10465), .ZN(n9081) );
  INV_X1 U10091 ( .A(n9077), .ZN(n9078) );
  AOI22_X1 U10092 ( .A1(n9079), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9078), .B2(
        n9157), .ZN(n9080) );
  OAI211_X1 U10093 ( .C1(n9082), .C2(n10461), .A(n9081), .B(n9080), .ZN(n9083)
         );
  AOI21_X1 U10094 ( .B1(n9215), .B2(n9100), .A(n9083), .ZN(n9084) );
  OAI21_X1 U10095 ( .B1(n9079), .B2(n9219), .A(n9084), .ZN(P2_U3275) );
  OAI211_X1 U10096 ( .C1(n9091), .C2(n9086), .A(n9085), .B(n10453), .ZN(n9088)
         );
  AOI21_X1 U10097 ( .B1(n9091), .B2(n9090), .A(n9089), .ZN(n9221) );
  INV_X1 U10098 ( .A(n9092), .ZN(n9093) );
  AOI21_X1 U10099 ( .B1(n9222), .B2(n9094), .A(n9093), .ZN(n9223) );
  NAND2_X1 U10100 ( .A1(n9223), .A2(n10465), .ZN(n9097) );
  AOI22_X1 U10101 ( .A1(n10466), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9095), 
        .B2(n9157), .ZN(n9096) );
  OAI211_X1 U10102 ( .C1(n9098), .C2(n10461), .A(n9097), .B(n9096), .ZN(n9099)
         );
  AOI21_X1 U10103 ( .B1(n9221), .B2(n9100), .A(n9099), .ZN(n9101) );
  OAI21_X1 U10104 ( .B1(n9079), .B2(n9225), .A(n9101), .ZN(P2_U3276) );
  XOR2_X1 U10105 ( .A(n9102), .B(n9110), .Z(n9230) );
  AOI22_X1 U10106 ( .A1(n6797), .A2(n9153), .B1(n10466), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n9115) );
  XNOR2_X1 U10107 ( .A(n9103), .B(n9118), .ZN(n9104) );
  NOR2_X1 U10108 ( .A1(n9104), .A2(n10613), .ZN(n9228) );
  INV_X1 U10109 ( .A(n9228), .ZN(n9107) );
  OAI22_X1 U10110 ( .A1(n9107), .A2(n9106), .B1(n10470), .B2(n9105), .ZN(n9113) );
  OAI211_X1 U10111 ( .C1(n9110), .C2(n9109), .A(n9108), .B(n10453), .ZN(n9112)
         );
  NAND2_X1 U10112 ( .A1(n9112), .A2(n9111), .ZN(n9227) );
  OAI21_X1 U10113 ( .B1(n9113), .B2(n9227), .A(n9164), .ZN(n9114) );
  OAI211_X1 U10114 ( .C1(n9230), .C2(n10460), .A(n9115), .B(n9114), .ZN(
        P2_U3277) );
  XNOR2_X1 U10115 ( .A(n9117), .B(n6831), .ZN(n9235) );
  AOI21_X1 U10116 ( .B1(n9231), .B2(n4899), .A(n9118), .ZN(n9232) );
  AOI22_X1 U10117 ( .A1(n10466), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9119), 
        .B2(n9157), .ZN(n9120) );
  OAI21_X1 U10118 ( .B1(n9121), .B2(n10461), .A(n9120), .ZN(n9129) );
  OAI211_X1 U10119 ( .C1(n6831), .C2(n9122), .A(n9123), .B(n10453), .ZN(n9127)
         );
  AOI22_X1 U10120 ( .A1(n9125), .A2(n10448), .B1(n10450), .B2(n9124), .ZN(
        n9126) );
  NOR2_X1 U10121 ( .A1(n9234), .A2(n10466), .ZN(n9128) );
  AOI211_X1 U10122 ( .C1(n9232), .C2(n10465), .A(n9129), .B(n9128), .ZN(n9130)
         );
  OAI21_X1 U10123 ( .B1(n9235), .B2(n10460), .A(n9130), .ZN(P2_U3278) );
  INV_X1 U10124 ( .A(n9131), .ZN(n9132) );
  XNOR2_X1 U10125 ( .A(n9133), .B(n9132), .ZN(n9135) );
  AOI21_X1 U10126 ( .B1(n9135), .B2(n10453), .A(n9134), .ZN(n9239) );
  OAI21_X1 U10127 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9139) );
  INV_X1 U10128 ( .A(n9139), .ZN(n9240) );
  NAND2_X1 U10129 ( .A1(n10466), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9140) );
  OAI21_X1 U10130 ( .B1(n10470), .B2(n9141), .A(n9140), .ZN(n9142) );
  AOI21_X1 U10131 ( .B1(n9237), .B2(n9153), .A(n9142), .ZN(n9147) );
  AOI21_X1 U10132 ( .B1(n9237), .B2(n9143), .A(n10613), .ZN(n9144) );
  AND2_X1 U10133 ( .A1(n9144), .A2(n4899), .ZN(n9236) );
  NAND2_X1 U10134 ( .A1(n9236), .A2(n9145), .ZN(n9146) );
  OAI211_X1 U10135 ( .C1(n9240), .C2(n10460), .A(n9147), .B(n9146), .ZN(n9148)
         );
  INV_X1 U10136 ( .A(n9148), .ZN(n9149) );
  OAI21_X1 U10137 ( .B1(n9079), .B2(n9239), .A(n9149), .ZN(P2_U3279) );
  INV_X1 U10138 ( .A(n9150), .ZN(n9152) );
  XNOR2_X1 U10139 ( .A(n9151), .B(n9159), .ZN(n10390) );
  AOI22_X1 U10140 ( .A1(n9153), .A2(n10374), .B1(n9152), .B2(n10390), .ZN(
        n9168) );
  INV_X1 U10141 ( .A(n9154), .ZN(n9155) );
  AOI21_X1 U10142 ( .B1(n10374), .B2(n9156), .A(n9155), .ZN(n10385) );
  AOI22_X1 U10143 ( .A1(n10465), .A2(n10385), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n9157), .ZN(n9167) );
  NAND2_X1 U10144 ( .A1(n10466), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9166) );
  NAND2_X1 U10145 ( .A1(n10390), .A2(n9160), .ZN(n9162) );
  AOI22_X1 U10146 ( .A1(n10448), .A2(n10451), .B1(n4868), .B2(n10450), .ZN(
        n9161) );
  NAND3_X1 U10147 ( .A1(n9163), .A2(n9162), .A3(n9161), .ZN(n10388) );
  NAND2_X1 U10148 ( .A1(n9164), .A2(n10388), .ZN(n9165) );
  NAND4_X1 U10149 ( .A1(n9168), .A2(n9167), .A3(n9166), .A4(n9165), .ZN(
        P2_U3294) );
  NAND3_X1 U10150 ( .A1(n9172), .A2(n10404), .A3(n9171), .ZN(n9174) );
  OAI211_X1 U10151 ( .C1(n9175), .C2(n10611), .A(n9174), .B(n9173), .ZN(n9251)
         );
  MUX2_X1 U10152 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9251), .S(n10620), .Z(
        P2_U3550) );
  AOI22_X1 U10153 ( .A1(n9177), .A2(n10404), .B1(n10403), .B2(n9176), .ZN(
        n9178) );
  OAI211_X1 U10154 ( .C1(n9180), .C2(n9245), .A(n9179), .B(n9178), .ZN(n9252)
         );
  MUX2_X1 U10155 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9252), .S(n10620), .Z(
        P2_U3548) );
  AOI22_X1 U10156 ( .A1(n9182), .A2(n10404), .B1(n10403), .B2(n9181), .ZN(
        n9183) );
  OAI211_X1 U10157 ( .C1(n9185), .C2(n9245), .A(n9184), .B(n9183), .ZN(n9253)
         );
  MUX2_X1 U10158 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9253), .S(n10620), .Z(
        P2_U3547) );
  AOI21_X1 U10159 ( .B1(n10403), .B2(n9187), .A(n9186), .ZN(n9188) );
  OAI211_X1 U10160 ( .C1(n9190), .C2(n9245), .A(n9189), .B(n9188), .ZN(n9254)
         );
  MUX2_X1 U10161 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9254), .S(n10620), .Z(
        P2_U3546) );
  AOI211_X1 U10162 ( .C1(n10403), .C2(n9193), .A(n9192), .B(n9191), .ZN(n9194)
         );
  OAI21_X1 U10163 ( .B1(n9195), .B2(n9245), .A(n9194), .ZN(n9255) );
  MUX2_X1 U10164 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9255), .S(n10620), .Z(
        P2_U3545) );
  INV_X1 U10165 ( .A(n9196), .ZN(n9201) );
  AOI22_X1 U10166 ( .A1(n9198), .A2(n10404), .B1(n10403), .B2(n9197), .ZN(
        n9199) );
  OAI211_X1 U10167 ( .C1(n9201), .C2(n9245), .A(n9200), .B(n9199), .ZN(n9256)
         );
  MUX2_X1 U10168 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9256), .S(n10620), .Z(
        P2_U3544) );
  NOR3_X1 U10169 ( .A1(n9203), .A2(n9202), .A3(n9245), .ZN(n9209) );
  INV_X1 U10170 ( .A(n9204), .ZN(n9205) );
  OAI22_X1 U10171 ( .A1(n9206), .A2(n10613), .B1(n9205), .B2(n10611), .ZN(
        n9207) );
  MUX2_X1 U10172 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9257), .S(n10620), .Z(
        P2_U3543) );
  AOI22_X1 U10173 ( .A1(n9211), .A2(n10404), .B1(n10403), .B2(n9210), .ZN(
        n9212) );
  OAI211_X1 U10174 ( .C1(n9214), .C2(n9245), .A(n9213), .B(n9212), .ZN(n9258)
         );
  MUX2_X1 U10175 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9258), .S(n10620), .Z(
        P2_U3542) );
  INV_X1 U10176 ( .A(n9215), .ZN(n9220) );
  AOI22_X1 U10177 ( .A1(n9217), .A2(n10404), .B1(n10403), .B2(n9216), .ZN(
        n9218) );
  OAI211_X1 U10178 ( .C1(n9220), .C2(n9245), .A(n9219), .B(n9218), .ZN(n9259)
         );
  MUX2_X1 U10179 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9259), .S(n10620), .Z(
        P2_U3541) );
  INV_X1 U10180 ( .A(n9221), .ZN(n9226) );
  AOI22_X1 U10181 ( .A1(n9223), .A2(n10404), .B1(n10403), .B2(n9222), .ZN(
        n9224) );
  OAI211_X1 U10182 ( .C1(n9226), .C2(n9245), .A(n9225), .B(n9224), .ZN(n9260)
         );
  MUX2_X1 U10183 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9260), .S(n10620), .Z(
        P2_U3540) );
  AOI211_X1 U10184 ( .C1(n10403), .C2(n6797), .A(n9228), .B(n9227), .ZN(n9229)
         );
  OAI21_X1 U10185 ( .B1(n9230), .B2(n9245), .A(n9229), .ZN(n9261) );
  MUX2_X1 U10186 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9261), .S(n10620), .Z(
        P2_U3539) );
  AOI22_X1 U10187 ( .A1(n9232), .A2(n10404), .B1(n10403), .B2(n9231), .ZN(
        n9233) );
  OAI211_X1 U10188 ( .C1(n9235), .C2(n9245), .A(n9234), .B(n9233), .ZN(n9262)
         );
  MUX2_X1 U10189 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9262), .S(n10620), .Z(
        P2_U3538) );
  AOI21_X1 U10190 ( .B1(n10403), .B2(n9237), .A(n9236), .ZN(n9238) );
  OAI211_X1 U10191 ( .C1(n9240), .C2(n9245), .A(n9239), .B(n9238), .ZN(n9263)
         );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9263), .S(n10620), .Z(
        P2_U3537) );
  AOI21_X1 U10193 ( .B1(n10403), .B2(n9242), .A(n9241), .ZN(n9243) );
  OAI211_X1 U10194 ( .C1(n9246), .C2(n9245), .A(n9244), .B(n9243), .ZN(n9264)
         );
  MUX2_X1 U10195 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9264), .S(n10620), .Z(
        P2_U3536) );
  MUX2_X1 U10196 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9247), .S(n10620), .Z(
        P2_U3533) );
  MUX2_X1 U10197 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9248), .S(n10620), .Z(
        P2_U3527) );
  MUX2_X1 U10198 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9249), .S(n10620), .Z(
        P2_U3525) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9250), .S(n10624), .Z(
        P2_U3519) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9251), .S(n10624), .Z(
        P2_U3518) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9252), .S(n10624), .Z(
        P2_U3516) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9253), .S(n10624), .Z(
        P2_U3515) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9254), .S(n10624), .Z(
        P2_U3514) );
  MUX2_X1 U10204 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9255), .S(n10624), .Z(
        P2_U3513) );
  MUX2_X1 U10205 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9256), .S(n10624), .Z(
        P2_U3512) );
  MUX2_X1 U10206 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9257), .S(n10624), .Z(
        P2_U3511) );
  MUX2_X1 U10207 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9258), .S(n10624), .Z(
        P2_U3510) );
  MUX2_X1 U10208 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9259), .S(n10624), .Z(
        P2_U3509) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9260), .S(n10624), .Z(
        P2_U3508) );
  MUX2_X1 U10210 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9261), .S(n10624), .Z(
        P2_U3507) );
  MUX2_X1 U10211 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9262), .S(n10624), .Z(
        P2_U3505) );
  MUX2_X1 U10212 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9263), .S(n10624), .Z(
        P2_U3502) );
  MUX2_X1 U10213 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9264), .S(n10624), .Z(
        P2_U3499) );
  NAND2_X1 U10214 ( .A1(n10189), .A2(n9265), .ZN(n9269) );
  NAND2_X1 U10215 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_STATE_REG_SCAN_IN), 
        .ZN(n9266) );
  OR3_X1 U10216 ( .A1(n9267), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9266), .ZN(
        n9268) );
  OAI211_X1 U10217 ( .C1(n9270), .C2(n9280), .A(n9269), .B(n9268), .ZN(
        P2_U3327) );
  INV_X1 U10218 ( .A(n9271), .ZN(n10193) );
  OAI222_X1 U10219 ( .A1(n8529), .A2(n10193), .B1(P2_U3152), .B2(n9273), .C1(
        n9272), .C2(n9280), .ZN(P2_U3329) );
  INV_X1 U10220 ( .A(n9274), .ZN(n10198) );
  OAI222_X1 U10221 ( .A1(n9280), .A2(n9276), .B1(n8529), .B2(n10198), .C1(
        n9275), .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U10222 ( .A(n10200), .ZN(n9277) );
  OAI222_X1 U10223 ( .A1(n9280), .A2(n9278), .B1(n8529), .B2(n9277), .C1(n6841), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U10224 ( .A(n10342), .ZN(n9282) );
  INV_X1 U10225 ( .A(n9279), .ZN(n10206) );
  OAI222_X1 U10226 ( .A1(P2_U3152), .A2(n9282), .B1(n8529), .B2(n10206), .C1(
        n9281), .C2(n9280), .ZN(P2_U3332) );
  INV_X1 U10227 ( .A(n9284), .ZN(n9285) );
  MUX2_X1 U10228 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9285), .S(P2_U3152), .Z(
        P2_U3358) );
  NAND2_X1 U10229 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  XOR2_X1 U10230 ( .A(n9289), .B(n9288), .Z(n9298) );
  NAND2_X1 U10231 ( .A1(n9401), .A2(n9672), .ZN(n9291) );
  OAI211_X1 U10232 ( .C1(n9292), .C2(n9405), .A(n9291), .B(n9290), .ZN(n9295)
         );
  NOR2_X1 U10233 ( .A1(n9293), .A2(n9388), .ZN(n9294) );
  AOI211_X1 U10234 ( .C1(n9296), .C2(n9402), .A(n9295), .B(n9294), .ZN(n9297)
         );
  OAI21_X1 U10235 ( .B1(n9298), .B2(n9410), .A(n9297), .ZN(P1_U3213) );
  INV_X1 U10236 ( .A(n9300), .ZN(n9302) );
  NAND2_X1 U10237 ( .A1(n9302), .A2(n9301), .ZN(n9304) );
  AOI22_X1 U10238 ( .A1(n6052), .A2(n9305), .B1(n9304), .B2(n9303), .ZN(n9310)
         );
  AOI22_X1 U10239 ( .A1(n9401), .A2(n9878), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9307) );
  NAND2_X1 U10240 ( .A1(n9402), .A2(n9883), .ZN(n9306) );
  OAI211_X1 U10241 ( .C1(n9919), .C2(n9405), .A(n9307), .B(n9306), .ZN(n9308)
         );
  AOI21_X1 U10242 ( .B1(n10094), .B2(n9408), .A(n9308), .ZN(n9309) );
  OAI21_X1 U10243 ( .B1(n9310), .B2(n9410), .A(n9309), .ZN(P1_U3214) );
  NAND2_X1 U10244 ( .A1(n9366), .A2(n9311), .ZN(n9313) );
  XOR2_X1 U10245 ( .A(n9313), .B(n9312), .Z(n9318) );
  NAND2_X1 U10246 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9774) );
  OAI21_X1 U10247 ( .B1(n9405), .B2(n9975), .A(n9774), .ZN(n9314) );
  AOI21_X1 U10248 ( .B1(n9401), .B2(n9944), .A(n9314), .ZN(n9315) );
  OAI21_X1 U10249 ( .B1(n9395), .B2(n9946), .A(n9315), .ZN(n9316) );
  AOI21_X1 U10250 ( .B1(n10117), .B2(n9408), .A(n9316), .ZN(n9317) );
  OAI21_X1 U10251 ( .B1(n9318), .B2(n9410), .A(n9317), .ZN(P1_U3217) );
  INV_X1 U10252 ( .A(n9319), .ZN(n9323) );
  NAND2_X1 U10253 ( .A1(n4896), .A2(n9322), .ZN(n9320) );
  AOI22_X1 U10254 ( .A1(n9323), .A2(n9322), .B1(n9321), .B2(n9320), .ZN(n9329)
         );
  NOR2_X1 U10255 ( .A1(n9395), .A2(n9918), .ZN(n9327) );
  AOI22_X1 U10256 ( .A1(n9879), .A2(n9401), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9324) );
  OAI21_X1 U10257 ( .B1(n9325), .B2(n9405), .A(n9324), .ZN(n9326) );
  AOI211_X1 U10258 ( .C1(n10108), .C2(n9408), .A(n9327), .B(n9326), .ZN(n9328)
         );
  OAI21_X1 U10259 ( .B1(n9329), .B2(n9410), .A(n9328), .ZN(P1_U3221) );
  XNOR2_X1 U10260 ( .A(n9332), .B(n9331), .ZN(n9333) );
  XNOR2_X1 U10261 ( .A(n9330), .B(n9333), .ZN(n9338) );
  AOI22_X1 U10262 ( .A1(n9401), .A2(n9844), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9335) );
  NAND2_X1 U10263 ( .A1(n9402), .A2(n9847), .ZN(n9334) );
  OAI211_X1 U10264 ( .C1(n9469), .C2(n9405), .A(n9335), .B(n9334), .ZN(n9336)
         );
  AOI21_X1 U10265 ( .B1(n10084), .B2(n9408), .A(n9336), .ZN(n9337) );
  OAI21_X1 U10266 ( .B1(n9338), .B2(n9410), .A(n9337), .ZN(P1_U3223) );
  OAI21_X1 U10267 ( .B1(n9340), .B2(n8544), .A(n9339), .ZN(n9341) );
  NAND2_X1 U10268 ( .A1(n9341), .A2(n9381), .ZN(n9346) );
  NOR2_X1 U10269 ( .A1(n9405), .A2(n9996), .ZN(n9344) );
  INV_X1 U10270 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9721) );
  OAI22_X1 U10271 ( .A1(n9342), .A2(n9999), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9721), .ZN(n9343) );
  AOI211_X1 U10272 ( .C1(n10004), .C2(n9402), .A(n9344), .B(n9343), .ZN(n9345)
         );
  OAI211_X1 U10273 ( .C1(n8630), .C2(n9388), .A(n9346), .B(n9345), .ZN(
        P1_U3224) );
  XNOR2_X1 U10274 ( .A(n9349), .B(n9348), .ZN(n9350) );
  XNOR2_X1 U10275 ( .A(n9347), .B(n9350), .ZN(n9356) );
  NOR2_X1 U10276 ( .A1(n9351), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9733) );
  AOI21_X1 U10277 ( .B1(n9401), .B2(n9943), .A(n9733), .ZN(n9353) );
  NAND2_X1 U10278 ( .A1(n9402), .A2(n9983), .ZN(n9352) );
  OAI211_X1 U10279 ( .C1(n10016), .C2(n9405), .A(n9353), .B(n9352), .ZN(n9354)
         );
  AOI21_X1 U10280 ( .B1(n10128), .B2(n9408), .A(n9354), .ZN(n9355) );
  OAI21_X1 U10281 ( .B1(n9356), .B2(n9410), .A(n9355), .ZN(P1_U3226) );
  INV_X1 U10282 ( .A(n9357), .ZN(n9358) );
  AOI21_X1 U10283 ( .B1(n9359), .B2(n9299), .A(n9358), .ZN(n9365) );
  AOI22_X1 U10284 ( .A1(n9401), .A2(n9863), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9361) );
  NAND2_X1 U10285 ( .A1(n9402), .A2(n9869), .ZN(n9360) );
  OAI211_X1 U10286 ( .C1(n9362), .C2(n9405), .A(n9361), .B(n9360), .ZN(n9363)
         );
  AOI21_X1 U10287 ( .B1(n10090), .B2(n9408), .A(n9363), .ZN(n9364) );
  OAI21_X1 U10288 ( .B1(n9365), .B2(n9410), .A(n9364), .ZN(P1_U3227) );
  NAND2_X1 U10289 ( .A1(n9367), .A2(n9366), .ZN(n9371) );
  XNOR2_X1 U10290 ( .A(n9369), .B(n9368), .ZN(n9370) );
  XNOR2_X1 U10291 ( .A(n9371), .B(n9370), .ZN(n9377) );
  NOR2_X1 U10292 ( .A1(n9395), .A2(n9931), .ZN(n9375) );
  AOI22_X1 U10293 ( .A1(n9928), .A2(n9401), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9372) );
  OAI21_X1 U10294 ( .B1(n9373), .B2(n9405), .A(n9372), .ZN(n9374) );
  AOI211_X1 U10295 ( .C1(n10112), .C2(n9408), .A(n9375), .B(n9374), .ZN(n9376)
         );
  OAI21_X1 U10296 ( .B1(n9377), .B2(n9410), .A(n9376), .ZN(P1_U3231) );
  INV_X1 U10297 ( .A(n10102), .ZN(n9905) );
  OAI21_X1 U10298 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9382) );
  NAND2_X1 U10299 ( .A1(n9382), .A2(n9381), .ZN(n9387) );
  AOI22_X1 U10300 ( .A1(n9401), .A2(n9897), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9383) );
  OAI21_X1 U10301 ( .B1(n9384), .B2(n9405), .A(n9383), .ZN(n9385) );
  AOI21_X1 U10302 ( .B1(n9903), .B2(n9402), .A(n9385), .ZN(n9386) );
  OAI211_X1 U10303 ( .C1(n9905), .C2(n9388), .A(n9387), .B(n9386), .ZN(
        P1_U3233) );
  XOR2_X1 U10304 ( .A(n9390), .B(n9389), .Z(n9391) );
  XNOR2_X1 U10305 ( .A(n9392), .B(n9391), .ZN(n9398) );
  NAND2_X1 U10306 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9746) );
  OAI21_X1 U10307 ( .B1(n9405), .B2(n9999), .A(n9746), .ZN(n9393) );
  AOI21_X1 U10308 ( .B1(n9401), .B2(n9956), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10309 ( .B1(n9395), .B2(n9966), .A(n9394), .ZN(n9396) );
  AOI21_X1 U10310 ( .B1(n10123), .B2(n9408), .A(n9396), .ZN(n9397) );
  OAI21_X1 U10311 ( .B1(n9398), .B2(n9410), .A(n9397), .ZN(P1_U3236) );
  XNOR2_X1 U10312 ( .A(n9399), .B(n9400), .ZN(n9411) );
  AOI22_X1 U10313 ( .A1(n9401), .A2(n9826), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9404) );
  NAND2_X1 U10314 ( .A1(n9402), .A2(n9832), .ZN(n9403) );
  OAI211_X1 U10315 ( .C1(n9406), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9407)
         );
  AOI21_X1 U10316 ( .B1(n10079), .B2(n9408), .A(n9407), .ZN(n9409) );
  OAI21_X1 U10317 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(P1_U3238) );
  INV_X1 U10318 ( .A(n9485), .ZN(n9504) );
  MUX2_X1 U10319 ( .A(n9539), .B(n9603), .S(n9504), .Z(n9479) );
  MUX2_X1 U10320 ( .A(n9537), .B(n9599), .S(n9485), .Z(n9476) );
  OAI21_X1 U10321 ( .B1(n9542), .B2(n9485), .A(n9855), .ZN(n9475) );
  MUX2_X1 U10322 ( .A(n9641), .B(n9592), .S(n9485), .Z(n9465) );
  NAND2_X1 U10323 ( .A1(n9415), .A2(n9412), .ZN(n9591) );
  NAND2_X1 U10324 ( .A1(n9591), .A2(n9416), .ZN(n9418) );
  INV_X1 U10325 ( .A(n9413), .ZN(n9414) );
  NAND2_X1 U10326 ( .A1(n9415), .A2(n9414), .ZN(n9417) );
  AND2_X1 U10327 ( .A1(n9417), .A2(n9416), .ZN(n9589) );
  MUX2_X1 U10328 ( .A(n9418), .B(n9589), .S(n9485), .Z(n9463) );
  MUX2_X1 U10329 ( .A(n9546), .B(n9580), .S(n9485), .Z(n9457) );
  XNOR2_X1 U10330 ( .A(n10510), .B(n9504), .ZN(n9419) );
  NAND2_X1 U10331 ( .A1(n9419), .A2(n10509), .ZN(n9421) );
  NAND2_X1 U10332 ( .A1(n9421), .A2(n9636), .ZN(n9420) );
  NAND2_X1 U10333 ( .A1(n9420), .A2(n9422), .ZN(n9426) );
  NAND2_X1 U10334 ( .A1(n9421), .A2(n9632), .ZN(n9424) );
  INV_X1 U10335 ( .A(n9422), .ZN(n10034) );
  AOI21_X1 U10336 ( .B1(n9424), .B2(n9423), .A(n10034), .ZN(n9425) );
  INV_X1 U10337 ( .A(n9427), .ZN(n9517) );
  MUX2_X1 U10338 ( .A(n9428), .B(n10033), .S(n9504), .Z(n9429) );
  MUX2_X1 U10339 ( .A(n9550), .B(n8040), .S(n9485), .Z(n9432) );
  NAND3_X1 U10340 ( .A1(n9433), .A2(n9518), .A3(n9432), .ZN(n9438) );
  AND2_X1 U10341 ( .A1(n9563), .A2(n9560), .ZN(n9436) );
  NOR2_X1 U10342 ( .A1(n9435), .A2(n5177), .ZN(n9549) );
  MUX2_X1 U10343 ( .A(n9436), .B(n9549), .S(n9485), .Z(n9437) );
  NAND2_X1 U10344 ( .A1(n9438), .A2(n9437), .ZN(n9443) );
  MUX2_X1 U10345 ( .A(n9674), .B(n9439), .S(n9504), .Z(n9440) );
  NAND2_X1 U10346 ( .A1(n9520), .A2(n9440), .ZN(n9441) );
  AND2_X1 U10347 ( .A1(n9522), .A2(n9441), .ZN(n9442) );
  NAND2_X1 U10348 ( .A1(n9443), .A2(n9442), .ZN(n9445) );
  AOI21_X1 U10349 ( .B1(n9445), .B2(n9564), .A(n9444), .ZN(n9451) );
  NAND3_X1 U10350 ( .A1(n9570), .A2(n9504), .A3(n9569), .ZN(n9450) );
  NAND2_X1 U10351 ( .A1(n9445), .A2(n9566), .ZN(n9446) );
  NAND2_X1 U10352 ( .A1(n9446), .A2(n9569), .ZN(n9447) );
  NAND4_X1 U10353 ( .A1(n9447), .A2(n9567), .A3(n9547), .A4(n9485), .ZN(n9449)
         );
  MUX2_X1 U10354 ( .A(n9547), .B(n9570), .S(n9485), .Z(n9448) );
  MUX2_X1 U10355 ( .A(n9548), .B(n9575), .S(n9485), .Z(n9452) );
  NAND3_X1 U10356 ( .A1(n9453), .A2(n9994), .A3(n9452), .ZN(n9455) );
  MUX2_X1 U10357 ( .A(n9545), .B(n9576), .S(n9504), .Z(n9454) );
  NAND3_X1 U10358 ( .A1(n9455), .A2(n9977), .A3(n9454), .ZN(n9456) );
  MUX2_X1 U10359 ( .A(n9583), .B(n9582), .S(n9485), .Z(n9458) );
  MUX2_X1 U10360 ( .A(n9586), .B(n9587), .S(n9504), .Z(n9459) );
  OAI21_X1 U10361 ( .B1(n9460), .B2(n9941), .A(n9459), .ZN(n9461) );
  NAND3_X1 U10362 ( .A1(n9915), .A2(n9935), .A3(n9461), .ZN(n9462) );
  NAND3_X1 U10363 ( .A1(n9901), .A2(n9463), .A3(n9462), .ZN(n9464) );
  NAND3_X1 U10364 ( .A1(n9876), .A2(n9465), .A3(n9464), .ZN(n9468) );
  NAND2_X1 U10365 ( .A1(n9542), .A2(n9594), .ZN(n9466) );
  NAND2_X1 U10366 ( .A1(n9466), .A2(n9485), .ZN(n9467) );
  NAND2_X1 U10367 ( .A1(n9468), .A2(n9467), .ZN(n9472) );
  OR2_X1 U10368 ( .A1(n10090), .A2(n9469), .ZN(n9471) );
  NAND2_X1 U10369 ( .A1(n9471), .A2(n9470), .ZN(n9597) );
  AOI22_X1 U10370 ( .A1(n9472), .A2(n9471), .B1(n9504), .B2(n9597), .ZN(n9474)
         );
  MUX2_X1 U10371 ( .A(n9543), .B(n9598), .S(n9504), .Z(n9473) );
  AND3_X1 U10372 ( .A1(n9791), .A2(n9479), .A3(n9478), .ZN(n9484) );
  INV_X1 U10373 ( .A(n9484), .ZN(n9480) );
  NAND3_X1 U10374 ( .A1(n9480), .A2(n9541), .A3(n9649), .ZN(n9481) );
  NAND2_X1 U10375 ( .A1(n9481), .A2(n9483), .ZN(n9487) );
  NAND2_X1 U10376 ( .A1(n9483), .A2(n9482), .ZN(n9646) );
  OAI21_X1 U10377 ( .B1(n9484), .B2(n9646), .A(n9649), .ZN(n9486) );
  MUX2_X1 U10378 ( .A(n9487), .B(n9486), .S(n9485), .Z(n9501) );
  NAND2_X1 U10379 ( .A1(n10189), .A2(n9493), .ZN(n9489) );
  INV_X1 U10380 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10186) );
  OR2_X1 U10381 ( .A1(n5548), .A2(n10186), .ZN(n9488) );
  NAND2_X1 U10382 ( .A1(n4867), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9492) );
  NAND2_X1 U10383 ( .A1(n4877), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U10384 ( .A1(n4873), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9490) );
  AND3_X1 U10385 ( .A1(n9492), .A2(n9491), .A3(n9490), .ZN(n9780) );
  NAND2_X1 U10386 ( .A1(n10056), .A2(n9780), .ZN(n9654) );
  NAND2_X1 U10387 ( .A1(n9494), .A2(n9493), .ZN(n9497) );
  OR2_X1 U10388 ( .A1(n5548), .A2(n9495), .ZN(n9496) );
  INV_X1 U10389 ( .A(n9651), .ZN(n9498) );
  NAND2_X1 U10390 ( .A1(n9498), .A2(n10056), .ZN(n9500) );
  INV_X1 U10391 ( .A(n9508), .ZN(n9670) );
  INV_X1 U10392 ( .A(n9780), .ZN(n9669) );
  NAND2_X1 U10393 ( .A1(n9670), .A2(n9669), .ZN(n9499) );
  NAND2_X1 U10394 ( .A1(n10060), .A2(n9499), .ZN(n9608) );
  INV_X1 U10395 ( .A(n10056), .ZN(n9782) );
  OAI21_X1 U10396 ( .B1(n9504), .B2(n9608), .A(n9656), .ZN(n9502) );
  NAND2_X1 U10397 ( .A1(n9502), .A2(n9654), .ZN(n9507) );
  OR2_X1 U10398 ( .A1(n9651), .A2(n9780), .ZN(n9503) );
  AND2_X1 U10399 ( .A1(n9654), .A2(n9503), .ZN(n9611) );
  INV_X1 U10400 ( .A(n9611), .ZN(n9505) );
  NAND2_X1 U10401 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NAND2_X1 U10402 ( .A1(n10060), .A2(n9508), .ZN(n9650) );
  AND2_X1 U10403 ( .A1(n9651), .A2(n9650), .ZN(n9534) );
  AND4_X1 U10404 ( .A1(n10476), .A2(n5159), .A3(n9510), .A4(n9509), .ZN(n9514)
         );
  NOR2_X1 U10405 ( .A1(n9511), .A2(n10413), .ZN(n9512) );
  NAND4_X1 U10406 ( .A1(n9514), .A2(n10509), .A3(n9513), .A4(n9512), .ZN(n9515) );
  NOR2_X1 U10407 ( .A1(n9515), .A2(n10046), .ZN(n9516) );
  NAND3_X1 U10408 ( .A1(n9518), .A2(n9517), .A3(n9516), .ZN(n9519) );
  NOR2_X1 U10409 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  NAND3_X1 U10410 ( .A1(n9523), .A2(n9522), .A3(n9521), .ZN(n9524) );
  OR4_X1 U10411 ( .A1(n8596), .A2(n9991), .A3(n9525), .A4(n9524), .ZN(n9526)
         );
  OR4_X1 U10412 ( .A1(n9954), .A2(n9526), .A3(n9941), .A4(n9973), .ZN(n9527)
         );
  NOR2_X1 U10413 ( .A1(n9910), .A2(n9527), .ZN(n9528) );
  NAND3_X1 U10414 ( .A1(n9901), .A2(n9935), .A3(n9528), .ZN(n9529) );
  NOR2_X1 U10415 ( .A1(n9881), .A2(n9529), .ZN(n9530) );
  NAND4_X1 U10416 ( .A1(n9837), .A2(n9855), .A3(n9530), .A4(n9868), .ZN(n9531)
         );
  NOR4_X1 U10417 ( .A1(n9796), .A2(n9532), .A3(n9815), .A4(n9531), .ZN(n9533)
         );
  NAND4_X1 U10418 ( .A1(n9656), .A2(n9534), .A3(n9654), .A4(n9533), .ZN(n9535)
         );
  AND2_X1 U10419 ( .A1(n9535), .A2(n9620), .ZN(n9612) );
  INV_X1 U10420 ( .A(n9612), .ZN(n9536) );
  OAI21_X1 U10421 ( .B1(n9618), .B2(n6163), .A(n9536), .ZN(n9615) );
  INV_X1 U10422 ( .A(n9537), .ZN(n9538) );
  NAND2_X1 U10423 ( .A1(n9603), .A2(n9538), .ZN(n9540) );
  NAND3_X1 U10424 ( .A1(n9541), .A2(n9540), .A3(n9539), .ZN(n9606) );
  NAND2_X1 U10425 ( .A1(n9543), .A2(n9542), .ZN(n9600) );
  NAND3_X1 U10426 ( .A1(n9594), .A2(n9589), .A3(n9586), .ZN(n9544) );
  OR3_X1 U10427 ( .A1(n9606), .A2(n9600), .A3(n9544), .ZN(n9642) );
  NAND3_X1 U10428 ( .A1(n9582), .A2(n9546), .A3(n9545), .ZN(n9578) );
  AND2_X1 U10429 ( .A1(n9548), .A2(n9547), .ZN(n9573) );
  INV_X1 U10430 ( .A(n9573), .ZN(n9558) );
  INV_X1 U10431 ( .A(n9560), .ZN(n9551) );
  OAI211_X1 U10432 ( .C1(n9551), .C2(n9550), .A(n9566), .B(n9549), .ZN(n9552)
         );
  INV_X1 U10433 ( .A(n9552), .ZN(n9553) );
  AND2_X1 U10434 ( .A1(n9553), .A2(n9567), .ZN(n9562) );
  INV_X1 U10435 ( .A(n9562), .ZN(n9556) );
  INV_X1 U10436 ( .A(n9554), .ZN(n9555) );
  OR2_X1 U10437 ( .A1(n9556), .A2(n9555), .ZN(n9557) );
  OR3_X1 U10438 ( .A1(n9578), .A2(n9558), .A3(n9557), .ZN(n9637) );
  INV_X1 U10439 ( .A(n9559), .ZN(n10035) );
  NAND3_X1 U10440 ( .A1(n9560), .A2(n10033), .A3(n8040), .ZN(n9561) );
  NAND2_X1 U10441 ( .A1(n9562), .A2(n9561), .ZN(n9571) );
  NAND2_X1 U10442 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  NAND3_X1 U10443 ( .A1(n9567), .A2(n9566), .A3(n9565), .ZN(n9568) );
  NAND4_X1 U10444 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9572)
         );
  NAND2_X1 U10445 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  AND3_X1 U10446 ( .A1(n9576), .A2(n9575), .A3(n9574), .ZN(n9577) );
  OR2_X1 U10447 ( .A1(n9578), .A2(n9577), .ZN(n9644) );
  OAI21_X1 U10448 ( .B1(n9637), .B2(n10035), .A(n9644), .ZN(n9579) );
  NAND2_X1 U10449 ( .A1(n9641), .A2(n9579), .ZN(n9607) );
  INV_X1 U10450 ( .A(n9580), .ZN(n9581) );
  NAND2_X1 U10451 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  NAND2_X1 U10452 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U10453 ( .A1(n9586), .A2(n9585), .ZN(n9588) );
  NAND2_X1 U10454 ( .A1(n9588), .A2(n9587), .ZN(n9590) );
  OAI211_X1 U10455 ( .C1(n9591), .C2(n9590), .A(n9589), .B(n9641), .ZN(n9593)
         );
  NAND2_X1 U10456 ( .A1(n9593), .A2(n9592), .ZN(n9595) );
  AND2_X1 U10457 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  NOR2_X1 U10458 ( .A1(n9597), .A2(n9596), .ZN(n9601) );
  OAI211_X1 U10459 ( .C1(n9601), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9602)
         );
  INV_X1 U10460 ( .A(n9602), .ZN(n9604) );
  AND2_X1 U10461 ( .A1(n9604), .A2(n9603), .ZN(n9605) );
  OR2_X1 U10462 ( .A1(n9606), .A2(n9605), .ZN(n9645) );
  OAI21_X1 U10463 ( .B1(n9642), .B2(n9607), .A(n9645), .ZN(n9609) );
  OAI211_X1 U10464 ( .C1(n9609), .C2(n9646), .A(n9608), .B(n9649), .ZN(n9610)
         );
  AOI211_X1 U10465 ( .C1(n9611), .C2(n9610), .A(n9620), .B(n9616), .ZN(n9613)
         );
  NOR2_X1 U10466 ( .A1(n9613), .A2(n9612), .ZN(n9614) );
  NOR3_X1 U10467 ( .A1(n9616), .A2(n7722), .A3(n9620), .ZN(n9617) );
  NAND2_X1 U10468 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U10469 ( .B1(n9679), .B2(n10364), .A(n9620), .ZN(n9623) );
  NAND3_X1 U10470 ( .A1(n9623), .A2(n9622), .A3(n9621), .ZN(n9625) );
  NAND2_X1 U10471 ( .A1(n9625), .A2(n9624), .ZN(n9628) );
  OAI211_X1 U10472 ( .C1(n7764), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9631)
         );
  NAND3_X1 U10473 ( .A1(n9631), .A2(n9630), .A3(n9629), .ZN(n9635) );
  INV_X1 U10474 ( .A(n9632), .ZN(n9633) );
  AOI21_X1 U10475 ( .B1(n9635), .B2(n9634), .A(n9633), .ZN(n9640) );
  INV_X1 U10476 ( .A(n9636), .ZN(n9639) );
  INV_X1 U10477 ( .A(n9637), .ZN(n9638) );
  OAI21_X1 U10478 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9643) );
  AOI211_X1 U10479 ( .C1(n9644), .C2(n9643), .A(n5183), .B(n9642), .ZN(n9648)
         );
  INV_X1 U10480 ( .A(n9645), .ZN(n9647) );
  NOR3_X1 U10481 ( .A1(n9648), .A2(n9647), .A3(n9646), .ZN(n9653) );
  NAND2_X1 U10482 ( .A1(n9650), .A2(n9649), .ZN(n9652) );
  OAI21_X1 U10483 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n9657) );
  INV_X1 U10484 ( .A(n9654), .ZN(n9655) );
  AOI21_X1 U10485 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9658) );
  XNOR2_X1 U10486 ( .A(n9658), .B(n10494), .ZN(n9660) );
  NOR3_X1 U10487 ( .A1(n9664), .A2(n6181), .A3(n10295), .ZN(n9666) );
  OAI21_X1 U10488 ( .B1(n7722), .B2(n9667), .A(P1_B_REG_SCAN_IN), .ZN(n9665)
         );
  OAI22_X1 U10489 ( .A1(n9668), .A2(n9667), .B1(n9666), .B2(n9665), .ZN(
        P1_U3240) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9669), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9670), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9795), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9826), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9844), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9863), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9878), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9897), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9879), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9928), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9956), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9943), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9671), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9672), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9673), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9674), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9675), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10039), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9676), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10513), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9677), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10516), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9678), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10513 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9679), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10514 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9680), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10515 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7714), .S(P1_U4006), .Z(
        P1_U3555) );
  AOI21_X1 U10516 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  NOR2_X1 U10517 ( .A1(n10332), .A2(n9684), .ZN(n9685) );
  AOI211_X1 U10518 ( .C1(n10311), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9692)
         );
  OAI21_X1 U10519 ( .B1(n9689), .B2(n4918), .A(n9688), .ZN(n9690) );
  AOI22_X1 U10520 ( .A1(n10336), .A2(n9690), .B1(n10324), .B2(
        P1_ADDR_REG_4__SCAN_IN), .ZN(n9691) );
  NAND3_X1 U10521 ( .A1(n9693), .A2(n9692), .A3(n9691), .ZN(P1_U3245) );
  NOR2_X1 U10522 ( .A1(n10316), .A2(n9694), .ZN(n9695) );
  AOI211_X1 U10523 ( .C1(n10324), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9696), .B(
        n9695), .ZN(n9707) );
  OAI21_X1 U10524 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9700) );
  NAND2_X1 U10525 ( .A1(n9700), .A2(n10315), .ZN(n9706) );
  OAI21_X1 U10526 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9704) );
  NAND2_X1 U10527 ( .A1(n9704), .A2(n10336), .ZN(n9705) );
  NAND3_X1 U10528 ( .A1(n9707), .A2(n9706), .A3(n9705), .ZN(P1_U3249) );
  NOR2_X1 U10529 ( .A1(n9709), .A2(n9708), .ZN(n9711) );
  NOR2_X1 U10530 ( .A1(n9711), .A2(n9710), .ZN(n9714) );
  NAND2_X1 U10531 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9738), .ZN(n9712) );
  OAI21_X1 U10532 ( .B1(n9738), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9712), .ZN(
        n9713) );
  NOR2_X1 U10533 ( .A1(n9714), .A2(n9713), .ZN(n9737) );
  AOI211_X1 U10534 ( .C1(n9714), .C2(n9713), .A(n9737), .B(n10305), .ZN(n9727)
         );
  NAND2_X1 U10535 ( .A1(n9716), .A2(n9715), .ZN(n9718) );
  NAND2_X1 U10536 ( .A1(n9718), .A2(n9717), .ZN(n9720) );
  XOR2_X1 U10537 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9738), .Z(n9719) );
  NAND2_X1 U10538 ( .A1(n9719), .A2(n9720), .ZN(n9728) );
  OAI211_X1 U10539 ( .C1(n9720), .C2(n9719), .A(n10315), .B(n9728), .ZN(n9724)
         );
  NOR2_X1 U10540 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9721), .ZN(n9722) );
  AOI21_X1 U10541 ( .B1(n10311), .B2(n9738), .A(n9722), .ZN(n9723) );
  OAI211_X1 U10542 ( .C1(n9725), .C2(n9776), .A(n9724), .B(n9723), .ZN(n9726)
         );
  OR2_X1 U10543 ( .A1(n9727), .A2(n9726), .ZN(P1_U3257) );
  INV_X1 U10544 ( .A(n9751), .ZN(n9758) );
  XNOR2_X1 U10545 ( .A(n9758), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9732) );
  INV_X1 U10546 ( .A(n9738), .ZN(n9730) );
  INV_X1 U10547 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9729) );
  OAI21_X1 U10548 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9731) );
  NAND2_X1 U10549 ( .A1(n9732), .A2(n9731), .ZN(n9756) );
  OAI211_X1 U10550 ( .C1(n9732), .C2(n9731), .A(n9756), .B(n10315), .ZN(n9735)
         );
  INV_X1 U10551 ( .A(n9733), .ZN(n9734) );
  OAI211_X1 U10552 ( .C1(n9776), .C2(n9736), .A(n9735), .B(n9734), .ZN(n9744)
         );
  AOI21_X1 U10553 ( .B1(n9738), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9737), .ZN(
        n9742) );
  INV_X1 U10554 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U10555 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n9739), .S(n9751), .Z(n9740) );
  INV_X1 U10556 ( .A(n9740), .ZN(n9741) );
  NOR2_X1 U10557 ( .A1(n9742), .A2(n9741), .ZN(n9750) );
  AOI211_X1 U10558 ( .C1(n9742), .C2(n9741), .A(n9750), .B(n10305), .ZN(n9743)
         );
  AOI211_X1 U10559 ( .C1(n10311), .C2(n9751), .A(n9744), .B(n9743), .ZN(n9745)
         );
  INV_X1 U10560 ( .A(n9745), .ZN(P1_U3258) );
  INV_X1 U10561 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10284) );
  NAND2_X1 U10562 ( .A1(n10311), .A2(n9772), .ZN(n9747) );
  OAI211_X1 U10563 ( .C1(n9776), .C2(n10284), .A(n9747), .B(n9746), .ZN(n9764)
         );
  INV_X1 U10564 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U10565 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9748), .S(n9772), .Z(n9749) );
  INV_X1 U10566 ( .A(n9749), .ZN(n9753) );
  AOI21_X1 U10567 ( .B1(n9751), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9750), .ZN(
        n9752) );
  NOR2_X1 U10568 ( .A1(n9752), .A2(n9753), .ZN(n9771) );
  AOI211_X1 U10569 ( .C1(n9753), .C2(n9752), .A(n9771), .B(n10305), .ZN(n9763)
         );
  INV_X1 U10570 ( .A(n9772), .ZN(n9755) );
  INV_X1 U10571 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U10572 ( .A1(n9755), .A2(n9754), .ZN(n9767) );
  OAI21_X1 U10573 ( .B1(n9755), .B2(n9754), .A(n9767), .ZN(n9760) );
  INV_X1 U10574 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9757) );
  OAI21_X1 U10575 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9759) );
  NOR2_X1 U10576 ( .A1(n9759), .A2(n9760), .ZN(n9765) );
  AOI21_X1 U10577 ( .B1(n9760), .B2(n9759), .A(n9765), .ZN(n9761) );
  NOR2_X1 U10578 ( .A1(n9761), .A2(n10332), .ZN(n9762) );
  OR3_X1 U10579 ( .A1(n9764), .A2(n9763), .A3(n9762), .ZN(P1_U3259) );
  INV_X1 U10580 ( .A(n9765), .ZN(n9766) );
  NAND2_X1 U10581 ( .A1(n9767), .A2(n9766), .ZN(n9769) );
  XNOR2_X1 U10582 ( .A(n10494), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9768) );
  XNOR2_X1 U10583 ( .A(n9769), .B(n9768), .ZN(n9778) );
  INV_X1 U10584 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U10585 ( .A(n9770), .B(P1_REG2_REG_19__SCAN_IN), .S(n10494), .Z(
        n9773) );
  NAND2_X1 U10586 ( .A1(n10311), .A2(n10494), .ZN(n9775) );
  OAI211_X1 U10587 ( .C1(n9776), .C2(n5300), .A(n9775), .B(n9774), .ZN(n9777)
         );
  NAND2_X1 U10588 ( .A1(n9787), .A2(n9786), .ZN(n9785) );
  XNOR2_X1 U10589 ( .A(n9785), .B(n10056), .ZN(n10058) );
  NOR2_X1 U10590 ( .A1(n9780), .A2(n9779), .ZN(n10059) );
  INV_X1 U10591 ( .A(n10059), .ZN(n9781) );
  NOR2_X1 U10592 ( .A1(n9781), .A2(n10502), .ZN(n9789) );
  NOR2_X1 U10593 ( .A1(n9782), .A2(n10530), .ZN(n9783) );
  AOI211_X1 U10594 ( .C1(n10502), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9789), .B(
        n9783), .ZN(n9784) );
  OAI21_X1 U10595 ( .B1(n10058), .B2(n10430), .A(n9784), .ZN(P1_U3261) );
  OAI21_X1 U10596 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n10062) );
  NOR2_X1 U10597 ( .A1(n9787), .A2(n10530), .ZN(n9788) );
  AOI211_X1 U10598 ( .C1(n10502), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9789), .B(
        n9788), .ZN(n9790) );
  OAI21_X1 U10599 ( .B1(n10430), .B2(n10062), .A(n9790), .ZN(P1_U3262) );
  AND2_X1 U10600 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  AOI22_X1 U10601 ( .A1(n9795), .A2(n10514), .B1(n10515), .B2(n9826), .ZN(
        n9801) );
  AND2_X1 U10602 ( .A1(n9797), .A2(n9796), .ZN(n9799) );
  OAI21_X1 U10603 ( .B1(n9799), .B2(n9798), .A(n10511), .ZN(n9800) );
  OAI211_X1 U10604 ( .C1(n10069), .C2(n10519), .A(n9801), .B(n9800), .ZN(
        n10071) );
  INV_X1 U10605 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9803) );
  OAI22_X1 U10606 ( .A1(n10536), .A2(n9803), .B1(n9802), .B2(n10531), .ZN(
        n9804) );
  AOI21_X1 U10607 ( .B1(n10066), .B2(n10045), .A(n9804), .ZN(n9807) );
  NAND2_X1 U10608 ( .A1(n10066), .A2(n9811), .ZN(n9805) );
  AND2_X1 U10609 ( .A1(n4902), .A2(n9805), .ZN(n10067) );
  NAND2_X1 U10610 ( .A1(n10067), .A2(n10526), .ZN(n9806) );
  OAI211_X1 U10611 ( .C1(n10069), .C2(n10431), .A(n9807), .B(n9806), .ZN(n9808) );
  AOI21_X1 U10612 ( .B1(n10071), .B2(n10536), .A(n9808), .ZN(n9809) );
  INV_X1 U10613 ( .A(n9809), .ZN(P1_U3263) );
  XNOR2_X1 U10614 ( .A(n9810), .B(n9815), .ZN(n10078) );
  INV_X1 U10615 ( .A(n9811), .ZN(n9812) );
  AOI21_X1 U10616 ( .B1(n10074), .B2(n9828), .A(n9812), .ZN(n10075) );
  AOI22_X1 U10617 ( .A1(n10502), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9813), 
        .B2(n10491), .ZN(n9814) );
  OAI21_X1 U10618 ( .B1(n5120), .B2(n10530), .A(n9814), .ZN(n9823) );
  AOI21_X1 U10619 ( .B1(n9816), .B2(n9815), .A(n10479), .ZN(n9821) );
  OAI22_X1 U10620 ( .A1(n9818), .A2(n10482), .B1(n9817), .B2(n10484), .ZN(
        n9819) );
  AOI21_X1 U10621 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n10077) );
  NOR2_X1 U10622 ( .A1(n10077), .A2(n10502), .ZN(n9822) );
  AOI211_X1 U10623 ( .C1(n10075), .C2(n10526), .A(n9823), .B(n9822), .ZN(n9824) );
  OAI21_X1 U10624 ( .B1(n10078), .B2(n10012), .A(n9824), .ZN(P1_U3264) );
  XNOR2_X1 U10625 ( .A(n9825), .B(n9837), .ZN(n9827) );
  AOI222_X1 U10626 ( .A1(n10511), .A2(n9827), .B1(n9826), .B2(n10514), .C1(
        n9863), .C2(n10515), .ZN(n10082) );
  INV_X1 U10627 ( .A(n9846), .ZN(n9830) );
  INV_X1 U10628 ( .A(n9828), .ZN(n9829) );
  AOI21_X1 U10629 ( .B1(n10079), .B2(n9830), .A(n9829), .ZN(n10080) );
  NOR2_X1 U10630 ( .A1(n9831), .A2(n10530), .ZN(n9836) );
  INV_X1 U10631 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9834) );
  INV_X1 U10632 ( .A(n9832), .ZN(n9833) );
  OAI22_X1 U10633 ( .A1(n10536), .A2(n9834), .B1(n9833), .B2(n10531), .ZN(
        n9835) );
  AOI211_X1 U10634 ( .C1(n10080), .C2(n10526), .A(n9836), .B(n9835), .ZN(n9842) );
  OAI21_X1 U10635 ( .B1(n9839), .B2(n8615), .A(n9838), .ZN(n10083) );
  INV_X1 U10636 ( .A(n10083), .ZN(n9840) );
  INV_X1 U10637 ( .A(n10012), .ZN(n10048) );
  NAND2_X1 U10638 ( .A1(n9840), .A2(n10048), .ZN(n9841) );
  OAI211_X1 U10639 ( .C1(n10082), .C2(n10502), .A(n9842), .B(n9841), .ZN(
        P1_U3265) );
  XNOR2_X1 U10640 ( .A(n9843), .B(n9855), .ZN(n9845) );
  AOI222_X1 U10641 ( .A1(n10511), .A2(n9845), .B1(n9878), .B2(n10515), .C1(
        n9844), .C2(n10514), .ZN(n10087) );
  AOI21_X1 U10642 ( .B1(n10084), .B2(n9859), .A(n9846), .ZN(n10085) );
  INV_X1 U10643 ( .A(n10084), .ZN(n9849) );
  AOI22_X1 U10644 ( .A1(n10502), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9847), 
        .B2(n10491), .ZN(n9848) );
  OAI21_X1 U10645 ( .B1(n9849), .B2(n10530), .A(n9848), .ZN(n9857) );
  NAND2_X1 U10646 ( .A1(n10096), .A2(n9851), .ZN(n9853) );
  AND2_X1 U10647 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  XOR2_X1 U10648 ( .A(n9855), .B(n9854), .Z(n10088) );
  NOR2_X1 U10649 ( .A1(n10088), .A2(n10012), .ZN(n9856) );
  AOI211_X1 U10650 ( .C1(n10085), .C2(n10526), .A(n9857), .B(n9856), .ZN(n9858) );
  OAI21_X1 U10651 ( .B1(n10502), .B2(n10087), .A(n9858), .ZN(P1_U3266) );
  INV_X1 U10652 ( .A(n9859), .ZN(n9860) );
  AOI211_X1 U10653 ( .C1(n10090), .C2(n9889), .A(n10583), .B(n9860), .ZN(
        n10089) );
  OAI21_X1 U10654 ( .B1(n9861), .B2(n9868), .A(n9862), .ZN(n9864) );
  AOI222_X1 U10655 ( .A1(n10511), .A2(n9864), .B1(n9897), .B2(n10515), .C1(
        n9863), .C2(n10514), .ZN(n10092) );
  INV_X1 U10656 ( .A(n10092), .ZN(n9865) );
  AOI21_X1 U10657 ( .B1(n10089), .B2(n9900), .A(n9865), .ZN(n9875) );
  NAND2_X1 U10658 ( .A1(n10096), .A2(n9866), .ZN(n9867) );
  XOR2_X1 U10659 ( .A(n9868), .B(n9867), .Z(n10093) );
  INV_X1 U10660 ( .A(n10093), .ZN(n9873) );
  INV_X1 U10661 ( .A(n10090), .ZN(n9871) );
  AOI22_X1 U10662 ( .A1(n10502), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9869), 
        .B2(n10491), .ZN(n9870) );
  OAI21_X1 U10663 ( .B1(n9871), .B2(n10530), .A(n9870), .ZN(n9872) );
  AOI21_X1 U10664 ( .B1(n9873), .B2(n10048), .A(n9872), .ZN(n9874) );
  OAI21_X1 U10665 ( .B1(n9875), .B2(n10502), .A(n9874), .ZN(P1_U3267) );
  XNOR2_X1 U10666 ( .A(n9877), .B(n9876), .ZN(n9880) );
  AOI222_X1 U10667 ( .A1(n10511), .A2(n9880), .B1(n9879), .B2(n10515), .C1(
        n9878), .C2(n10514), .ZN(n10100) );
  OR2_X1 U10668 ( .A1(n9882), .A2(n9881), .ZN(n10097) );
  NAND3_X1 U10669 ( .A1(n10097), .A2(n10096), .A3(n10048), .ZN(n9892) );
  INV_X1 U10670 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9885) );
  INV_X1 U10671 ( .A(n9883), .ZN(n9884) );
  OAI22_X1 U10672 ( .A1(n10536), .A2(n9885), .B1(n9884), .B2(n10531), .ZN(
        n9886) );
  AOI21_X1 U10673 ( .B1(n10094), .B2(n10045), .A(n9886), .ZN(n9891) );
  NAND2_X1 U10674 ( .A1(n10094), .A2(n9894), .ZN(n9888) );
  AND2_X1 U10675 ( .A1(n9889), .A2(n9888), .ZN(n10095) );
  NAND2_X1 U10676 ( .A1(n10095), .A2(n10526), .ZN(n9890) );
  AND3_X1 U10677 ( .A1(n9892), .A2(n9891), .A3(n9890), .ZN(n9893) );
  OAI21_X1 U10678 ( .B1(n10100), .B2(n10502), .A(n9893), .ZN(P1_U3268) );
  AOI211_X1 U10679 ( .C1(n10102), .C2(n9912), .A(n10583), .B(n9887), .ZN(
        n10101) );
  OAI21_X1 U10680 ( .B1(n9901), .B2(n9895), .A(n9896), .ZN(n9898) );
  AOI222_X1 U10681 ( .A1(n10511), .A2(n9898), .B1(n9897), .B2(n10514), .C1(
        n9928), .C2(n10515), .ZN(n10104) );
  INV_X1 U10682 ( .A(n10104), .ZN(n9899) );
  AOI21_X1 U10683 ( .B1(n10101), .B2(n9900), .A(n9899), .ZN(n9909) );
  XNOR2_X1 U10684 ( .A(n9902), .B(n9901), .ZN(n10105) );
  INV_X1 U10685 ( .A(n10105), .ZN(n9907) );
  AOI22_X1 U10686 ( .A1(n9903), .A2(n10491), .B1(n10502), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9904) );
  OAI21_X1 U10687 ( .B1(n9905), .B2(n10530), .A(n9904), .ZN(n9906) );
  AOI21_X1 U10688 ( .B1(n9907), .B2(n10048), .A(n9906), .ZN(n9908) );
  OAI21_X1 U10689 ( .B1(n9909), .B2(n10502), .A(n9908), .ZN(P1_U3269) );
  XNOR2_X1 U10690 ( .A(n9911), .B(n9910), .ZN(n10111) );
  INV_X1 U10691 ( .A(n9930), .ZN(n9914) );
  INV_X1 U10692 ( .A(n9912), .ZN(n9913) );
  AOI211_X1 U10693 ( .C1(n10108), .C2(n9914), .A(n10583), .B(n9913), .ZN(
        n10106) );
  INV_X1 U10694 ( .A(n10106), .ZN(n9922) );
  XNOR2_X1 U10695 ( .A(n9916), .B(n9915), .ZN(n9917) );
  AOI22_X1 U10696 ( .A1(n9917), .A2(n10511), .B1(n10515), .B2(n9944), .ZN(
        n10109) );
  INV_X1 U10697 ( .A(n9918), .ZN(n9920) );
  NOR2_X1 U10698 ( .A1(n9919), .A2(n10484), .ZN(n10107) );
  AOI21_X1 U10699 ( .B1(n10491), .B2(n9920), .A(n10107), .ZN(n9921) );
  OAI211_X1 U10700 ( .C1(n10494), .C2(n9922), .A(n10109), .B(n9921), .ZN(n9923) );
  NAND2_X1 U10701 ( .A1(n9923), .A2(n10536), .ZN(n9925) );
  AOI22_X1 U10702 ( .A1(n10108), .A2(n10045), .B1(n10502), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9924) );
  OAI211_X1 U10703 ( .C1(n10111), .C2(n10012), .A(n9925), .B(n9924), .ZN(
        P1_U3270) );
  OAI21_X1 U10704 ( .B1(n9935), .B2(n9927), .A(n9926), .ZN(n9929) );
  AOI222_X1 U10705 ( .A1(n10511), .A2(n9929), .B1(n9928), .B2(n10514), .C1(
        n9956), .C2(n10515), .ZN(n10115) );
  AOI21_X1 U10706 ( .B1(n10112), .B2(n9948), .A(n9930), .ZN(n10113) );
  INV_X1 U10707 ( .A(n10112), .ZN(n9934) );
  INV_X1 U10708 ( .A(n9931), .ZN(n9932) );
  AOI22_X1 U10709 ( .A1(n10502), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9932), 
        .B2(n10491), .ZN(n9933) );
  OAI21_X1 U10710 ( .B1(n9934), .B2(n10530), .A(n9933), .ZN(n9938) );
  XNOR2_X1 U10711 ( .A(n9936), .B(n9935), .ZN(n10116) );
  NOR2_X1 U10712 ( .A1(n10116), .A2(n10012), .ZN(n9937) );
  AOI211_X1 U10713 ( .C1(n10113), .C2(n10526), .A(n9938), .B(n9937), .ZN(n9939) );
  OAI21_X1 U10714 ( .B1(n10502), .B2(n10115), .A(n9939), .ZN(P1_U3271) );
  XNOR2_X1 U10715 ( .A(n9940), .B(n9941), .ZN(n10121) );
  OAI21_X1 U10716 ( .B1(n4951), .B2(n8585), .A(n9942), .ZN(n9945) );
  AOI222_X1 U10717 ( .A1(n10511), .A2(n9945), .B1(n9944), .B2(n10514), .C1(
        n9943), .C2(n10515), .ZN(n10120) );
  OAI21_X1 U10718 ( .B1(n9946), .B2(n10531), .A(n10120), .ZN(n9947) );
  NAND2_X1 U10719 ( .A1(n9947), .A2(n10536), .ZN(n9952) );
  AOI21_X1 U10720 ( .B1(n10117), .B2(n9964), .A(n5115), .ZN(n10118) );
  INV_X1 U10721 ( .A(n10117), .ZN(n9949) );
  OAI22_X1 U10722 ( .A1(n9949), .A2(n10530), .B1(n9770), .B2(n10536), .ZN(
        n9950) );
  AOI21_X1 U10723 ( .B1(n10118), .B2(n10526), .A(n9950), .ZN(n9951) );
  OAI211_X1 U10724 ( .C1(n10121), .C2(n10012), .A(n9952), .B(n9951), .ZN(
        P1_U3272) );
  OAI21_X1 U10725 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n10127) );
  AOI22_X1 U10726 ( .A1(n9957), .A2(n10515), .B1(n9956), .B2(n10514), .ZN(
        n9962) );
  OAI211_X1 U10727 ( .C1(n9960), .C2(n9959), .A(n9958), .B(n10511), .ZN(n9961)
         );
  OAI211_X1 U10728 ( .C1(n10127), .C2(n10519), .A(n9962), .B(n9961), .ZN(
        n10122) );
  NAND2_X1 U10729 ( .A1(n10122), .A2(n10536), .ZN(n9971) );
  INV_X1 U10730 ( .A(n9982), .ZN(n9963) );
  NAND2_X1 U10731 ( .A1(n9963), .A2(n10123), .ZN(n9965) );
  AND2_X1 U10732 ( .A1(n9965), .A2(n9964), .ZN(n10124) );
  OAI22_X1 U10733 ( .A1(n10536), .A2(n9748), .B1(n9966), .B2(n10531), .ZN(
        n9969) );
  NOR2_X1 U10734 ( .A1(n9967), .A2(n10530), .ZN(n9968) );
  AOI211_X1 U10735 ( .C1(n10124), .C2(n10526), .A(n9969), .B(n9968), .ZN(n9970) );
  OAI211_X1 U10736 ( .C1(n10127), .C2(n10431), .A(n9971), .B(n9970), .ZN(
        P1_U3273) );
  OAI21_X1 U10737 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n9986) );
  OAI22_X1 U10738 ( .A1(n9975), .A2(n10484), .B1(n10016), .B2(n10482), .ZN(
        n9981) );
  OAI211_X1 U10739 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n10511), .ZN(n9979)
         );
  INV_X1 U10740 ( .A(n9979), .ZN(n9980) );
  AOI211_X1 U10741 ( .C1(n10555), .C2(n9986), .A(n9981), .B(n9980), .ZN(n10131) );
  AOI21_X1 U10742 ( .B1(n10128), .B2(n10001), .A(n9982), .ZN(n10129) );
  INV_X1 U10743 ( .A(n10128), .ZN(n9985) );
  AOI22_X1 U10744 ( .A1(n10502), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9983), 
        .B2(n10491), .ZN(n9984) );
  OAI21_X1 U10745 ( .B1(n9985), .B2(n10530), .A(n9984), .ZN(n9988) );
  INV_X1 U10746 ( .A(n9986), .ZN(n10132) );
  NOR2_X1 U10747 ( .A1(n10132), .A2(n10431), .ZN(n9987) );
  AOI211_X1 U10748 ( .C1(n10129), .C2(n10526), .A(n9988), .B(n9987), .ZN(n9989) );
  OAI21_X1 U10749 ( .B1(n10502), .B2(n10131), .A(n9989), .ZN(P1_U3274) );
  NAND2_X1 U10750 ( .A1(n10015), .A2(n9990), .ZN(n9992) );
  XNOR2_X1 U10751 ( .A(n9992), .B(n9991), .ZN(n10137) );
  OAI211_X1 U10752 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n10511), .ZN(n9998)
         );
  OR2_X1 U10753 ( .A1(n9996), .A2(n10482), .ZN(n9997) );
  OAI211_X1 U10754 ( .C1(n9999), .C2(n10484), .A(n9998), .B(n9997), .ZN(n10133) );
  INV_X1 U10755 ( .A(n10000), .ZN(n10026) );
  AOI21_X1 U10756 ( .B1(n10135), .B2(n10026), .A(n10583), .ZN(n10002) );
  AND2_X1 U10757 ( .A1(n10002), .A2(n10001), .ZN(n10134) );
  NAND2_X1 U10758 ( .A1(n10134), .A2(n10003), .ZN(n10009) );
  INV_X1 U10759 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10006) );
  INV_X1 U10760 ( .A(n10004), .ZN(n10005) );
  OAI22_X1 U10761 ( .A1(n10536), .A2(n10006), .B1(n10005), .B2(n10531), .ZN(
        n10007) );
  AOI21_X1 U10762 ( .B1(n10135), .B2(n10045), .A(n10007), .ZN(n10008) );
  NAND2_X1 U10763 ( .A1(n10009), .A2(n10008), .ZN(n10010) );
  AOI21_X1 U10764 ( .B1(n10133), .B2(n10536), .A(n10010), .ZN(n10011) );
  OAI21_X1 U10765 ( .B1(n10012), .B2(n10137), .A(n10011), .ZN(P1_U3275) );
  NAND2_X1 U10766 ( .A1(n10013), .A2(n10019), .ZN(n10014) );
  OAI22_X1 U10767 ( .A1(n10017), .A2(n10482), .B1(n10016), .B2(n10484), .ZN(
        n10023) );
  OAI211_X1 U10768 ( .C1(n10020), .C2(n10019), .A(n10018), .B(n10511), .ZN(
        n10021) );
  INV_X1 U10769 ( .A(n10021), .ZN(n10022) );
  AOI211_X1 U10770 ( .C1(n10138), .C2(n10555), .A(n10023), .B(n10022), .ZN(
        n10142) );
  NAND2_X1 U10771 ( .A1(n10139), .A2(n10024), .ZN(n10025) );
  AND2_X1 U10772 ( .A1(n10026), .A2(n10025), .ZN(n10140) );
  NAND2_X1 U10773 ( .A1(n10140), .A2(n10526), .ZN(n10030) );
  OAI22_X1 U10774 ( .A1(n10536), .A2(n8004), .B1(n10027), .B2(n10531), .ZN(
        n10028) );
  AOI21_X1 U10775 ( .B1(n10139), .B2(n10045), .A(n10028), .ZN(n10029) );
  NAND2_X1 U10776 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  AOI21_X1 U10777 ( .B1(n10138), .B2(n10527), .A(n10031), .ZN(n10032) );
  OAI21_X1 U10778 ( .B1(n10142), .B2(n10502), .A(n10032), .ZN(P1_U3276) );
  INV_X1 U10779 ( .A(n10033), .ZN(n10038) );
  OAI21_X1 U10780 ( .B1(n10035), .B2(n10034), .A(n10046), .ZN(n10036) );
  OAI211_X1 U10781 ( .C1(n10038), .C2(n10037), .A(n10036), .B(n10511), .ZN(
        n10041) );
  AOI22_X1 U10782 ( .A1(n10515), .A2(n10513), .B1(n10039), .B2(n10514), .ZN(
        n10040) );
  NAND2_X1 U10783 ( .A1(n10041), .A2(n10040), .ZN(n10559) );
  NAND2_X1 U10784 ( .A1(n10559), .A2(n10536), .ZN(n10055) );
  INV_X1 U10785 ( .A(n10042), .ZN(n10043) );
  OAI22_X1 U10786 ( .A1(n10536), .A2(n7397), .B1(n10043), .B2(n10531), .ZN(
        n10044) );
  AOI21_X1 U10787 ( .B1(n10560), .B2(n10045), .A(n10044), .ZN(n10054) );
  OR2_X1 U10788 ( .A1(n10047), .A2(n10046), .ZN(n10566) );
  NAND3_X1 U10789 ( .A1(n10565), .A2(n10566), .A3(n10048), .ZN(n10053) );
  AND2_X1 U10790 ( .A1(n10049), .A2(n10560), .ZN(n10050) );
  NOR2_X1 U10791 ( .A1(n10051), .A2(n10050), .ZN(n10563) );
  NAND2_X1 U10792 ( .A1(n10563), .A2(n10526), .ZN(n10052) );
  NAND4_X1 U10793 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        P1_U3283) );
  AOI21_X1 U10794 ( .B1(n10056), .B2(n10561), .A(n10059), .ZN(n10057) );
  OAI21_X1 U10795 ( .B1(n10058), .B2(n10583), .A(n10057), .ZN(n10163) );
  MUX2_X1 U10796 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10163), .S(n10591), .Z(
        P1_U3554) );
  AOI21_X1 U10797 ( .B1(n10060), .B2(n10561), .A(n10059), .ZN(n10061) );
  OAI21_X1 U10798 ( .B1(n10062), .B2(n10583), .A(n10061), .ZN(n10164) );
  MUX2_X1 U10799 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10164), .S(n10591), .Z(
        P1_U3553) );
  MUX2_X1 U10800 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10165), .S(n10591), .Z(
        P1_U3552) );
  INV_X1 U10801 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U10802 ( .A1(n10067), .A2(n10562), .B1(n10561), .B2(n10066), .ZN(
        n10068) );
  OAI21_X1 U10803 ( .B1(n10069), .B2(n10550), .A(n10068), .ZN(n10070) );
  NOR2_X1 U10804 ( .A1(n10071), .A2(n10070), .ZN(n10166) );
  MUX2_X1 U10805 ( .A(n10072), .B(n10166), .S(n10591), .Z(n10073) );
  INV_X1 U10806 ( .A(n10073), .ZN(P1_U3551) );
  AOI22_X1 U10807 ( .A1(n10075), .A2(n10562), .B1(n10561), .B2(n10074), .ZN(
        n10076) );
  OAI211_X1 U10808 ( .C1(n10078), .C2(n10162), .A(n10077), .B(n10076), .ZN(
        n10169) );
  MUX2_X1 U10809 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10169), .S(n10591), .Z(
        P1_U3550) );
  AOI22_X1 U10810 ( .A1(n10080), .A2(n10562), .B1(n10561), .B2(n10079), .ZN(
        n10081) );
  OAI211_X1 U10811 ( .C1(n10162), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10170) );
  MUX2_X1 U10812 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10170), .S(n10591), .Z(
        P1_U3549) );
  AOI22_X1 U10813 ( .A1(n10085), .A2(n10562), .B1(n10561), .B2(n10084), .ZN(
        n10086) );
  OAI211_X1 U10814 ( .C1(n10088), .C2(n10162), .A(n10087), .B(n10086), .ZN(
        n10171) );
  MUX2_X1 U10815 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10171), .S(n10591), .Z(
        P1_U3548) );
  AOI21_X1 U10816 ( .B1(n10561), .B2(n10090), .A(n10089), .ZN(n10091) );
  OAI211_X1 U10817 ( .C1(n10093), .C2(n10162), .A(n10092), .B(n10091), .ZN(
        n10172) );
  MUX2_X1 U10818 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10172), .S(n10591), .Z(
        P1_U3547) );
  AOI22_X1 U10819 ( .A1(n10095), .A2(n10562), .B1(n10561), .B2(n10094), .ZN(
        n10099) );
  INV_X1 U10820 ( .A(n10162), .ZN(n10564) );
  NAND3_X1 U10821 ( .A1(n10097), .A2(n10096), .A3(n10564), .ZN(n10098) );
  NAND3_X1 U10822 ( .A1(n10100), .A2(n10099), .A3(n10098), .ZN(n10173) );
  MUX2_X1 U10823 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10173), .S(n10591), .Z(
        P1_U3546) );
  AOI21_X1 U10824 ( .B1(n10561), .B2(n10102), .A(n10101), .ZN(n10103) );
  OAI211_X1 U10825 ( .C1(n10162), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10174) );
  MUX2_X1 U10826 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10174), .S(n10591), .Z(
        P1_U3545) );
  AOI211_X1 U10827 ( .C1(n10561), .C2(n10108), .A(n10107), .B(n10106), .ZN(
        n10110) );
  OAI211_X1 U10828 ( .C1(n10162), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10175) );
  MUX2_X1 U10829 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10175), .S(n10591), .Z(
        P1_U3544) );
  AOI22_X1 U10830 ( .A1(n10113), .A2(n10562), .B1(n10561), .B2(n10112), .ZN(
        n10114) );
  OAI211_X1 U10831 ( .C1(n10162), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10176) );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10176), .S(n10591), .Z(
        P1_U3543) );
  AOI22_X1 U10833 ( .A1(n10118), .A2(n10562), .B1(n10561), .B2(n10117), .ZN(
        n10119) );
  OAI211_X1 U10834 ( .C1(n10162), .C2(n10121), .A(n10120), .B(n10119), .ZN(
        n10177) );
  MUX2_X1 U10835 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10177), .S(n10591), .Z(
        P1_U3542) );
  INV_X1 U10836 ( .A(n10122), .ZN(n10126) );
  AOI22_X1 U10837 ( .A1(n10124), .A2(n10562), .B1(n10561), .B2(n10123), .ZN(
        n10125) );
  OAI211_X1 U10838 ( .C1(n10550), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        n10178) );
  MUX2_X1 U10839 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10178), .S(n10591), .Z(
        P1_U3541) );
  AOI22_X1 U10840 ( .A1(n10129), .A2(n10562), .B1(n10561), .B2(n10128), .ZN(
        n10130) );
  OAI211_X1 U10841 ( .C1(n10132), .C2(n10550), .A(n10131), .B(n10130), .ZN(
        n10179) );
  MUX2_X1 U10842 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10179), .S(n10591), .Z(
        P1_U3540) );
  AOI211_X1 U10843 ( .C1(n10561), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10136) );
  OAI21_X1 U10844 ( .B1(n10162), .B2(n10137), .A(n10136), .ZN(n10180) );
  MUX2_X1 U10845 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10180), .S(n10591), .Z(
        P1_U3539) );
  INV_X1 U10846 ( .A(n10138), .ZN(n10143) );
  AOI22_X1 U10847 ( .A1(n10140), .A2(n10562), .B1(n10561), .B2(n10139), .ZN(
        n10141) );
  OAI211_X1 U10848 ( .C1(n10550), .C2(n10143), .A(n10142), .B(n10141), .ZN(
        n10181) );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10181), .S(n10591), .Z(
        P1_U3538) );
  AOI211_X1 U10850 ( .C1(n10561), .C2(n10146), .A(n10145), .B(n10144), .ZN(
        n10147) );
  OAI21_X1 U10851 ( .B1(n10162), .B2(n10148), .A(n10147), .ZN(n10182) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10182), .S(n10591), .Z(
        P1_U3537) );
  INV_X1 U10853 ( .A(n10550), .ZN(n10588) );
  NAND2_X1 U10854 ( .A1(n10149), .A2(n10588), .ZN(n10154) );
  OAI22_X1 U10855 ( .A1(n10151), .A2(n10583), .B1(n10150), .B2(n10581), .ZN(
        n10152) );
  INV_X1 U10856 ( .A(n10152), .ZN(n10153) );
  NAND2_X1 U10857 ( .A1(n10154), .A2(n10153), .ZN(n10155) );
  MUX2_X1 U10858 ( .A(n10183), .B(P1_REG1_REG_13__SCAN_IN), .S(n10589), .Z(
        P1_U3536) );
  AOI211_X1 U10859 ( .C1(n10561), .C2(n10159), .A(n10158), .B(n10157), .ZN(
        n10160) );
  OAI21_X1 U10860 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(n10184) );
  MUX2_X1 U10861 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10184), .S(n10591), .Z(
        P1_U3535) );
  MUX2_X1 U10862 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10163), .S(n10595), .Z(
        P1_U3522) );
  MUX2_X1 U10863 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10164), .S(n10595), .Z(
        P1_U3521) );
  MUX2_X1 U10864 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10165), .S(n10595), .Z(
        P1_U3520) );
  INV_X1 U10865 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10167) );
  MUX2_X1 U10866 ( .A(n10167), .B(n10166), .S(n10595), .Z(n10168) );
  INV_X1 U10867 ( .A(n10168), .ZN(P1_U3519) );
  MUX2_X1 U10868 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10169), .S(n10595), .Z(
        P1_U3518) );
  MUX2_X1 U10869 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10170), .S(n10595), .Z(
        P1_U3517) );
  MUX2_X1 U10870 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10171), .S(n10595), .Z(
        P1_U3516) );
  MUX2_X1 U10871 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10172), .S(n10595), .Z(
        P1_U3515) );
  MUX2_X1 U10872 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10173), .S(n10595), .Z(
        P1_U3514) );
  MUX2_X1 U10873 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10174), .S(n10595), .Z(
        P1_U3513) );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10175), .S(n10595), .Z(
        P1_U3512) );
  MUX2_X1 U10875 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10176), .S(n10595), .Z(
        P1_U3511) );
  MUX2_X1 U10876 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10177), .S(n10595), .Z(
        P1_U3510) );
  MUX2_X1 U10877 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10178), .S(n10595), .Z(
        P1_U3508) );
  MUX2_X1 U10878 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10179), .S(n10595), .Z(
        P1_U3505) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10180), .S(n10595), .Z(
        P1_U3502) );
  MUX2_X1 U10880 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10181), .S(n10595), .Z(
        P1_U3499) );
  MUX2_X1 U10881 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10182), .S(n10595), .Z(
        P1_U3496) );
  MUX2_X1 U10882 ( .A(n10183), .B(P1_REG0_REG_13__SCAN_IN), .S(n10592), .Z(
        P1_U3493) );
  MUX2_X1 U10883 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10184), .S(n10595), .Z(
        P1_U3490) );
  INV_X1 U10884 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10185) );
  NAND3_X1 U10885 ( .A1(n10185), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10187) );
  OAI22_X1 U10886 ( .A1(n5465), .A2(n10187), .B1(n10186), .B2(n10204), .ZN(
        n10188) );
  AOI21_X1 U10887 ( .B1(n10189), .B2(n10199), .A(n10188), .ZN(n10190) );
  INV_X1 U10888 ( .A(n10190), .ZN(P1_U3322) );
  OAI222_X1 U10889 ( .A1(n10197), .A2(n10193), .B1(n10192), .B2(P1_U3084), 
        .C1(n10191), .C2(n10204), .ZN(P1_U3324) );
  AOI21_X1 U10890 ( .B1(n10195), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n10194), 
        .ZN(n10196) );
  OAI21_X1 U10891 ( .B1(n10198), .B2(n10197), .A(n10196), .ZN(P1_U3325) );
  NAND2_X1 U10892 ( .A1(n10200), .A2(n10199), .ZN(n10202) );
  OAI211_X1 U10893 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10201), .ZN(
        P1_U3326) );
  OAI222_X1 U10894 ( .A1(n10207), .A2(P1_U3084), .B1(n10197), .B2(n10206), 
        .C1(n10205), .C2(n10204), .ZN(P1_U3327) );
  MUX2_X1 U10895 ( .A(n10208), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X2 U10896 ( .A(n10210), .ZN(n10228) );
  INV_X1 U10897 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U10898 ( .A1(n10228), .A2(n10209), .ZN(P1_U3321) );
  INV_X1 U10899 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U10900 ( .A1(n10228), .A2(n10211), .ZN(P1_U3320) );
  INV_X1 U10901 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U10902 ( .A1(n10228), .A2(n10212), .ZN(P1_U3319) );
  INV_X1 U10903 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U10904 ( .A1(n10228), .A2(n10213), .ZN(P1_U3318) );
  INV_X1 U10905 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U10906 ( .A1(n10228), .A2(n10214), .ZN(P1_U3317) );
  INV_X1 U10907 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U10908 ( .A1(n10228), .A2(n10215), .ZN(P1_U3316) );
  INV_X1 U10909 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U10910 ( .A1(n10228), .A2(n10216), .ZN(P1_U3315) );
  INV_X1 U10911 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U10912 ( .A1(n10228), .A2(n10217), .ZN(P1_U3314) );
  INV_X1 U10913 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U10914 ( .A1(n10228), .A2(n10218), .ZN(P1_U3313) );
  INV_X1 U10915 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U10916 ( .A1(n10228), .A2(n10219), .ZN(P1_U3312) );
  INV_X1 U10917 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U10918 ( .A1(n10228), .A2(n10220), .ZN(P1_U3311) );
  INV_X1 U10919 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U10920 ( .A1(n10228), .A2(n10221), .ZN(P1_U3310) );
  INV_X1 U10921 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U10922 ( .A1(n10228), .A2(n10222), .ZN(P1_U3309) );
  INV_X1 U10923 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U10924 ( .A1(n10228), .A2(n10223), .ZN(P1_U3308) );
  INV_X1 U10925 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U10926 ( .A1(n10228), .A2(n10224), .ZN(P1_U3307) );
  INV_X1 U10927 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U10928 ( .A1(n10228), .A2(n10225), .ZN(P1_U3306) );
  INV_X1 U10929 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U10930 ( .A1(n10228), .A2(n10226), .ZN(P1_U3305) );
  INV_X1 U10931 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U10932 ( .A1(n10228), .A2(n10227), .ZN(P1_U3304) );
  INV_X1 U10933 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U10934 ( .A1(n10228), .A2(n10229), .ZN(P1_U3303) );
  INV_X1 U10935 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U10936 ( .A1(n10228), .A2(n10230), .ZN(P1_U3302) );
  INV_X1 U10937 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10231) );
  NOR2_X1 U10938 ( .A1(n10228), .A2(n10231), .ZN(P1_U3301) );
  INV_X1 U10939 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U10940 ( .A1(n10228), .A2(n10232), .ZN(P1_U3300) );
  INV_X1 U10941 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U10942 ( .A1(n10228), .A2(n10233), .ZN(P1_U3299) );
  INV_X1 U10943 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U10944 ( .A1(n10228), .A2(n10234), .ZN(P1_U3298) );
  INV_X1 U10945 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U10946 ( .A1(n10228), .A2(n10235), .ZN(P1_U3297) );
  INV_X1 U10947 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U10948 ( .A1(n10228), .A2(n10236), .ZN(P1_U3296) );
  INV_X1 U10949 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10237) );
  NOR2_X1 U10950 ( .A1(n10228), .A2(n10237), .ZN(P1_U3295) );
  INV_X1 U10951 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U10952 ( .A1(n10228), .A2(n10238), .ZN(P1_U3294) );
  INV_X1 U10953 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10239) );
  NOR2_X1 U10954 ( .A1(n10228), .A2(n10239), .ZN(P1_U3293) );
  INV_X1 U10955 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U10956 ( .A1(n10228), .A2(n10240), .ZN(P1_U3292) );
  NOR2_X1 U10957 ( .A1(n10342), .A2(n10241), .ZN(n10246) );
  INV_X1 U10958 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10245) );
  INV_X1 U10959 ( .A(n10242), .ZN(n10244) );
  AOI22_X1 U10960 ( .A1(n10347), .A2(n10246), .B1(n10245), .B2(n10344), .ZN(
        P2_U3438) );
  AND2_X1 U10961 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10344), .ZN(P2_U3326) );
  AND2_X1 U10962 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10344), .ZN(P2_U3325) );
  AND2_X1 U10963 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10344), .ZN(P2_U3324) );
  AND2_X1 U10964 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10344), .ZN(P2_U3323) );
  AND2_X1 U10965 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10344), .ZN(P2_U3322) );
  AND2_X1 U10966 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10344), .ZN(P2_U3321) );
  AND2_X1 U10967 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10344), .ZN(P2_U3320) );
  AND2_X1 U10968 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10344), .ZN(P2_U3319) );
  AND2_X1 U10969 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10344), .ZN(P2_U3318) );
  AND2_X1 U10970 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10344), .ZN(P2_U3317) );
  AND2_X1 U10971 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10344), .ZN(P2_U3316) );
  AND2_X1 U10972 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10344), .ZN(P2_U3315) );
  AND2_X1 U10973 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10344), .ZN(P2_U3314) );
  AND2_X1 U10974 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10344), .ZN(P2_U3313) );
  AND2_X1 U10975 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10344), .ZN(P2_U3312) );
  AND2_X1 U10976 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10344), .ZN(P2_U3311) );
  AND2_X1 U10977 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10344), .ZN(P2_U3310) );
  AND2_X1 U10978 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10344), .ZN(P2_U3309) );
  AND2_X1 U10979 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10344), .ZN(P2_U3308) );
  AND2_X1 U10980 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10344), .ZN(P2_U3307) );
  AND2_X1 U10981 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10344), .ZN(P2_U3306) );
  AND2_X1 U10982 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10344), .ZN(P2_U3305) );
  AND2_X1 U10983 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10344), .ZN(P2_U3304) );
  AND2_X1 U10984 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10344), .ZN(P2_U3303) );
  AND2_X1 U10985 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10344), .ZN(P2_U3302) );
  AND2_X1 U10986 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10344), .ZN(P2_U3301) );
  AND2_X1 U10987 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10344), .ZN(P2_U3300) );
  AND2_X1 U10988 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10344), .ZN(P2_U3299) );
  AND2_X1 U10989 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10344), .ZN(P2_U3298) );
  AND2_X1 U10990 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10344), .ZN(P2_U3297) );
  XOR2_X1 U10991 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U10992 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U10993 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  XOR2_X1 U10994 ( .A(n10251), .B(n10250), .Z(ADD_1071_U5) );
  XOR2_X1 U10995 ( .A(n10253), .B(n10252), .Z(ADD_1071_U54) );
  XOR2_X1 U10996 ( .A(n10255), .B(n10254), .Z(ADD_1071_U53) );
  XNOR2_X1 U10997 ( .A(n10257), .B(n10256), .ZN(ADD_1071_U52) );
  NOR2_X1 U10998 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  XOR2_X1 U10999 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10260), .Z(ADD_1071_U51) );
  XOR2_X1 U11000 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10261), .Z(ADD_1071_U50) );
  XOR2_X1 U11001 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10262), .Z(ADD_1071_U49) );
  XOR2_X1 U11002 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10263), .Z(ADD_1071_U48) );
  XOR2_X1 U11003 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10264), .Z(ADD_1071_U47) );
  XOR2_X1 U11004 ( .A(n10266), .B(n10265), .Z(ADD_1071_U63) );
  XOR2_X1 U11005 ( .A(n10268), .B(n10267), .Z(ADD_1071_U62) );
  XNOR2_X1 U11006 ( .A(n10270), .B(n10269), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11007 ( .A(n10272), .B(n10271), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11008 ( .A(n10274), .B(n10273), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11009 ( .A(n10276), .B(n10275), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11010 ( .A(n10278), .B(n10277), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11011 ( .A(n10280), .B(n10279), .ZN(ADD_1071_U56) );
  NOR2_X1 U11012 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  XNOR2_X1 U11013 ( .A(n10284), .B(n10283), .ZN(ADD_1071_U55) );
  INV_X1 U11014 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10286) );
  AOI21_X1 U11015 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(P1_U3441) );
  INV_X1 U11016 ( .A(n10288), .ZN(n10292) );
  OAI211_X1 U11017 ( .C1(n10290), .C2(n10294), .A(P1_STATE_REG_SCAN_IN), .B(
        n4872), .ZN(n10291) );
  OAI22_X1 U11018 ( .A1(n10332), .A2(P1_REG1_REG_0__SCAN_IN), .B1(n10292), 
        .B2(n10291), .ZN(n10297) );
  NAND3_X1 U11019 ( .A1(n10295), .A2(n10294), .A3(n10293), .ZN(n10296) );
  NAND2_X1 U11020 ( .A1(n10297), .A2(n10296), .ZN(n10299) );
  AOI22_X1 U11021 ( .A1(n10324), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10298) );
  OAI21_X1 U11022 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(P1_U3241) );
  OAI21_X1 U11023 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(n10304) );
  AOI22_X1 U11024 ( .A1(n10304), .A2(n10315), .B1(n10324), .B2(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n10314) );
  AOI211_X1 U11025 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        n10309) );
  AOI211_X1 U11026 ( .C1(n10312), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10313) );
  NAND2_X1 U11027 ( .A1(n10314), .A2(n10313), .ZN(P1_U3251) );
  NAND2_X1 U11028 ( .A1(n10315), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10317) );
  OAI21_X1 U11029 ( .B1(n10333), .B2(n10317), .A(n10316), .ZN(n10318) );
  INV_X1 U11030 ( .A(n10318), .ZN(n10341) );
  INV_X1 U11031 ( .A(n10319), .ZN(n10321) );
  INV_X1 U11032 ( .A(n10327), .ZN(n10320) );
  NOR3_X1 U11033 ( .A1(n10321), .A2(n10329), .A3(n10320), .ZN(n10322) );
  AOI211_X1 U11034 ( .C1(n10324), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10323), 
        .B(n10322), .ZN(n10339) );
  NOR2_X1 U11035 ( .A1(n10325), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10328) );
  AOI211_X1 U11036 ( .C1(n10329), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10337) );
  INV_X1 U11037 ( .A(n10330), .ZN(n10334) );
  AOI211_X1 U11038 ( .C1(n10334), .C2(n10333), .A(n10332), .B(n10331), .ZN(
        n10335) );
  AOI21_X1 U11039 ( .B1(n10337), .B2(n10336), .A(n10335), .ZN(n10338) );
  OAI211_X1 U11040 ( .C1(n10341), .C2(n10340), .A(n10339), .B(n10338), .ZN(
        P1_U3252) );
  NOR2_X1 U11041 ( .A1(n10343), .A2(n10342), .ZN(n10346) );
  INV_X1 U11042 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U11043 ( .A1(n10347), .A2(n10346), .B1(n10345), .B2(n10344), .ZN(
        P2_U3437) );
  XOR2_X1 U11044 ( .A(n5297), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11045 ( .A(n10348), .ZN(n10352) );
  OAI21_X1 U11046 ( .B1(n7736), .B2(n10581), .A(n10349), .ZN(n10351) );
  AOI211_X1 U11047 ( .C1(n10588), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10355) );
  INV_X1 U11048 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U11049 ( .A1(n10591), .A2(n10355), .B1(n10353), .B2(n10589), .ZN(
        P1_U3524) );
  INV_X1 U11050 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U11051 ( .A1(n10595), .A2(n10355), .B1(n10354), .B2(n10592), .ZN(
        P1_U3457) );
  OAI22_X1 U11052 ( .A1(n10356), .A2(n10613), .B1(n6847), .B2(n10611), .ZN(
        n10359) );
  INV_X1 U11053 ( .A(n10357), .ZN(n10358) );
  AOI211_X1 U11054 ( .C1(n10617), .C2(n10360), .A(n10359), .B(n10358), .ZN(
        n10362) );
  AOI22_X1 U11055 ( .A1(n10620), .A2(n10362), .B1(n8168), .B2(n10619), .ZN(
        P2_U3521) );
  INV_X1 U11056 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U11057 ( .A1(n10624), .A2(n10362), .B1(n10361), .B2(n10621), .ZN(
        P2_U3454) );
  INV_X1 U11058 ( .A(n10363), .ZN(n10368) );
  OAI22_X1 U11059 ( .A1(n10365), .A2(n10583), .B1(n10364), .B2(n10581), .ZN(
        n10367) );
  AOI211_X1 U11060 ( .C1(n10588), .C2(n10368), .A(n10367), .B(n10366), .ZN(
        n10371) );
  INV_X1 U11061 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U11062 ( .A1(n10591), .A2(n10371), .B1(n10369), .B2(n10589), .ZN(
        P1_U3525) );
  INV_X1 U11063 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U11064 ( .A1(n10595), .A2(n10371), .B1(n10370), .B2(n10592), .ZN(
        P1_U3460) );
  NAND2_X1 U11065 ( .A1(n10372), .A2(n4868), .ZN(n10381) );
  NAND2_X1 U11066 ( .A1(n10373), .A2(n10451), .ZN(n10380) );
  NAND2_X1 U11067 ( .A1(n6759), .A2(n10374), .ZN(n10379) );
  OAI211_X1 U11068 ( .C1(n10377), .C2(n10376), .A(n10375), .B(n8665), .ZN(
        n10378) );
  AND4_X1 U11069 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  OAI21_X1 U11070 ( .B1(n10384), .B2(n10383), .A(n10382), .ZN(P2_U3239) );
  INV_X1 U11071 ( .A(n10385), .ZN(n10387) );
  OAI22_X1 U11072 ( .A1(n10387), .A2(n10613), .B1(n10386), .B2(n10611), .ZN(
        n10389) );
  AOI211_X1 U11073 ( .C1(n10391), .C2(n10390), .A(n10389), .B(n10388), .ZN(
        n10392) );
  AOI22_X1 U11074 ( .A1(n10620), .A2(n10392), .B1(n8166), .B2(n10619), .ZN(
        P2_U3522) );
  AOI22_X1 U11075 ( .A1(n10624), .A2(n10392), .B1(n6294), .B2(n10621), .ZN(
        P2_U3457) );
  INV_X1 U11076 ( .A(n10393), .ZN(n10394) );
  AND2_X1 U11077 ( .A1(n10394), .A2(n10588), .ZN(n10397) );
  OAI22_X1 U11078 ( .A1(n10395), .A2(n10583), .B1(n7846), .B2(n10581), .ZN(
        n10396) );
  NOR3_X1 U11079 ( .A1(n10398), .A2(n10397), .A3(n10396), .ZN(n10401) );
  INV_X1 U11080 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U11081 ( .A1(n10591), .A2(n10401), .B1(n10399), .B2(n10589), .ZN(
        P1_U3526) );
  INV_X1 U11082 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U11083 ( .A1(n10595), .A2(n10401), .B1(n10400), .B2(n10592), .ZN(
        P1_U3463) );
  AOI22_X1 U11084 ( .A1(n10405), .A2(n10404), .B1(n10403), .B2(n10402), .ZN(
        n10406) );
  OAI211_X1 U11085 ( .C1(n10408), .C2(n10596), .A(n10407), .B(n10406), .ZN(
        n10409) );
  INV_X1 U11086 ( .A(n10409), .ZN(n10411) );
  AOI22_X1 U11087 ( .A1(n10620), .A2(n10411), .B1(n8165), .B2(n10619), .ZN(
        P2_U3523) );
  INV_X1 U11088 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U11089 ( .A1(n10624), .A2(n10411), .B1(n10410), .B2(n10621), .ZN(
        P2_U3460) );
  INV_X1 U11090 ( .A(n10413), .ZN(n10414) );
  XNOR2_X1 U11091 ( .A(n10412), .B(n10414), .ZN(n10432) );
  XNOR2_X1 U11092 ( .A(n10415), .B(n10414), .ZN(n10416) );
  NAND2_X1 U11093 ( .A1(n10416), .A2(n10511), .ZN(n10421) );
  OAI22_X1 U11094 ( .A1(n10418), .A2(n10482), .B1(n10417), .B2(n10484), .ZN(
        n10419) );
  INV_X1 U11095 ( .A(n10419), .ZN(n10420) );
  OAI211_X1 U11096 ( .C1(n10432), .C2(n10519), .A(n10421), .B(n10420), .ZN(
        n10439) );
  INV_X1 U11097 ( .A(n10432), .ZN(n10422) );
  AND2_X1 U11098 ( .A1(n10422), .A2(n10588), .ZN(n10426) );
  NOR2_X1 U11099 ( .A1(n10423), .A2(n10434), .ZN(n10424) );
  OR2_X1 U11100 ( .A1(n10477), .A2(n10424), .ZN(n10429) );
  OAI22_X1 U11101 ( .A1(n10429), .A2(n10583), .B1(n10434), .B2(n10581), .ZN(
        n10425) );
  NOR3_X1 U11102 ( .A1(n10439), .A2(n10426), .A3(n10425), .ZN(n10428) );
  AOI22_X1 U11103 ( .A1(n10591), .A2(n10428), .B1(n7328), .B2(n10589), .ZN(
        P1_U3527) );
  INV_X1 U11104 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U11105 ( .A1(n10595), .A2(n10428), .B1(n10427), .B2(n10592), .ZN(
        P1_U3466) );
  OAI22_X1 U11106 ( .A1(n10432), .A2(n10431), .B1(n10430), .B2(n10429), .ZN(
        n10433) );
  INV_X1 U11107 ( .A(n10433), .ZN(n10441) );
  NOR2_X1 U11108 ( .A1(n10530), .A2(n10434), .ZN(n10438) );
  INV_X1 U11109 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10436) );
  OAI22_X1 U11110 ( .A1(n10536), .A2(n10436), .B1(n10435), .B2(n10531), .ZN(
        n10437) );
  AOI211_X1 U11111 ( .C1(n10439), .C2(n10536), .A(n10438), .B(n10437), .ZN(
        n10440) );
  NAND2_X1 U11112 ( .A1(n10441), .A2(n10440), .ZN(P1_U3287) );
  XNOR2_X1 U11113 ( .A(n10447), .B(n10442), .ZN(n10458) );
  OR2_X1 U11114 ( .A1(n10443), .A2(n10462), .ZN(n10444) );
  NAND2_X1 U11115 ( .A1(n10445), .A2(n10444), .ZN(n10463) );
  OAI22_X1 U11116 ( .A1(n10463), .A2(n10613), .B1(n10462), .B2(n10611), .ZN(
        n10455) );
  XOR2_X1 U11117 ( .A(n10447), .B(n10446), .Z(n10452) );
  AOI222_X1 U11118 ( .A1(n10453), .A2(n10452), .B1(n10451), .B2(n10450), .C1(
        n10449), .C2(n10448), .ZN(n10474) );
  INV_X1 U11119 ( .A(n10474), .ZN(n10454) );
  AOI211_X1 U11120 ( .C1(n10458), .C2(n10617), .A(n10455), .B(n10454), .ZN(
        n10457) );
  AOI22_X1 U11121 ( .A1(n10620), .A2(n10457), .B1(n8163), .B2(n10619), .ZN(
        P2_U3524) );
  INV_X1 U11122 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U11123 ( .A1(n10624), .A2(n10457), .B1(n10456), .B2(n10621), .ZN(
        P2_U3463) );
  INV_X1 U11124 ( .A(n10458), .ZN(n10459) );
  OAI22_X1 U11125 ( .A1(n10462), .A2(n10461), .B1(n10460), .B2(n10459), .ZN(
        n10472) );
  INV_X1 U11126 ( .A(n10463), .ZN(n10464) );
  NAND2_X1 U11127 ( .A1(n10465), .A2(n10464), .ZN(n10468) );
  NAND2_X1 U11128 ( .A1(n10466), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10467) );
  OAI211_X1 U11129 ( .C1(n10470), .C2(n10469), .A(n10468), .B(n10467), .ZN(
        n10471) );
  NOR2_X1 U11130 ( .A1(n10472), .A2(n10471), .ZN(n10473) );
  OAI21_X1 U11131 ( .B1(n9079), .B2(n10474), .A(n10473), .ZN(P2_U3292) );
  XNOR2_X1 U11132 ( .A(n10475), .B(n7859), .ZN(n10498) );
  OAI211_X1 U11133 ( .C1(n10477), .C2(n7851), .A(n10562), .B(n10506), .ZN(
        n10495) );
  OAI21_X1 U11134 ( .B1(n7851), .B2(n10581), .A(n10495), .ZN(n10485) );
  XNOR2_X1 U11135 ( .A(n7859), .B(n10478), .ZN(n10480) );
  OAI222_X1 U11136 ( .A1(n10484), .A2(n10483), .B1(n10482), .B2(n10481), .C1(
        n10480), .C2(n10479), .ZN(n10496) );
  AOI211_X1 U11137 ( .C1(n10564), .C2(n10498), .A(n10485), .B(n10496), .ZN(
        n10488) );
  INV_X1 U11138 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11139 ( .A1(n10591), .A2(n10488), .B1(n10486), .B2(n10589), .ZN(
        P1_U3528) );
  INV_X1 U11140 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U11141 ( .A1(n10595), .A2(n10488), .B1(n10487), .B2(n10592), .ZN(
        P1_U3469) );
  INV_X1 U11142 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U11143 ( .A1(n10492), .A2(n10491), .B1(n10490), .B2(n10489), .ZN(
        n10493) );
  OAI21_X1 U11144 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10497) );
  AOI211_X1 U11145 ( .C1(n10499), .C2(n10498), .A(n10497), .B(n10496), .ZN(
        n10500) );
  AOI22_X1 U11146 ( .A1(n10502), .A2(n10501), .B1(n10500), .B2(n10536), .ZN(
        P1_U3286) );
  INV_X1 U11147 ( .A(n10503), .ZN(n10504) );
  AOI21_X1 U11148 ( .B1(n10509), .B2(n10505), .A(n10504), .ZN(n10520) );
  INV_X1 U11149 ( .A(n10520), .ZN(n10528) );
  INV_X1 U11150 ( .A(n10506), .ZN(n10508) );
  OAI21_X1 U11151 ( .B1(n10508), .B2(n10529), .A(n10507), .ZN(n10524) );
  OAI22_X1 U11152 ( .A1(n10524), .A2(n10583), .B1(n10529), .B2(n10581), .ZN(
        n10521) );
  XOR2_X1 U11153 ( .A(n10510), .B(n10509), .Z(n10512) );
  NAND2_X1 U11154 ( .A1(n10512), .A2(n10511), .ZN(n10518) );
  AOI22_X1 U11155 ( .A1(n10516), .A2(n10515), .B1(n10514), .B2(n10513), .ZN(
        n10517) );
  OAI211_X1 U11156 ( .C1(n10520), .C2(n10519), .A(n10518), .B(n10517), .ZN(
        n10537) );
  AOI211_X1 U11157 ( .C1(n10588), .C2(n10528), .A(n10521), .B(n10537), .ZN(
        n10523) );
  AOI22_X1 U11158 ( .A1(n10591), .A2(n10523), .B1(n7333), .B2(n10589), .ZN(
        P1_U3529) );
  INV_X1 U11159 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U11160 ( .A1(n10595), .A2(n10523), .B1(n10522), .B2(n10592), .ZN(
        P1_U3472) );
  INV_X1 U11161 ( .A(n10524), .ZN(n10525) );
  AOI22_X1 U11162 ( .A1(n10528), .A2(n10527), .B1(n10526), .B2(n10525), .ZN(
        n10539) );
  NOR2_X1 U11163 ( .A1(n10530), .A2(n10529), .ZN(n10535) );
  INV_X1 U11164 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10533) );
  OAI22_X1 U11165 ( .A1(n10536), .A2(n10533), .B1(n10532), .B2(n10531), .ZN(
        n10534) );
  AOI211_X1 U11166 ( .C1(n10537), .C2(n10536), .A(n10535), .B(n10534), .ZN(
        n10538) );
  NAND2_X1 U11167 ( .A1(n10539), .A2(n10538), .ZN(P1_U3285) );
  OAI22_X1 U11168 ( .A1(n10540), .A2(n10613), .B1(n5227), .B2(n10611), .ZN(
        n10541) );
  AOI21_X1 U11169 ( .B1(n10542), .B2(n10617), .A(n10541), .ZN(n10543) );
  AND2_X1 U11170 ( .A1(n10544), .A2(n10543), .ZN(n10546) );
  AOI22_X1 U11171 ( .A1(n10620), .A2(n10546), .B1(n8173), .B2(n10619), .ZN(
        P2_U3526) );
  INV_X1 U11172 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U11173 ( .A1(n10624), .A2(n10546), .B1(n10545), .B2(n10621), .ZN(
        P2_U3469) );
  INV_X1 U11174 ( .A(n10551), .ZN(n10554) );
  AOI21_X1 U11175 ( .B1(n10561), .B2(n10548), .A(n10547), .ZN(n10549) );
  OAI21_X1 U11176 ( .B1(n10551), .B2(n10550), .A(n10549), .ZN(n10553) );
  AOI211_X1 U11177 ( .C1(n10555), .C2(n10554), .A(n10553), .B(n10552), .ZN(
        n10558) );
  INV_X1 U11178 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U11179 ( .A1(n10591), .A2(n10558), .B1(n10556), .B2(n10589), .ZN(
        P1_U3530) );
  INV_X1 U11180 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U11181 ( .A1(n10595), .A2(n10558), .B1(n10557), .B2(n10592), .ZN(
        P1_U3475) );
  INV_X1 U11182 ( .A(n10559), .ZN(n10569) );
  AOI22_X1 U11183 ( .A1(n10563), .A2(n10562), .B1(n10561), .B2(n10560), .ZN(
        n10568) );
  NAND3_X1 U11184 ( .A1(n10566), .A2(n10565), .A3(n10564), .ZN(n10567) );
  AOI22_X1 U11185 ( .A1(n10591), .A2(n10572), .B1(n10570), .B2(n10589), .ZN(
        P1_U3531) );
  INV_X1 U11186 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U11187 ( .A1(n10595), .A2(n10572), .B1(n10571), .B2(n10592), .ZN(
        P1_U3478) );
  OAI21_X1 U11188 ( .B1(n10574), .B2(n10611), .A(n10573), .ZN(n10577) );
  INV_X1 U11189 ( .A(n10575), .ZN(n10576) );
  AOI211_X1 U11190 ( .C1(n10578), .C2(n10617), .A(n10577), .B(n10576), .ZN(
        n10580) );
  AOI22_X1 U11191 ( .A1(n10620), .A2(n10580), .B1(n8218), .B2(n10619), .ZN(
        P2_U3528) );
  INV_X1 U11192 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U11193 ( .A1(n10624), .A2(n10580), .B1(n10579), .B2(n10621), .ZN(
        P2_U3475) );
  OAI22_X1 U11194 ( .A1(n10584), .A2(n10583), .B1(n10582), .B2(n10581), .ZN(
        n10586) );
  AOI211_X1 U11195 ( .C1(n10588), .C2(n10587), .A(n10586), .B(n10585), .ZN(
        n10594) );
  INV_X1 U11196 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10590) );
  AOI22_X1 U11197 ( .A1(n10591), .A2(n10594), .B1(n10590), .B2(n10589), .ZN(
        P1_U3532) );
  INV_X1 U11198 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11199 ( .A1(n10595), .A2(n10594), .B1(n10593), .B2(n10592), .ZN(
        P1_U3481) );
  NOR2_X1 U11200 ( .A1(n10597), .A2(n10596), .ZN(n10601) );
  OAI22_X1 U11201 ( .A1(n10599), .A2(n10613), .B1(n10598), .B2(n10611), .ZN(
        n10600) );
  NOR3_X1 U11202 ( .A1(n10602), .A2(n10601), .A3(n10600), .ZN(n10604) );
  AOI22_X1 U11203 ( .A1(n10620), .A2(n10604), .B1(n8248), .B2(n10619), .ZN(
        P2_U3530) );
  INV_X1 U11204 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U11205 ( .A1(n10624), .A2(n10604), .B1(n10603), .B2(n10621), .ZN(
        P2_U3481) );
  OAI22_X1 U11206 ( .A1(n10605), .A2(n10613), .B1(n5212), .B2(n10611), .ZN(
        n10607) );
  AOI211_X1 U11207 ( .C1(n10608), .C2(n10617), .A(n10607), .B(n10606), .ZN(
        n10610) );
  AOI22_X1 U11208 ( .A1(n10620), .A2(n10610), .B1(n8806), .B2(n10619), .ZN(
        P2_U3532) );
  INV_X1 U11209 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U11210 ( .A1(n10624), .A2(n10610), .B1(n10609), .B2(n10621), .ZN(
        P2_U3487) );
  OAI22_X1 U11211 ( .A1(n10614), .A2(n10613), .B1(n10612), .B2(n10611), .ZN(
        n10615) );
  AOI211_X1 U11212 ( .C1(n10618), .C2(n10617), .A(n10616), .B(n10615), .ZN(
        n10623) );
  AOI22_X1 U11213 ( .A1(n10620), .A2(n10623), .B1(n8842), .B2(n10619), .ZN(
        P2_U3534) );
  INV_X1 U11214 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U11215 ( .A1(n10624), .A2(n10623), .B1(n10622), .B2(n10621), .ZN(
        P2_U3493) );
  XNOR2_X1 U11216 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI22_X1 U11217 ( .A1(n10655), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10635) );
  AOI211_X1 U11218 ( .C1(n10627), .C2(n10626), .A(n10625), .B(n10636), .ZN(
        n10628) );
  AOI21_X1 U11219 ( .B1(n10642), .B2(n10629), .A(n10628), .ZN(n10634) );
  OAI211_X1 U11220 ( .C1(n10632), .C2(n10631), .A(n10653), .B(n10630), .ZN(
        n10633) );
  NAND3_X1 U11221 ( .A1(n10635), .A2(n10634), .A3(n10633), .ZN(P2_U3247) );
  AOI22_X1 U11222 ( .A1(n10655), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10649) );
  AOI211_X1 U11223 ( .C1(n10639), .C2(n10638), .A(n10637), .B(n10636), .ZN(
        n10640) );
  AOI21_X1 U11224 ( .B1(n10642), .B2(n10641), .A(n10640), .ZN(n10648) );
  NOR2_X1 U11225 ( .A1(n10657), .A2(n10643), .ZN(n10646) );
  OAI211_X1 U11226 ( .C1(n10646), .C2(n10645), .A(n10653), .B(n10644), .ZN(
        n10647) );
  NAND3_X1 U11227 ( .A1(n10649), .A2(n10648), .A3(n10647), .ZN(P2_U3246) );
  OAI211_X1 U11228 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10651), .A(n10650), .B(
        P2_IR_REG_0__SCAN_IN), .ZN(n10652) );
  AOI21_X1 U11229 ( .B1(n10654), .B2(n6266), .A(n10652), .ZN(n10659) );
  AOI22_X1 U11230 ( .A1(n10654), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10653), .ZN(n10658) );
  AOI22_X1 U11231 ( .A1(n10655), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10656) );
  OAI221_X1 U11232 ( .B1(n10659), .B2(n10658), .C1(n10659), .C2(n10657), .A(
        n10656), .ZN(P2_U3245) );
  CLKBUF_X1 U4930 ( .A(n5618), .Z(n6090) );
  CLKBUF_X1 U4939 ( .A(n6279), .Z(n6883) );
  OR2_X1 U4943 ( .A1(n4864), .A2(n9106), .ZN(n6302) );
  CLKBUF_X1 U5130 ( .A(n6796), .Z(n9231) );
endmodule

