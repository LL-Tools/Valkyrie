

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
         n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
         n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
         n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
         n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
         n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
         n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125,
         n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
         n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
         n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
         n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
         n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
         n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
         n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
         n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
         n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
         n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269,
         n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277,
         n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
         n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293,
         n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
         n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
         n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
         n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
         n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
         n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341,
         n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
         n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
         n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
         n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
         n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
         n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397,
         n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
         n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413,
         n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
         n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
         n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
         n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
         n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461,
         n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469,
         n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
         n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485,
         n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
         n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
         n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509,
         n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
         n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
         n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533,
         n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541,
         n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
         n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557,
         n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
         n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
         n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581,
         n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
         n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
         n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
         n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613,
         n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
         n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
         n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
         n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
         n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
         n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751;

  AOI211_X1 U11262 ( .C1(n19003), .C2(n18947), .A(n16911), .B(n16910), .ZN(
        n16912) );
  AOI211_X1 U11263 ( .C1(n17457), .C2(n18948), .A(n16710), .B(n16709), .ZN(
        n16711) );
  INV_X1 U11264 ( .A(n18532), .ZN(n18520) );
  NAND2_X1 U11265 ( .A1(n13077), .A2(n11337), .ZN(n13115) );
  INV_X1 U11267 ( .A(n12043), .ZN(n16012) );
  AND2_X1 U11268 ( .A1(n12499), .A2(n12495), .ZN(n12533) );
  NOR2_X1 U11269 ( .A1(n12494), .A2(n12485), .ZN(n19615) );
  NOR2_X1 U11270 ( .A1(n17274), .A2(n17273), .ZN(n19425) );
  NAND2_X1 U11271 ( .A1(n12976), .A2(n12975), .ZN(n14843) );
  NAND2_X1 U11272 ( .A1(n12943), .A2(n12944), .ZN(n12988) );
  CLKBUF_X2 U11273 ( .A(n17233), .Z(n18029) );
  CLKBUF_X2 U11274 ( .A(n12874), .Z(n13710) );
  CLKBUF_X2 U11275 ( .A(n12847), .Z(n12903) );
  BUF_X1 U11277 ( .A(n14268), .Z(n22386) );
  CLKBUF_X2 U11278 ( .A(n17806), .Z(n11170) );
  INV_X1 U11279 ( .A(n11158), .ZN(n11168) );
  NOR2_X1 U11280 ( .A1(n12977), .A2(n14459), .ZN(n17364) );
  INV_X2 U11281 ( .A(n13924), .ZN(n13906) );
  AND2_X1 U11282 ( .A1(n15837), .A2(n14477), .ZN(n14471) );
  INV_X1 U11283 ( .A(n12977), .ZN(n22457) );
  AND2_X1 U11284 ( .A1(n11209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12144) );
  AND2_X1 U11285 ( .A1(n13943), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13911) );
  AND2_X1 U11286 ( .A1(n13938), .A2(n12086), .ZN(n13929) );
  INV_X1 U11287 ( .A(n11918), .ZN(n11902) );
  AND2_X1 U11288 ( .A1(n12811), .A2(n17370), .ZN(n13089) );
  NAND2_X1 U11289 ( .A1(n11798), .A2(n11797), .ZN(n11866) );
  AND2_X1 U11290 ( .A1(n12085), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11210) );
  INV_X2 U11291 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14755) );
  INV_X2 U11292 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14722) );
  CLKBUF_X1 U11293 ( .A(n19389), .Z(n11155) );
  NOR2_X1 U11294 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19120), .ZN(
        n19389) );
  CLKBUF_X1 U11295 ( .A(n21928), .Z(n11156) );
  NOR2_X1 U11296 ( .A1(n15907), .A2(n15840), .ZN(n21928) );
  NAND2_X2 U11297 ( .A1(n20342), .A2(n13149), .ZN(n20348) );
  BUF_X4 U11298 ( .A(n13544), .Z(n13693) );
  OAI22_X1 U11300 ( .A1(n17054), .A2(n19015), .B1(n17074), .B2(n17069), .ZN(
        n17059) );
  AND2_X1 U11301 ( .A1(n13938), .A2(n12074), .ZN(n13913) );
  OR2_X1 U11302 ( .A1(n12672), .A2(n12667), .ZN(n12669) );
  AND2_X1 U11303 ( .A1(n12085), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11209) );
  INV_X1 U11304 ( .A(n13926), .ZN(n12365) );
  AND2_X1 U11305 ( .A1(n13940), .A2(n14755), .ZN(n13930) );
  AND2_X1 U11306 ( .A1(n13940), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13928) );
  NAND2_X1 U11307 ( .A1(n11823), .A2(n11822), .ZN(n11888) );
  NAND2_X1 U11308 ( .A1(n21633), .A2(n21191), .ZN(n21183) );
  NOR2_X1 U11309 ( .A1(n21183), .A2(n17191), .ZN(n18023) );
  INV_X1 U11310 ( .A(n15881), .ZN(n15841) );
  INV_X1 U11311 ( .A(n15878), .ZN(n15886) );
  AND2_X1 U11312 ( .A1(n12650), .A2(n12651), .ZN(n12646) );
  AND2_X1 U11313 ( .A1(n11209), .A2(n14755), .ZN(n13918) );
  AND2_X1 U11314 ( .A1(n11162), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13914) );
  CLKBUF_X2 U11317 ( .A(n16024), .Z(n11166) );
  CLKBUF_X3 U11319 ( .A(n18023), .Z(n17997) );
  BUF_X1 U11320 ( .A(n16300), .Z(n20391) );
  INV_X1 U11321 ( .A(n16004), .ZN(n12574) );
  OR2_X1 U11322 ( .A1(n12835), .A2(n12834), .ZN(n14636) );
  NOR2_X2 U11323 ( .A1(n16106), .A2(n16107), .ZN(n16094) );
  NAND2_X1 U11324 ( .A1(n11855), .A2(n11893), .ZN(n14151) );
  NAND2_X1 U11325 ( .A1(n18901), .A2(n18900), .ZN(n18906) );
  AND2_X1 U11326 ( .A1(n14662), .A2(n11300), .ZN(n15061) );
  NOR2_X1 U11327 ( .A1(n11716), .A2(n15793), .ZN(n11720) );
  INV_X2 U11328 ( .A(n18830), .ZN(n11167) );
  NOR2_X1 U11329 ( .A1(n21218), .A2(n19211), .ZN(n21153) );
  INV_X1 U11330 ( .A(n20723), .ZN(n20932) );
  AOI211_X1 U11332 ( .C1(n17457), .C2(n11600), .A(n16022), .B(n16021), .ZN(
        n16023) );
  AOI211_X1 U11333 ( .C1(n19003), .C2(n19524), .A(n16037), .B(n16036), .ZN(
        n16038) );
  INV_X1 U11334 ( .A(n17221), .ZN(n17238) );
  OR2_X1 U11335 ( .A1(n17190), .A2(n21183), .ZN(n11158) );
  BUF_X1 U11336 ( .A(n17806), .Z(n11203) );
  AND2_X2 U11337 ( .A1(n12085), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11205) );
  AND2_X2 U11338 ( .A1(n12793), .A2(n11326), .ZN(n16723) );
  NAND4_X1 U11339 ( .A1(n14270), .A2(n14636), .A3(n14271), .A4(n22528), .ZN(
        n17413) );
  NAND2_X2 U11340 ( .A1(n16874), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16860) );
  NOR2_X4 U11341 ( .A1(n17468), .A2(n17099), .ZN(n16874) );
  AND2_X1 U11342 ( .A1(n17370), .A2(n14598), .ZN(n12847) );
  OR2_X1 U11343 ( .A1(n22236), .A2(n14268), .ZN(n15881) );
  NAND2_X4 U11344 ( .A1(n12068), .A2(n11854), .ZN(n11893) );
  INV_X4 U11345 ( .A(n11861), .ZN(n11854) );
  AND2_X4 U11346 ( .A1(n12809), .A2(n17368), .ZN(n11160) );
  AND2_X2 U11347 ( .A1(n12809), .A2(n17368), .ZN(n13363) );
  BUF_X4 U11348 ( .A(n18014), .Z(n18041) );
  CLKBUF_X1 U11349 ( .A(n14060), .Z(n11161) );
  CLKBUF_X3 U11350 ( .A(n14060), .Z(n11162) );
  CLKBUF_X3 U11351 ( .A(n14060), .Z(n11163) );
  AND2_X2 U11352 ( .A1(n14724), .A2(n11741), .ZN(n14060) );
  OAI22_X1 U11355 ( .A1(n11739), .A2(n11698), .B1(n16018), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11707) );
  NAND2_X2 U11356 ( .A1(n16723), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16717) );
  AOI21_X2 U11357 ( .B1(n17024), .B2(n16818), .A(n16811), .ZN(n17027) );
  AND2_X4 U11358 ( .A1(n14080), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12176) );
  AND2_X1 U11359 ( .A1(n12069), .A2(n19593), .ZN(n16024) );
  AND2_X1 U11360 ( .A1(n12810), .A2(n14597), .ZN(n12874) );
  INV_X2 U11361 ( .A(n18515), .ZN(n18527) );
  AND2_X4 U11362 ( .A1(n17369), .A2(n17368), .ZN(n13646) );
  NAND2_X2 U11363 ( .A1(n11851), .A2(n11850), .ZN(n11877) );
  INV_X1 U11364 ( .A(n17465), .ZN(n11172) );
  NOR2_X2 U11365 ( .A1(n15551), .A2(n11313), .ZN(n15767) );
  AND2_X1 U11367 ( .A1(n11336), .A2(n13179), .ZN(n11495) );
  NAND2_X1 U11368 ( .A1(n14655), .A2(n13795), .ZN(n14654) );
  AOI21_X1 U11369 ( .B1(n11677), .B2(n12558), .A(n11294), .ZN(n11349) );
  INV_X4 U11370 ( .A(n13169), .ZN(n20353) );
  NAND2_X1 U11372 ( .A1(n12491), .A2(n12476), .ZN(n18648) );
  NAND2_X1 U11373 ( .A1(n15841), .A2(n16057), .ZN(n15878) );
  INV_X4 U11374 ( .A(n15821), .ZN(n22236) );
  INV_X2 U11375 ( .A(n21211), .ZN(n20529) );
  INV_X2 U11376 ( .A(n21063), .ZN(n20997) );
  CLKBUF_X2 U11377 ( .A(n11869), .Z(n12609) );
  CLKBUF_X2 U11378 ( .A(n11890), .Z(n15617) );
  NAND2_X1 U11379 ( .A1(n11810), .A2(n11809), .ZN(n14352) );
  CLKBUF_X3 U11380 ( .A(n17232), .Z(n17991) );
  CLKBUF_X2 U11381 ( .A(n13089), .Z(n13712) );
  CLKBUF_X2 U11382 ( .A(n12945), .Z(n13720) );
  CLKBUF_X2 U11383 ( .A(n13390), .Z(n13707) );
  BUF_X2 U11384 ( .A(n12082), .Z(n12083) );
  BUF_X4 U11385 ( .A(n17264), .Z(n11169) );
  OR2_X1 U11386 ( .A1(n21182), .A2(n20535), .ZN(n11246) );
  CLKBUF_X2 U11387 ( .A(n12950), .Z(n13721) );
  INV_X2 U11388 ( .A(n17686), .ZN(n11171) );
  INV_X2 U11389 ( .A(n17363), .ZN(n13722) );
  AND2_X1 U11390 ( .A1(n14483), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12811) );
  INV_X2 U11391 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21190) );
  AND2_X1 U11393 ( .A1(n11180), .A2(n11181), .ZN(n15968) );
  NAND2_X1 U11394 ( .A1(n16713), .A2(n16712), .ZN(n16714) );
  NAND2_X1 U11395 ( .A1(n12735), .A2(n16702), .ZN(n15963) );
  OAI21_X1 U11396 ( .B1(n16002), .B2(n16001), .A(n16000), .ZN(n16009) );
  NOR2_X1 U11397 ( .A1(n16800), .A2(n17012), .ZN(n16799) );
  AND2_X1 U11398 ( .A1(n11250), .A2(n16533), .ZN(n16535) );
  NAND2_X1 U11399 ( .A1(n12712), .A2(n16746), .ZN(n11670) );
  AND2_X1 U11400 ( .A1(n16838), .A2(n16776), .ZN(n16830) );
  NOR2_X1 U11401 ( .A1(n14055), .A2(n14054), .ZN(n16539) );
  NAND2_X1 U11402 ( .A1(n11661), .A2(n11662), .ZN(n16752) );
  NOR2_X1 U11403 ( .A1(n16885), .A2(n16884), .ZN(n17146) );
  NAND3_X1 U11404 ( .A1(n11332), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n16330), .ZN(n13181) );
  NAND2_X1 U11405 ( .A1(n16564), .A2(n11251), .ZN(n14015) );
  NAND2_X1 U11406 ( .A1(n16566), .A2(n16565), .ZN(n16564) );
  NAND2_X1 U11407 ( .A1(n11333), .A2(n13169), .ZN(n16330) );
  NAND2_X1 U11408 ( .A1(n11221), .A2(n12773), .ZN(n12783) );
  NOR2_X1 U11409 ( .A1(n11647), .A2(n15787), .ZN(n11646) );
  NAND2_X1 U11410 ( .A1(n15731), .A2(n15730), .ZN(n15729) );
  OAI21_X1 U11411 ( .B1(n12773), .B2(n12779), .A(n12778), .ZN(n12780) );
  AND2_X1 U11412 ( .A1(n16610), .A2(n16609), .ZN(n18956) );
  NAND2_X1 U11413 ( .A1(n15069), .A2(n11637), .ZN(n12775) );
  INV_X1 U11414 ( .A(n15999), .ZN(n11173) );
  CLKBUF_X1 U11415 ( .A(n12771), .Z(n12776) );
  NOR2_X1 U11416 ( .A1(n21495), .A2(n21476), .ZN(n18331) );
  AND2_X1 U11417 ( .A1(n16653), .A2(n16638), .ZN(n16640) );
  OR2_X1 U11418 ( .A1(n11347), .A2(n11349), .ZN(n11346) );
  NOR2_X1 U11419 ( .A1(n16659), .A2(n16652), .ZN(n16653) );
  NAND2_X1 U11420 ( .A1(n11347), .A2(n11349), .ZN(n12614) );
  INV_X1 U11421 ( .A(n14654), .ZN(n13796) );
  NAND2_X1 U11422 ( .A1(n11353), .A2(n12769), .ZN(n11640) );
  OR2_X1 U11423 ( .A1(n16673), .A2(n16661), .ZN(n16659) );
  AND2_X1 U11424 ( .A1(n12708), .A2(n16964), .ZN(n16753) );
  NAND2_X1 U11425 ( .A1(n12612), .A2(n12611), .ZN(n12777) );
  NOR2_X1 U11426 ( .A1(n19552), .A2(n19657), .ZN(n19966) );
  AND2_X1 U11427 ( .A1(n12734), .A2(n16725), .ZN(n16702) );
  OR2_X1 U11428 ( .A1(n18263), .A2(n11538), .ZN(n18287) );
  OR2_X1 U11429 ( .A1(n12607), .A2(n12606), .ZN(n12612) );
  AND2_X1 U11430 ( .A1(n18258), .A2(n11536), .ZN(n18263) );
  AOI221_X1 U11431 ( .B1(n18515), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19421), .C2(n20553), .A(n18514), .ZN(n18516) );
  AND2_X1 U11432 ( .A1(n12444), .A2(n12714), .ZN(n12719) );
  AND4_X1 U11433 ( .A1(n12557), .A2(n12556), .A3(n12555), .A4(n12554), .ZN(
        n12558) );
  NAND2_X1 U11434 ( .A1(n11335), .A2(n11334), .ZN(n16404) );
  INV_X1 U11435 ( .A(n18513), .ZN(n18521) );
  AND2_X1 U11436 ( .A1(n18257), .A2(n18242), .ZN(n11536) );
  NAND2_X1 U11437 ( .A1(n16764), .A2(n11663), .ZN(n11662) );
  OR2_X1 U11438 ( .A1(n18845), .A2(n16849), .ZN(n12691) );
  NOR2_X1 U11439 ( .A1(n21372), .A2(n18385), .ZN(n21378) );
  NAND2_X1 U11440 ( .A1(n18258), .A2(n18132), .ZN(n18186) );
  OAI22_X1 U11441 ( .A1(n12550), .A2(n12471), .B1(n12551), .B2(n13850), .ZN(
        n12483) );
  OAI22_X1 U11442 ( .A1(n12535), .A2(n12481), .B1(n12534), .B2(n12480), .ZN(
        n12482) );
  AND2_X1 U11443 ( .A1(n12443), .A2(n12701), .ZN(n12703) );
  NAND2_X2 U11444 ( .A1(n12479), .A2(n12478), .ZN(n12534) );
  AND2_X1 U11445 ( .A1(n12660), .A2(n16776), .ZN(n16836) );
  AND2_X1 U11446 ( .A1(n12499), .A2(n12498), .ZN(n12538) );
  NAND2_X1 U11447 ( .A1(n13120), .A2(n11236), .ZN(n13162) );
  NOR2_X1 U11448 ( .A1(n12502), .A2(n12485), .ZN(n12548) );
  OR2_X1 U11449 ( .A1(n18806), .A2(n12659), .ZN(n16776) );
  INV_X1 U11450 ( .A(n15615), .ZN(n12395) );
  NOR2_X2 U11451 ( .A1(n21225), .A2(n18531), .ZN(n18443) );
  NAND2_X1 U11452 ( .A1(n13078), .A2(n13115), .ZN(n15517) );
  NAND3_X1 U11453 ( .A1(n11385), .A2(n18122), .A3(n11277), .ZN(n18434) );
  NOR2_X1 U11454 ( .A1(n14536), .A2(n14526), .ZN(n14572) );
  AND2_X1 U11455 ( .A1(n12655), .A2(n12661), .ZN(n12650) );
  AND2_X1 U11456 ( .A1(n21690), .A2(n21630), .ZN(n21692) );
  NAND2_X1 U11457 ( .A1(n18441), .A2(n18442), .ZN(n18440) );
  NOR2_X1 U11458 ( .A1(n22634), .A2(n15825), .ZN(n22451) );
  NOR2_X1 U11459 ( .A1(n12669), .A2(n12656), .ZN(n12655) );
  NAND2_X1 U11460 ( .A1(n16279), .A2(n14638), .ZN(n16281) );
  INV_X2 U11461 ( .A(n21491), .ZN(n21658) );
  INV_X1 U11462 ( .A(n12495), .ZN(n12497) );
  AND2_X1 U11463 ( .A1(n11462), .A2(n11298), .ZN(n14624) );
  NAND2_X1 U11464 ( .A1(n18448), .A2(n18085), .ZN(n18441) );
  AND2_X1 U11465 ( .A1(n12493), .A2(n12492), .ZN(n12495) );
  NAND2_X1 U11466 ( .A1(n18648), .A2(n18992), .ZN(n12485) );
  NAND2_X1 U11467 ( .A1(n11581), .A2(n11292), .ZN(n12672) );
  CLKBUF_X1 U11468 ( .A(n14843), .Z(n14970) );
  INV_X1 U11469 ( .A(n12645), .ZN(n11581) );
  NAND2_X1 U11470 ( .A1(n18460), .A2(n18081), .ZN(n18148) );
  CLKBUF_X1 U11471 ( .A(n12472), .Z(n12491) );
  NOR2_X2 U11472 ( .A1(n21652), .A2(n21600), .ZN(n21603) );
  INV_X2 U11473 ( .A(n16571), .ZN(n16604) );
  OR2_X1 U11474 ( .A1(n13023), .A2(n13022), .ZN(n13024) );
  NAND2_X1 U11475 ( .A1(n13023), .A2(n13022), .ZN(n17321) );
  OR2_X2 U11476 ( .A1(n13241), .A2(n13240), .ZN(n15830) );
  AND2_X1 U11477 ( .A1(n11935), .A2(n11936), .ZN(n12461) );
  AND2_X1 U11478 ( .A1(n12492), .A2(n12473), .ZN(n18637) );
  NAND2_X1 U11479 ( .A1(n18474), .A2(n18117), .ZN(n18119) );
  NAND2_X1 U11480 ( .A1(n11944), .A2(n11943), .ZN(n11949) );
  AOI21_X2 U11481 ( .B1(n17978), .B2(n21155), .A(n21167), .ZN(n21611) );
  NOR2_X1 U11482 ( .A1(n12167), .A2(n12166), .ZN(n14690) );
  NAND2_X1 U11483 ( .A1(n18481), .A2(n18073), .ZN(n18076) );
  NAND2_X1 U11484 ( .A1(n11354), .A2(n12465), .ZN(n12473) );
  AND2_X1 U11485 ( .A1(n11703), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11700) );
  AND3_X1 U11486 ( .A1(n11929), .A2(n11931), .A3(n11930), .ZN(n11659) );
  NAND2_X1 U11487 ( .A1(n11223), .A2(n11916), .ZN(n11354) );
  OAI211_X1 U11488 ( .C1(n12037), .C2(n19030), .A(n11939), .B(n11938), .ZN(
        n11945) );
  NAND2_X1 U11489 ( .A1(n12623), .A2(n12624), .ZN(n12631) );
  NAND2_X1 U11490 ( .A1(n18482), .A2(n18483), .ZN(n18481) );
  NAND2_X1 U11491 ( .A1(n17334), .A2(n20472), .ZN(n17335) );
  CLKBUF_X1 U11492 ( .A(n13018), .Z(n13059) );
  NAND2_X1 U11493 ( .A1(n18498), .A2(n18072), .ZN(n18482) );
  INV_X1 U11494 ( .A(n17299), .ZN(n20472) );
  OR2_X1 U11495 ( .A1(n12167), .A2(n12162), .ZN(n14368) );
  AND2_X1 U11496 ( .A1(n12437), .A2(n12620), .ZN(n12623) );
  NAND2_X1 U11497 ( .A1(n18500), .A2(n18499), .ZN(n18498) );
  NAND2_X1 U11498 ( .A1(n18495), .A2(n18113), .ZN(n18115) );
  AOI21_X1 U11499 ( .B1(n14407), .B2(n12161), .A(n12160), .ZN(n12167) );
  NOR2_X1 U11500 ( .A1(n17289), .A2(n21211), .ZN(n21666) );
  OR2_X1 U11501 ( .A1(n17294), .A2(n11503), .ZN(n17289) );
  AND2_X1 U11502 ( .A1(n14399), .A2(n14400), .ZN(n12141) );
  AND2_X1 U11503 ( .A1(n12937), .A2(n12938), .ZN(n11328) );
  CLKBUF_X1 U11504 ( .A(n11920), .Z(n11921) );
  NAND2_X1 U11505 ( .A1(n13038), .A2(n13036), .ZN(n13239) );
  NOR2_X1 U11506 ( .A1(n11579), .A2(n11577), .ZN(n11576) );
  AND2_X1 U11507 ( .A1(n12577), .A2(n12432), .ZN(n12566) );
  OAI211_X1 U11508 ( .C1(n12372), .C2(n12758), .A(n12158), .B(n12114), .ZN(
        n14400) );
  INV_X2 U11509 ( .A(n16057), .ZN(n15889) );
  NAND2_X1 U11510 ( .A1(n11891), .A2(n14322), .ZN(n14350) );
  NAND2_X2 U11511 ( .A1(n12936), .A2(n15883), .ZN(n15897) );
  INV_X2 U11512 ( .A(n12936), .ZN(n16057) );
  AND2_X1 U11513 ( .A1(n14320), .A2(n15617), .ZN(n11891) );
  AND3_X1 U11514 ( .A1(n15892), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15821), 
        .ZN(n13220) );
  AND2_X2 U11515 ( .A1(n11856), .A2(n12070), .ZN(n12093) );
  OR2_X1 U11516 ( .A1(n12182), .A2(n12181), .ZN(n12507) );
  NAND3_X1 U11517 ( .A1(n17284), .A2(n17283), .A3(n17282), .ZN(n21211) );
  AND2_X1 U11518 ( .A1(n12137), .A2(n12136), .ZN(n12759) );
  AND2_X1 U11519 ( .A1(n12113), .A2(n12112), .ZN(n12758) );
  AND2_X2 U11521 ( .A1(n15825), .A2(n12977), .ZN(n14271) );
  AND2_X1 U11522 ( .A1(n12069), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13762) );
  NAND3_X1 U11523 ( .A1(n11867), .A2(n11881), .A3(n19528), .ZN(n11892) );
  NAND2_X1 U11524 ( .A1(n13247), .A2(n14477), .ZN(n14637) );
  INV_X1 U11525 ( .A(n19425), .ZN(n11507) );
  AND2_X1 U11526 ( .A1(n11877), .A2(n14352), .ZN(n11875) );
  OR2_X1 U11527 ( .A1(n12157), .A2(n12156), .ZN(n12764) );
  NOR2_X1 U11528 ( .A1(n15524), .A2(n15892), .ZN(n14270) );
  NAND3_X1 U11529 ( .A1(n17231), .A2(n17230), .A3(n17229), .ZN(n21063) );
  AND2_X1 U11530 ( .A1(n13761), .A2(n11860), .ZN(n11853) );
  INV_X1 U11531 ( .A(n14352), .ZN(n14921) );
  INV_X2 U11532 ( .A(U212), .ZN(n11174) );
  INV_X2 U11533 ( .A(n11869), .ZN(n12069) );
  AND2_X1 U11534 ( .A1(n11769), .A2(n11768), .ZN(n11869) );
  INV_X1 U11535 ( .A(n11888), .ZN(n11860) );
  NAND2_X2 U11536 ( .A1(n11220), .A2(n11675), .ZN(n14477) );
  INV_X1 U11538 ( .A(n11866), .ZN(n11355) );
  AND4_X1 U11539 ( .A1(n12860), .A2(n12859), .A3(n12858), .A4(n12857), .ZN(
        n12866) );
  NAND2_X2 U11540 ( .A1(U214), .A2(n20401), .ZN(n20456) );
  NAND2_X1 U11541 ( .A1(n11836), .A2(n11835), .ZN(n11890) );
  INV_X2 U11542 ( .A(U214), .ZN(n20446) );
  INV_X1 U11544 ( .A(n11158), .ZN(n11207) );
  NAND3_X1 U11545 ( .A1(n11796), .A2(n11795), .A3(n11794), .ZN(n11797) );
  OAI21_X1 U11546 ( .B1(n11834), .B2(n11833), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11835) );
  AND3_X1 U11547 ( .A1(n11843), .A2(n11842), .A3(n14755), .ZN(n11844) );
  AND2_X2 U11548 ( .A1(n14083), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12241) );
  NAND2_X2 U11549 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20459), .ZN(n20260) );
  OR2_X2 U11550 ( .A1(n20459), .A2(n17426), .ZN(n17357) );
  OR2_X2 U11551 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14149), .ZN(n18830) );
  AND2_X1 U11552 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  AND2_X1 U11553 ( .A1(n11841), .A2(n11840), .ZN(n11843) );
  AND2_X1 U11554 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  AND3_X1 U11555 ( .A1(n11793), .A2(n11792), .A3(n11791), .ZN(n11796) );
  INV_X2 U11556 ( .A(n19293), .ZN(U215) );
  NAND2_X1 U11557 ( .A1(n12083), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13924) );
  INV_X4 U11558 ( .A(n11246), .ZN(n18043) );
  CLKBUF_X2 U11559 ( .A(n12896), .Z(n13647) );
  INV_X1 U11560 ( .A(n17686), .ZN(n17901) );
  INV_X4 U11561 ( .A(n11245), .ZN(n18028) );
  CLKBUF_X3 U11562 ( .A(n13544), .Z(n13718) );
  CLKBUF_X2 U11563 ( .A(n12852), .Z(n13686) );
  INV_X2 U11564 ( .A(n21620), .ZN(n11176) );
  INV_X2 U11565 ( .A(n22749), .ZN(n20459) );
  INV_X2 U11566 ( .A(n20119), .ZN(n20179) );
  AND2_X1 U11567 ( .A1(n12810), .A2(n17370), .ZN(n12896) );
  OR2_X1 U11568 ( .A1(n21182), .A2(n17190), .ZN(n17686) );
  NAND2_X1 U11569 ( .A1(n21184), .A2(n21191), .ZN(n21173) );
  NOR2_X1 U11570 ( .A1(n17192), .A2(n17191), .ZN(n18014) );
  BUF_X4 U11571 ( .A(n18015), .Z(n11177) );
  OR2_X1 U11572 ( .A1(n21182), .A2(n17191), .ZN(n11245) );
  AND2_X1 U11573 ( .A1(n17369), .A2(n14598), .ZN(n12852) );
  AND2_X1 U11574 ( .A1(n12981), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12810) );
  AND2_X1 U11575 ( .A1(n13019), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17369) );
  AND2_X1 U11576 ( .A1(n13058), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17370) );
  NAND2_X2 U11577 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21190), .ZN(
        n17191) );
  NOR2_X2 U11578 ( .A1(n21181), .A2(n21190), .ZN(n21184) );
  INV_X1 U11579 ( .A(n11204), .ZN(n11178) );
  NAND2_X1 U11580 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21181), .ZN(
        n17190) );
  NAND2_X1 U11581 ( .A1(n21633), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n21194) );
  NAND2_X1 U11582 ( .A1(n21181), .A2(n21190), .ZN(n20535) );
  NOR2_X4 U11583 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14785) );
  AND2_X1 U11584 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12745) );
  INV_X2 U11585 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21181) );
  INV_X2 U11586 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U11587 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11718) );
  NOR2_X1 U11588 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12809) );
  NOR2_X2 U11589 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14598) );
  AND2_X2 U11590 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U11591 ( .B1(n16772), .B2(n12685), .A(n12684), .ZN(n12695) );
  AND2_X1 U11592 ( .A1(n11186), .A2(n16702), .ZN(n11179) );
  AND2_X1 U11593 ( .A1(n11186), .A2(n16702), .ZN(n16703) );
  NAND2_X1 U11594 ( .A1(n15070), .A2(n15643), .ZN(n15069) );
  XNOR2_X1 U11595 ( .A(n11640), .B(n11639), .ZN(n15070) );
  NAND2_X1 U11596 ( .A1(n12735), .A2(n11182), .ZN(n11180) );
  OR2_X1 U11597 ( .A1(n11173), .A2(n15962), .ZN(n11181) );
  AND2_X1 U11598 ( .A1(n16702), .A2(n15999), .ZN(n11182) );
  CLKBUF_X1 U11599 ( .A(n19585), .Z(n11183) );
  XNOR2_X1 U11600 ( .A(n15968), .B(n15967), .ZN(n11184) );
  CLKBUF_X1 U11601 ( .A(n15069), .Z(n11185) );
  NAND3_X1 U11602 ( .A1(n11670), .A2(n11669), .A3(n11290), .ZN(n11186) );
  NOR2_X2 U11603 ( .A1(n16717), .A2(n11654), .ZN(n16019) );
  OAI21_X1 U11604 ( .B1(n11197), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16712), .ZN(n16706) );
  NAND2_X1 U11605 ( .A1(n12730), .A2(n11190), .ZN(n11187) );
  NAND2_X1 U11606 ( .A1(n11187), .A2(n11188), .ZN(n16002) );
  OR2_X1 U11607 ( .A1(n11189), .A2(n11195), .ZN(n11188) );
  INV_X1 U11608 ( .A(n11193), .ZN(n11189) );
  AND2_X1 U11609 ( .A1(n12729), .A2(n11193), .ZN(n11190) );
  NAND2_X1 U11610 ( .A1(n12730), .A2(n12729), .ZN(n11191) );
  OR2_X1 U11611 ( .A1(n12775), .A2(n12774), .ZN(n12779) );
  OAI21_X1 U11612 ( .B1(n11221), .B2(n12782), .A(n12781), .ZN(n11192) );
  AND2_X2 U11613 ( .A1(n11378), .A2(n11377), .ZN(n11221) );
  OAI21_X1 U11614 ( .B1(n11221), .B2(n12782), .A(n12781), .ZN(n15738) );
  XNOR2_X2 U11615 ( .A(n16719), .B(n16907), .ZN(n16909) );
  OR2_X1 U11616 ( .A1(n11194), .A2(n16702), .ZN(n11193) );
  INV_X1 U11617 ( .A(n15962), .ZN(n11194) );
  AND2_X1 U11618 ( .A1(n12732), .A2(n15962), .ZN(n11195) );
  INV_X1 U11619 ( .A(n11741), .ZN(n11196) );
  NOR2_X1 U11620 ( .A1(n11179), .A2(n11279), .ZN(n11197) );
  CLKBUF_X1 U11621 ( .A(n14375), .Z(n11198) );
  AND2_X1 U11622 ( .A1(n13937), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13912) );
  AOI21_X1 U11623 ( .B1(n11917), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11932), .ZN(n11934) );
  AND2_X2 U11624 ( .A1(n11890), .A2(n11866), .ZN(n11856) );
  NAND2_X1 U11625 ( .A1(n11659), .A2(n11934), .ZN(n11936) );
  AND2_X2 U11626 ( .A1(n11376), .A2(n11909), .ZN(n12468) );
  NAND2_X1 U11627 ( .A1(n11339), .A2(n11936), .ZN(n12457) );
  NAND2_X1 U11628 ( .A1(n11267), .A2(n11439), .ZN(n12494) );
  AND2_X1 U11629 ( .A1(n14318), .A2(n11854), .ZN(n12065) );
  OAI21_X2 U11630 ( .B1(n14342), .B2(n14349), .A(n11885), .ZN(n11886) );
  INV_X2 U11631 ( .A(n21619), .ZN(n21600) );
  AND2_X1 U11632 ( .A1(n12745), .A2(n11741), .ZN(n11199) );
  AND2_X1 U11633 ( .A1(n12745), .A2(n11741), .ZN(n11200) );
  INV_X1 U11634 ( .A(n12083), .ZN(n11201) );
  AND2_X2 U11635 ( .A1(n12745), .A2(n11741), .ZN(n12082) );
  AND2_X2 U11636 ( .A1(n12085), .A2(n14722), .ZN(n11202) );
  AND2_X2 U11637 ( .A1(n12085), .A2(n14722), .ZN(n12072) );
  INV_X2 U11638 ( .A(n13944), .ZN(n14083) );
  NOR2_X1 U11639 ( .A1(n17190), .A2(n17192), .ZN(n17806) );
  AND2_X1 U11640 ( .A1(n12085), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11204) );
  INV_X4 U11641 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11741) );
  NAND2_X2 U11642 ( .A1(n11914), .A2(n11895), .ZN(n11917) );
  NOR2_X1 U11643 ( .A1(n17190), .A2(n21194), .ZN(n17264) );
  AOI21_X2 U11644 ( .B1(n12694), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11681), .ZN(n12700) );
  NAND2_X2 U11645 ( .A1(n12459), .A2(n12458), .ZN(n11439) );
  NOR2_X1 U11646 ( .A1(n21194), .A2(n20541), .ZN(n11208) );
  NOR2_X1 U11647 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21173), .ZN(
        n11211) );
  NOR2_X2 U11648 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21173), .ZN(
        n11212) );
  NOR2_X1 U11649 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21173), .ZN(
        n18017) );
  NOR2_X4 U11650 ( .A1(n20535), .A2(n21183), .ZN(n17221) );
  NAND2_X2 U11651 ( .A1(n11441), .A2(n11440), .ZN(n16772) );
  NOR2_X1 U11652 ( .A1(n21633), .A2(n21173), .ZN(n11213) );
  AND2_X4 U11653 ( .A1(n14724), .A2(n11741), .ZN(n11214) );
  OAI21_X2 U11654 ( .B1(n16752), .B2(n16753), .A(n16754), .ZN(n16745) );
  NOR2_X2 U11655 ( .A1(n21208), .A2(n21582), .ZN(n21491) );
  NAND2_X2 U11656 ( .A1(n21603), .A2(n21611), .ZN(n21582) );
  NOR2_X1 U11657 ( .A1(n21183), .A2(n17191), .ZN(n11215) );
  NAND2_X1 U11658 ( .A1(n12941), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13018) );
  AND3_X1 U11659 ( .A1(n12934), .A2(n14886), .A3(n12933), .ZN(n12939) );
  INV_X1 U11660 ( .A(n15524), .ZN(n13247) );
  XNOR2_X1 U11661 ( .A(n12986), .B(n13009), .ZN(n14847) );
  OAI21_X1 U11662 ( .B1(n13018), .B2(n12981), .A(n12983), .ZN(n12986) );
  INV_X2 U11663 ( .A(n11937), .ZN(n12037) );
  XNOR2_X1 U11664 ( .A(n15632), .B(n13782), .ZN(n14294) );
  INV_X1 U11665 ( .A(n17438), .ZN(n11450) );
  NAND2_X1 U11666 ( .A1(n13761), .A2(n11866), .ZN(n11431) );
  AND2_X1 U11667 ( .A1(n17369), .A2(n12811), .ZN(n12945) );
  OR2_X1 U11668 ( .A1(n14636), .A2(n22253), .ZN(n13734) );
  NAND2_X1 U11669 ( .A1(n14684), .A2(n11533), .ZN(n14685) );
  NAND2_X1 U11670 ( .A1(n11534), .A2(n15841), .ZN(n11533) );
  INV_X1 U11671 ( .A(n14630), .ZN(n11534) );
  NAND2_X1 U11672 ( .A1(n11502), .A2(n14979), .ZN(n11501) );
  AND2_X1 U11673 ( .A1(n13014), .A2(n22122), .ZN(n11502) );
  NAND2_X1 U11674 ( .A1(n12985), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13009) );
  NOR2_X1 U11675 ( .A1(n12069), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12070) );
  AND2_X1 U11676 ( .A1(n12683), .A2(n16786), .ZN(n12684) );
  NOR2_X1 U11677 ( .A1(n17435), .A2(n11364), .ZN(n11363) );
  NAND2_X1 U11678 ( .A1(n11645), .A2(n11269), .ZN(n11362) );
  AND2_X1 U11679 ( .A1(n11253), .A2(n12789), .ZN(n11365) );
  INV_X1 U11680 ( .A(n15614), .ZN(n12394) );
  AND2_X1 U11681 ( .A1(n11664), .A2(n11444), .ZN(n11443) );
  NAND2_X1 U11682 ( .A1(n11448), .A2(n11446), .ZN(n11444) );
  NOR2_X1 U11683 ( .A1(n11665), .A2(n16880), .ZN(n11664) );
  INV_X1 U11684 ( .A(n11666), .ZN(n11665) );
  AOI21_X1 U11685 ( .B1(n14499), .B2(n11466), .A(n11465), .ZN(n11464) );
  INV_X1 U11686 ( .A(n14496), .ZN(n11465) );
  OAI21_X1 U11687 ( .B1(n12775), .B2(n12776), .A(n15642), .ZN(n11378) );
  OR2_X1 U11688 ( .A1(n12092), .A2(n12091), .ZN(n12608) );
  NAND2_X1 U11689 ( .A1(n11949), .A2(n11947), .ZN(n12458) );
  NAND2_X1 U11690 ( .A1(n11587), .A2(n13771), .ZN(n13774) );
  NAND2_X1 U11691 ( .A1(n12484), .A2(n13781), .ZN(n11587) );
  NAND2_X1 U11692 ( .A1(n13756), .A2(n14730), .ZN(n12477) );
  NOR2_X1 U11693 ( .A1(n21208), .A2(n17289), .ZN(n17299) );
  INV_X1 U11694 ( .A(n21221), .ZN(n17285) );
  OR2_X1 U11695 ( .A1(n12916), .A2(n12919), .ZN(n12922) );
  AND4_X1 U11696 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n12870), .ZN(
        n12889) );
  NOR2_X1 U11697 ( .A1(n11263), .A2(n11330), .ZN(n11329) );
  OAI21_X1 U11698 ( .B1(n13181), .B2(n16433), .A(n13169), .ZN(n16284) );
  AND2_X1 U11699 ( .A1(n16284), .A2(n16283), .ZN(n16294) );
  NAND2_X1 U11700 ( .A1(n13064), .A2(n13063), .ZN(n14988) );
  NOR2_X1 U11701 ( .A1(n11173), .A2(n11284), .ZN(n16000) );
  AND2_X1 U11702 ( .A1(n11306), .A2(n11634), .ZN(n11633) );
  INV_X1 U11703 ( .A(n16557), .ZN(n11634) );
  AOI21_X1 U11704 ( .B1(n18648), .B2(n13781), .A(n13780), .ZN(n14293) );
  NAND2_X1 U11705 ( .A1(n13777), .A2(n13776), .ZN(n15632) );
  NAND2_X1 U11706 ( .A1(n18352), .A2(n11415), .ZN(n11414) );
  OR2_X1 U11707 ( .A1(n18352), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11417) );
  NOR2_X1 U11708 ( .A1(n11416), .A2(n18318), .ZN(n11415) );
  XNOR2_X1 U11709 ( .A(n18076), .B(n11535), .ZN(n18471) );
  INV_X1 U11710 ( .A(n18077), .ZN(n11535) );
  OR2_X1 U11711 ( .A1(n21418), .A2(n21441), .ZN(n18347) );
  AND2_X1 U11712 ( .A1(n13058), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11499) );
  NOR2_X1 U11713 ( .A1(n13244), .A2(n15892), .ZN(n12869) );
  BUF_X4 U11714 ( .A(n12852), .Z(n13708) );
  NOR2_X1 U11715 ( .A1(n11583), .A2(n11308), .ZN(n11582) );
  NAND2_X1 U11716 ( .A1(n12564), .A2(n12426), .ZN(n11348) );
  AND2_X1 U11717 ( .A1(n11358), .A2(n11276), .ZN(n11359) );
  NAND2_X1 U11718 ( .A1(n11631), .A2(n16095), .ZN(n11630) );
  INV_X1 U11719 ( .A(n16087), .ZN(n11631) );
  AND2_X1 U11720 ( .A1(n13171), .A2(n11498), .ZN(n11497) );
  INV_X1 U11721 ( .A(n13178), .ZN(n11498) );
  NAND2_X1 U11722 ( .A1(n14650), .A2(n13008), .ZN(n13056) );
  NAND2_X1 U11723 ( .A1(n16348), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U11724 ( .A1(n11333), .A2(n16349), .ZN(n16300) );
  OR2_X1 U11725 ( .A1(n11497), .A2(n11496), .ZN(n11336) );
  INV_X1 U11726 ( .A(n13177), .ZN(n11496) );
  INV_X1 U11727 ( .A(n20373), .ZN(n13171) );
  NOR2_X1 U11728 ( .A1(n16149), .A2(n11521), .ZN(n11520) );
  INV_X1 U11729 ( .A(n16214), .ZN(n11521) );
  INV_X1 U11730 ( .A(n13139), .ZN(n11331) );
  INV_X1 U11731 ( .A(n14957), .ZN(n11525) );
  INV_X1 U11732 ( .A(n14947), .ZN(n14953) );
  AND2_X1 U11733 ( .A1(n14683), .A2(n14682), .ZN(n14686) );
  OAI21_X1 U11734 ( .B1(n15878), .B2(P1_EBX_REG_1__SCAN_IN), .A(n14594), .ZN(
        n14684) );
  INV_X1 U11735 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13019) );
  AND4_X2 U11736 ( .A1(n12868), .A2(n12867), .A3(n12866), .A4(n12865), .ZN(
        n14268) );
  AND4_X1 U11737 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n12853), .ZN(
        n12867) );
  AND4_X1 U11738 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12865) );
  OR2_X1 U11739 ( .A1(n14971), .A2(n14970), .ZN(n15519) );
  AND2_X1 U11740 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14597) );
  INV_X1 U11741 ( .A(n15830), .ZN(n15824) );
  NAND2_X1 U11742 ( .A1(n12710), .A2(n12704), .ZN(n11574) );
  INV_X1 U11743 ( .A(n12702), .ZN(n12443) );
  NOR2_X1 U11744 ( .A1(n16600), .A2(n15770), .ZN(n11617) );
  NAND2_X1 U11745 ( .A1(n11981), .A2(n11615), .ZN(n11614) );
  INV_X1 U11746 ( .A(n14932), .ZN(n11615) );
  NOR2_X1 U11747 ( .A1(n17453), .A2(n11555), .ZN(n11554) );
  INV_X1 U11748 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11555) );
  INV_X1 U11749 ( .A(n14613), .ZN(n11620) );
  NOR2_X1 U11750 ( .A1(n11455), .A2(n11454), .ZN(n11453) );
  OAI21_X1 U11751 ( .B1(n11455), .B2(n16829), .A(n11456), .ZN(n11452) );
  INV_X1 U11752 ( .A(n16828), .ZN(n11454) );
  INV_X1 U11753 ( .A(n14809), .ZN(n11981) );
  INV_X1 U11754 ( .A(n11363), .ZN(n11360) );
  NAND2_X1 U11755 ( .A1(n11297), .A2(n11450), .ZN(n11446) );
  XNOR2_X1 U11756 ( .A(n12784), .B(n16849), .ZN(n12785) );
  XNOR2_X1 U11757 ( .A(n11352), .B(n12770), .ZN(n11639) );
  INV_X1 U11758 ( .A(n12563), .ZN(n12530) );
  AND2_X1 U11759 ( .A1(n11940), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U11760 ( .A1(n11892), .A2(n14921), .ZN(n11374) );
  NAND2_X1 U11761 ( .A1(n14350), .A2(n14352), .ZN(n11375) );
  NAND2_X1 U11762 ( .A1(n13756), .A2(n13781), .ZN(n13760) );
  NAND2_X1 U11763 ( .A1(n11837), .A2(n11261), .ZN(n11859) );
  AOI22_X1 U11764 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11838) );
  AOI21_X1 U11765 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19563), .A(
        n12056), .ZN(n12052) );
  NAND2_X1 U11766 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21191), .ZN(
        n17192) );
  NOR2_X1 U11767 ( .A1(n20535), .A2(n21194), .ZN(n18015) );
  NOR2_X1 U11768 ( .A1(n11419), .A2(n11422), .ZN(n11418) );
  INV_X1 U11769 ( .A(n11420), .ZN(n11419) );
  NAND2_X1 U11770 ( .A1(n11686), .A2(n11412), .ZN(n11411) );
  NOR2_X1 U11771 ( .A1(n18232), .A2(n20877), .ZN(n11412) );
  AND2_X1 U11772 ( .A1(n21390), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11539) );
  NOR2_X1 U11773 ( .A1(n20997), .A2(n20970), .ZN(n17290) );
  OR2_X1 U11774 ( .A1(n21002), .A2(n18079), .ZN(n18082) );
  AND2_X1 U11775 ( .A1(n18086), .A2(n18089), .ZN(n11549) );
  INV_X1 U11776 ( .A(n18125), .ZN(n11383) );
  NAND2_X1 U11777 ( .A1(n11390), .A2(n11389), .ZN(n18108) );
  NAND2_X1 U11778 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U11779 ( .A1(n11504), .A2(n17288), .ZN(n17294) );
  INV_X1 U11780 ( .A(n13159), .ZN(n11491) );
  AND2_X1 U11781 ( .A1(n15696), .A2(n11489), .ZN(n11488) );
  NAND2_X1 U11782 ( .A1(n11490), .A2(n13159), .ZN(n11489) );
  INV_X1 U11783 ( .A(n20347), .ZN(n11490) );
  NAND2_X1 U11784 ( .A1(n13300), .A2(n13299), .ZN(n15109) );
  OAI21_X1 U11785 ( .B1(n14971), .B2(n13398), .A(n13269), .ZN(n14585) );
  OR2_X1 U11786 ( .A1(n15684), .A2(n15683), .ZN(n15690) );
  NAND2_X1 U11787 ( .A1(n20348), .A2(n20347), .ZN(n20346) );
  INV_X1 U11788 ( .A(n15892), .ZN(n15837) );
  NAND2_X1 U11789 ( .A1(n12987), .A2(n12988), .ZN(n14979) );
  NAND2_X1 U11790 ( .A1(n11501), .A2(n13000), .ZN(n13261) );
  OAI21_X1 U11791 ( .B1(n16514), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13035), 
        .ZN(n13046) );
  NAND2_X1 U11792 ( .A1(n13046), .A2(n13045), .ZN(n13076) );
  INV_X1 U11793 ( .A(n13265), .ZN(n13045) );
  INV_X1 U11794 ( .A(n13075), .ZN(n11338) );
  AND2_X1 U11795 ( .A1(n15892), .A2(n14636), .ZN(n12846) );
  NAND2_X1 U11796 ( .A1(n11255), .A2(n13058), .ZN(n17363) );
  AND2_X1 U11797 ( .A1(n22356), .A2(n22632), .ZN(n22314) );
  INV_X1 U11798 ( .A(n22632), .ZN(n22285) );
  NOR2_X1 U11799 ( .A1(n22325), .A2(n22285), .ZN(n22362) );
  NOR2_X1 U11800 ( .A1(n14971), .A2(n16503), .ZN(n15027) );
  AND2_X1 U11801 ( .A1(n11561), .A2(n11164), .ZN(n11558) );
  NAND2_X1 U11802 ( .A1(n18917), .A2(n11564), .ZN(n11563) );
  INV_X1 U11803 ( .A(n18908), .ZN(n11564) );
  AND2_X1 U11804 ( .A1(n12002), .A2(n12001), .ZN(n15714) );
  NAND2_X1 U11805 ( .A1(n11252), .A2(n15578), .ZN(n15713) );
  INV_X1 U11806 ( .A(n11460), .ZN(n11459) );
  NAND2_X1 U11807 ( .A1(n16010), .A2(n11607), .ZN(n11606) );
  INV_X1 U11808 ( .A(n12796), .ZN(n11607) );
  NAND2_X1 U11809 ( .A1(n11605), .A2(n11604), .ZN(n11603) );
  INV_X1 U11810 ( .A(n16546), .ZN(n11604) );
  INV_X1 U11811 ( .A(n16016), .ZN(n11605) );
  NOR3_X1 U11812 ( .A1(n16543), .A2(n16546), .A3(n12796), .ZN(n16011) );
  OR2_X1 U11813 ( .A1(n16543), .A2(n16546), .ZN(n16544) );
  AND2_X1 U11814 ( .A1(n11995), .A2(n11994), .ZN(n15553) );
  XNOR2_X1 U11815 ( .A(n12787), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17435) );
  NAND2_X1 U11816 ( .A1(n12788), .A2(n11468), .ZN(n12787) );
  AND2_X1 U11817 ( .A1(n14572), .A2(n11288), .ZN(n14615) );
  NOR2_X1 U11818 ( .A1(n16849), .A2(n15965), .ZN(n11571) );
  AOI21_X1 U11819 ( .B1(n15964), .B2(n11468), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U11820 ( .A1(n18944), .A2(n16849), .ZN(n16704) );
  NAND2_X1 U11821 ( .A1(n12695), .A2(n17012), .ZN(n12698) );
  INV_X1 U11822 ( .A(n15720), .ZN(n11478) );
  NOR2_X1 U11823 ( .A1(n17004), .A2(n17018), .ZN(n11380) );
  NOR2_X1 U11824 ( .A1(n16860), .A2(n17004), .ZN(n16832) );
  INV_X1 U11825 ( .A(n16797), .ZN(n16885) );
  NAND2_X1 U11826 ( .A1(n11468), .A2(n11467), .ZN(n11466) );
  NAND2_X1 U11827 ( .A1(n11462), .A2(n11464), .ZN(n14582) );
  NAND2_X1 U11828 ( .A1(n11351), .A2(n12594), .ZN(n15740) );
  INV_X1 U11829 ( .A(n12780), .ZN(n12781) );
  AOI21_X1 U11830 ( .B1(n11467), .B2(n12608), .A(n12224), .ZN(n14498) );
  AND2_X1 U11831 ( .A1(n12226), .A2(n12225), .ZN(n14499) );
  INV_X1 U11832 ( .A(n11946), .ZN(n11943) );
  INV_X1 U11833 ( .A(n11945), .ZN(n11944) );
  OR2_X1 U11834 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  AOI21_X1 U11835 ( .B1(n14294), .B2(n14293), .A(n13784), .ZN(n14416) );
  NOR2_X1 U11836 ( .A1(n11874), .A2(n11877), .ZN(n11880) );
  NOR2_X1 U11837 ( .A1(n19660), .A2(n19642), .ZN(n19695) );
  NAND2_X1 U11838 ( .A1(n19715), .A2(n19708), .ZN(n19648) );
  NAND2_X1 U11839 ( .A1(n19660), .A2(n19642), .ZN(n19552) );
  INV_X1 U11840 ( .A(n19715), .ZN(n20005) );
  INV_X1 U11841 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19593) );
  AOI21_X1 U11842 ( .B1(n20932), .B2(n11402), .A(n11401), .ZN(n11400) );
  INV_X1 U11843 ( .A(n20919), .ZN(n11401) );
  INV_X1 U11844 ( .A(n20908), .ZN(n11402) );
  NOR2_X1 U11845 ( .A1(n17299), .A2(n21163), .ZN(n20972) );
  NOR2_X1 U11846 ( .A1(n11278), .A2(n20901), .ZN(n18352) );
  INV_X1 U11847 ( .A(n18280), .ZN(n18319) );
  NAND2_X1 U11848 ( .A1(n18276), .A2(n21425), .ZN(n21418) );
  NAND2_X1 U11849 ( .A1(n18369), .A2(n21505), .ZN(n18258) );
  AOI21_X1 U11850 ( .B1(n18078), .B2(n21293), .A(n11368), .ZN(n11366) );
  INV_X1 U11851 ( .A(n18078), .ZN(n11367) );
  INV_X1 U11852 ( .A(n18462), .ZN(n11368) );
  NAND2_X1 U11853 ( .A1(n18471), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18470) );
  NAND2_X1 U11854 ( .A1(n18525), .A2(n18518), .ZN(n18517) );
  INV_X1 U11855 ( .A(n21184), .ZN(n20541) );
  INV_X1 U11856 ( .A(n21167), .ZN(n21187) );
  OAI22_X1 U11857 ( .A1(n21658), .A2(n21650), .B1(n21219), .B2(n21579), .ZN(
        n21630) );
  OR2_X1 U11858 ( .A1(n13749), .A2(n16289), .ZN(n13751) );
  XNOR2_X1 U11859 ( .A(n13744), .B(n13743), .ZN(n16044) );
  INV_X1 U11860 ( .A(n16407), .ZN(n20388) );
  INV_X1 U11861 ( .A(n20379), .ZN(n20395) );
  AND2_X1 U11862 ( .A1(n13745), .A2(n22292), .ZN(n20385) );
  AND2_X1 U11863 ( .A1(n14305), .A2(n17399), .ZN(n20392) );
  INV_X1 U11864 ( .A(n11484), .ZN(n11483) );
  AOI21_X1 U11865 ( .B1(n11484), .B2(n11280), .A(n11482), .ZN(n11481) );
  NAND2_X1 U11866 ( .A1(n14979), .A2(n13014), .ZN(n22339) );
  OR2_X1 U11867 ( .A1(n22275), .A2(n22274), .ZN(n22577) );
  NAND2_X1 U11868 ( .A1(n11560), .A2(n11164), .ZN(n18918) );
  OR2_X1 U11869 ( .A1(n18906), .A2(n18908), .ZN(n11560) );
  OR2_X1 U11870 ( .A1(n18906), .A2(n11563), .ZN(n11559) );
  OR2_X1 U11871 ( .A1(n11164), .A2(n11562), .ZN(n11561) );
  AND2_X1 U11872 ( .A1(n14122), .A2(n18631), .ZN(n16571) );
  INV_X1 U11873 ( .A(n19642), .ZN(n17481) );
  INV_X1 U11874 ( .A(n17477), .ZN(n19550) );
  OR2_X1 U11875 ( .A1(n16558), .A2(n16553), .ZN(n18924) );
  NAND2_X1 U11876 ( .A1(n16841), .A2(n17055), .ZN(n11345) );
  NOR2_X1 U11877 ( .A1(n16832), .A2(n17446), .ZN(n11344) );
  NAND2_X1 U11878 ( .A1(n14378), .A2(n14760), .ZN(n19015) );
  INV_X1 U11879 ( .A(n19694), .ZN(n19708) );
  INV_X1 U11880 ( .A(n20069), .ZN(n20079) );
  NOR2_X1 U11881 ( .A1(n19623), .A2(n19675), .ZN(n20069) );
  AOI21_X1 U11882 ( .B1(n20932), .B2(n11405), .A(n18138), .ZN(n11404) );
  INV_X1 U11883 ( .A(n20771), .ZN(n11405) );
  NAND2_X1 U11884 ( .A1(n20772), .A2(n20771), .ZN(n20782) );
  CLKBUF_X1 U11885 ( .A(n20792), .Z(n20934) );
  INV_X1 U11886 ( .A(n11393), .ZN(n11392) );
  OAI21_X1 U11887 ( .B1(n21475), .B2(n18388), .A(n11394), .ZN(n11393) );
  NAND2_X1 U11888 ( .A1(n18360), .A2(n18343), .ZN(n11394) );
  NAND2_X1 U11889 ( .A1(n18341), .A2(n21468), .ZN(n11395) );
  NOR2_X1 U11890 ( .A1(n18337), .A2(n11516), .ZN(n18284) );
  NAND2_X1 U11891 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11517), .ZN(
        n11516) );
  INV_X1 U11892 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11517) );
  NOR3_X2 U11893 ( .A1(P3_STATEBS16_REG_SCAN_IN), .A2(n18515), .A3(n21158), 
        .ZN(n18360) );
  AND2_X1 U11894 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18489) );
  AOI21_X2 U11895 ( .B1(n20467), .B2(n21688), .A(n21692), .ZN(n18515) );
  NOR2_X2 U11896 ( .A1(n18216), .A2(n18360), .ZN(n18513) );
  AND2_X1 U11897 ( .A1(n21500), .A2(n11545), .ZN(n11544) );
  OR2_X1 U11898 ( .A1(n21499), .A2(n21556), .ZN(n21500) );
  OAI21_X1 U11899 ( .B1(n22528), .B2(n14467), .A(n14881), .ZN(n13221) );
  AOI22_X1 U11900 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n12538), .B1(
        n12539), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12540) );
  NOR2_X1 U11901 ( .A1(n11912), .A2(n11739), .ZN(n11357) );
  AOI22_X1 U11902 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11820) );
  CLKBUF_X1 U11903 ( .A(n13358), .Z(n13711) );
  AND2_X1 U11904 ( .A1(n15679), .A2(n15763), .ZN(n11609) );
  CLKBUF_X2 U11905 ( .A(n13088), .Z(n13717) );
  NAND2_X1 U11906 ( .A1(n13120), .A2(n13119), .ZN(n13140) );
  AOI21_X1 U11907 ( .B1(n13358), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11500), .ZN(n12812) );
  AND2_X1 U11908 ( .A1(n11255), .A2(n11499), .ZN(n11500) );
  INV_X1 U11909 ( .A(n13911), .ZN(n13894) );
  INV_X1 U11910 ( .A(n13912), .ZN(n13896) );
  NOR2_X1 U11911 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13938) );
  INV_X1 U11912 ( .A(n12621), .ZN(n12437) );
  NAND3_X1 U11913 ( .A1(n12788), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n11468), .ZN(n12789) );
  INV_X1 U11914 ( .A(n16779), .ZN(n11456) );
  NAND2_X1 U11915 ( .A1(n16807), .A2(n16820), .ZN(n11455) );
  NAND2_X1 U11916 ( .A1(n14498), .A2(n11466), .ZN(n11462) );
  INV_X1 U11917 ( .A(n12777), .ZN(n12613) );
  INV_X1 U11918 ( .A(n12614), .ZN(n11340) );
  NAND2_X1 U11919 ( .A1(n12614), .A2(n12777), .ZN(n11668) );
  AOI22_X1 U11920 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12548), .B1(
        n19585), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12524) );
  AND2_X1 U11921 ( .A1(n12533), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12517) );
  AOI22_X1 U11922 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19615), .B1(
        n12549), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12523) );
  INV_X1 U11923 ( .A(n14318), .ZN(n14316) );
  XNOR2_X1 U11924 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12053) );
  AND2_X1 U11925 ( .A1(n12054), .A2(n12053), .ZN(n12056) );
  NOR2_X1 U11926 ( .A1(n18108), .A2(n21015), .ZN(n18054) );
  AND2_X1 U11927 ( .A1(n18099), .A2(n18054), .ZN(n18075) );
  NOR2_X1 U11928 ( .A1(n11507), .A2(n20529), .ZN(n17291) );
  INV_X1 U11929 ( .A(n14471), .ZN(n12919) );
  AND2_X1 U11930 ( .A1(n13190), .A2(n13220), .ZN(n13238) );
  AND2_X1 U11931 ( .A1(n13201), .A2(n13228), .ZN(n14262) );
  NAND2_X1 U11932 ( .A1(n12888), .A2(n12887), .ZN(n11330) );
  AND4_X1 U11933 ( .A1(n12886), .A2(n12885), .A3(n12884), .A4(n12883), .ZN(
        n12887) );
  AND4_X1 U11934 ( .A1(n12878), .A2(n12877), .A3(n12876), .A4(n12875), .ZN(
        n12888) );
  NOR2_X1 U11935 ( .A1(n11632), .A2(n11630), .ZN(n11629) );
  INV_X1 U11936 ( .A(n16074), .ZN(n11632) );
  AND2_X1 U11937 ( .A1(n11625), .A2(n11624), .ZN(n11623) );
  INV_X1 U11938 ( .A(n16173), .ZN(n11624) );
  AND2_X1 U11939 ( .A1(n16355), .A2(n16186), .ZN(n11625) );
  OR2_X1 U11940 ( .A1(n11609), .A2(n11610), .ZN(n11608) );
  AND2_X1 U11941 ( .A1(n15679), .A2(n16144), .ZN(n11610) );
  XNOR2_X1 U11942 ( .A(n13162), .B(n13152), .ZN(n13305) );
  NAND2_X1 U11943 ( .A1(n13005), .A2(n13004), .ZN(n13006) );
  NAND2_X1 U11944 ( .A1(n11501), .A2(n11225), .ZN(n13005) );
  AND2_X1 U11945 ( .A1(n11530), .A2(n11529), .ZN(n11528) );
  INV_X1 U11946 ( .A(n16181), .ZN(n11529) );
  AND2_X1 U11947 ( .A1(n20308), .A2(n16187), .ZN(n11530) );
  NAND2_X1 U11948 ( .A1(n14671), .A2(n13057), .ZN(n13082) );
  NOR2_X1 U11949 ( .A1(n22528), .A2(n22386), .ZN(n13190) );
  NAND2_X1 U11950 ( .A1(n15837), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13038) );
  OR2_X1 U11951 ( .A1(n12912), .A2(n12913), .ZN(n14459) );
  AOI21_X1 U11952 ( .B1(n17421), .B2(n14875), .A(n22129), .ZN(n14846) );
  INV_X1 U11953 ( .A(n12725), .ZN(n11584) );
  NOR2_X1 U11954 ( .A1(n11574), .A2(n11575), .ZN(n11573) );
  INV_X1 U11955 ( .A(n12717), .ZN(n11575) );
  INV_X1 U11956 ( .A(n12670), .ZN(n11580) );
  INV_X1 U11957 ( .A(n12644), .ZN(n11583) );
  NAND2_X1 U11958 ( .A1(n11581), .A2(n11582), .ZN(n12675) );
  NAND2_X1 U11959 ( .A1(n12635), .A2(n12636), .ZN(n12645) );
  AND2_X1 U11960 ( .A1(n12438), .A2(n12633), .ZN(n12635) );
  INV_X1 U11961 ( .A(n12634), .ZN(n12438) );
  NAND2_X1 U11962 ( .A1(n11570), .A2(n12630), .ZN(n12634) );
  INV_X1 U11963 ( .A(n12631), .ZN(n11570) );
  NAND2_X1 U11964 ( .A1(n12574), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12624) );
  CLKBUF_X1 U11965 ( .A(n13943), .Z(n14078) );
  CLKBUF_X1 U11966 ( .A(n13937), .Z(n14079) );
  CLKBUF_X1 U11967 ( .A(n13940), .Z(n14084) );
  OAI211_X1 U11968 ( .C1(n16539), .C2(n16552), .A(n16541), .B(n16549), .ZN(
        n14071) );
  NOR2_X1 U11969 ( .A1(n16559), .A2(n14016), .ZN(n14055) );
  AND2_X1 U11970 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  NOR2_X1 U11971 ( .A1(n11597), .A2(n11596), .ZN(n11595) );
  INV_X1 U11972 ( .A(n16587), .ZN(n11596) );
  INV_X1 U11973 ( .A(n13914), .ZN(n13877) );
  NAND2_X1 U11974 ( .A1(n11598), .A2(n13873), .ZN(n11597) );
  INV_X1 U11975 ( .A(n16595), .ZN(n11598) );
  INV_X1 U11976 ( .A(n15768), .ZN(n11590) );
  NAND2_X1 U11977 ( .A1(n13812), .A2(n11593), .ZN(n11592) );
  INV_X1 U11978 ( .A(n15716), .ZN(n11593) );
  OAI21_X1 U11979 ( .B1(n15617), .B2(n17511), .A(n19593), .ZN(n11460) );
  INV_X1 U11980 ( .A(n12784), .ZN(n12788) );
  NOR2_X1 U11981 ( .A1(n16624), .A2(n11477), .ZN(n11476) );
  NAND2_X1 U11982 ( .A1(n16608), .A2(n16628), .ZN(n11477) );
  OAI21_X1 U11983 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n16704), .ZN(n12729) );
  INV_X1 U11984 ( .A(n16570), .ZN(n11635) );
  AND2_X1 U11985 ( .A1(n16580), .A2(n16577), .ZN(n11636) );
  NOR2_X1 U11986 ( .A1(n11651), .A2(n16952), .ZN(n11649) );
  INV_X1 U11987 ( .A(n15063), .ZN(n11469) );
  AND2_X1 U11988 ( .A1(n11312), .A2(n17150), .ZN(n11666) );
  INV_X1 U11989 ( .A(n14583), .ZN(n11461) );
  NAND2_X1 U11990 ( .A1(n12614), .A2(n11346), .ZN(n12771) );
  NAND2_X1 U11991 ( .A1(n11641), .A2(n12508), .ZN(n12564) );
  OAI21_X1 U11992 ( .B1(n11643), .B2(n11642), .A(n12069), .ZN(n11641) );
  AOI22_X1 U11993 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U11994 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11782) );
  INV_X1 U11995 ( .A(n11354), .ZN(n12467) );
  NAND3_X1 U11996 ( .A1(n11892), .A2(n12609), .A3(n11889), .ZN(n14349) );
  NAND2_X1 U11997 ( .A1(n11803), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U11998 ( .A1(n11808), .A2(n14755), .ZN(n11809) );
  INV_X1 U11999 ( .A(n12485), .ZN(n12478) );
  NOR2_X1 U12000 ( .A1(n17306), .A2(n21165), .ZN(n17580) );
  INV_X1 U12001 ( .A(n11418), .ZN(n11416) );
  NOR2_X1 U12002 ( .A1(n20543), .A2(n11421), .ZN(n11420) );
  INV_X1 U12003 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11421) );
  NOR2_X1 U12004 ( .A1(n18227), .A2(n18232), .ZN(n18246) );
  NOR2_X1 U12005 ( .A1(n20758), .A2(n11408), .ZN(n11407) );
  NOR2_X1 U12006 ( .A1(n18095), .A2(n11427), .ZN(n11426) );
  NAND2_X1 U12007 ( .A1(n18094), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18095) );
  INV_X1 U12008 ( .A(n11429), .ZN(n11427) );
  INV_X1 U12009 ( .A(n18410), .ZN(n18094) );
  AND2_X1 U12010 ( .A1(n11426), .A2(n11428), .ZN(n20680) );
  NOR2_X1 U12011 ( .A1(n18472), .A2(n11430), .ZN(n11429) );
  INV_X1 U12012 ( .A(n20574), .ZN(n11428) );
  NAND2_X1 U12013 ( .A1(n18186), .A2(n11322), .ZN(n11538) );
  INV_X1 U12014 ( .A(n21525), .ZN(n11537) );
  OR2_X1 U12015 ( .A1(n18441), .A2(n18329), .ZN(n11369) );
  INV_X1 U12016 ( .A(n11369), .ZN(n18401) );
  INV_X1 U12017 ( .A(n18124), .ZN(n11386) );
  XNOR2_X1 U12018 ( .A(n18115), .B(n11388), .ZN(n18485) );
  INV_X1 U12019 ( .A(n18114), .ZN(n11388) );
  AND2_X1 U12020 ( .A1(n11272), .A2(n18108), .ZN(n18056) );
  NOR2_X1 U12021 ( .A1(n21153), .A2(n11505), .ZN(n17314) );
  NOR2_X1 U12022 ( .A1(n11507), .A2(n11506), .ZN(n11505) );
  OR2_X1 U12023 ( .A1(n11506), .A2(n17291), .ZN(n17310) );
  NAND2_X1 U12024 ( .A1(n17285), .A2(n21027), .ZN(n21166) );
  NAND2_X1 U12025 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21182) );
  NAND2_X1 U12026 ( .A1(n14467), .A2(n12977), .ZN(n12936) );
  AOI21_X1 U12027 ( .B1(n13286), .B2(n13463), .A(n13285), .ZN(n14716) );
  AND2_X1 U12028 ( .A1(n14870), .A2(n22161), .ZN(n20183) );
  INV_X1 U12029 ( .A(n14580), .ZN(n14521) );
  AND2_X1 U12030 ( .A1(n16094), .A2(n11626), .ZN(n16065) );
  AND2_X1 U12031 ( .A1(n11627), .A2(n11629), .ZN(n11626) );
  INV_X1 U12032 ( .A(n16066), .ZN(n11627) );
  INV_X1 U12033 ( .A(n11630), .ZN(n11628) );
  AND2_X1 U12034 ( .A1(n16183), .A2(n11621), .ZN(n20297) );
  AND2_X1 U12035 ( .A1(n11622), .A2(n11623), .ZN(n11621) );
  INV_X1 U12036 ( .A(n20295), .ZN(n11622) );
  NAND2_X1 U12037 ( .A1(n16183), .A2(n11623), .ZN(n20296) );
  NAND2_X1 U12038 ( .A1(n16183), .A2(n11625), .ZN(n16354) );
  NOR2_X1 U12039 ( .A1(n13487), .A2(n22027), .ZN(n13488) );
  AND2_X1 U12040 ( .A1(n13421), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13469) );
  AND2_X1 U12041 ( .A1(n13439), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13421) );
  AND2_X1 U12042 ( .A1(n13454), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13439) );
  AND2_X1 U12043 ( .A1(n13403), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13454) );
  INV_X1 U12044 ( .A(n15120), .ZN(n11586) );
  INV_X1 U12045 ( .A(n15109), .ZN(n11585) );
  NOR2_X1 U12046 ( .A1(n13289), .A2(n13288), .ZN(n13294) );
  NAND2_X1 U12047 ( .A1(n14674), .A2(n13272), .ZN(n14814) );
  AND2_X1 U12048 ( .A1(n13259), .A2(n13258), .ZN(n14484) );
  NOR2_X1 U12049 ( .A1(n13189), .A2(n11280), .ZN(n11480) );
  INV_X1 U12050 ( .A(n13188), .ZN(n11482) );
  AND2_X1 U12051 ( .A1(n13187), .A2(n13186), .ZN(n11484) );
  NOR2_X1 U12052 ( .A1(n11219), .A2(n16076), .ZN(n16075) );
  OR2_X1 U12053 ( .A1(n16172), .A2(n11522), .ZN(n11219) );
  OR3_X1 U12054 ( .A1(n16114), .A2(n16083), .A3(n11523), .ZN(n11522) );
  NAND2_X1 U12055 ( .A1(n16300), .A2(n16301), .ZN(n11332) );
  OR2_X1 U12056 ( .A1(n20299), .A2(n16170), .ZN(n16172) );
  NAND2_X1 U12057 ( .A1(n16175), .A2(n20300), .ZN(n20299) );
  NAND2_X1 U12058 ( .A1(n11495), .A2(n11496), .ZN(n11492) );
  AND2_X1 U12059 ( .A1(n16122), .A2(n11526), .ZN(n16477) );
  AND2_X1 U12060 ( .A1(n11528), .A2(n11527), .ZN(n11526) );
  INV_X1 U12061 ( .A(n16479), .ZN(n11527) );
  NAND2_X1 U12062 ( .A1(n16122), .A2(n11528), .ZN(n16478) );
  NAND2_X1 U12063 ( .A1(n16122), .A2(n11530), .ZN(n20311) );
  AND2_X1 U12064 ( .A1(n16122), .A2(n16187), .ZN(n20309) );
  NAND2_X1 U12065 ( .A1(n16388), .A2(n13171), .ZN(n16379) );
  OR2_X1 U12066 ( .A1(n13169), .A2(n21729), .ZN(n11335) );
  NOR2_X1 U12067 ( .A1(n11519), .A2(n16204), .ZN(n11518) );
  INV_X1 U12068 ( .A(n11520), .ZN(n11519) );
  NAND2_X1 U12069 ( .A1(n20287), .A2(n16214), .ZN(n16215) );
  NAND2_X1 U12070 ( .A1(n20287), .A2(n11520), .ZN(n16203) );
  BUF_X1 U12071 ( .A(n16388), .Z(n16389) );
  NAND2_X1 U12072 ( .A1(n11487), .A2(n11486), .ZN(n15731) );
  AOI21_X1 U12073 ( .B1(n11488), .B2(n11491), .A(n11265), .ZN(n11486) );
  AND2_X1 U12074 ( .A1(n11259), .A2(n15124), .ZN(n11524) );
  AND2_X1 U12075 ( .A1(n14953), .A2(n11259), .ZN(n15125) );
  AND2_X1 U12076 ( .A1(n14956), .A2(n14955), .ZN(n14957) );
  NAND2_X1 U12077 ( .A1(n20327), .A2(n13103), .ZN(n20335) );
  NAND2_X1 U12078 ( .A1(n14953), .A2(n11676), .ZN(n20316) );
  INV_X1 U12079 ( .A(n14685), .ZN(n11532) );
  XNOR2_X1 U12080 ( .A(n14684), .B(n14630), .ZN(n15558) );
  NAND2_X1 U12081 ( .A1(n13014), .A2(n13013), .ZN(n13023) );
  OAI211_X1 U12082 ( .C1(n15528), .C2(n13752), .A(n13021), .B(n13020), .ZN(
        n13022) );
  OR2_X1 U12083 ( .A1(n13059), .A2(n13019), .ZN(n13021) );
  INV_X1 U12084 ( .A(n14641), .ZN(n11337) );
  INV_X1 U12085 ( .A(n13076), .ZN(n13077) );
  OR2_X1 U12086 ( .A1(n14256), .A2(n12928), .ZN(n14476) );
  OR2_X2 U12087 ( .A1(n12845), .A2(n12844), .ZN(n15892) );
  OR2_X1 U12088 ( .A1(n15517), .A2(n14842), .ZN(n14972) );
  INV_X2 U12089 ( .A(n14459), .ZN(n15825) );
  OR2_X2 U12090 ( .A1(n12825), .A2(n12824), .ZN(n15524) );
  INV_X1 U12091 ( .A(n15519), .ZN(n15026) );
  NOR2_X1 U12092 ( .A1(n13253), .A2(n14641), .ZN(n15028) );
  AOI21_X1 U12093 ( .B1(n22251), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22285), 
        .ZN(n22268) );
  NAND2_X1 U12094 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15824), .ZN(n16509) );
  NAND2_X1 U12095 ( .A1(n12719), .A2(n11243), .ZN(n12728) );
  INV_X1 U12096 ( .A(n11557), .ZN(n11556) );
  AOI21_X1 U12097 ( .B1(n11558), .B2(n11563), .A(n18931), .ZN(n11557) );
  INV_X1 U12098 ( .A(n11574), .ZN(n11572) );
  NAND2_X1 U12099 ( .A1(n12703), .A2(n12704), .ZN(n12711) );
  NAND2_X1 U12100 ( .A1(n12646), .A2(n11311), .ZN(n12702) );
  NAND2_X1 U12101 ( .A1(n12646), .A2(n12647), .ZN(n12696) );
  NAND2_X1 U12102 ( .A1(n11708), .A2(n11233), .ZN(n11726) );
  NAND2_X1 U12103 ( .A1(n11432), .A2(n11933), .ZN(n11935) );
  INV_X1 U12104 ( .A(n11659), .ZN(n11432) );
  NAND2_X1 U12105 ( .A1(n16533), .A2(n16534), .ZN(n14073) );
  XNOR2_X1 U12106 ( .A(n14015), .B(n14014), .ZN(n16561) );
  XNOR2_X1 U12107 ( .A(n13997), .B(n13994), .ZN(n16566) );
  INV_X1 U12108 ( .A(n15551), .ZN(n11591) );
  NAND2_X1 U12109 ( .A1(n14662), .A2(n14708), .ZN(n14721) );
  CLKBUF_X1 U12110 ( .A(n14211), .Z(n15622) );
  NAND2_X1 U12111 ( .A1(n11700), .A2(n11242), .ZN(n11737) );
  AND2_X1 U12112 ( .A1(n11700), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11702) );
  NOR2_X1 U12113 ( .A1(n11734), .A2(n18885), .ZN(n11733) );
  NAND2_X1 U12114 ( .A1(n11566), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11734) );
  NOR2_X1 U12115 ( .A1(n16592), .A2(n16589), .ZN(n16588) );
  NAND2_X1 U12116 ( .A1(n15712), .A2(n11616), .ZN(n16592) );
  AND2_X1 U12117 ( .A1(n11286), .A2(n11618), .ZN(n11616) );
  INV_X1 U12118 ( .A(n16594), .ZN(n11618) );
  AND2_X1 U12119 ( .A1(n12011), .A2(n12010), .ZN(n16600) );
  NAND2_X1 U12120 ( .A1(n15712), .A2(n12006), .ZN(n16601) );
  NAND2_X1 U12121 ( .A1(n11435), .A2(n11433), .ZN(n16837) );
  NAND2_X1 U12122 ( .A1(n11438), .A2(n11434), .ZN(n11433) );
  INV_X1 U12123 ( .A(n16775), .ZN(n11434) );
  AND2_X1 U12124 ( .A1(n11708), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11725) );
  INV_X1 U12125 ( .A(n15553), .ZN(n11996) );
  AND2_X1 U12126 ( .A1(n11992), .A2(n11991), .ZN(n15097) );
  AND2_X1 U12127 ( .A1(n11613), .A2(n14940), .ZN(n11612) );
  INV_X1 U12128 ( .A(n11614), .ZN(n11613) );
  AND2_X1 U12129 ( .A1(n11986), .A2(n11985), .ZN(n14932) );
  NOR2_X1 U12130 ( .A1(n14710), .A2(n11614), .ZN(n14941) );
  AND2_X1 U12131 ( .A1(n11224), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11553) );
  AND2_X1 U12132 ( .A1(n11291), .A2(n14656), .ZN(n11619) );
  AND2_X1 U12133 ( .A1(n14572), .A2(n11291), .ZN(n14657) );
  INV_X1 U12134 ( .A(n12783), .ZN(n11341) );
  NAND2_X1 U12135 ( .A1(n11655), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11654) );
  INV_X1 U12136 ( .A(n15974), .ZN(n11655) );
  AND2_X1 U12137 ( .A1(n16640), .A2(n11472), .ZN(n16027) );
  AND2_X1 U12138 ( .A1(n11476), .A2(n11473), .ZN(n11472) );
  INV_X1 U12139 ( .A(n12420), .ZN(n11473) );
  NOR2_X1 U12140 ( .A1(n16624), .A2(n11475), .ZN(n11474) );
  INV_X1 U12141 ( .A(n16628), .ZN(n11475) );
  NAND2_X1 U12142 ( .A1(n16588), .A2(n11306), .ZN(n16568) );
  NAND2_X1 U12143 ( .A1(n18896), .A2(n11468), .ZN(n16746) );
  NAND2_X1 U12144 ( .A1(n16976), .A2(n16671), .ZN(n16673) );
  NOR2_X1 U12145 ( .A1(n16977), .A2(n16978), .ZN(n16976) );
  NAND2_X1 U12146 ( .A1(n18873), .A2(n11468), .ZN(n16764) );
  NOR2_X1 U12147 ( .A1(n11363), .A2(n11244), .ZN(n11361) );
  INV_X1 U12148 ( .A(n17003), .ZN(n12404) );
  INV_X1 U12149 ( .A(n17002), .ZN(n12405) );
  NAND2_X1 U12150 ( .A1(n11458), .A2(n11457), .ZN(n16977) );
  INV_X1 U12151 ( .A(n16682), .ZN(n11457) );
  NAND2_X1 U12152 ( .A1(n16783), .A2(n16782), .ZN(n16800) );
  OR2_X1 U12153 ( .A1(n18823), .A2(n12689), .ZN(n16828) );
  NAND2_X1 U12154 ( .A1(n12395), .A2(n12394), .ZN(n15719) );
  NOR2_X1 U12155 ( .A1(n14720), .A2(n11471), .ZN(n11470) );
  INV_X1 U12156 ( .A(n14708), .ZN(n11471) );
  NAND2_X1 U12157 ( .A1(n14662), .A2(n11282), .ZN(n15062) );
  AOI21_X1 U12158 ( .B1(n11443), .B2(n11445), .A(n11295), .ZN(n11440) );
  INV_X1 U12159 ( .A(n11446), .ZN(n11445) );
  NAND2_X1 U12160 ( .A1(n11611), .A2(n11981), .ZN(n14933) );
  AND2_X1 U12161 ( .A1(n12640), .A2(n17123), .ZN(n16880) );
  INV_X1 U12162 ( .A(n14709), .ZN(n11976) );
  NAND2_X1 U12163 ( .A1(n11442), .A2(n11446), .ZN(n17152) );
  NAND2_X1 U12164 ( .A1(n15777), .A2(n11447), .ZN(n11442) );
  AND2_X1 U12165 ( .A1(n19010), .A2(n15981), .ZN(n17156) );
  NAND2_X1 U12166 ( .A1(n14572), .A2(n14573), .ZN(n14614) );
  NAND2_X1 U12167 ( .A1(n12775), .A2(n12776), .ZN(n11377) );
  AND3_X1 U12168 ( .A1(n12206), .A2(n12205), .A3(n12204), .ZN(n14831) );
  AND2_X1 U12169 ( .A1(n14534), .A2(n11949), .ZN(n11589) );
  AND2_X1 U12170 ( .A1(n14378), .A2(n14758), .ZN(n17047) );
  CLKBUF_X1 U12171 ( .A(n12421), .Z(n12422) );
  XNOR2_X1 U12172 ( .A(n12141), .B(n12118), .ZN(n14406) );
  CLKBUF_X1 U12173 ( .A(n14373), .Z(n14374) );
  NAND2_X1 U12174 ( .A1(n13786), .A2(n13785), .ZN(n14696) );
  INV_X1 U12175 ( .A(n13766), .ZN(n14695) );
  OR2_X1 U12177 ( .A1(n19551), .A2(n19550), .ZN(n19633) );
  NAND2_X1 U12178 ( .A1(n11688), .A2(n11844), .ZN(n11851) );
  NOR3_X2 U12179 ( .A1(n15619), .A2(n22141), .A3(n19648), .ZN(n20011) );
  NOR3_X2 U12180 ( .A1(n22141), .A2(n15622), .A3(n19648), .ZN(n20010) );
  INV_X1 U12181 ( .A(n20011), .ZN(n19961) );
  NAND2_X1 U12182 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19715), .ZN(n20007) );
  NAND2_X1 U12183 ( .A1(n17307), .A2(n19211), .ZN(n11503) );
  AOI21_X1 U12184 ( .B1(n17304), .B2(n17303), .A(n17302), .ZN(n21656) );
  AOI211_X1 U12185 ( .C1(n11168), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17228), .B(n17227), .ZN(n17229) );
  NAND2_X1 U12186 ( .A1(n20529), .A2(n19425), .ZN(n20970) );
  INV_X1 U12187 ( .A(n20527), .ZN(n20479) );
  NAND2_X1 U12188 ( .A1(n18352), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18322) );
  NAND2_X1 U12189 ( .A1(n11410), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11409) );
  INV_X1 U12190 ( .A(n11411), .ZN(n11410) );
  NOR2_X1 U12191 ( .A1(n18227), .A2(n11411), .ZN(n18298) );
  NOR2_X1 U12192 ( .A1(n21233), .A2(n18251), .ZN(n18275) );
  NAND3_X1 U12193 ( .A1(n18188), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18227) );
  NAND2_X1 U12194 ( .A1(n18135), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18214) );
  NAND2_X1 U12195 ( .A1(n18379), .A2(n11235), .ZN(n18096) );
  NAND2_X1 U12196 ( .A1(n18379), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18146) );
  NOR2_X1 U12197 ( .A1(n18166), .A2(n20701), .ZN(n18379) );
  NAND2_X1 U12198 ( .A1(n11426), .A2(n11424), .ZN(n18166) );
  NOR2_X1 U12199 ( .A1(n20574), .A2(n11425), .ZN(n11424) );
  INV_X1 U12200 ( .A(n21343), .ZN(n18168) );
  NAND2_X1 U12201 ( .A1(n11428), .A2(n11429), .ZN(n18454) );
  NAND2_X1 U12202 ( .A1(n21490), .A2(n21491), .ZN(n21504) );
  INV_X1 U12203 ( .A(n18347), .ZN(n21499) );
  AOI21_X1 U12204 ( .B1(n21495), .B2(n21651), .A(n11546), .ZN(n11545) );
  INV_X1 U12205 ( .A(n21501), .ZN(n11546) );
  INV_X1 U12206 ( .A(n18287), .ZN(n18306) );
  NAND2_X1 U12207 ( .A1(n18186), .A2(n11539), .ZN(n18259) );
  NOR2_X1 U12208 ( .A1(n17335), .A2(n11512), .ZN(n17978) );
  OR2_X1 U12209 ( .A1(n11511), .A2(n17335), .ZN(n21188) );
  NAND2_X1 U12210 ( .A1(n21187), .A2(n11513), .ZN(n11511) );
  AOI21_X1 U12211 ( .B1(n18440), .B2(n11226), .A(n11296), .ZN(n11548) );
  AND2_X1 U12212 ( .A1(n18383), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21373) );
  NAND2_X1 U12213 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18168), .ZN(
        n18384) );
  NOR2_X1 U12214 ( .A1(n18384), .A2(n21372), .ZN(n18383) );
  NAND2_X1 U12215 ( .A1(n21557), .A2(n21356), .ZN(n21343) );
  NAND2_X1 U12216 ( .A1(n11384), .A2(n11382), .ZN(n21346) );
  NAND2_X1 U12217 ( .A1(n18434), .A2(n11307), .ZN(n11384) );
  NAND2_X1 U12218 ( .A1(n11383), .A2(n21356), .ZN(n11382) );
  AND2_X1 U12219 ( .A1(n11369), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21557) );
  NAND2_X1 U12220 ( .A1(n18433), .A2(n18125), .ZN(n21331) );
  AOI211_X1 U12221 ( .C1(n17901), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17281), .B(n17280), .ZN(n17282) );
  NAND2_X1 U12222 ( .A1(n18434), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18433) );
  OR2_X1 U12223 ( .A1(n21316), .A2(n21315), .ZN(n21328) );
  XNOR2_X1 U12224 ( .A(n18148), .B(n18083), .ZN(n18449) );
  NAND2_X1 U12225 ( .A1(n18463), .A2(n18120), .ZN(n18451) );
  XNOR2_X1 U12226 ( .A(n18119), .B(n11387), .ZN(n18464) );
  INV_X1 U12227 ( .A(n18118), .ZN(n11387) );
  NAND2_X1 U12228 ( .A1(n18464), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18463) );
  XNOR2_X1 U12229 ( .A(n18070), .B(n21274), .ZN(n18500) );
  INV_X1 U12230 ( .A(n18108), .ZN(n18071) );
  NAND2_X1 U12231 ( .A1(n18507), .A2(n18112), .ZN(n18496) );
  NAND2_X1 U12232 ( .A1(n18496), .A2(n18497), .ZN(n18495) );
  INV_X1 U12233 ( .A(n21579), .ZN(n21651) );
  INV_X1 U12234 ( .A(n21214), .ZN(n17975) );
  XNOR2_X1 U12235 ( .A(n18056), .B(n11370), .ZN(n18512) );
  INV_X1 U12236 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U12237 ( .A1(n18511), .A2(n18512), .ZN(n18510) );
  NOR2_X1 U12238 ( .A1(n19211), .A2(n11506), .ZN(n21214) );
  NAND2_X1 U12239 ( .A1(n21212), .A2(n21211), .ZN(n21208) );
  OR3_X1 U12240 ( .A1(n17261), .A2(n17260), .A3(n11508), .ZN(n21218) );
  NOR2_X1 U12241 ( .A1(n18067), .A2(n18066), .ZN(n18526) );
  XNOR2_X1 U12242 ( .A(n21145), .B(n11550), .ZN(n18518) );
  NOR2_X1 U12243 ( .A1(n17335), .A2(n11264), .ZN(n21163) );
  NOR2_X1 U12244 ( .A1(n11512), .A2(n17298), .ZN(n11510) );
  NOR2_X1 U12245 ( .A1(n17254), .A2(n17253), .ZN(n21221) );
  INV_X1 U12246 ( .A(n21218), .ZN(n21027) );
  NOR2_X1 U12247 ( .A1(n20231), .A2(n22011), .ZN(n22021) );
  INV_X1 U12248 ( .A(n22079), .ZN(n22100) );
  AND2_X1 U12249 ( .A1(n22050), .A2(n14880), .ZN(n22108) );
  INV_X1 U12250 ( .A(n22107), .ZN(n22096) );
  AND2_X1 U12251 ( .A1(n22050), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22061) );
  INV_X1 U12252 ( .A(n16219), .ZN(n20323) );
  INV_X1 U12253 ( .A(n16281), .ZN(n22379) );
  NAND2_X2 U12254 ( .A1(n14635), .A2(n15833), .ZN(n22375) );
  OR2_X1 U12255 ( .A1(n14634), .A2(n14633), .ZN(n14635) );
  INV_X1 U12256 ( .A(n22375), .ZN(n16279) );
  BUF_X1 U12257 ( .A(n20199), .Z(n20208) );
  CLKBUF_X1 U12258 ( .A(n20194), .Z(n21698) );
  CLKBUF_X1 U12259 ( .A(n14519), .Z(n14869) );
  NOR2_X1 U12260 ( .A1(n16183), .A2(n20307), .ZN(n22217) );
  AND2_X1 U12261 ( .A1(n16121), .A2(n16191), .ZN(n22214) );
  OR2_X1 U12262 ( .A1(n16194), .A2(n16119), .ZN(n16121) );
  AOI21_X1 U12263 ( .B1(n16133), .B2(n16132), .A(n16131), .ZN(n20367) );
  NAND2_X1 U12264 ( .A1(n20346), .A2(n13159), .ZN(n15697) );
  NAND2_X1 U12265 ( .A1(n11485), .A2(n11488), .ZN(n15695) );
  OR2_X1 U12266 ( .A1(n20348), .A2(n11491), .ZN(n11485) );
  CLKBUF_X1 U12267 ( .A(n14650), .Z(n21927) );
  INV_X1 U12268 ( .A(n14970), .ZN(n16503) );
  NAND2_X1 U12269 ( .A1(n13266), .A2(n13265), .ZN(n14971) );
  INV_X1 U12270 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22237) );
  CLKBUF_X1 U12271 ( .A(n14476), .Z(n17404) );
  OAI21_X1 U12272 ( .B1(n22286), .B2(n22666), .A(n22362), .ZN(n22668) );
  OAI211_X1 U12273 ( .C1(n22691), .C2(n22316), .A(n22315), .B(n22314), .ZN(
        n22694) );
  INV_X1 U12274 ( .A(n22729), .ZN(n22717) );
  AND2_X1 U12275 ( .A1(n15028), .A2(n14997), .ZN(n22733) );
  INV_X1 U12276 ( .A(n22417), .ZN(n22424) );
  INV_X1 U12277 ( .A(n22743), .ZN(n22232) );
  INV_X1 U12278 ( .A(n14984), .ZN(n22521) );
  INV_X1 U12279 ( .A(n22559), .ZN(n22566) );
  NAND2_X1 U12280 ( .A1(n15028), .A2(n15026), .ZN(n22747) );
  INV_X1 U12281 ( .A(n22722), .ZN(n22738) );
  INV_X1 U12282 ( .A(n15964), .ZN(n15966) );
  NAND2_X1 U12283 ( .A1(n12646), .A2(n11241), .ZN(n12681) );
  NAND2_X1 U12284 ( .A1(n11552), .A2(n18850), .ZN(n18849) );
  NAND2_X1 U12285 ( .A1(n12621), .A2(n12617), .ZN(n18688) );
  AND2_X1 U12286 ( .A1(n14221), .A2(n22141), .ZN(n18957) );
  OR2_X1 U12287 ( .A1(n12797), .A2(n16011), .ZN(n16536) );
  INV_X1 U12288 ( .A(n14808), .ZN(n11588) );
  INV_X1 U12289 ( .A(n19660), .ZN(n19573) );
  AND2_X1 U12290 ( .A1(n15623), .A2(n15619), .ZN(n19908) );
  INV_X1 U12291 ( .A(n19822), .ZN(n19912) );
  CLKBUF_X1 U12293 ( .A(n17530), .Z(n17542) );
  XNOR2_X1 U12294 ( .A(n11697), .B(n18974), .ZN(n16018) );
  INV_X1 U12295 ( .A(n11602), .ZN(n11601) );
  NOR3_X1 U12296 ( .A1(n16543), .A2(n11606), .A3(n11603), .ZN(n11599) );
  OAI21_X1 U12297 ( .B1(n11606), .B2(n16546), .A(n16016), .ZN(n11602) );
  XOR2_X1 U12298 ( .A(n16010), .B(n16011), .Z(n15977) );
  INV_X1 U12299 ( .A(n16536), .ZN(n18958) );
  INV_X1 U12300 ( .A(n18637), .ZN(n18992) );
  XNOR2_X1 U12301 ( .A(n16020), .B(n11698), .ZN(n16035) );
  NAND2_X1 U12302 ( .A1(n11653), .A2(n11652), .ZN(n16020) );
  NOR2_X1 U12303 ( .A1(n11654), .A2(n15965), .ZN(n11652) );
  XNOR2_X1 U12304 ( .A(n16007), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16008) );
  XNOR2_X1 U12305 ( .A(n15963), .B(n11682), .ZN(n16901) );
  AND2_X1 U12306 ( .A1(n12395), .A2(n11289), .ZN(n17031) );
  NAND2_X1 U12307 ( .A1(n17147), .A2(n11379), .ZN(n17447) );
  NAND2_X1 U12308 ( .A1(n16885), .A2(n16884), .ZN(n11379) );
  NAND2_X1 U12309 ( .A1(n11463), .A2(n11466), .ZN(n14497) );
  OR2_X1 U12310 ( .A1(n14498), .A2(n14499), .ZN(n11463) );
  NAND2_X1 U12311 ( .A1(n11192), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11648) );
  CLKBUF_X1 U12312 ( .A(n15740), .Z(n15741) );
  AND2_X1 U12313 ( .A1(n14378), .A2(n14357), .ZN(n17048) );
  INV_X1 U12314 ( .A(n17166), .ZN(n19024) );
  OR2_X1 U12315 ( .A1(n15632), .A2(n14253), .ZN(n17477) );
  INV_X1 U12316 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19592) );
  XNOR2_X1 U12317 ( .A(n14415), .B(n14417), .ZN(n19642) );
  AND2_X1 U12318 ( .A1(n14694), .A2(n14697), .ZN(n19660) );
  OR2_X1 U12319 ( .A1(n14696), .A2(n14695), .ZN(n14697) );
  INV_X1 U12320 ( .A(n20086), .ZN(n20088) );
  INV_X1 U12321 ( .A(n19751), .ZN(n20076) );
  OAI21_X1 U12322 ( .B1(n19620), .B2(n19619), .A(n19618), .ZN(n20070) );
  NOR2_X1 U12323 ( .A1(n19581), .A2(n19633), .ZN(n20055) );
  OAI21_X1 U12324 ( .B1(n15667), .B2(n15666), .A(n15665), .ZN(n20042) );
  INV_X1 U12325 ( .A(n19895), .ZN(n19900) );
  INV_X1 U12326 ( .A(n19818), .ZN(n19808) );
  INV_X1 U12327 ( .A(n20016), .ZN(n20027) );
  NOR2_X1 U12328 ( .A1(n19552), .A2(n19675), .ZN(n20016) );
  NOR2_X1 U12329 ( .A1(n19552), .A2(n19643), .ZN(n20109) );
  AND2_X1 U12330 ( .A1(n12749), .A2(n17476), .ZN(n19043) );
  CLKBUF_X1 U12331 ( .A(n17572), .Z(n17568) );
  AND2_X1 U12332 ( .A1(n20970), .A2(n17583), .ZN(n20462) );
  NAND2_X1 U12333 ( .A1(n11399), .A2(n11398), .ZN(n20947) );
  AOI21_X1 U12334 ( .B1(n11400), .B2(n20723), .A(n20723), .ZN(n11398) );
  NAND2_X1 U12335 ( .A1(n20917), .A2(n20932), .ZN(n20918) );
  NAND2_X1 U12336 ( .A1(n11397), .A2(n11400), .ZN(n20931) );
  OR2_X1 U12337 ( .A1(n20907), .A2(n20723), .ZN(n11397) );
  NAND2_X1 U12338 ( .A1(n20907), .A2(n20908), .ZN(n20917) );
  AOI21_X1 U12339 ( .B1(n20932), .B2(n20758), .A(n20757), .ZN(n20760) );
  INV_X1 U12340 ( .A(n20941), .ZN(n20900) );
  INV_X1 U12341 ( .A(n20912), .ZN(n20962) );
  NOR2_X1 U12342 ( .A1(n17583), .A2(n20969), .ZN(n17952) );
  INV_X1 U12343 ( .A(n21082), .ZN(n21078) );
  NOR2_X1 U12344 ( .A1(n21094), .A2(n21088), .ZN(n21087) );
  NOR2_X1 U12345 ( .A1(n21069), .A2(n21070), .ZN(n21095) );
  INV_X1 U12346 ( .A(n21100), .ZN(n21064) );
  NAND2_X1 U12347 ( .A1(n21064), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21069) );
  NOR3_X1 U12348 ( .A1(n21113), .A2(n21062), .A3(n21061), .ZN(n21107) );
  NOR2_X1 U12349 ( .A1(n21119), .A2(n21130), .ZN(n21114) );
  NOR2_X1 U12350 ( .A1(n17990), .A2(n17989), .ZN(n21002) );
  INV_X1 U12351 ( .A(n18098), .ZN(n21015) );
  OAI22_X1 U12352 ( .A1(n20972), .A2(n20971), .B1(n20970), .B2(n20969), .ZN(
        n21150) );
  INV_X1 U12353 ( .A(n21144), .ZN(n21147) );
  INV_X1 U12354 ( .A(n21018), .ZN(n21148) );
  CLKBUF_X1 U12355 ( .A(n18593), .Z(n21627) );
  CLKBUF_X1 U12356 ( .A(n18597), .Z(n18601) );
  CLKBUF_X1 U12357 ( .A(n20525), .Z(n20507) );
  CLKBUF_X1 U12358 ( .A(n20524), .Z(n20521) );
  NOR2_X1 U12359 ( .A1(n20472), .A2(n20971), .ZN(n20525) );
  NOR2_X1 U12360 ( .A1(n20507), .A2(n20479), .ZN(n20524) );
  INV_X1 U12361 ( .A(n18443), .ZN(n18389) );
  NAND2_X1 U12362 ( .A1(n18202), .A2(n11325), .ZN(n18337) );
  NOR2_X1 U12363 ( .A1(n21414), .A2(n21415), .ZN(n11515) );
  INV_X1 U12364 ( .A(n21414), .ZN(n11514) );
  NAND2_X1 U12365 ( .A1(n21580), .A2(n18252), .ZN(n21233) );
  NAND2_X1 U12366 ( .A1(n21373), .A2(n18252), .ZN(n21236) );
  NAND2_X1 U12367 ( .A1(n18202), .A2(n21390), .ZN(n18278) );
  NOR2_X1 U12368 ( .A1(n18432), .A2(n21224), .ZN(n18202) );
  OAI21_X1 U12369 ( .B1(n20543), .B2(n18320), .A(n19252), .ZN(n18280) );
  AND2_X1 U12370 ( .A1(n18379), .A2(n11406), .ZN(n18135) );
  AND2_X1 U12371 ( .A1(n11235), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11406) );
  INV_X1 U12372 ( .A(n18360), .ZN(n18310) );
  INV_X1 U12373 ( .A(n21580), .ZN(n21377) );
  AOI22_X1 U12374 ( .A1(n21557), .A2(n18443), .B1(n18520), .B2(n21331), .ZN(
        n18432) );
  NOR2_X2 U12375 ( .A1(n21492), .A2(n18531), .ZN(n18444) );
  NAND2_X1 U12376 ( .A1(n18489), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20574) );
  INV_X1 U12377 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20553) );
  NAND2_X1 U12378 ( .A1(n20529), .A2(n21692), .ZN(n18532) );
  NAND2_X1 U12379 ( .A1(n21211), .A2(n21692), .ZN(n18531) );
  OR2_X1 U12380 ( .A1(n18347), .A2(n21476), .ZN(n18317) );
  INV_X1 U12381 ( .A(n21536), .ZN(n21556) );
  NAND2_X1 U12382 ( .A1(n18258), .A2(n18257), .ZN(n18264) );
  AND2_X1 U12383 ( .A1(n21378), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21580) );
  INV_X1 U12384 ( .A(n18383), .ZN(n21383) );
  NOR2_X2 U12385 ( .A1(n21163), .A2(n21168), .ZN(n21619) );
  NOR2_X1 U12386 ( .A1(n21658), .A2(n21225), .ZN(n21536) );
  NAND2_X1 U12387 ( .A1(n18470), .A2(n18078), .ZN(n18461) );
  NOR3_X2 U12388 ( .A1(n20462), .A2(n17976), .A3(n17975), .ZN(n21652) );
  INV_X1 U12389 ( .A(n21602), .ZN(n21470) );
  INV_X1 U12390 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21646) );
  CLKBUF_X1 U12391 ( .A(n19419), .Z(n19293) );
  AOI21_X1 U12392 ( .B1(n16044), .B2(n20385), .A(n13754), .ZN(n13755) );
  NAND2_X1 U12393 ( .A1(n11559), .A2(n11561), .ZN(n18929) );
  AND2_X1 U12394 ( .A1(n14532), .A2(n11234), .ZN(n14609) );
  OR2_X1 U12395 ( .A1(n17029), .A2(n17445), .ZN(n11373) );
  NAND2_X1 U12396 ( .A1(n11343), .A2(n11342), .ZN(P2_U2997) );
  AOI21_X1 U12397 ( .B1(n17046), .B2(n17462), .A(n16835), .ZN(n11342) );
  NAND2_X1 U12398 ( .A1(n11345), .A2(n11344), .ZN(n11343) );
  OR2_X1 U12399 ( .A1(n17029), .A2(n17166), .ZN(n11372) );
  NAND2_X1 U12400 ( .A1(n20782), .A2(n20932), .ZN(n20783) );
  OR2_X1 U12401 ( .A1(n11391), .A2(n18342), .ZN(P3_U2800) );
  OR2_X1 U12402 ( .A1(n18346), .A2(n21468), .ZN(n11396) );
  INV_X1 U12403 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18503) );
  NOR2_X1 U12404 ( .A1(n11257), .A2(n11541), .ZN(n11540) );
  NOR2_X1 U12405 ( .A1(n21620), .A2(n21511), .ZN(n11541) );
  NOR2_X1 U12406 ( .A1(n17191), .A2(n21194), .ZN(n17593) );
  BUF_X1 U12407 ( .A(n17593), .Z(n18044) );
  NAND2_X1 U12408 ( .A1(n12793), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16760) );
  NAND2_X1 U12409 ( .A1(n13796), .A2(n11216), .ZN(n14935) );
  NAND2_X1 U12410 ( .A1(n11362), .A2(n11361), .ZN(n16768) );
  INV_X1 U12411 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U12412 ( .A1(n14921), .A2(n11877), .ZN(n11923) );
  AND3_X1 U12413 ( .A1(n11270), .A2(n11551), .A3(n11227), .ZN(n21145) );
  INV_X1 U12414 ( .A(n21145), .ZN(n11389) );
  AND2_X1 U12415 ( .A1(n11304), .A2(n14936), .ZN(n11216) );
  AND4_X1 U12416 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11569), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11217) );
  AND2_X2 U12417 ( .A1(n13938), .A2(n12085), .ZN(n12101) );
  OR3_X1 U12418 ( .A1(n21182), .A2(n21181), .A3(n21190), .ZN(n11218) );
  NOR2_X1 U12419 ( .A1(n20535), .A2(n17192), .ZN(n17233) );
  AND2_X1 U12420 ( .A1(n12810), .A2(n12809), .ZN(n13390) );
  AND2_X1 U12421 ( .A1(n12809), .A2(n14598), .ZN(n12950) );
  AND3_X1 U12422 ( .A1(n12815), .A2(n12814), .A3(n11260), .ZN(n11220) );
  NAND2_X1 U12423 ( .A1(n16553), .A2(n16554), .ZN(n16543) );
  NAND2_X1 U12424 ( .A1(n16588), .A2(n11636), .ZN(n16567) );
  NAND2_X1 U12425 ( .A1(n15712), .A2(n11286), .ZN(n15804) );
  AND2_X1 U12426 ( .A1(n16852), .A2(n16868), .ZN(n11222) );
  AND3_X1 U12427 ( .A1(n11915), .A2(n11275), .A3(n11914), .ZN(n11223) );
  AND2_X1 U12428 ( .A1(n11554), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11224) );
  NOR2_X2 U12429 ( .A1(n17208), .A2(n17207), .ZN(n21212) );
  INV_X1 U12430 ( .A(n21212), .ZN(n11506) );
  AND2_X1 U12431 ( .A1(n15571), .A2(n15679), .ZN(n15680) );
  INV_X1 U12432 ( .A(n19211), .ZN(n21026) );
  NOR2_X1 U12433 ( .A1(n17198), .A2(n17197), .ZN(n19211) );
  AND2_X1 U12434 ( .A1(n13000), .A2(n14467), .ZN(n11225) );
  AND2_X1 U12435 ( .A1(n11549), .A2(n11283), .ZN(n11226) );
  AND4_X1 U12436 ( .A1(n18022), .A2(n18021), .A3(n18020), .A4(n18019), .ZN(
        n11227) );
  AND2_X1 U12437 ( .A1(n18202), .A2(n11324), .ZN(n11228) );
  AND2_X1 U12438 ( .A1(n13299), .A2(n11586), .ZN(n11229) );
  OR2_X1 U12439 ( .A1(n16764), .A2(n11663), .ZN(n11230) );
  AND2_X1 U12440 ( .A1(n11290), .A2(n12724), .ZN(n11231) );
  AND2_X1 U12441 ( .A1(n11222), .A2(n11438), .ZN(n11232) );
  NAND2_X1 U12443 ( .A1(n11720), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11714) );
  AND3_X1 U12444 ( .A1(n13306), .A2(n13300), .A3(n11229), .ZN(n15119) );
  NAND2_X1 U12445 ( .A1(n11720), .A2(n11224), .ZN(n11712) );
  AND2_X1 U12446 ( .A1(n11462), .A2(n11287), .ZN(n14581) );
  NOR2_X1 U12447 ( .A1(n15807), .A2(n11597), .ZN(n16586) );
  NAND2_X1 U12448 ( .A1(n11591), .A2(n13812), .ZN(n15575) );
  INV_X1 U12449 ( .A(n11718), .ZN(n11569) );
  AND2_X1 U12450 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11233) );
  NOR2_X1 U12451 ( .A1(n11735), .A2(n16729), .ZN(n11703) );
  AND2_X1 U12452 ( .A1(n14531), .A2(n11310), .ZN(n11234) );
  AND2_X1 U12453 ( .A1(n11407), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11235) );
  INV_X1 U12454 ( .A(n12561), .ZN(n11577) );
  AND2_X1 U12455 ( .A1(n11331), .A2(n13119), .ZN(n11236) );
  AND2_X1 U12456 ( .A1(n11289), .A2(n17030), .ZN(n11237) );
  AND2_X1 U12457 ( .A1(n11233), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11238) );
  AND2_X1 U12458 ( .A1(n11234), .A2(n14608), .ZN(n11239) );
  NAND2_X1 U12459 ( .A1(n14532), .A2(n14531), .ZN(n14525) );
  NAND2_X1 U12460 ( .A1(n11868), .A2(n14344), .ZN(n11240) );
  NAND2_X1 U12461 ( .A1(n11733), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11705) );
  AND2_X1 U12462 ( .A1(n12647), .A2(n11320), .ZN(n11241) );
  AND2_X1 U12463 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11242) );
  AND2_X1 U12464 ( .A1(n12720), .A2(n11584), .ZN(n11243) );
  NAND2_X1 U12465 ( .A1(n16961), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11244) );
  CLKBUF_X1 U12466 ( .A(n18018), .Z(n17934) );
  NAND2_X4 U12467 ( .A1(n13162), .A2(n13161), .ZN(n13169) );
  NOR2_X2 U12468 ( .A1(n18082), .A2(n21492), .ZN(n18329) );
  INV_X1 U12469 ( .A(n18329), .ZN(n21505) );
  INV_X1 U12470 ( .A(n12096), .ZN(n13892) );
  NAND2_X1 U12472 ( .A1(n11340), .A2(n12613), .ZN(n12784) );
  OR2_X1 U12473 ( .A1(n16198), .A2(n16197), .ZN(n11247) );
  AND2_X1 U12474 ( .A1(n11437), .A2(n11436), .ZN(n16847) );
  NAND2_X1 U12475 ( .A1(n16797), .A2(n16961), .ZN(n16792) );
  NOR2_X1 U12476 ( .A1(n20298), .A2(n20297), .ZN(n11248) );
  NAND2_X1 U12477 ( .A1(n11494), .A2(n13177), .ZN(n16356) );
  AND2_X1 U12478 ( .A1(n12793), .A2(n11649), .ZN(n16734) );
  AND2_X1 U12479 ( .A1(n12793), .A2(n11650), .ZN(n16743) );
  OR3_X1 U12480 ( .A1(n16172), .A2(n16114), .A3(n11523), .ZN(n11249) );
  NAND2_X1 U12481 ( .A1(n11375), .A2(n11374), .ZN(n11910) );
  OR2_X1 U12482 ( .A1(n14071), .A2(n14070), .ZN(n11250) );
  INV_X1 U12483 ( .A(n11869), .ZN(n12068) );
  NAND2_X1 U12484 ( .A1(n17290), .A2(n17580), .ZN(n11513) );
  OR2_X1 U12485 ( .A1(n13997), .A2(n13998), .ZN(n11251) );
  NAND2_X1 U12486 ( .A1(n17152), .A2(n17150), .ZN(n17134) );
  AND2_X1 U12487 ( .A1(n15095), .A2(n11996), .ZN(n11252) );
  NAND2_X1 U12488 ( .A1(n12786), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U12489 ( .A1(n12700), .A2(n12699), .ZN(n16763) );
  AND2_X1 U12490 ( .A1(n11676), .A2(n11525), .ZN(n11254) );
  AND3_X1 U12491 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U12492 ( .A1(n12703), .A2(n11572), .ZN(n11256) );
  AND2_X1 U12493 ( .A1(n16117), .A2(n13505), .ZN(n16183) );
  NOR3_X1 U12494 ( .A1(n21510), .A2(n21569), .A3(n21509), .ZN(n11257) );
  NOR2_X1 U12495 ( .A1(n16819), .A2(n16778), .ZN(n11258) );
  NAND2_X1 U12496 ( .A1(n18231), .A2(n18527), .ZN(n18320) );
  NOR2_X1 U12497 ( .A1(n16561), .A2(n16560), .ZN(n16559) );
  AND2_X1 U12498 ( .A1(n11254), .A2(n15114), .ZN(n11259) );
  NAND2_X1 U12499 ( .A1(n14295), .A2(n18992), .ZN(n12501) );
  OAI21_X1 U12500 ( .B1(n12771), .B2(n11468), .A(n18677), .ZN(n12593) );
  INV_X1 U12501 ( .A(n16860), .ZN(n11381) );
  NAND2_X1 U12502 ( .A1(n18637), .A2(n12475), .ZN(n12500) );
  INV_X1 U12503 ( .A(n12500), .ZN(n12469) );
  AND2_X1 U12504 ( .A1(n12813), .A2(n12812), .ZN(n11260) );
  AND2_X1 U12505 ( .A1(n11888), .A2(n11890), .ZN(n11261) );
  AND3_X1 U12506 ( .A1(n11788), .A2(n11787), .A3(n11786), .ZN(n11262) );
  NAND4_X1 U12507 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n11263) );
  INV_X1 U12508 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12073) );
  INV_X1 U12509 ( .A(n11513), .ZN(n11512) );
  AOI21_X1 U12510 ( .B1(n16830), .B2(n11453), .A(n11452), .ZN(n11451) );
  NOR2_X1 U12511 ( .A1(n18450), .A2(n21316), .ZN(n18121) );
  NAND2_X1 U12512 ( .A1(n21187), .A2(n11510), .ZN(n11264) );
  NAND2_X1 U12513 ( .A1(n20297), .A2(n16169), .ZN(n16106) );
  AND2_X1 U12514 ( .A1(n13167), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11265) );
  AND2_X1 U12515 ( .A1(n12510), .A2(n12509), .ZN(n11266) );
  AND2_X1 U12516 ( .A1(n11371), .A2(n12484), .ZN(n11267) );
  OR2_X1 U12517 ( .A1(n12645), .A2(n11583), .ZN(n11268) );
  NOR2_X1 U12518 ( .A1(n20997), .A2(n19295), .ZN(n17307) );
  AND2_X1 U12519 ( .A1(n16183), .A2(n16186), .ZN(n16184) );
  NAND2_X1 U12520 ( .A1(n15571), .A2(n11609), .ZN(n15762) );
  AND2_X1 U12521 ( .A1(n11644), .A2(n11365), .ZN(n11269) );
  NAND2_X1 U12522 ( .A1(n16837), .A2(n16836), .ZN(n16838) );
  AND2_X1 U12523 ( .A1(n18024), .A2(n18025), .ZN(n11270) );
  AND2_X1 U12524 ( .A1(n11644), .A2(n11253), .ZN(n11271) );
  NAND2_X1 U12525 ( .A1(n21020), .A2(n21145), .ZN(n11272) );
  AND2_X1 U12526 ( .A1(n15571), .A2(n11608), .ZN(n11273) );
  AND2_X1 U12527 ( .A1(n11854), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11274) );
  NAND2_X1 U12528 ( .A1(n11667), .A2(n18688), .ZN(n12618) );
  AND2_X1 U12529 ( .A1(n11359), .A2(n11356), .ZN(n11275) );
  AND2_X1 U12530 ( .A1(n11911), .A2(n19032), .ZN(n11276) );
  NAND2_X1 U12531 ( .A1(n18452), .A2(n18451), .ZN(n11277) );
  AND2_X1 U12532 ( .A1(n12065), .A2(n13762), .ZN(n11913) );
  INV_X1 U12533 ( .A(n11600), .ZN(n16034) );
  OR2_X1 U12534 ( .A1(n18227), .A2(n11409), .ZN(n11278) );
  AND2_X1 U12535 ( .A1(n13785), .A2(n13775), .ZN(n14415) );
  NOR2_X1 U12536 ( .A1(n11247), .A2(n16123), .ZN(n16122) );
  NOR2_X1 U12537 ( .A1(n15551), .A2(n11592), .ZN(n15715) );
  NOR2_X1 U12538 ( .A1(n11710), .A2(n11694), .ZN(n11711) );
  OR2_X1 U12539 ( .A1(n18933), .A2(n16849), .ZN(n11279) );
  NOR2_X1 U12540 ( .A1(n11718), .A2(n15946), .ZN(n11717) );
  AND2_X1 U12541 ( .A1(n11720), .A2(n11553), .ZN(n11713) );
  AND2_X1 U12542 ( .A1(n11720), .A2(n11554), .ZN(n11715) );
  NAND2_X1 U12543 ( .A1(n12989), .A2(n14847), .ZN(n13014) );
  AND2_X1 U12544 ( .A1(n13169), .A2(n16432), .ZN(n11280) );
  OR2_X1 U12545 ( .A1(n12583), .A2(n12433), .ZN(n11281) );
  AND2_X1 U12546 ( .A1(n11470), .A2(n14874), .ZN(n11282) );
  NAND2_X1 U12547 ( .A1(n18329), .A2(n21584), .ZN(n11283) );
  AND2_X1 U12548 ( .A1(n15119), .A2(n15572), .ZN(n15571) );
  AND2_X1 U12549 ( .A1(n16477), .A2(n16176), .ZN(n16175) );
  AND2_X1 U12550 ( .A1(n16588), .A2(n16580), .ZN(n16576) );
  NAND2_X1 U12551 ( .A1(n11585), .A2(n13306), .ZN(n15107) );
  AND2_X1 U12552 ( .A1(n15964), .A2(n11571), .ZN(n11284) );
  AND2_X1 U12553 ( .A1(n15712), .A2(n11617), .ZN(n11285) );
  AND2_X1 U12554 ( .A1(n11617), .A2(n15805), .ZN(n11286) );
  XNOR2_X1 U12555 ( .A(n12618), .B(n15787), .ZN(n15739) );
  OAI21_X1 U12556 ( .B1(n12775), .B2(n12776), .A(n11377), .ZN(n15638) );
  AND2_X1 U12557 ( .A1(n11464), .A2(n11461), .ZN(n11287) );
  AND2_X1 U12558 ( .A1(n11620), .A2(n14573), .ZN(n11288) );
  NOR2_X1 U12559 ( .A1(n14717), .A2(n14716), .ZN(n14718) );
  AND2_X1 U12560 ( .A1(n12394), .A2(n11478), .ZN(n11289) );
  AND2_X1 U12561 ( .A1(n11711), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11708) );
  AND2_X1 U12562 ( .A1(n12395), .A2(n11237), .ZN(n16690) );
  AND2_X1 U12563 ( .A1(n14624), .A2(n14661), .ZN(n14662) );
  AND2_X1 U12564 ( .A1(n16726), .A2(n16727), .ZN(n11290) );
  OAI21_X1 U12565 ( .B1(n16582), .B2(n16583), .A(n11679), .ZN(n16574) );
  AND2_X1 U12566 ( .A1(n11288), .A2(n14606), .ZN(n11291) );
  NAND2_X1 U12567 ( .A1(n17152), .A2(n11666), .ZN(n16877) );
  AND2_X1 U12568 ( .A1(n11582), .A2(n11580), .ZN(n11292) );
  AND2_X1 U12569 ( .A1(n11559), .A2(n11558), .ZN(n11293) );
  INV_X1 U12570 ( .A(n15712), .ZN(n15771) );
  NOR2_X1 U12571 ( .A1(n15713), .A2(n15714), .ZN(n15712) );
  NAND2_X1 U12572 ( .A1(n12405), .A2(n12404), .ZN(n17001) );
  INV_X1 U12573 ( .A(n17001), .ZN(n11458) );
  NAND2_X1 U12574 ( .A1(n11594), .A2(n13873), .ZN(n15806) );
  INV_X1 U12575 ( .A(n12426), .ZN(n12770) );
  OR2_X1 U12576 ( .A1(n12203), .A2(n12202), .ZN(n12426) );
  INV_X1 U12577 ( .A(n15770), .ZN(n12006) );
  NAND2_X1 U12578 ( .A1(n15767), .A2(n16599), .ZN(n15807) );
  XNOR2_X1 U12579 ( .A(n13761), .B(n11355), .ZN(n14325) );
  AND2_X1 U12580 ( .A1(n12559), .A2(n12609), .ZN(n11294) );
  NAND2_X1 U12581 ( .A1(n16879), .A2(n16878), .ZN(n11295) );
  AND2_X1 U12582 ( .A1(n16588), .A2(n11633), .ZN(n16553) );
  AND2_X1 U12583 ( .A1(n11283), .A2(n18329), .ZN(n11296) );
  NAND2_X1 U12584 ( .A1(n17437), .A2(n11449), .ZN(n11297) );
  INV_X1 U12585 ( .A(n11448), .ZN(n11447) );
  NAND2_X1 U12586 ( .A1(n11450), .A2(n15779), .ZN(n11448) );
  NAND2_X1 U12587 ( .A1(n14695), .A2(n14696), .ZN(n14694) );
  NAND2_X1 U12588 ( .A1(n12565), .A2(n12566), .ZN(n12583) );
  INV_X1 U12589 ( .A(n12583), .ZN(n11578) );
  AND2_X1 U12590 ( .A1(n11287), .A2(n14625), .ZN(n11298) );
  AND2_X1 U12591 ( .A1(n11237), .A2(n16691), .ZN(n11299) );
  AND2_X1 U12592 ( .A1(n11282), .A2(n11469), .ZN(n11300) );
  AND2_X1 U12593 ( .A1(n11238), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11301) );
  AND2_X1 U12594 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11302) );
  BUF_X1 U12595 ( .A(n12084), .Z(n14080) );
  NAND2_X1 U12596 ( .A1(n12070), .A2(n16004), .ZN(n12372) );
  INV_X1 U12597 ( .A(n12372), .ZN(n11467) );
  NAND2_X1 U12598 ( .A1(n14694), .A2(n13791), .ZN(n14532) );
  NOR2_X1 U12599 ( .A1(n14691), .A2(n14831), .ZN(n14832) );
  AND2_X1 U12600 ( .A1(n11708), .A2(n11238), .ZN(n11303) );
  INV_X1 U12601 ( .A(n16845), .ZN(n11438) );
  AND2_X1 U12602 ( .A1(n14713), .A2(n11588), .ZN(n11304) );
  AND2_X1 U12603 ( .A1(n14953), .A2(n11254), .ZN(n15113) );
  NOR2_X1 U12604 ( .A1(n11727), .A2(n16812), .ZN(n11728) );
  NOR2_X1 U12605 ( .A1(n14685), .A2(n14686), .ZN(n14817) );
  AND2_X1 U12606 ( .A1(n18379), .A2(n11407), .ZN(n11305) );
  AND2_X1 U12607 ( .A1(n11636), .A2(n11635), .ZN(n11306) );
  NAND2_X1 U12608 ( .A1(n13796), .A2(n14713), .ZN(n14712) );
  NOR2_X1 U12609 ( .A1(n18214), .A2(n18213), .ZN(n18188) );
  AND2_X1 U12610 ( .A1(n21356), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11307) );
  AND2_X1 U12611 ( .A1(n12574), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11308) );
  AND2_X1 U12612 ( .A1(n20287), .A2(n11518), .ZN(n16136) );
  NOR2_X1 U12613 ( .A1(n15099), .A2(n15100), .ZN(n11309) );
  NOR2_X1 U12614 ( .A1(n13794), .A2(n14570), .ZN(n11310) );
  INV_X1 U12615 ( .A(n11566), .ZN(n11731) );
  NOR2_X1 U12616 ( .A1(n11729), .A2(n16791), .ZN(n11566) );
  AND2_X1 U12617 ( .A1(n11241), .A2(n12680), .ZN(n11311) );
  NOR2_X1 U12618 ( .A1(n11705), .A2(n16739), .ZN(n11696) );
  NOR2_X1 U12619 ( .A1(n15096), .A2(n15097), .ZN(n15095) );
  NAND2_X1 U12620 ( .A1(n12642), .A2(n17140), .ZN(n11312) );
  OR2_X1 U12621 ( .A1(n11592), .A2(n11590), .ZN(n11313) );
  NAND2_X1 U12622 ( .A1(n11976), .A2(n11684), .ZN(n14710) );
  INV_X1 U12623 ( .A(n11686), .ZN(n11413) );
  AND2_X1 U12624 ( .A1(n14662), .A2(n11470), .ZN(n11314) );
  AND2_X1 U12625 ( .A1(n13796), .A2(n11304), .ZN(n11315) );
  AND2_X1 U12626 ( .A1(n11608), .A2(n15800), .ZN(n11316) );
  AND2_X1 U12627 ( .A1(n11216), .A2(n11309), .ZN(n11317) );
  AND2_X1 U12628 ( .A1(n11242), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11318) );
  INV_X1 U12629 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22122) );
  INV_X1 U12630 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11565) );
  NAND2_X1 U12631 ( .A1(n14636), .A2(n22528), .ZN(n11319) );
  OR2_X1 U12632 ( .A1(n16004), .A2(n12442), .ZN(n11320) );
  INV_X1 U12633 ( .A(n18917), .ZN(n11562) );
  OR3_X1 U12634 ( .A1(n18227), .A2(n11413), .A3(n18232), .ZN(n11321) );
  NAND2_X1 U12635 ( .A1(n11859), .A2(n11858), .ZN(n14774) );
  NAND2_X1 U12636 ( .A1(n18352), .A2(n11420), .ZN(n11423) );
  AND2_X1 U12637 ( .A1(n11539), .A2(n11537), .ZN(n11322) );
  AND2_X1 U12638 ( .A1(n11243), .A2(n12737), .ZN(n11323) );
  BUF_X1 U12639 ( .A(n11860), .Z(n19828) );
  NOR2_X1 U12640 ( .A1(n20574), .A2(n18472), .ZN(n18409) );
  NOR2_X1 U12641 ( .A1(n18013), .A2(n18012), .ZN(n21020) );
  INV_X1 U12642 ( .A(n21020), .ZN(n11390) );
  AND2_X1 U12643 ( .A1(n21390), .A2(n11514), .ZN(n11324) );
  AND2_X1 U12644 ( .A1(n21390), .A2(n11515), .ZN(n11325) );
  INV_X1 U12645 ( .A(n11651), .ZN(n11650) );
  NAND2_X1 U12646 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11651) );
  INV_X1 U12647 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11663) );
  AND2_X1 U12648 ( .A1(n11649), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11326) );
  INV_X1 U12649 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11550) );
  INV_X1 U12650 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11430) );
  INV_X1 U12651 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11408) );
  INV_X1 U12652 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11425) );
  INV_X1 U12653 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11422) );
  CLKBUF_X1 U12654 ( .A(n20959), .Z(n11327) );
  NOR4_X1 U12655 ( .A1(n11176), .A2(n20530), .A3(n20934), .A4(n21683), .ZN(
        n20959) );
  OR2_X1 U12656 ( .A1(n14846), .A2(n22126), .ZN(n22634) );
  OR3_X2 U12657 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), 
        .A3(n20463), .ZN(n21620) );
  NOR2_X1 U12658 ( .A1(n21655), .A2(n20470), .ZN(n20530) );
  NOR2_X1 U12659 ( .A1(n21627), .A2(n18584), .ZN(n18597) );
  OAI22_X2 U12660 ( .A1(n22390), .A2(n22640), .B1(n22639), .B2(n22389), .ZN(
        n22426) );
  OAI22_X2 U12661 ( .A1(n22384), .A2(n22640), .B1(n22639), .B2(n22239), .ZN(
        n22365) );
  OAI22_X2 U12662 ( .A1(n22641), .A2(n22640), .B1(n22639), .B2(n22638), .ZN(
        n22742) );
  OAI22_X2 U12663 ( .A1(n22247), .A2(n22640), .B1(n22639), .B2(n22246), .ZN(
        n22371) );
  OAI22_X2 U12664 ( .A1(n22388), .A2(n22640), .B1(n22639), .B2(n22387), .ZN(
        n22420) );
  OAI22_X2 U12665 ( .A1(n22459), .A2(n22640), .B1(n22639), .B2(n22458), .ZN(
        n22491) );
  NAND2_X2 U12666 ( .A1(n14226), .A2(n14297), .ZN(n14227) );
  INV_X2 U12667 ( .A(n18611), .ZN(n18615) );
  OAI22_X2 U12668 ( .A1(n22530), .A2(n22639), .B1(n22529), .B2(n22640), .ZN(
        n22562) );
  NAND3_X1 U12669 ( .A1(n17404), .A2(n11328), .A3(n14477), .ZN(n14478) );
  NAND4_X1 U12670 ( .A1(n12984), .A2(n12940), .A3(n11328), .A4(n12939), .ZN(
        n12941) );
  NAND2_X4 U12671 ( .A1(n22457), .A2(n15821), .ZN(n15883) );
  NAND2_X4 U12672 ( .A1(n11329), .A2(n12889), .ZN(n15821) );
  OR2_X2 U12673 ( .A1(n20353), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11334) );
  NAND2_X1 U12674 ( .A1(n13173), .A2(n11335), .ZN(n20370) );
  OAI21_X1 U12675 ( .B1(n20374), .B2(n16392), .A(n11335), .ZN(n16394) );
  INV_X2 U12676 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13058) );
  AOI21_X2 U12677 ( .B1(n17360), .B2(n22122), .A(n11338), .ZN(n14641) );
  NAND2_X1 U12678 ( .A1(n12464), .A2(n11339), .ZN(n12484) );
  NAND2_X1 U12679 ( .A1(n12461), .A2(n12460), .ZN(n11339) );
  NOR2_X2 U12680 ( .A1(n11348), .A2(n12563), .ZN(n11347) );
  INV_X1 U12681 ( .A(n15776), .ZN(n11647) );
  NAND2_X1 U12682 ( .A1(n11341), .A2(n15776), .ZN(n11644) );
  NAND2_X1 U12683 ( .A1(n17052), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16841) );
  NAND2_X2 U12684 ( .A1(n11172), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17468) );
  NAND2_X2 U12685 ( .A1(n16797), .A2(n17082), .ZN(n17465) );
  AND2_X2 U12686 ( .A1(n11362), .A2(n11360), .ZN(n16797) );
  NAND2_X2 U12687 ( .A1(n11350), .A2(n12619), .ZN(n15777) );
  NAND2_X1 U12688 ( .A1(n15740), .A2(n15739), .ZN(n11350) );
  NAND2_X1 U12689 ( .A1(n15639), .A2(n15640), .ZN(n11351) );
  OR2_X2 U12690 ( .A1(n16703), .A2(n11279), .ZN(n16713) );
  NAND2_X1 U12691 ( .A1(n12530), .A2(n12564), .ZN(n11352) );
  NAND2_X1 U12692 ( .A1(n12767), .A2(n15085), .ZN(n11353) );
  AND2_X1 U12693 ( .A1(n11860), .A2(n11866), .ZN(n11867) );
  NAND2_X1 U12694 ( .A1(n11881), .A2(n11355), .ZN(n11882) );
  NAND3_X1 U12695 ( .A1(n11868), .A2(n14344), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11918) );
  NAND3_X1 U12696 ( .A1(n11868), .A2(n14344), .A3(n11357), .ZN(n11356) );
  NAND3_X1 U12697 ( .A1(n13762), .A2(n14318), .A3(n11274), .ZN(n11358) );
  INV_X1 U12698 ( .A(n11913), .ZN(n16014) );
  OR2_X2 U12699 ( .A1(n16717), .A2(n16893), .ZN(n16719) );
  NAND2_X1 U12700 ( .A1(n11271), .A2(n11645), .ZN(n17434) );
  INV_X1 U12701 ( .A(n12789), .ZN(n11364) );
  OAI21_X1 U12702 ( .B1(n18471), .B2(n11367), .A(n11366), .ZN(n18460) );
  INV_X2 U12703 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21191) );
  AND2_X1 U12704 ( .A1(n11371), .A2(n11949), .ZN(n14535) );
  NAND2_X1 U12705 ( .A1(n11371), .A2(n11589), .ZN(n14536) );
  NAND2_X2 U12706 ( .A1(n11439), .A2(n11371), .ZN(n13756) );
  NAND2_X2 U12707 ( .A1(n12457), .A2(n11948), .ZN(n11371) );
  AND2_X4 U12708 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U12709 ( .A1(n17028), .A2(n11372), .ZN(P2_U3027) );
  NAND2_X1 U12710 ( .A1(n16817), .A2(n11373), .ZN(P2_U2995) );
  NAND2_X1 U12711 ( .A1(n12472), .A2(n11157), .ZN(n12460) );
  NAND2_X1 U12712 ( .A1(n11906), .A2(n11905), .ZN(n11376) );
  NOR2_X2 U12713 ( .A1(n16818), .A2(n17024), .ZN(n16811) );
  NAND2_X2 U12714 ( .A1(n11381), .A2(n11380), .ZN(n16818) );
  NAND2_X1 U12715 ( .A1(n18121), .A2(n11386), .ZN(n11385) );
  NAND3_X1 U12716 ( .A1(n11396), .A2(n11395), .A3(n11392), .ZN(n11391) );
  NAND2_X1 U12717 ( .A1(n20907), .A2(n11400), .ZN(n11399) );
  NAND2_X1 U12718 ( .A1(n11403), .A2(n11404), .ZN(n20791) );
  NAND2_X1 U12720 ( .A1(n20770), .A2(n20932), .ZN(n20772) );
  OAI211_X2 U12721 ( .C1(n11418), .C2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n11417), .B(n11414), .ZN(n20723) );
  INV_X1 U12722 ( .A(n11423), .ZN(n18349) );
  NAND2_X1 U12723 ( .A1(n11861), .A2(n11869), .ZN(n11855) );
  OAI21_X1 U12724 ( .B1(n11855), .B2(n11431), .A(n14921), .ZN(n11658) );
  AND2_X2 U12725 ( .A1(n11785), .A2(n11784), .ZN(n13761) );
  AND2_X2 U12726 ( .A1(n11754), .A2(n11755), .ZN(n11861) );
  INV_X1 U12727 ( .A(n16773), .ZN(n11437) );
  NAND2_X1 U12728 ( .A1(n16774), .A2(n17464), .ZN(n11436) );
  NAND3_X1 U12729 ( .A1(n11436), .A2(n11437), .A3(n11232), .ZN(n11435) );
  INV_X1 U12730 ( .A(n12484), .ZN(n14730) );
  NAND2_X1 U12732 ( .A1(n15777), .A2(n11443), .ZN(n11441) );
  OAI21_X1 U12733 ( .B1(n15777), .B2(n15778), .A(n15779), .ZN(n17436) );
  NAND2_X1 U12734 ( .A1(n15778), .A2(n15779), .ZN(n11449) );
  AOI21_X1 U12735 ( .B1(n16830), .B2(n16828), .A(n16777), .ZN(n16819) );
  INV_X1 U12736 ( .A(n11451), .ZN(n16781) );
  NAND3_X1 U12737 ( .A1(n12094), .A2(n12095), .A3(n11459), .ZN(n14399) );
  INV_X2 U12738 ( .A(n16849), .ZN(n11468) );
  AND2_X1 U12739 ( .A1(n16640), .A2(n11474), .ZN(n16607) );
  NAND2_X1 U12740 ( .A1(n16640), .A2(n11476), .ZN(n16610) );
  NAND2_X1 U12741 ( .A1(n16640), .A2(n16628), .ZN(n16623) );
  NAND2_X1 U12742 ( .A1(n12395), .A2(n11299), .ZN(n17002) );
  INV_X2 U12743 ( .A(n14477), .ZN(n22528) );
  NAND2_X1 U12744 ( .A1(n16294), .A2(n11480), .ZN(n11479) );
  OAI211_X1 U12745 ( .C1(n16294), .C2(n11483), .A(n11481), .B(n11479), .ZN(
        n15934) );
  NAND2_X1 U12746 ( .A1(n20348), .A2(n11488), .ZN(n11487) );
  NAND2_X1 U12747 ( .A1(n16388), .A2(n11495), .ZN(n11493) );
  NAND2_X1 U12748 ( .A1(n16388), .A2(n11497), .ZN(n11494) );
  NAND3_X1 U12749 ( .A1(n11493), .A2(n13169), .A3(n11492), .ZN(n16348) );
  INV_X2 U12750 ( .A(n17363), .ZN(n13691) );
  NAND3_X1 U12751 ( .A1(n17286), .A2(n21166), .A3(n17306), .ZN(n11504) );
  OR2_X2 U12752 ( .A1(n21582), .A2(n21211), .ZN(n21579) );
  NAND3_X1 U12753 ( .A1(n17263), .A2(n17262), .A3(n11509), .ZN(n11508) );
  NOR2_X1 U12754 ( .A1(n16172), .A2(n16114), .ZN(n16113) );
  INV_X1 U12755 ( .A(n16099), .ZN(n11523) );
  NAND2_X1 U12756 ( .A1(n14953), .A2(n11524), .ZN(n15684) );
  INV_X1 U12757 ( .A(n14686), .ZN(n11531) );
  NAND3_X1 U12758 ( .A1(n11532), .A2(n14818), .A3(n11531), .ZN(n14947) );
  NAND2_X1 U12759 ( .A1(n18291), .A2(n21509), .ZN(n21490) );
  NAND2_X1 U12760 ( .A1(n18295), .A2(n21510), .ZN(n18291) );
  NAND2_X1 U12761 ( .A1(n18296), .A2(n18329), .ZN(n18295) );
  NAND2_X1 U12762 ( .A1(n11542), .A2(n11540), .ZN(P3_U2834) );
  NAND3_X1 U12763 ( .A1(n21508), .A2(n21620), .A3(n11543), .ZN(n11542) );
  NAND2_X1 U12764 ( .A1(n11547), .A2(n11544), .ZN(n11543) );
  NAND2_X1 U12765 ( .A1(n21493), .A2(n21494), .ZN(n11547) );
  AOI21_X1 U12766 ( .B1(n18440), .B2(n11549), .A(n18329), .ZN(n18090) );
  AOI21_X1 U12767 ( .B1(n18091), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11548), .ZN(n18370) );
  NAND2_X1 U12768 ( .A1(n18440), .A2(n18086), .ZN(n18403) );
  AND2_X1 U12769 ( .A1(n18026), .A2(n18027), .ZN(n11551) );
  INV_X2 U12770 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21633) );
  OAI211_X1 U12771 ( .C1(n11552), .C2(n18850), .A(n18849), .B(n18980), .ZN(
        n18851) );
  NAND2_X1 U12772 ( .A1(n18838), .A2(n11164), .ZN(n11552) );
  AOI21_X1 U12773 ( .B1(n18906), .B2(n11558), .A(n11556), .ZN(n18930) );
  NAND2_X1 U12774 ( .A1(n11708), .A2(n11301), .ZN(n11727) );
  NAND2_X1 U12775 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11568) );
  NAND3_X1 U12776 ( .A1(n11569), .A2(n11567), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11716) );
  NOR2_X1 U12777 ( .A1(n18676), .A2(n11568), .ZN(n11567) );
  NAND3_X1 U12778 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11569), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U12779 ( .A1(n11700), .A2(n11318), .ZN(n11697) );
  NAND2_X1 U12780 ( .A1(n12703), .A2(n11573), .ZN(n12715) );
  NAND3_X1 U12781 ( .A1(n11578), .A2(n12584), .A3(n12561), .ZN(n12616) );
  NAND3_X1 U12782 ( .A1(n11578), .A2(n12584), .A3(n11576), .ZN(n12621) );
  INV_X1 U12783 ( .A(n12615), .ZN(n11579) );
  NAND2_X1 U12784 ( .A1(n12719), .A2(n11323), .ZN(n16003) );
  NAND2_X1 U12785 ( .A1(n12719), .A2(n12720), .ZN(n12726) );
  INV_X1 U12786 ( .A(n12728), .ZN(n12736) );
  INV_X1 U12787 ( .A(n15807), .ZN(n11594) );
  NAND2_X1 U12788 ( .A1(n11594), .A2(n11595), .ZN(n16582) );
  NAND2_X1 U12789 ( .A1(n14532), .A2(n11239), .ZN(n14607) );
  AOI211_X1 U12790 ( .C1(n16543), .C2(n16016), .A(n11599), .B(n11601), .ZN(
        n11600) );
  AND2_X2 U12791 ( .A1(n15571), .A2(n11316), .ZN(n16117) );
  INV_X1 U12792 ( .A(n14710), .ZN(n11611) );
  NAND2_X1 U12793 ( .A1(n11611), .A2(n11612), .ZN(n15096) );
  NAND2_X1 U12794 ( .A1(n14572), .A2(n11619), .ZN(n14709) );
  AND2_X1 U12795 ( .A1(n16094), .A2(n11628), .ZN(n16086) );
  NAND2_X1 U12796 ( .A1(n16094), .A2(n11629), .ZN(n16073) );
  NAND2_X1 U12797 ( .A1(n16094), .A2(n16095), .ZN(n16085) );
  NAND2_X1 U12798 ( .A1(n11638), .A2(n11639), .ZN(n11637) );
  INV_X1 U12799 ( .A(n11640), .ZN(n11638) );
  NAND3_X1 U12800 ( .A1(n12489), .A2(n12504), .A3(n12505), .ZN(n11642) );
  NAND4_X1 U12801 ( .A1(n12488), .A2(n12503), .A3(n12506), .A4(n12487), .ZN(
        n11643) );
  NAND2_X1 U12802 ( .A1(n11646), .A2(n15738), .ZN(n11645) );
  NAND2_X1 U12803 ( .A1(n11648), .A2(n12783), .ZN(n15775) );
  INV_X1 U12804 ( .A(n16717), .ZN(n11653) );
  NAND2_X1 U12805 ( .A1(n11656), .A2(n11852), .ZN(n14375) );
  INV_X1 U12806 ( .A(n11920), .ZN(n11656) );
  NAND3_X1 U12807 ( .A1(n11658), .A2(n14151), .A3(n11657), .ZN(n11920) );
  INV_X1 U12808 ( .A(n11859), .ZN(n11657) );
  AND3_X2 U12809 ( .A1(n11853), .A2(n11856), .A3(n11875), .ZN(n14318) );
  NAND3_X1 U12810 ( .A1(n11903), .A2(n11904), .A3(n11660), .ZN(n11907) );
  NAND2_X1 U12811 ( .A1(n11864), .A2(n11302), .ZN(n11660) );
  AND2_X2 U12812 ( .A1(n11864), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11937) );
  NAND3_X1 U12813 ( .A1(n12700), .A2(n12699), .A3(n11230), .ZN(n11661) );
  NAND3_X1 U12814 ( .A1(n12784), .A2(n16849), .A3(n11668), .ZN(n11667) );
  AND2_X1 U12815 ( .A1(n12784), .A2(n11668), .ZN(n12773) );
  NAND2_X1 U12816 ( .A1(n12713), .A2(n16952), .ZN(n11669) );
  NAND2_X1 U12817 ( .A1(n11670), .A2(n11669), .ZN(n16724) );
  NAND3_X1 U12818 ( .A1(n11670), .A2(n11669), .A3(n11231), .ZN(n12730) );
  AND2_X1 U12819 ( .A1(n13787), .A2(n13790), .ZN(n13791) );
  AND2_X1 U12820 ( .A1(n19612), .A2(n11196), .ZN(n12059) );
  NAND2_X1 U12821 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U12822 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U12823 ( .A1(n12468), .A2(n12473), .ZN(n12472) );
  INV_X1 U12824 ( .A(n15095), .ZN(n15554) );
  AOI22_X1 U12825 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U12826 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U12827 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U12828 ( .A1(n12082), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U12829 ( .A1(n11199), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U12830 ( .A1(n12082), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11756) );
  AOI21_X1 U12831 ( .B1(n11200), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n14755), .ZN(n11846) );
  AOI21_X1 U12832 ( .B1(n12082), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11787) );
  NAND2_X1 U12833 ( .A1(n12082), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11770) );
  AOI21_X1 U12834 ( .B1(n12082), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14755), .ZN(n11792) );
  AOI22_X1 U12835 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11818) );
  OR2_X1 U12836 ( .A1(n18819), .A2(n18821), .ZN(n11671) );
  INV_X1 U12837 ( .A(n12115), .ZN(n12398) );
  AOI21_X1 U12838 ( .B1(n13298), .B2(n13463), .A(n13297), .ZN(n14946) );
  INV_X1 U12839 ( .A(n14946), .ZN(n13299) );
  AND2_X1 U12840 ( .A1(n15977), .A2(n16571), .ZN(n11672) );
  AND2_X1 U12841 ( .A1(n12804), .A2(n12803), .ZN(n11673) );
  INV_X1 U12842 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11694) );
  OR2_X1 U12843 ( .A1(n16161), .A2(n22111), .ZN(n11674) );
  AND4_X1 U12844 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n11675) );
  AND2_X1 U12845 ( .A1(n20313), .A2(n20321), .ZN(n11676) );
  AND4_X1 U12846 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n11677) );
  OR2_X1 U12847 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11678) );
  OR2_X1 U12848 ( .A1(n13976), .A2(n12069), .ZN(n11679) );
  AND2_X1 U12849 ( .A1(n16604), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11680) );
  NAND3_X1 U12850 ( .A1(n16785), .A2(n12693), .A3(n16807), .ZN(n11681) );
  AND2_X1 U12851 ( .A1(n15962), .A2(n15999), .ZN(n11682) );
  AND3_X1 U12852 ( .A1(n11847), .A2(n11846), .A3(n11845), .ZN(n11683) );
  NAND2_X1 U12853 ( .A1(n11975), .A2(n11974), .ZN(n11684) );
  INV_X1 U12854 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11695) );
  XNOR2_X1 U12855 ( .A(P1_REIP_REG_30__SCAN_IN), .B(n16067), .ZN(n11685) );
  AND2_X1 U12856 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11686) );
  INV_X1 U12857 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18318) );
  OR2_X1 U12858 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11687) );
  INV_X1 U12859 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18087) );
  AND2_X1 U12860 ( .A1(n11839), .A2(n11838), .ZN(n11688) );
  OR2_X1 U12861 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11689) );
  OR2_X1 U12862 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11690) );
  OR2_X1 U12863 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11691) );
  INV_X1 U12864 ( .A(n16389), .ZN(n16401) );
  OR2_X1 U12865 ( .A1(n18255), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11692) );
  INV_X1 U12866 ( .A(n14935), .ZN(n14939) );
  OR2_X1 U12867 ( .A1(n18329), .A2(n18263), .ZN(n11693) );
  INV_X1 U12868 ( .A(n13239), .ZN(n13219) );
  NOR2_X1 U12869 ( .A1(n13219), .A2(n14257), .ZN(n13222) );
  OR2_X1 U12870 ( .A1(n13203), .A2(n13207), .ZN(n13193) );
  NAND2_X1 U12871 ( .A1(n11209), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U12872 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11771) );
  AND2_X1 U12873 ( .A1(n11940), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11899) );
  AND2_X1 U12874 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  AOI22_X1 U12875 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11209), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11761) );
  INV_X1 U12876 ( .A(n11923), .ZN(n11852) );
  NAND2_X1 U12877 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11845) );
  AND2_X1 U12878 ( .A1(n13118), .A2(n13117), .ZN(n13119) );
  INV_X1 U12879 ( .A(n13115), .ZN(n13120) );
  INV_X1 U12880 ( .A(n13220), .ZN(n13232) );
  OAI21_X1 U12881 ( .B1(n14894), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12974), 
        .ZN(n12969) );
  NOR2_X1 U12882 ( .A1(n12517), .A2(n12516), .ZN(n12522) );
  AOI21_X1 U12883 ( .B1(n15895), .B2(n12930), .A(n12929), .ZN(n12984) );
  OR2_X1 U12884 ( .A1(n12220), .A2(n12219), .ZN(n12434) );
  NAND2_X1 U12885 ( .A1(n12507), .A2(n12609), .ZN(n12508) );
  INV_X1 U12886 ( .A(n12773), .ZN(n12782) );
  NAND2_X1 U12887 ( .A1(n13765), .A2(n13764), .ZN(n13787) );
  NAND2_X1 U12888 ( .A1(n18377), .A2(n18087), .ZN(n18088) );
  AOI21_X1 U12889 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n22122), .A(
        n13236), .ZN(n13237) );
  NAND2_X1 U12890 ( .A1(n22528), .A2(n15524), .ZN(n14588) );
  AND2_X1 U12891 ( .A1(n13679), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13680) );
  OR2_X1 U12892 ( .A1(n12956), .A2(n12955), .ZN(n13165) );
  INV_X1 U12893 ( .A(n14676), .ZN(n13270) );
  OR2_X1 U12894 ( .A1(n13169), .A2(n21811), .ZN(n13168) );
  NAND2_X1 U12895 ( .A1(n13043), .A2(n13042), .ZN(n13262) );
  INV_X1 U12896 ( .A(n14653), .ZN(n13795) );
  INV_X1 U12897 ( .A(n15808), .ZN(n13873) );
  OR2_X1 U12898 ( .A1(n12141), .A2(n12140), .ZN(n12161) );
  NAND2_X1 U12899 ( .A1(n12731), .A2(n16907), .ZN(n12732) );
  INV_X1 U12900 ( .A(n12093), .ZN(n12163) );
  AND2_X1 U12902 ( .A1(n13239), .A2(n14262), .ZN(n13240) );
  AOI21_X1 U12903 ( .B1(n13238), .B2(n14262), .A(n13237), .ZN(n13241) );
  NOR2_X1 U12904 ( .A1(n21964), .A2(n22253), .ZN(n14889) );
  AND4_X1 U12905 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12868) );
  AND2_X1 U12906 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n13605), .ZN(
        n13606) );
  INV_X1 U12907 ( .A(n13734), .ZN(n13741) );
  INV_X1 U12908 ( .A(n13398), .ZN(n13463) );
  AOI21_X1 U12909 ( .B1(n13305), .B2(n13463), .A(n13304), .ZN(n15108) );
  OAI21_X1 U12910 ( .B1(n13253), .B2(n13398), .A(n13252), .ZN(n13254) );
  OR2_X1 U12911 ( .A1(n20370), .A2(n16390), .ZN(n16377) );
  NAND2_X1 U12912 ( .A1(n13261), .A2(n13262), .ZN(n13265) );
  INV_X1 U12913 ( .A(n15576), .ZN(n13812) );
  AND2_X1 U12914 ( .A1(n11958), .A2(n11957), .ZN(n14526) );
  INV_X1 U12915 ( .A(n15647), .ZN(n12224) );
  INV_X1 U12916 ( .A(n11218), .ZN(n17671) );
  INV_X1 U12917 ( .A(n17307), .ZN(n17977) );
  NAND2_X1 U12918 ( .A1(n18075), .A2(n18074), .ZN(n18079) );
  NOR2_X1 U12919 ( .A1(n18452), .A2(n18451), .ZN(n18450) );
  INV_X1 U12920 ( .A(n17978), .ZN(n21168) );
  OR2_X1 U12921 ( .A1(n17977), .A2(n21166), .ZN(n17976) );
  INV_X1 U12922 ( .A(n17413), .ZN(n12925) );
  NOR2_X1 U12923 ( .A1(n13322), .A2(n13317), .ZN(n13346) );
  INV_X1 U12924 ( .A(n22050), .ZN(n21964) );
  NOR2_X1 U12925 ( .A1(n13399), .A2(n13371), .ZN(n13403) );
  NOR2_X1 U12926 ( .A1(n13351), .A2(n13347), .ZN(n13352) );
  OR2_X1 U12927 ( .A1(n20392), .A2(n13746), .ZN(n16407) );
  AND2_X1 U12928 ( .A1(n21707), .A2(n21878), .ZN(n21826) );
  OR2_X1 U12929 ( .A1(n22275), .A2(n22231), .ZN(n22245) );
  INV_X1 U12930 ( .A(n14844), .ZN(n22265) );
  INV_X1 U12931 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22238) );
  AND2_X1 U12932 ( .A1(n14842), .A2(n14641), .ZN(n15016) );
  INV_X1 U12933 ( .A(n15027), .ZN(n22274) );
  INV_X1 U12934 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22251) );
  INV_X1 U12935 ( .A(n16509), .ZN(n22129) );
  AND2_X1 U12936 ( .A1(n11980), .A2(n11979), .ZN(n14809) );
  AND2_X1 U12937 ( .A1(n11967), .A2(n11966), .ZN(n14613) );
  NAND2_X1 U12938 ( .A1(n14071), .A2(n14070), .ZN(n16533) );
  INV_X1 U12939 ( .A(n11166), .ZN(n12355) );
  OR2_X1 U12940 ( .A1(n18886), .A2(n12709), .ZN(n16754) );
  INV_X1 U12941 ( .A(n12750), .ZN(n14314) );
  AND2_X1 U12942 ( .A1(n14360), .A2(n14359), .ZN(n14758) );
  INV_X1 U12943 ( .A(n11165), .ZN(n18809) );
  NAND2_X1 U12944 ( .A1(n19573), .A2(n19642), .ZN(n19623) );
  AND2_X1 U12945 ( .A1(n15656), .A2(n19709), .ZN(n15667) );
  NAND2_X1 U12946 ( .A1(n19660), .A2(n17481), .ZN(n19581) );
  OR2_X1 U12947 ( .A1(n19551), .A2(n17477), .ZN(n19675) );
  INV_X1 U12948 ( .A(n20010), .ZN(n19960) );
  CLKBUF_X1 U12949 ( .A(n14318), .Z(n14804) );
  NOR2_X1 U12950 ( .A1(n21134), .A2(n21133), .ZN(n21132) );
  INV_X1 U12951 ( .A(n18084), .ZN(n18083) );
  INV_X1 U12952 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18472) );
  AOI21_X1 U12953 ( .B1(n21506), .B2(n21602), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21507) );
  AND2_X1 U12954 ( .A1(n18256), .A2(n11692), .ZN(n18257) );
  NAND2_X1 U12955 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21346), .ZN(
        n18385) );
  NOR2_X1 U12956 ( .A1(n21207), .A2(n17976), .ZN(n17582) );
  NOR2_X1 U12957 ( .A1(n17244), .A2(n17243), .ZN(n19295) );
  OAI211_X1 U12958 ( .C1(n11685), .C2(n22085), .A(n16061), .B(n11674), .ZN(
        n16062) );
  AND2_X1 U12959 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n13536), .ZN(
        n13537) );
  AND2_X1 U12960 ( .A1(n14892), .A2(n14891), .ZN(n22079) );
  AND2_X1 U12961 ( .A1(n22050), .A2(n14897), .ZN(n22107) );
  INV_X1 U12962 ( .A(n16217), .ZN(n20322) );
  AND2_X1 U12963 ( .A1(n15814), .A2(n15813), .ZN(n22378) );
  OR2_X1 U12964 ( .A1(n16147), .A2(n15801), .ZN(n16132) );
  AND2_X1 U12965 ( .A1(n13294), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13301) );
  XNOR2_X1 U12966 ( .A(n13082), .B(n15909), .ZN(n14826) );
  AND2_X1 U12967 ( .A1(n16407), .A2(n13748), .ZN(n20379) );
  INV_X1 U12968 ( .A(n21734), .ZN(n21819) );
  NAND2_X1 U12969 ( .A1(n15834), .A2(n15833), .ZN(n15907) );
  INV_X1 U12970 ( .A(n21705), .ZN(n21821) );
  INV_X1 U12971 ( .A(n22245), .ZN(n22648) );
  INV_X1 U12972 ( .A(n22652), .ZN(n22654) );
  INV_X1 U12973 ( .A(n15526), .ZN(n22660) );
  INV_X1 U12974 ( .A(n22577), .ZN(n22667) );
  AND2_X1 U12975 ( .A1(n15016), .A2(n22230), .ZN(n22674) );
  AND2_X1 U12976 ( .A1(n15016), .A2(n14997), .ZN(n22583) );
  AND2_X1 U12977 ( .A1(n15016), .A2(n15026), .ZN(n22686) );
  AND2_X1 U12978 ( .A1(n15016), .A2(n15027), .ZN(n22693) );
  INV_X1 U12979 ( .A(n22715), .ZN(n22704) );
  INV_X1 U12980 ( .A(n14972), .ZN(n14969) );
  NOR2_X1 U12981 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14846), .ZN(n22632) );
  AND2_X1 U12982 ( .A1(n14971), .A2(n16503), .ZN(n22230) );
  INV_X1 U12983 ( .A(n22625), .ZN(n22617) );
  INV_X1 U12984 ( .A(n22350), .ZN(n22369) );
  INV_X1 U12985 ( .A(n22488), .ZN(n22495) );
  AND2_X1 U12986 ( .A1(n15028), .A2(n15027), .ZN(n22743) );
  OR2_X1 U12987 ( .A1(n14311), .A2(n14119), .ZN(n14912) );
  NAND2_X1 U12988 ( .A1(n11165), .A2(n11671), .ZN(n18839) );
  INV_X1 U12989 ( .A(n18973), .ZN(n18955) );
  INV_X1 U12990 ( .A(n16606), .ZN(n16596) );
  XNOR2_X1 U12991 ( .A(n14294), .B(n14293), .ZN(n19551) );
  AND2_X1 U12992 ( .A1(n14397), .A2(n14396), .ZN(n19905) );
  AND2_X1 U12993 ( .A1(n14299), .A2(n22182), .ZN(n17509) );
  AND2_X1 U12994 ( .A1(n17452), .A2(n14290), .ZN(n17443) );
  AND2_X1 U12995 ( .A1(n17452), .A2(n17340), .ZN(n17457) );
  XNOR2_X1 U12996 ( .A(n12785), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15776) );
  AND2_X1 U12997 ( .A1(n14339), .A2(n18631), .ZN(n14378) );
  AND2_X1 U12998 ( .A1(n14378), .A2(n14365), .ZN(n19003) );
  OAI21_X2 U12999 ( .B1(n17179), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14915), 
        .ZN(n19715) );
  NAND2_X1 U13000 ( .A1(n14912), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17179) );
  AND3_X1 U13001 ( .A1(n14740), .A2(n14739), .A3(n14738), .ZN(n15630) );
  AND2_X1 U13002 ( .A1(n19695), .A2(n19688), .ZN(n19899) );
  AND2_X1 U13003 ( .A1(n19695), .A2(n19676), .ZN(n20102) );
  OAI21_X1 U13004 ( .B1(n19654), .B2(n19653), .A(n19652), .ZN(n20082) );
  OAI21_X1 U13005 ( .B1(n19654), .B2(n19651), .A(n19650), .ZN(n20083) );
  INV_X1 U13006 ( .A(n19943), .ZN(n20081) );
  NOR2_X1 U13007 ( .A1(n19623), .A2(n19657), .ZN(n20062) );
  NOR2_X1 U13008 ( .A1(n19623), .A2(n19643), .ZN(n19980) );
  NOR2_X1 U13009 ( .A1(n19581), .A2(n19675), .ZN(n20048) );
  INV_X1 U13010 ( .A(n19959), .ZN(n19950) );
  AOI21_X1 U13011 ( .B1(n20015), .B2(n19715), .A(n19537), .ZN(n20018) );
  INV_X1 U13012 ( .A(n19732), .ZN(n19764) );
  NAND2_X1 U13013 ( .A1(n21690), .A2(n21656), .ZN(n20470) );
  NOR2_X1 U13014 ( .A1(n21163), .A2(n17335), .ZN(n21655) );
  INV_X1 U13015 ( .A(n20531), .ZN(n20534) );
  NAND2_X1 U13016 ( .A1(n21667), .A2(n20534), .ZN(n20957) );
  INV_X1 U13017 ( .A(n20957), .ZN(n20915) );
  INV_X1 U13018 ( .A(n17952), .ZN(n17953) );
  NAND2_X1 U13019 ( .A1(n21095), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21094) );
  NOR2_X1 U13020 ( .A1(n21063), .A2(n21106), .ZN(n21101) );
  NAND2_X1 U13021 ( .A1(n21114), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21113) );
  NAND4_X1 U13022 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(n20996), .A4(n21150), .ZN(n21134) );
  INV_X1 U13023 ( .A(n21139), .ZN(n21120) );
  OAI21_X1 U13024 ( .B1(n17582), .B2(n17581), .A(n21690), .ZN(n20969) );
  NAND2_X1 U13025 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18449), .ZN(
        n18448) );
  INV_X1 U13026 ( .A(n21507), .ZN(n21508) );
  NOR2_X2 U13027 ( .A1(n21470), .A2(n21321), .ZN(n21623) );
  NOR3_X1 U13028 ( .A1(n17582), .A2(n17315), .A3(n21215), .ZN(n21644) );
  INV_X1 U13029 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21637) );
  NAND2_X1 U13030 ( .A1(n14305), .A2(n15895), .ZN(n16043) );
  OAI211_X1 U13031 ( .C1(n14453), .C2(n22135), .A(n16043), .B(n14868), .ZN(
        n21696) );
  INV_X1 U13032 ( .A(n22093), .ZN(n22111) );
  INV_X1 U13033 ( .A(n22108), .ZN(n22052) );
  INV_X1 U13034 ( .A(n22061), .ZN(n22098) );
  NAND2_X1 U13035 ( .A1(n20326), .A2(n22633), .ZN(n16217) );
  INV_X1 U13036 ( .A(n16274), .ZN(n16278) );
  OR2_X1 U13037 ( .A1(n16043), .A2(n14467), .ZN(n14519) );
  OAI21_X1 U13038 ( .B1(n16117), .B2(n15802), .A(n16132), .ZN(n22008) );
  INV_X1 U13039 ( .A(n20392), .ZN(n22113) );
  INV_X1 U13040 ( .A(n11156), .ZN(n21862) );
  INV_X1 U13041 ( .A(n21925), .ZN(n21906) );
  OR2_X1 U13042 ( .A1(n22275), .A2(n15518), .ZN(n22652) );
  INV_X1 U13043 ( .A(n22674), .ZN(n22671) );
  INV_X1 U13044 ( .A(n22583), .ZN(n22683) );
  INV_X1 U13045 ( .A(n22686), .ZN(n22593) );
  NAND2_X1 U13046 ( .A1(n14969), .A2(n22230), .ZN(n22702) );
  AOI22_X1 U13047 ( .A1(n22326), .A2(n22331), .B1(n22325), .B2(n22324), .ZN(
        n22709) );
  NAND2_X1 U13048 ( .A1(n14969), .A2(n15026), .ZN(n22715) );
  AOI22_X1 U13049 ( .A1(n22342), .A2(n22346), .B1(n22341), .B2(n22340), .ZN(
        n22723) );
  INV_X1 U13050 ( .A(n22522), .ZN(n22520) );
  INV_X1 U13051 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22253) );
  OR2_X1 U13052 ( .A1(n18954), .A2(n19593), .ZN(n18973) );
  NOR2_X1 U13053 ( .A1(n11672), .A2(n11680), .ZN(n14123) );
  XNOR2_X1 U13054 ( .A(n14095), .B(n14094), .ZN(n15961) );
  INV_X1 U13055 ( .A(n19905), .ZN(n19770) );
  AND2_X1 U13056 ( .A1(n19912), .A2(n19911), .ZN(n19781) );
  NOR2_X1 U13057 ( .A1(n17509), .A2(n17542), .ZN(n17529) );
  INV_X1 U13058 ( .A(n17509), .ZN(n17544) );
  INV_X1 U13059 ( .A(n17443), .ZN(n17475) );
  NAND2_X1 U13060 ( .A1(n19057), .A2(n12798), .ZN(n17452) );
  INV_X1 U13061 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19612) );
  INV_X1 U13062 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19689) );
  INV_X1 U13063 ( .A(n19899), .ZN(n20116) );
  NAND2_X1 U13064 ( .A1(n19695), .A2(n19658), .ZN(n20098) );
  NAND2_X1 U13065 ( .A1(n19695), .A2(n19644), .ZN(n20086) );
  AND2_X1 U13066 ( .A1(n19632), .A2(n19631), .ZN(n19751) );
  INV_X1 U13067 ( .A(n20062), .ZN(n20073) );
  INV_X1 U13068 ( .A(n19980), .ZN(n20066) );
  INV_X1 U13069 ( .A(n20048), .ZN(n19979) );
  AND2_X1 U13070 ( .A1(n15660), .A2(n15659), .ZN(n20046) );
  INV_X1 U13071 ( .A(n19561), .ZN(n20039) );
  INV_X1 U13072 ( .A(n19955), .ZN(n19953) );
  INV_X1 U13073 ( .A(n19814), .ZN(n19812) );
  INV_X1 U13074 ( .A(n19966), .ZN(n20021) );
  NAND4_X1 U13075 ( .A1(n20534), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n21211), 
        .A4(n20533), .ZN(n20912) );
  INV_X1 U13076 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20664) );
  INV_X1 U13077 ( .A(n20963), .ZN(n20903) );
  AND2_X1 U13078 ( .A1(n21063), .A2(n21150), .ZN(n21139) );
  INV_X1 U13079 ( .A(n21225), .ZN(n21492) );
  NOR2_X1 U13080 ( .A1(n18003), .A2(n18002), .ZN(n21012) );
  INV_X1 U13081 ( .A(n20479), .ZN(n20523) );
  INV_X1 U13082 ( .A(n18444), .ZN(n18388) );
  INV_X1 U13083 ( .A(n21623), .ZN(n21569) );
  INV_X1 U13084 ( .A(n21615), .ZN(n21591) );
  INV_X1 U13085 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21640) );
  OR2_X1 U13086 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18564), .ZN(n22205) );
  OAI21_X1 U13087 ( .B1(n16901), .B2(n17445), .A(n11673), .ZN(P2_U2985) );
  INV_X1 U13088 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11698) );
  INV_X1 U13089 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18676) );
  INV_X1 U13090 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15793) );
  INV_X1 U13091 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17453) );
  INV_X1 U13092 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18747) );
  NAND2_X1 U13093 ( .A1(n11713), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11710) );
  INV_X1 U13094 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16812) );
  NAND2_X1 U13095 ( .A1(n11728), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11729) );
  INV_X1 U13096 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16791) );
  INV_X1 U13097 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12018) );
  INV_X1 U13098 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18885) );
  INV_X1 U13099 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16739) );
  INV_X1 U13100 ( .A(n11696), .ZN(n11735) );
  INV_X1 U13101 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16729) );
  INV_X1 U13102 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18974) );
  OAI21_X1 U13103 ( .B1(n11702), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n11737), .ZN(n11699) );
  INV_X1 U13104 ( .A(n11699), .ZN(n18960) );
  NOR2_X1 U13105 ( .A1(n11700), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11701) );
  OR2_X1 U13106 ( .A1(n11702), .A2(n11701), .ZN(n16708) );
  INV_X1 U13107 ( .A(n16708), .ZN(n18942) );
  NOR2_X1 U13108 ( .A1(n11703), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11704) );
  OR2_X1 U13109 ( .A1(n11700), .A2(n11704), .ZN(n16716) );
  INV_X1 U13110 ( .A(n16716), .ZN(n18931) );
  AOI21_X1 U13111 ( .B1(n16739), .B2(n11705), .A(n11696), .ZN(n18908) );
  OR2_X1 U13112 ( .A1(n11733), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11706) );
  NAND2_X1 U13113 ( .A1(n11705), .A2(n11706), .ZN(n18901) );
  NOR2_X1 U13114 ( .A1(n11708), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11709) );
  NOR2_X1 U13115 ( .A1(n11725), .A2(n11709), .ZN(n18799) );
  AOI21_X1 U13116 ( .B1(n11710), .B2(n11694), .A(n11711), .ZN(n18775) );
  AOI21_X1 U13117 ( .B1(n11712), .B2(n18747), .A(n11713), .ZN(n18753) );
  AOI21_X1 U13118 ( .B1(n17453), .B2(n11714), .A(n11715), .ZN(n18722) );
  AOI21_X1 U13119 ( .B1(n15793), .B2(n11716), .A(n11720), .ZN(n18700) );
  AOI21_X1 U13120 ( .B1(n18676), .B2(n11719), .A(n11217), .ZN(n18682) );
  AOI21_X1 U13121 ( .B1(n15946), .B2(n11718), .A(n11717), .ZN(n15944) );
  OAI22_X1 U13122 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15673) );
  OAI22_X1 U13123 ( .A1(n11739), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14249), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15672) );
  AND2_X1 U13124 ( .A1(n15673), .A2(n15672), .ZN(n15538) );
  OAI21_X1 U13125 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11718), .ZN(n15539) );
  NAND2_X1 U13126 ( .A1(n15538), .A2(n15539), .ZN(n15942) );
  NOR2_X1 U13127 ( .A1(n15944), .A2(n15942), .ZN(n18669) );
  OAI21_X1 U13128 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11717), .A(
        n11719), .ZN(n18668) );
  NAND2_X1 U13129 ( .A1(n18669), .A2(n18668), .ZN(n18680) );
  NOR2_X1 U13130 ( .A1(n18682), .A2(n18680), .ZN(n18691) );
  OAI21_X1 U13131 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11217), .A(
        n11716), .ZN(n18692) );
  NAND2_X1 U13132 ( .A1(n18691), .A2(n18692), .ZN(n18699) );
  NOR2_X1 U13133 ( .A1(n18700), .A2(n18699), .ZN(n18714) );
  OAI21_X1 U13134 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11720), .A(
        n11714), .ZN(n18715) );
  NAND2_X1 U13135 ( .A1(n18714), .A2(n18715), .ZN(n18721) );
  NOR2_X1 U13136 ( .A1(n18722), .A2(n18721), .ZN(n18737) );
  OAI21_X1 U13137 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11715), .A(
        n11712), .ZN(n18738) );
  NAND2_X1 U13138 ( .A1(n18737), .A2(n18738), .ZN(n18754) );
  NOR2_X1 U13139 ( .A1(n18753), .A2(n18754), .ZN(n18752) );
  OAI21_X1 U13140 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11713), .A(
        n11710), .ZN(n18760) );
  NAND2_X1 U13141 ( .A1(n18752), .A2(n18760), .ZN(n18773) );
  NOR2_X1 U13142 ( .A1(n18775), .A2(n18773), .ZN(n18781) );
  INV_X1 U13143 ( .A(n11708), .ZN(n11724) );
  INV_X1 U13144 ( .A(n11711), .ZN(n11722) );
  INV_X1 U13145 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U13146 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  NAND2_X1 U13147 ( .A1(n11724), .A2(n11723), .ZN(n18782) );
  NAND2_X1 U13148 ( .A1(n18781), .A2(n18782), .ZN(n18797) );
  NOR2_X1 U13149 ( .A1(n18799), .A2(n18797), .ZN(n18808) );
  OAI21_X1 U13150 ( .B1(n11725), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n11726), .ZN(n18811) );
  NAND2_X1 U13151 ( .A1(n18808), .A2(n18811), .ZN(n18819) );
  AOI21_X1 U13152 ( .B1(n11726), .B2(n11695), .A(n11303), .ZN(n18821) );
  OAI21_X1 U13153 ( .B1(n11303), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11727), .ZN(n18840) );
  NAND2_X1 U13154 ( .A1(n18839), .A2(n18840), .ZN(n18838) );
  AOI21_X1 U13155 ( .B1(n16812), .B2(n11727), .A(n11728), .ZN(n16814) );
  INV_X1 U13156 ( .A(n16814), .ZN(n18850) );
  NAND2_X1 U13157 ( .A1(n18849), .A2(n11164), .ZN(n18857) );
  OR2_X1 U13158 ( .A1(n11728), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11730) );
  NAND2_X1 U13159 ( .A1(n11729), .A2(n11730), .ZN(n18858) );
  NAND2_X1 U13160 ( .A1(n18857), .A2(n18858), .ZN(n18856) );
  NAND2_X1 U13161 ( .A1(n11165), .A2(n18856), .ZN(n18867) );
  AOI21_X1 U13162 ( .B1(n16791), .B2(n11729), .A(n11566), .ZN(n16789) );
  INV_X1 U13163 ( .A(n16789), .ZN(n18868) );
  NAND2_X1 U13164 ( .A1(n18867), .A2(n18868), .ZN(n18866) );
  NAND2_X1 U13165 ( .A1(n18866), .A2(n11165), .ZN(n18876) );
  NAND2_X1 U13166 ( .A1(n11731), .A2(n12018), .ZN(n11732) );
  NAND2_X1 U13167 ( .A1(n11734), .A2(n11732), .ZN(n18877) );
  NAND2_X1 U13168 ( .A1(n18876), .A2(n18877), .ZN(n18875) );
  NAND2_X1 U13169 ( .A1(n18875), .A2(n11164), .ZN(n18891) );
  AOI21_X1 U13170 ( .B1(n18885), .B2(n11734), .A(n11733), .ZN(n16757) );
  INV_X1 U13171 ( .A(n16757), .ZN(n18892) );
  NAND2_X1 U13172 ( .A1(n18891), .A2(n18892), .ZN(n18890) );
  NAND2_X1 U13173 ( .A1(n11164), .A2(n18890), .ZN(n18900) );
  AND2_X1 U13174 ( .A1(n11735), .A2(n16729), .ZN(n11736) );
  OR2_X1 U13175 ( .A1(n11736), .A2(n11703), .ZN(n18917) );
  NOR2_X1 U13176 ( .A1(n18809), .A2(n18930), .ZN(n18941) );
  NOR2_X1 U13177 ( .A1(n18942), .A2(n18941), .ZN(n18940) );
  NOR2_X1 U13178 ( .A1(n18809), .A2(n18940), .ZN(n18959) );
  NOR2_X1 U13179 ( .A1(n18960), .A2(n18959), .ZN(n18979) );
  NOR2_X1 U13180 ( .A1(n18809), .A2(n18979), .ZN(n11738) );
  XOR2_X1 U13181 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n11737), .Z(
        n18978) );
  XNOR2_X1 U13182 ( .A(n11738), .B(n18978), .ZN(n11740) );
  INV_X1 U13183 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11739) );
  INV_X1 U13184 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19594) );
  INV_X1 U13185 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22141) );
  NAND4_X1 U13186 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n11739), .A3(n19594), 
        .A4(n22141), .ZN(n19039) );
  NAND2_X1 U13187 ( .A1(n11740), .A2(n18980), .ZN(n12456) );
  NOR2_X4 U13188 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14724) );
  AND2_X4 U13189 ( .A1(n14724), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13937) );
  AOI22_X1 U13190 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11745) );
  AND3_X4 U13191 ( .A1(n14722), .A2(n11741), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12084) );
  AND3_X4 U13192 ( .A1(n12073), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U13193 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11744) );
  AND2_X4 U13194 ( .A1(n14785), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13943) );
  AOI22_X1 U13195 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U13196 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U13197 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  NAND2_X1 U13198 ( .A1(n11746), .A2(n14755), .ZN(n11755) );
  AOI22_X1 U13199 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U13200 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U13201 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U13202 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U13203 ( .A1(n11199), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11747) );
  AND2_X1 U13204 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND4_X1 U13205 ( .A1(n11752), .A2(n11751), .A3(n11750), .A4(n11749), .ZN(
        n11753) );
  NAND2_X1 U13206 ( .A1(n11753), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11754) );
  AOI22_X1 U13207 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U13208 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11759) );
  NAND2_X1 U13209 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11757) );
  NAND4_X1 U13210 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11762) );
  NAND2_X1 U13211 ( .A1(n11762), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11769) );
  AOI22_X1 U13212 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U13213 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U13214 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U13215 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11199), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U13216 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11767) );
  NAND2_X1 U13217 ( .A1(n11767), .A2(n14755), .ZN(n11768) );
  AOI22_X1 U13218 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13219 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U13220 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11776) );
  NAND2_X1 U13221 ( .A1(n11776), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11785) );
  AOI22_X1 U13222 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11781) );
  NAND2_X1 U13223 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U13224 ( .A1(n12082), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11777) );
  NAND4_X1 U13225 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  NAND2_X1 U13226 ( .A1(n11783), .A2(n14755), .ZN(n11784) );
  AOI22_X1 U13227 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U13228 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11789) );
  NAND3_X1 U13229 ( .A1(n11262), .A2(n11790), .A3(n11789), .ZN(n11798) );
  AOI22_X1 U13230 ( .A1(n11214), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12072), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U13231 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13943), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U13232 ( .A1(n11163), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12072), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U13233 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13234 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13943), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U13235 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  AOI22_X1 U13236 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13237 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U13238 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11161), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U13239 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11199), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11804) );
  NAND4_X1 U13240 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11808) );
  INV_X1 U13241 ( .A(n11866), .ZN(n11811) );
  NAND2_X2 U13242 ( .A1(n13761), .A2(n11811), .ZN(n11889) );
  NAND2_X1 U13243 ( .A1(n11889), .A2(n14352), .ZN(n11837) );
  AOI22_X1 U13244 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U13245 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U13246 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U13247 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11200), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U13248 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11816) );
  NAND2_X1 U13249 ( .A1(n11816), .A2(n14755), .ZN(n11823) );
  AOI22_X1 U13250 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U13251 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11817) );
  NAND4_X1 U13252 ( .A1(n11820), .A2(n11819), .A3(n11818), .A4(n11817), .ZN(
        n11821) );
  NAND2_X1 U13253 ( .A1(n11821), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11822) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13943), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U13255 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U13256 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11205), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U13257 ( .A1(n12072), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12082), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11824) );
  NAND4_X1 U13258 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11828) );
  NAND2_X1 U13259 ( .A1(n11828), .A2(n14755), .ZN(n11836) );
  AOI22_X1 U13260 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U13261 ( .A1(n11202), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12082), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U13262 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11829) );
  NAND3_X1 U13263 ( .A1(n11831), .A2(n11830), .A3(n11829), .ZN(n11834) );
  AOI22_X1 U13264 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n13943), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11832) );
  INV_X1 U13265 ( .A(n11832), .ZN(n11833) );
  AOI22_X1 U13266 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11214), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U13267 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U13268 ( .A1(n12084), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13940), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U13269 ( .A1(n13943), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U13270 ( .A1(n13937), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11210), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11848) );
  NAND3_X1 U13271 ( .A1(n11683), .A2(n11849), .A3(n11848), .ZN(n11850) );
  NAND2_X1 U13272 ( .A1(n12065), .A2(n12609), .ZN(n11863) );
  INV_X1 U13273 ( .A(n11855), .ZN(n11857) );
  INV_X2 U13274 ( .A(n13761), .ZN(n11881) );
  NAND4_X1 U13275 ( .A1(n11852), .A2(n11857), .A3(n11856), .A4(n11881), .ZN(
        n11897) );
  NAND3_X1 U13276 ( .A1(n19828), .A2(n11881), .A3(n14921), .ZN(n11858) );
  NAND3_X1 U13277 ( .A1(n11860), .A2(n11811), .A3(n11890), .ZN(n11874) );
  AND2_X1 U13278 ( .A1(n11880), .A2(n11861), .ZN(n11862) );
  NAND2_X1 U13279 ( .A1(n14774), .A2(n11862), .ZN(n14148) );
  NAND4_X1 U13280 ( .A1(n14375), .A2(n11863), .A3(n11897), .A4(n14148), .ZN(
        n11864) );
  NAND2_X1 U13281 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11873) );
  NOR2_X1 U13282 ( .A1(n11923), .A2(n11893), .ZN(n11868) );
  INV_X1 U13283 ( .A(n11890), .ZN(n19528) );
  INV_X1 U13284 ( .A(n11892), .ZN(n14344) );
  INV_X1 U13285 ( .A(n11902), .ZN(n12043) );
  AOI22_X1 U13286 ( .A1(n16012), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11871) );
  NAND2_X1 U13287 ( .A1(n12045), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11870) );
  AND2_X1 U13288 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  NAND2_X1 U13289 ( .A1(n11873), .A2(n11872), .ZN(n16010) );
  INV_X1 U13290 ( .A(n11874), .ZN(n11876) );
  NAND3_X1 U13291 ( .A1(n11876), .A2(n11875), .A3(n11881), .ZN(n12750) );
  NAND3_X1 U13292 ( .A1(n12750), .A2(n12069), .A3(n11877), .ZN(n11878) );
  NAND2_X1 U13293 ( .A1(n11878), .A2(n14316), .ZN(n14120) );
  INV_X1 U13294 ( .A(n14120), .ZN(n11879) );
  NAND2_X1 U13295 ( .A1(n11854), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14117) );
  NAND2_X1 U13296 ( .A1(n11879), .A2(n14300), .ZN(n11887) );
  INV_X1 U13297 ( .A(n11880), .ZN(n14776) );
  NAND2_X1 U13298 ( .A1(n11882), .A2(n11877), .ZN(n11883) );
  NAND2_X1 U13299 ( .A1(n14776), .A2(n11883), .ZN(n11884) );
  NAND2_X1 U13300 ( .A1(n11884), .A2(n14774), .ZN(n14342) );
  NOR2_X1 U13301 ( .A1(n11854), .A2(n11739), .ZN(n11885) );
  AND2_X2 U13302 ( .A1(n11887), .A2(n11886), .ZN(n11914) );
  NAND2_X1 U13303 ( .A1(n14325), .A2(n19828), .ZN(n14322) );
  NAND2_X1 U13304 ( .A1(n11889), .A2(n11888), .ZN(n14320) );
  NOR2_X1 U13305 ( .A1(n11893), .A2(n11739), .ZN(n11894) );
  NAND2_X1 U13306 ( .A1(n11910), .A2(n11894), .ZN(n11895) );
  NAND2_X1 U13307 ( .A1(n11917), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11901) );
  INV_X1 U13308 ( .A(n12065), .ZN(n11896) );
  NAND2_X1 U13309 ( .A1(n11896), .A2(n14148), .ZN(n12421) );
  INV_X1 U13310 ( .A(n12421), .ZN(n11898) );
  NAND2_X1 U13311 ( .A1(n11898), .A2(n11897), .ZN(n14373) );
  NOR2_X1 U13312 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11940) );
  AOI21_X1 U13313 ( .B1(n14373), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11899), 
        .ZN(n11900) );
  NAND2_X1 U13314 ( .A1(n11901), .A2(n11900), .ZN(n11908) );
  INV_X1 U13315 ( .A(n11908), .ZN(n11906) );
  NAND2_X1 U13316 ( .A1(n11913), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U13317 ( .A1(n11902), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11903) );
  INV_X1 U13318 ( .A(n11907), .ZN(n11905) );
  NAND2_X1 U13319 ( .A1(n11908), .A2(n11907), .ZN(n11909) );
  NAND2_X1 U13320 ( .A1(n11937), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11916) );
  NAND3_X1 U13321 ( .A1(n11910), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14349), 
        .ZN(n11915) );
  INV_X1 U13322 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U13323 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11911) );
  INV_X1 U13324 ( .A(n11940), .ZN(n19032) );
  NAND2_X1 U13325 ( .A1(n11918), .A2(n11741), .ZN(n11919) );
  NAND2_X1 U13326 ( .A1(n11917), .A2(n11919), .ZN(n11928) );
  INV_X1 U13327 ( .A(n11893), .ZN(n14102) );
  NAND2_X1 U13328 ( .A1(n11919), .A2(n14102), .ZN(n11922) );
  NAND2_X1 U13329 ( .A1(n11922), .A2(n11921), .ZN(n11926) );
  NOR2_X1 U13330 ( .A1(n11923), .A2(n11739), .ZN(n11925) );
  AOI21_X1 U13331 ( .B1(n11926), .B2(n11925), .A(n11924), .ZN(n11927) );
  NAND2_X1 U13332 ( .A1(n11928), .A2(n11927), .ZN(n12465) );
  NAND2_X1 U13333 ( .A1(n11937), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U13334 ( .A1(n11913), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U13335 ( .A1(n11902), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11929) );
  OAI21_X1 U13336 ( .B1(n19592), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14913), 
        .ZN(n11932) );
  INV_X1 U13337 ( .A(n11934), .ZN(n11933) );
  INV_X1 U13338 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19030) );
  AOI22_X1 U13339 ( .A1(n11902), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U13340 ( .A1(n11913), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11938) );
  NAND2_X1 U13341 ( .A1(n11917), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U13342 ( .A1(n11940), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U13343 ( .A1(n11942), .A2(n11941), .ZN(n11946) );
  NAND2_X1 U13344 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  INV_X1 U13345 ( .A(n12458), .ZN(n11948) );
  INV_X1 U13346 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U13347 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11951) );
  AOI22_X1 U13348 ( .A1(n16012), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11950) );
  OAI211_X1 U13349 ( .C1(n16014), .C2(n11952), .A(n11951), .B(n11950), .ZN(
        n14534) );
  NAND2_X1 U13350 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11958) );
  INV_X1 U13351 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U13352 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11954) );
  NAND2_X1 U13353 ( .A1(n11902), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11953) );
  OAI211_X1 U13354 ( .C1(n16014), .C2(n11955), .A(n11954), .B(n11953), .ZN(
        n11956) );
  INV_X1 U13355 ( .A(n11956), .ZN(n11957) );
  NAND2_X1 U13356 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11964) );
  INV_X1 U13357 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U13358 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U13359 ( .A1(n16012), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11959) );
  OAI211_X1 U13360 ( .C1(n16014), .C2(n11961), .A(n11960), .B(n11959), .ZN(
        n11962) );
  INV_X1 U13361 ( .A(n11962), .ZN(n11963) );
  NAND2_X1 U13362 ( .A1(n11964), .A2(n11963), .ZN(n14573) );
  NAND2_X1 U13363 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11967) );
  INV_X1 U13364 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12436) );
  INV_X1 U13365 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14913) );
  OAI22_X1 U13366 ( .A1(n12043), .A2(n12436), .B1(n14913), .B2(n15793), .ZN(
        n11965) );
  AOI21_X1 U13367 ( .B1(n12045), .B2(P2_REIP_REG_7__SCAN_IN), .A(n11965), .ZN(
        n11966) );
  INV_X1 U13368 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U13369 ( .A1(n16012), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U13370 ( .A1(n12045), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11968) );
  OAI211_X1 U13371 ( .C1(n12037), .C2(n12628), .A(n11969), .B(n11968), .ZN(
        n14606) );
  INV_X1 U13372 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U13373 ( .A1(n16012), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11971) );
  NAND2_X1 U13374 ( .A1(n12045), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11970) );
  OAI211_X1 U13375 ( .C1(n12037), .C2(n16884), .A(n11971), .B(n11970), .ZN(
        n14656) );
  NAND2_X1 U13376 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11975) );
  AOI22_X1 U13377 ( .A1(n16012), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11973) );
  NAND2_X1 U13378 ( .A1(n12045), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11972) );
  AND2_X1 U13379 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  NAND2_X1 U13380 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11980) );
  INV_X1 U13381 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11977) );
  OAI22_X1 U13382 ( .A1(n12043), .A2(n11977), .B1(n14913), .B2(n18747), .ZN(
        n11978) );
  AOI21_X1 U13383 ( .B1(n12045), .B2(P2_REIP_REG_11__SCAN_IN), .A(n11978), 
        .ZN(n11979) );
  NAND2_X1 U13384 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11986) );
  INV_X1 U13385 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11983) );
  INV_X1 U13386 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11982) );
  OAI22_X1 U13387 ( .A1(n12043), .A2(n11983), .B1(n14913), .B2(n11982), .ZN(
        n11984) );
  AOI21_X1 U13388 ( .B1(n12045), .B2(P2_REIP_REG_12__SCAN_IN), .A(n11984), 
        .ZN(n11985) );
  INV_X1 U13389 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U13390 ( .A1(n16012), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11988) );
  NAND2_X1 U13391 ( .A1(n12045), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11987) );
  OAI211_X1 U13392 ( .C1(n12037), .C2(n17099), .A(n11988), .B(n11987), .ZN(
        n14940) );
  NAND2_X1 U13393 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11992) );
  AOI22_X1 U13394 ( .A1(n16012), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11990) );
  NAND2_X1 U13395 ( .A1(n12045), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11989) );
  AND2_X1 U13396 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  NAND2_X1 U13397 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11995) );
  INV_X1 U13398 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12440) );
  INV_X1 U13399 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18793) );
  OAI22_X1 U13400 ( .A1(n12043), .A2(n12440), .B1(n14913), .B2(n18793), .ZN(
        n11993) );
  AOI21_X1 U13401 ( .B1(n12045), .B2(P2_REIP_REG_15__SCAN_IN), .A(n11993), 
        .ZN(n11994) );
  INV_X1 U13402 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U13403 ( .A1(n16012), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11998) );
  NAND2_X1 U13404 ( .A1(n12045), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11997) );
  OAI211_X1 U13405 ( .C1(n12037), .C2(n12658), .A(n11998), .B(n11997), .ZN(
        n15578) );
  NAND2_X1 U13406 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12002) );
  AOI22_X1 U13407 ( .A1(n16012), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12000) );
  NAND2_X1 U13408 ( .A1(n12045), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11999) );
  AND2_X1 U13409 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  NAND2_X1 U13410 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12005) );
  INV_X1 U13411 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18832) );
  OAI22_X1 U13412 ( .A1(n12043), .A2(n18832), .B1(n14913), .B2(n11565), .ZN(
        n12003) );
  AOI21_X1 U13413 ( .B1(n12045), .B2(P2_REIP_REG_18__SCAN_IN), .A(n12003), 
        .ZN(n12004) );
  AND2_X1 U13414 ( .A1(n12005), .A2(n12004), .ZN(n15770) );
  NAND2_X1 U13415 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12011) );
  INV_X1 U13416 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17560) );
  NAND2_X1 U13417 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U13418 ( .A1(n16012), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12007) );
  OAI211_X1 U13419 ( .C1(n16014), .C2(n17560), .A(n12008), .B(n12007), .ZN(
        n12009) );
  INV_X1 U13420 ( .A(n12009), .ZN(n12010) );
  INV_X1 U13421 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U13422 ( .A1(n16012), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12013) );
  NAND2_X1 U13423 ( .A1(n12045), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12012) );
  OAI211_X1 U13424 ( .C1(n12037), .C2(n17012), .A(n12013), .B(n12012), .ZN(
        n15805) );
  NAND2_X1 U13425 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12017) );
  INV_X1 U13426 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12014) );
  OAI22_X1 U13427 ( .A1(n12043), .A2(n12014), .B1(n14913), .B2(n16791), .ZN(
        n12015) );
  AOI21_X1 U13428 ( .B1(n12045), .B2(P2_REIP_REG_21__SCAN_IN), .A(n12015), 
        .ZN(n12016) );
  AND2_X1 U13429 ( .A1(n12017), .A2(n12016), .ZN(n16594) );
  NAND2_X1 U13430 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12022) );
  INV_X1 U13431 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12019) );
  OAI22_X1 U13432 ( .A1(n12043), .A2(n12019), .B1(n14913), .B2(n12018), .ZN(
        n12020) );
  AOI21_X1 U13433 ( .B1(n12045), .B2(P2_REIP_REG_22__SCAN_IN), .A(n12020), 
        .ZN(n12021) );
  AND2_X1 U13434 ( .A1(n12022), .A2(n12021), .ZN(n16589) );
  INV_X1 U13435 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U13436 ( .A1(n16012), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12024) );
  NAND2_X1 U13437 ( .A1(n12045), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12023) );
  OAI211_X1 U13438 ( .C1(n12037), .C2(n16964), .A(n12024), .B(n12023), .ZN(
        n16580) );
  INV_X1 U13439 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U13440 ( .A1(n16012), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12026) );
  NAND2_X1 U13441 ( .A1(n12045), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U13442 ( .C1(n12037), .C2(n16952), .A(n12026), .B(n12025), .ZN(
        n16577) );
  NAND2_X1 U13443 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12030) );
  INV_X1 U13444 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12027) );
  OAI22_X1 U13445 ( .A1(n12043), .A2(n12027), .B1(n14913), .B2(n16739), .ZN(
        n12028) );
  AOI21_X1 U13446 ( .B1(n12045), .B2(P2_REIP_REG_25__SCAN_IN), .A(n12028), 
        .ZN(n12029) );
  AND2_X1 U13447 ( .A1(n12030), .A2(n12029), .ZN(n16570) );
  NAND2_X1 U13448 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12034) );
  INV_X1 U13449 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12031) );
  OAI22_X1 U13450 ( .A1(n12043), .A2(n12031), .B1(n14913), .B2(n16729), .ZN(
        n12032) );
  AOI21_X1 U13451 ( .B1(n12045), .B2(P2_REIP_REG_26__SCAN_IN), .A(n12032), 
        .ZN(n12033) );
  AND2_X1 U13452 ( .A1(n12034), .A2(n12033), .ZN(n16557) );
  INV_X1 U13453 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U13454 ( .A1(n16012), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12036) );
  NAND2_X1 U13455 ( .A1(n12045), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12035) );
  OAI211_X1 U13456 ( .C1(n12037), .C2(n16893), .A(n12036), .B(n12035), .ZN(
        n16554) );
  NAND2_X1 U13457 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12041) );
  AOI22_X1 U13458 ( .A1(n16012), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12039) );
  NAND2_X1 U13459 ( .A1(n12045), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12038) );
  AND2_X1 U13460 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  AND2_X1 U13461 ( .A1(n12041), .A2(n12040), .ZN(n16546) );
  NAND2_X1 U13462 ( .A1(n11865), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12047) );
  INV_X1 U13463 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12042) );
  INV_X1 U13464 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12801) );
  OAI22_X1 U13465 ( .A1(n12043), .A2(n12042), .B1(n14913), .B2(n12801), .ZN(
        n12044) );
  AOI21_X1 U13466 ( .B1(n12045), .B2(P2_REIP_REG_29__SCAN_IN), .A(n12044), 
        .ZN(n12046) );
  AND2_X1 U13467 ( .A1(n12047), .A2(n12046), .ZN(n12796) );
  INV_X1 U13468 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19563) );
  XNOR2_X1 U13469 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U13470 ( .A1(n12753), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U13471 ( .A1(n19689), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U13472 ( .A1(n12061), .A2(n12048), .ZN(n12058) );
  XNOR2_X1 U13473 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U13474 ( .A1(n12058), .A2(n12057), .ZN(n12050) );
  NAND2_X1 U13475 ( .A1(n19592), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12049) );
  NAND2_X1 U13476 ( .A1(n12050), .A2(n12049), .ZN(n12054) );
  INV_X1 U13477 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18987) );
  INV_X1 U13478 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17343) );
  NOR2_X1 U13479 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17343), .ZN(
        n12051) );
  AOI221_X1 U13480 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12052), 
        .C1(n18987), .C2(n12052), .A(n12051), .ZN(n14118) );
  NAND3_X1 U13481 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12052), .A3(
        n18987), .ZN(n14096) );
  NOR2_X1 U13482 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  OR2_X1 U13483 ( .A1(n12056), .A2(n12055), .ZN(n14109) );
  XNOR2_X1 U13484 ( .A(n12058), .B(n12057), .ZN(n14108) );
  INV_X1 U13485 ( .A(n12753), .ZN(n12060) );
  INV_X1 U13486 ( .A(n12059), .ZN(n12571) );
  NAND2_X1 U13487 ( .A1(n12060), .A2(n12571), .ZN(n12062) );
  NAND2_X1 U13488 ( .A1(n12062), .A2(n12061), .ZN(n14103) );
  NOR3_X1 U13489 ( .A1(n14109), .A2(n14108), .A3(n14103), .ZN(n12063) );
  AND2_X1 U13490 ( .A1(n14096), .A2(n12063), .ZN(n12064) );
  OR2_X1 U13491 ( .A1(n14118), .A2(n12064), .ZN(n14759) );
  AND3_X1 U13492 ( .A1(n14913), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18631) );
  NAND2_X1 U13493 ( .A1(n12065), .A2(n18631), .ZN(n12066) );
  NOR2_X1 U13494 ( .A1(n14759), .A2(n12066), .ZN(n14152) );
  NAND2_X1 U13495 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n22174) );
  AND2_X1 U13496 ( .A1(n12069), .A2(n22174), .ZN(n12067) );
  AND2_X1 U13497 ( .A1(n14152), .A2(n12067), .ZN(n14221) );
  NOR2_X1 U13498 ( .A1(n15617), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12115) );
  INV_X2 U13499 ( .A(n12398), .ZN(n16025) );
  AOI222_X1 U13500 ( .A1(n12093), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n16025), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n11166), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12420) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15670) );
  INV_X1 U13502 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13899) );
  OAI22_X1 U13503 ( .A1(n13896), .A2(n15670), .B1(n13877), .B2(n13899), .ZN(
        n12071) );
  INV_X1 U13504 ( .A(n12071), .ZN(n12081) );
  AND2_X2 U13505 ( .A1(n13943), .A2(n14755), .ZN(n13917) );
  AOI22_X1 U13506 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12080) );
  INV_X1 U13507 ( .A(n12072), .ZN(n13944) );
  AOI22_X1 U13508 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12079) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U13510 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12076) );
  AND2_X1 U13511 ( .A1(n12073), .A2(n11196), .ZN(n12074) );
  NAND2_X1 U13512 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12075) );
  OAI211_X1 U13513 ( .C1(n13894), .C2(n12599), .A(n12076), .B(n12075), .ZN(
        n12077) );
  INV_X1 U13514 ( .A(n12077), .ZN(n12078) );
  NAND4_X1 U13515 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n12092) );
  NAND2_X2 U13516 ( .A1(n12083), .A2(n14755), .ZN(n13926) );
  AOI22_X1 U13517 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13906), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U13518 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12089) );
  AND2_X1 U13519 ( .A1(n11741), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12086) );
  AOI22_X1 U13520 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U13521 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12087) );
  NAND4_X1 U13522 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n12087), .ZN(
        n12091) );
  NAND2_X1 U13523 ( .A1(n12093), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12095) );
  INV_X1 U13524 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n17511) );
  NAND2_X1 U13525 ( .A1(n12069), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12094) );
  AOI22_X1 U13526 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13527 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U13528 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U13529 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12097) );
  AND4_X1 U13530 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12113) );
  AOI22_X1 U13531 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12105) );
  NAND2_X1 U13532 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U13533 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U13534 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12102) );
  NAND4_X1 U13535 ( .A1(n12105), .A2(n12104), .A3(n12103), .A4(n12102), .ZN(
        n12111) );
  NAND2_X1 U13536 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12109) );
  NAND2_X1 U13537 ( .A1(n13906), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12108) );
  NAND2_X1 U13538 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12107) );
  NAND2_X1 U13539 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12106) );
  NAND4_X1 U13540 ( .A1(n12109), .A2(n12108), .A3(n12107), .A4(n12106), .ZN(
        n12110) );
  NOR2_X1 U13541 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  INV_X1 U13542 ( .A(n11889), .ZN(n14401) );
  NAND2_X1 U13543 ( .A1(n14401), .A2(n16024), .ZN(n12158) );
  MUX2_X1 U13544 ( .A(n15617), .B(n19612), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12114) );
  INV_X1 U13545 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17548) );
  NAND2_X1 U13546 ( .A1(n12093), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12117) );
  INV_X1 U13547 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U13548 ( .A1(n12115), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n16024), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12116) );
  NAND2_X1 U13549 ( .A1(n12117), .A2(n12116), .ZN(n12140) );
  INV_X1 U13550 ( .A(n12140), .ZN(n12118) );
  AND2_X1 U13551 ( .A1(n11889), .A2(n15617), .ZN(n14398) );
  MUX2_X1 U13552 ( .A(n14398), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n12139) );
  AOI22_X1 U13553 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U13554 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U13555 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12120) );
  NAND2_X1 U13556 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12119) );
  NAND4_X1 U13557 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12119), .ZN(
        n12128) );
  NAND2_X1 U13558 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U13559 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12125) );
  NAND2_X1 U13560 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U13561 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12123) );
  NAND4_X1 U13562 ( .A1(n12126), .A2(n12125), .A3(n12124), .A4(n12123), .ZN(
        n12127) );
  NOR2_X1 U13563 ( .A1(n12128), .A2(n12127), .ZN(n12137) );
  AOI22_X1 U13564 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U13565 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U13566 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U13567 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12129) );
  NAND4_X1 U13568 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12135) );
  INV_X1 U13569 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12133) );
  INV_X1 U13570 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12514) );
  OAI22_X1 U13571 ( .A1(n13926), .A2(n12133), .B1(n13924), .B2(n12514), .ZN(
        n12134) );
  NOR2_X1 U13572 ( .A1(n12135), .A2(n12134), .ZN(n12136) );
  NOR2_X1 U13573 ( .A1(n12372), .A2(n12759), .ZN(n12138) );
  NOR2_X1 U13574 ( .A1(n12139), .A2(n12138), .ZN(n14405) );
  NAND2_X1 U13575 ( .A1(n14406), .A2(n14405), .ZN(n14407) );
  AOI22_X1 U13576 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U13577 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U13578 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12142) );
  AND2_X1 U13579 ( .A1(n12143), .A2(n12142), .ZN(n12147) );
  AOI22_X1 U13580 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U13581 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U13582 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12157) );
  INV_X1 U13583 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12150) );
  INV_X1 U13584 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12149) );
  OAI22_X1 U13585 ( .A1(n13926), .A2(n12150), .B1(n13924), .B2(n12149), .ZN(
        n12151) );
  INV_X1 U13586 ( .A(n12151), .ZN(n12155) );
  AOI22_X1 U13587 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13588 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12153) );
  NAND2_X1 U13589 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12152) );
  NAND4_X1 U13590 ( .A1(n12155), .A2(n12154), .A3(n12153), .A4(n12152), .ZN(
        n12156) );
  INV_X1 U13591 ( .A(n12764), .ZN(n12526) );
  OR2_X1 U13592 ( .A1(n12372), .A2(n12526), .ZN(n12159) );
  OAI211_X1 U13593 ( .C1(n19593), .C2(n19592), .A(n12159), .B(n12158), .ZN(
        n12160) );
  AND3_X1 U13594 ( .A1(n14407), .A2(n12161), .A3(n12160), .ZN(n12162) );
  NAND2_X1 U13595 ( .A1(n12093), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U13596 ( .A1(n16025), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11166), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U13597 ( .A1(n12165), .A2(n12164), .ZN(n14366) );
  NOR2_X1 U13598 ( .A1(n14368), .A2(n14366), .ZN(n12166) );
  NAND2_X1 U13599 ( .A1(n12093), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13600 ( .A1(n16025), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12186) );
  INV_X1 U13601 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12480) );
  INV_X1 U13602 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12471) );
  OAI22_X1 U13603 ( .A1(n13896), .A2(n12480), .B1(n13894), .B2(n12471), .ZN(
        n12168) );
  INV_X1 U13604 ( .A(n12168), .ZN(n12175) );
  AOI22_X1 U13605 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U13606 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12173) );
  INV_X1 U13607 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13850) );
  NAND2_X1 U13608 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12170) );
  NAND2_X1 U13609 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12169) );
  OAI211_X1 U13610 ( .C1(n13877), .C2(n13850), .A(n12170), .B(n12169), .ZN(
        n12171) );
  INV_X1 U13611 ( .A(n12171), .ZN(n12172) );
  NAND4_X1 U13612 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n12182) );
  AOI22_X1 U13613 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13906), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U13614 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U13615 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12178) );
  NAND2_X1 U13616 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12177) );
  NAND4_X1 U13617 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12181) );
  INV_X1 U13618 ( .A(n12507), .ZN(n12183) );
  OR2_X1 U13619 ( .A1(n12372), .A2(n12183), .ZN(n12185) );
  NAND2_X1 U13620 ( .A1(n11166), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12184) );
  NAND4_X1 U13621 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n14689) );
  NAND2_X1 U13622 ( .A1(n14690), .A2(n14689), .ZN(n14691) );
  NAND2_X1 U13623 ( .A1(n12093), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U13624 ( .A1(n16025), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11166), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12205) );
  INV_X1 U13625 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12189) );
  INV_X1 U13626 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12188) );
  OAI22_X1 U13627 ( .A1(n13896), .A2(n12189), .B1(n13894), .B2(n12188), .ZN(
        n12190) );
  INV_X1 U13628 ( .A(n12190), .ZN(n12197) );
  AOI22_X1 U13629 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U13630 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12195) );
  INV_X1 U13631 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13865) );
  NAND2_X1 U13632 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U13633 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12191) );
  OAI211_X1 U13634 ( .C1(n13877), .C2(n13865), .A(n12192), .B(n12191), .ZN(
        n12193) );
  INV_X1 U13635 ( .A(n12193), .ZN(n12194) );
  NAND4_X1 U13636 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12203) );
  AOI22_X1 U13637 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13906), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13638 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U13639 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U13640 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12198) );
  NAND4_X1 U13641 ( .A1(n12201), .A2(n12200), .A3(n12199), .A4(n12198), .ZN(
        n12202) );
  OR2_X1 U13642 ( .A1(n12372), .A2(n12770), .ZN(n12204) );
  AOI22_X1 U13643 ( .A1(n12093), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n16025), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12223) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12536) );
  INV_X1 U13645 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12552) );
  OAI22_X1 U13646 ( .A1(n13896), .A2(n12536), .B1(n13894), .B2(n12552), .ZN(
        n12207) );
  INV_X1 U13647 ( .A(n12207), .ZN(n12214) );
  AOI22_X1 U13648 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U13649 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12212) );
  INV_X1 U13650 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13884) );
  NAND2_X1 U13651 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12209) );
  NAND2_X1 U13652 ( .A1(n13913), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12208) );
  OAI211_X1 U13653 ( .C1(n13877), .C2(n13884), .A(n12209), .B(n12208), .ZN(
        n12210) );
  INV_X1 U13654 ( .A(n12210), .ZN(n12211) );
  NAND4_X1 U13655 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12220) );
  AOI22_X1 U13656 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13906), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U13657 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U13658 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U13659 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12215) );
  NAND4_X1 U13660 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  INV_X1 U13661 ( .A(n12434), .ZN(n12559) );
  INV_X1 U13662 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15642) );
  OAI22_X1 U13663 ( .A1(n12372), .A2(n12559), .B1(n12355), .B2(n15642), .ZN(
        n12221) );
  INV_X1 U13664 ( .A(n12221), .ZN(n12222) );
  NAND2_X1 U13665 ( .A1(n12223), .A2(n12222), .ZN(n15648) );
  NAND2_X1 U13666 ( .A1(n14832), .A2(n15648), .ZN(n15647) );
  NAND2_X1 U13667 ( .A1(n12093), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U13668 ( .A1(n16025), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11166), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U13669 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12096), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U13670 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12229) );
  NAND2_X1 U13671 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12228) );
  NAND2_X1 U13672 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12227) );
  NAND4_X1 U13673 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12236) );
  NAND2_X1 U13674 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12234) );
  NAND2_X1 U13675 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12233) );
  NAND2_X1 U13676 ( .A1(n13906), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12232) );
  NAND2_X1 U13677 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12231) );
  NAND4_X1 U13678 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12235) );
  NOR2_X1 U13679 ( .A1(n12236), .A2(n12235), .ZN(n12248) );
  AOI22_X1 U13680 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12101), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U13681 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U13682 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12238) );
  NAND2_X1 U13683 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12237) );
  NAND4_X1 U13684 ( .A1(n12240), .A2(n12239), .A3(n12238), .A4(n12237), .ZN(
        n12246) );
  INV_X1 U13685 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12244) );
  INV_X1 U13686 ( .A(n12241), .ZN(n12243) );
  INV_X1 U13687 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12242) );
  OAI22_X1 U13688 ( .A1(n12244), .A2(n12243), .B1(n13926), .B2(n12242), .ZN(
        n12245) );
  NOR2_X1 U13689 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  INV_X1 U13690 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15788) );
  INV_X1 U13691 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17524) );
  INV_X1 U13692 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17551) );
  OAI222_X1 U13693 ( .A1(n12355), .A2(n15788), .B1(n12398), .B2(n17524), .C1(
        n12163), .C2(n17551), .ZN(n14496) );
  AOI22_X1 U13694 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13914), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13695 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12365), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U13696 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U13697 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12249) );
  AND2_X1 U13698 ( .A1(n12250), .A2(n12249), .ZN(n12252) );
  AOI22_X1 U13699 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U13700 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12260) );
  AOI22_X1 U13701 ( .A1(n13906), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U13702 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U13703 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U13704 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12255) );
  NAND4_X1 U13705 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12259) );
  OR2_X1 U13706 ( .A1(n12260), .A2(n12259), .ZN(n14608) );
  INV_X1 U13707 ( .A(n14608), .ZN(n12262) );
  AOI22_X1 U13708 ( .A1(n16025), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11166), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12261) );
  OAI21_X1 U13709 ( .B1(n12262), .B2(n12372), .A(n12261), .ZN(n12263) );
  AOI21_X1 U13710 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(n12093), .A(n12263), .ZN(
        n14583) );
  AOI22_X1 U13711 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U13712 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12266) );
  NAND2_X1 U13713 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12265) );
  NAND2_X1 U13714 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12264) );
  NAND4_X1 U13715 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12273) );
  NAND2_X1 U13716 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12271) );
  NAND2_X1 U13717 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U13718 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U13719 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12268) );
  NAND4_X1 U13720 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  NOR2_X1 U13721 ( .A1(n12273), .A2(n12272), .ZN(n12282) );
  AOI22_X1 U13722 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U13723 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12276) );
  NAND2_X1 U13724 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12275) );
  NAND2_X1 U13725 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12274) );
  NAND4_X1 U13726 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12280) );
  INV_X1 U13727 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12518) );
  INV_X1 U13728 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12278) );
  OAI22_X1 U13729 ( .A1(n13926), .A2(n12518), .B1(n13924), .B2(n12278), .ZN(
        n12279) );
  NOR2_X1 U13730 ( .A1(n12280), .A2(n12279), .ZN(n12281) );
  AND2_X1 U13731 ( .A1(n12282), .A2(n12281), .ZN(n14653) );
  NAND2_X1 U13732 ( .A1(n12093), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U13733 ( .A1(n16025), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11166), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12283) );
  OAI211_X1 U13734 ( .C1(n14653), .C2(n12372), .A(n12284), .B(n12283), .ZN(
        n14625) );
  AOI22_X1 U13735 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13914), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U13736 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13906), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U13737 ( .A1(n13929), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U13738 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12285) );
  AND2_X1 U13739 ( .A1(n12286), .A2(n12285), .ZN(n12288) );
  AOI22_X1 U13740 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U13741 ( .A1(n12290), .A2(n12289), .A3(n12288), .A4(n12287), .ZN(
        n12296) );
  AOI22_X1 U13742 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U13743 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U13744 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12096), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U13745 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12291) );
  NAND4_X1 U13746 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12295) );
  NOR2_X1 U13747 ( .A1(n12296), .A2(n12295), .ZN(n14711) );
  NAND2_X1 U13748 ( .A1(n12093), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U13749 ( .A1(n16025), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12297) );
  OAI211_X1 U13750 ( .C1(n14711), .C2(n12372), .A(n12298), .B(n12297), .ZN(
        n14661) );
  AOI22_X1 U13751 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U13752 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12301) );
  NAND2_X1 U13753 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12300) );
  NAND2_X1 U13754 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12299) );
  NAND4_X1 U13755 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12308) );
  NAND2_X1 U13756 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12306) );
  NAND2_X1 U13757 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12305) );
  NAND2_X1 U13758 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U13759 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12303) );
  NAND4_X1 U13760 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12307) );
  NOR2_X1 U13761 ( .A1(n12308), .A2(n12307), .ZN(n12316) );
  AOI22_X1 U13762 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U13763 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12311) );
  NAND2_X1 U13764 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12310) );
  NAND2_X1 U13765 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12309) );
  NAND4_X1 U13766 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12314) );
  INV_X1 U13767 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12481) );
  INV_X1 U13768 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13763) );
  OAI22_X1 U13769 ( .A1(n13926), .A2(n12481), .B1(n13924), .B2(n13763), .ZN(
        n12313) );
  NOR2_X1 U13770 ( .A1(n12314), .A2(n12313), .ZN(n12315) );
  AND2_X1 U13771 ( .A1(n12316), .A2(n12315), .ZN(n14808) );
  NAND2_X1 U13772 ( .A1(n12093), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U13773 ( .A1(n16025), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12317) );
  OAI211_X1 U13774 ( .C1(n14808), .C2(n12372), .A(n12318), .B(n12317), .ZN(
        n14708) );
  NAND2_X1 U13775 ( .A1(n12093), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U13776 ( .A1(n16025), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U13777 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U13778 ( .A1(n13929), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U13779 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12319) );
  AND2_X1 U13780 ( .A1(n12320), .A2(n12319), .ZN(n12323) );
  AOI22_X1 U13781 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U13782 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12321) );
  NAND4_X1 U13783 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .ZN(
        n12332) );
  INV_X1 U13784 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12325) );
  INV_X1 U13785 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13792) );
  OAI22_X1 U13786 ( .A1(n13926), .A2(n12325), .B1(n13924), .B2(n13792), .ZN(
        n12326) );
  INV_X1 U13787 ( .A(n12326), .ZN(n12330) );
  AOI22_X1 U13788 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U13789 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12096), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U13790 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12327) );
  NAND4_X1 U13791 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12331) );
  OR2_X1 U13792 ( .A1(n12332), .A2(n12331), .ZN(n14936) );
  INV_X1 U13793 ( .A(n14936), .ZN(n12333) );
  OR2_X1 U13794 ( .A1(n12372), .A2(n12333), .ZN(n12334) );
  AND3_X1 U13795 ( .A1(n12336), .A2(n12335), .A3(n12334), .ZN(n14720) );
  AOI22_X1 U13796 ( .A1(n12093), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n16025), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U13797 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U13798 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12339) );
  NAND2_X1 U13799 ( .A1(n13911), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U13800 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12337) );
  NAND4_X1 U13801 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12346) );
  NAND2_X1 U13802 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12344) );
  NAND2_X1 U13803 ( .A1(n12241), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12343) );
  NAND2_X1 U13804 ( .A1(n13918), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12342) );
  NAND2_X1 U13805 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12341) );
  NAND4_X1 U13806 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12345) );
  NOR2_X1 U13807 ( .A1(n12346), .A2(n12345), .ZN(n12354) );
  AOI22_X1 U13808 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12350) );
  NAND2_X1 U13809 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12349) );
  NAND2_X1 U13810 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12348) );
  NAND2_X1 U13811 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12347) );
  NAND4_X1 U13812 ( .A1(n12350), .A2(n12349), .A3(n12348), .A4(n12347), .ZN(
        n12352) );
  INV_X1 U13813 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13880) );
  INV_X1 U13814 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14569) );
  OAI22_X1 U13815 ( .A1(n13926), .A2(n13880), .B1(n13924), .B2(n14569), .ZN(
        n12351) );
  NOR2_X1 U13816 ( .A1(n12352), .A2(n12351), .ZN(n12353) );
  AND2_X1 U13817 ( .A1(n12354), .A2(n12353), .ZN(n15100) );
  OAI22_X1 U13818 ( .A1(n12372), .A2(n15100), .B1(n12355), .B2(n17099), .ZN(
        n12356) );
  INV_X1 U13819 ( .A(n12356), .ZN(n12357) );
  NAND2_X1 U13820 ( .A1(n12358), .A2(n12357), .ZN(n14874) );
  NAND2_X1 U13821 ( .A1(n12093), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U13822 ( .A1(n16025), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U13823 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U13824 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12360) );
  NAND2_X1 U13825 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12359) );
  AND2_X1 U13826 ( .A1(n12360), .A2(n12359), .ZN(n12363) );
  AOI22_X1 U13827 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U13828 ( .A1(n13906), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U13829 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12371) );
  AOI22_X1 U13830 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U13831 ( .A1(n13928), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13930), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U13832 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U13833 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12366) );
  NAND4_X1 U13834 ( .A1(n12369), .A2(n12368), .A3(n12367), .A4(n12366), .ZN(
        n12370) );
  NOR2_X1 U13835 ( .A1(n12371), .A2(n12370), .ZN(n15099) );
  OR2_X1 U13836 ( .A1(n12372), .A2(n15099), .ZN(n12373) );
  AND3_X1 U13837 ( .A1(n12375), .A2(n12374), .A3(n12373), .ZN(n15063) );
  INV_X1 U13838 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17558) );
  AOI22_X1 U13839 ( .A1(n16025), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U13840 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13911), .B1(
        n13912), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U13841 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13913), .B1(
        n12096), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U13842 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12376) );
  AND2_X1 U13843 ( .A1(n12377), .A2(n12376), .ZN(n12380) );
  AOI22_X1 U13844 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U13845 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12144), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U13846 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12389) );
  INV_X1 U13847 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12382) );
  INV_X1 U13848 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13794) );
  OAI22_X1 U13849 ( .A1(n13926), .A2(n12382), .B1(n13924), .B2(n13794), .ZN(
        n12383) );
  INV_X1 U13850 ( .A(n12383), .ZN(n12387) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12176), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U13852 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13929), .B1(
        n12101), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U13853 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12384) );
  NAND4_X1 U13854 ( .A1(n12387), .A2(n12386), .A3(n12385), .A4(n12384), .ZN(
        n12388) );
  OR2_X1 U13855 ( .A1(n12389), .A2(n12388), .ZN(n15552) );
  NAND2_X1 U13856 ( .A1(n11467), .A2(n15552), .ZN(n12390) );
  OAI211_X1 U13857 ( .C1(n12163), .C2(n17558), .A(n12391), .B(n12390), .ZN(
        n15105) );
  NAND2_X1 U13858 ( .A1(n15061), .A2(n15105), .ZN(n15615) );
  NAND2_X1 U13859 ( .A1(n12093), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U13860 ( .A1(n16025), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12392) );
  AND2_X1 U13861 ( .A1(n12393), .A2(n12392), .ZN(n15614) );
  NAND2_X1 U13862 ( .A1(n12093), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U13863 ( .A1(n16025), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12396) );
  AND2_X1 U13864 ( .A1(n12397), .A2(n12396), .ZN(n15720) );
  INV_X1 U13865 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U13866 ( .A1(n16025), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12399) );
  OAI21_X1 U13867 ( .B1(n12163), .B2(n12400), .A(n12399), .ZN(n17030) );
  AOI22_X1 U13868 ( .A1(n16025), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12401) );
  OAI21_X1 U13869 ( .B1(n12163), .B2(n17560), .A(n12401), .ZN(n16691) );
  NAND2_X1 U13870 ( .A1(n12093), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U13871 ( .A1(n16025), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12402) );
  AND2_X1 U13872 ( .A1(n12403), .A2(n12402), .ZN(n17003) );
  NAND2_X1 U13873 ( .A1(n12093), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U13874 ( .A1(n16025), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12406) );
  AND2_X1 U13875 ( .A1(n12407), .A2(n12406), .ZN(n16682) );
  NAND2_X1 U13876 ( .A1(n12093), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U13877 ( .A1(n16025), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12408) );
  AND2_X1 U13878 ( .A1(n12409), .A2(n12408), .ZN(n16978) );
  INV_X1 U13879 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18882) );
  AOI22_X1 U13880 ( .A1(n16025), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12410) );
  OAI21_X1 U13881 ( .B1(n12163), .B2(n18882), .A(n12410), .ZN(n16671) );
  NAND2_X1 U13882 ( .A1(n12093), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U13883 ( .A1(n16025), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12411) );
  AND2_X1 U13884 ( .A1(n12412), .A2(n12411), .ZN(n16661) );
  NAND2_X1 U13885 ( .A1(n12093), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U13886 ( .A1(n16025), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12413) );
  AND2_X1 U13887 ( .A1(n12414), .A2(n12413), .ZN(n16652) );
  INV_X1 U13888 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18921) );
  AOI22_X1 U13889 ( .A1(n16025), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12415) );
  OAI21_X1 U13890 ( .B1(n12163), .B2(n18921), .A(n12415), .ZN(n16638) );
  INV_X1 U13891 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U13892 ( .A1(n16025), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12416) );
  OAI21_X1 U13893 ( .B1(n12163), .B2(n17566), .A(n12416), .ZN(n16628) );
  NAND2_X1 U13894 ( .A1(n12093), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U13895 ( .A1(n16025), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12417) );
  AND2_X1 U13896 ( .A1(n12418), .A2(n12417), .ZN(n16624) );
  INV_X1 U13897 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U13898 ( .A1(n16025), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11166), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12419) );
  OAI21_X1 U13899 ( .B1(n12163), .B2(n17569), .A(n12419), .ZN(n16608) );
  AOI21_X1 U13900 ( .B1(n12420), .B2(n16610), .A(n16027), .ZN(n15997) );
  NOR2_X1 U13901 ( .A1(n14759), .A2(n11898), .ZN(n14734) );
  NAND2_X1 U13902 ( .A1(n14734), .A2(n18631), .ZN(n18628) );
  AND2_X1 U13903 ( .A1(n12609), .A2(n11854), .ZN(n14327) );
  NAND2_X1 U13904 ( .A1(n14327), .A2(n22141), .ZN(n12423) );
  INV_X1 U13905 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n22173) );
  OR2_X1 U13906 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22173), .ZN(n17577) );
  INV_X2 U13907 ( .A(n17577), .ZN(n22172) );
  INV_X1 U13908 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22181) );
  NAND2_X1 U13909 ( .A1(n22172), .A2(n22181), .ZN(n17572) );
  NOR2_X1 U13910 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17338) );
  NAND2_X1 U13911 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17338), .ZN(n17546) );
  NAND2_X1 U13912 ( .A1(n17568), .A2(n17546), .ZN(n22182) );
  NAND2_X1 U13913 ( .A1(n22174), .A2(n22182), .ZN(n14310) );
  NOR2_X1 U13914 ( .A1(n12423), .A2(n14310), .ZN(n14803) );
  INV_X1 U13915 ( .A(n14803), .ZN(n12424) );
  OR2_X1 U13916 ( .A1(n18628), .A2(n12424), .ZN(n18922) );
  INV_X1 U13917 ( .A(n18922), .ZN(n18977) );
  AOI22_X1 U13918 ( .A1(n15977), .A2(n18957), .B1(n15997), .B2(n18977), .ZN(
        n12454) );
  NAND2_X1 U13919 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19594), .ZN(n19041) );
  NOR3_X1 U13920 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19593), .A3(n19041), 
        .ZN(n19045) );
  INV_X1 U13921 ( .A(n19039), .ZN(n18980) );
  NOR2_X1 U13922 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15936) );
  INV_X1 U13923 ( .A(n15936), .ZN(n19034) );
  NOR2_X1 U13924 ( .A1(n19034), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n17427) );
  INV_X1 U13925 ( .A(n17427), .ZN(n14149) );
  NOR3_X1 U13926 ( .A1(n19045), .A2(n18980), .A3(n11167), .ZN(n12425) );
  AND2_X2 U13927 ( .A1(n18628), .A2(n12425), .ZN(n18954) );
  MUX2_X1 U13928 ( .A(n14096), .B(n12426), .S(n14102), .Z(n12752) );
  INV_X1 U13929 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18662) );
  MUX2_X1 U13930 ( .A(n12752), .B(n18662), .S(n12574), .Z(n12584) );
  INV_X1 U13931 ( .A(n12584), .ZN(n12433) );
  INV_X1 U13932 ( .A(n14109), .ZN(n12427) );
  MUX2_X1 U13933 ( .A(n12507), .B(n12427), .S(n11893), .Z(n12751) );
  INV_X1 U13934 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12428) );
  MUX2_X1 U13935 ( .A(n12751), .B(n12428), .S(n12574), .Z(n12565) );
  INV_X1 U13936 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12429) );
  MUX2_X1 U13937 ( .A(n12429), .B(n12764), .S(n16004), .Z(n12577) );
  INV_X1 U13938 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n12430) );
  NAND2_X1 U13939 ( .A1(n12430), .A2(n11912), .ZN(n12431) );
  MUX2_X1 U13940 ( .A(n12431), .B(n12759), .S(n16004), .Z(n12578) );
  INV_X1 U13941 ( .A(n12578), .ZN(n12432) );
  INV_X1 U13942 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12435) );
  MUX2_X1 U13943 ( .A(n12435), .B(n12434), .S(n16004), .Z(n12561) );
  INV_X1 U13944 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18687) );
  MUX2_X1 U13945 ( .A(n18687), .B(n12608), .S(n16004), .Z(n12615) );
  MUX2_X1 U13946 ( .A(n12436), .B(n11468), .S(n16004), .Z(n12620) );
  NAND2_X1 U13947 ( .A1(n12574), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12630) );
  NAND2_X1 U13948 ( .A1(n12574), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12633) );
  NAND2_X1 U13949 ( .A1(n12574), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12636) );
  NAND2_X1 U13950 ( .A1(n12574), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12644) );
  INV_X1 U13951 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12439) );
  NOR2_X1 U13952 ( .A1(n16004), .A2(n12439), .ZN(n12670) );
  NOR2_X1 U13953 ( .A1(n16004), .A2(n12440), .ZN(n12667) );
  INV_X1 U13954 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12441) );
  NOR2_X1 U13955 ( .A1(n16004), .A2(n12441), .ZN(n12656) );
  NAND2_X1 U13956 ( .A1(n12574), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U13957 ( .A1(n12574), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U13958 ( .A1(n12574), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12647) );
  INV_X1 U13959 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U13960 ( .A1(n12574), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U13961 ( .A1(n12574), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12701) );
  NAND2_X1 U13962 ( .A1(n12574), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U13963 ( .A1(n12574), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U13964 ( .A1(n12574), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12717) );
  INV_X1 U13965 ( .A(n12715), .ZN(n12444) );
  NAND2_X1 U13966 ( .A1(n12574), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U13967 ( .A1(n12574), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12720) );
  INV_X1 U13968 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12445) );
  NOR2_X1 U13969 ( .A1(n16004), .A2(n12445), .ZN(n12725) );
  NAND2_X1 U13970 ( .A1(n12574), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U13971 ( .A1(n12574), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12446) );
  XNOR2_X1 U13972 ( .A(n16003), .B(n12446), .ZN(n15964) );
  NAND2_X1 U13973 ( .A1(n22141), .A2(n22174), .ZN(n12447) );
  NAND2_X1 U13974 ( .A1(n14152), .A2(n12447), .ZN(n12449) );
  INV_X1 U13975 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n18972) );
  OR3_X1 U13976 ( .A1(n12449), .A2(n12609), .A3(n18972), .ZN(n18969) );
  NAND2_X1 U13977 ( .A1(n14152), .A2(n12609), .ZN(n14297) );
  NOR2_X1 U13978 ( .A1(n14310), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12448) );
  OR2_X1 U13979 ( .A1(n14297), .A2(n12448), .ZN(n18971) );
  OR2_X1 U13980 ( .A1(n12449), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U13981 ( .A1(n18971), .A2(n12450), .ZN(n18951) );
  AOI22_X1 U13982 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18954), .ZN(n12451) );
  OAI21_X1 U13983 ( .B1(n15966), .B2(n18969), .A(n12451), .ZN(n12452) );
  AOI21_X1 U13984 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18955), .A(
        n12452), .ZN(n12453) );
  AND2_X1 U13985 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  NAND2_X1 U13986 ( .A1(n12456), .A2(n12455), .ZN(P2_U2825) );
  INV_X1 U13987 ( .A(n12457), .ZN(n12459) );
  INV_X1 U13988 ( .A(n12460), .ZN(n12463) );
  INV_X1 U13989 ( .A(n12461), .ZN(n12462) );
  NAND2_X1 U13990 ( .A1(n12463), .A2(n12462), .ZN(n12464) );
  NAND2_X1 U13991 ( .A1(n13756), .A2(n12484), .ZN(n12490) );
  INV_X1 U13992 ( .A(n12490), .ZN(n12486) );
  INV_X1 U13993 ( .A(n12465), .ZN(n12466) );
  NAND2_X1 U13994 ( .A1(n12467), .A2(n12466), .ZN(n12492) );
  INV_X1 U13995 ( .A(n12468), .ZN(n12475) );
  NAND2_X2 U13996 ( .A1(n12486), .A2(n12469), .ZN(n12550) );
  INV_X1 U13997 ( .A(n12477), .ZN(n12470) );
  NAND2_X2 U13998 ( .A1(n12470), .A2(n12469), .ZN(n12551) );
  INV_X1 U13999 ( .A(n12477), .ZN(n12496) );
  INV_X1 U14000 ( .A(n12473), .ZN(n12474) );
  NAND2_X1 U14001 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  INV_X1 U14002 ( .A(n18648), .ZN(n14295) );
  NAND2_X2 U14003 ( .A1(n12496), .A2(n12498), .ZN(n12535) );
  INV_X1 U14004 ( .A(n12477), .ZN(n12479) );
  NOR2_X1 U14005 ( .A1(n12483), .A2(n12482), .ZN(n12489) );
  OR2_X2 U14006 ( .A1(n13756), .A2(n12484), .ZN(n12502) );
  AOI22_X1 U14007 ( .A1(n19615), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12548), .ZN(n12488) );
  AND2_X2 U14009 ( .A1(n12486), .A2(n12478), .ZN(n12549) );
  AOI22_X1 U14010 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12531), .B1(
        n12549), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12487) );
  INV_X1 U14011 ( .A(n12490), .ZN(n12499) );
  INV_X1 U14012 ( .A(n12491), .ZN(n12493) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12545), .B1(
        n12533), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12506) );
  AND2_X2 U14014 ( .A1(n12496), .A2(n12495), .ZN(n12539) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12546), .B1(
        n12539), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12505) );
  NOR2_X2 U14016 ( .A1(n12502), .A2(n12497), .ZN(n12547) );
  INV_X1 U14017 ( .A(n12501), .ZN(n12498) );
  AOI22_X1 U14018 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12547), .B1(
        n12538), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12504) );
  NOR2_X2 U14019 ( .A1(n12502), .A2(n12500), .ZN(n12532) );
  NOR2_X2 U14020 ( .A1(n12502), .A2(n12501), .ZN(n12544) );
  AOI22_X1 U14021 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12532), .B1(
        n12544), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12503) );
  AOI21_X1 U14022 ( .B1(n12531), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n12609), .ZN(n12510) );
  NAND2_X1 U14023 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12509) );
  AOI22_X1 U14024 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12546), .B1(
        n12547), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U14025 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12545), .B1(
        n12544), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U14026 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12532), .B1(
        n12538), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12511) );
  NAND4_X1 U14027 ( .A1(n11266), .A2(n12513), .A3(n12512), .A4(n12511), .ZN(
        n12529) );
  INV_X1 U14028 ( .A(n12551), .ZN(n19585) );
  INV_X1 U14029 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12515) );
  NOR2_X1 U14030 ( .A1(n12534), .A2(n12515), .ZN(n12516) );
  INV_X1 U14031 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12519) );
  OAI22_X1 U14032 ( .A1(n12519), .A2(n12550), .B1(n12535), .B2(n12518), .ZN(
        n12520) );
  INV_X1 U14033 ( .A(n12520), .ZN(n12521) );
  NAND4_X1 U14034 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12528) );
  NOR2_X1 U14035 ( .A1(n12758), .A2(n12069), .ZN(n14285) );
  INV_X1 U14036 ( .A(n12759), .ZN(n12525) );
  NAND2_X1 U14037 ( .A1(n14285), .A2(n12525), .ZN(n12763) );
  NAND2_X1 U14038 ( .A1(n12763), .A2(n12526), .ZN(n12527) );
  OAI21_X2 U14039 ( .B1(n12529), .B2(n12528), .A(n12527), .ZN(n12563) );
  AOI22_X1 U14040 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12531), .B1(
        n19615), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U14041 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12532), .B1(
        n12533), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12542) );
  OAI22_X1 U14042 ( .A1(n12536), .A2(n12534), .B1(n12535), .B2(n13880), .ZN(
        n12537) );
  INV_X1 U14043 ( .A(n12537), .ZN(n12541) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12544), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U14045 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12546), .B1(
        n12547), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U14046 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19678), .B1(
        n12549), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12555) );
  OAI22_X1 U14047 ( .A1(n12552), .A2(n12550), .B1(n12551), .B2(n13884), .ZN(
        n12553) );
  INV_X1 U14048 ( .A(n12553), .ZN(n12554) );
  NAND2_X1 U14049 ( .A1(n11281), .A2(n11577), .ZN(n12562) );
  NAND2_X1 U14050 ( .A1(n12616), .A2(n12562), .ZN(n18677) );
  XNOR2_X1 U14051 ( .A(n12593), .B(n15642), .ZN(n15639) );
  XNOR2_X1 U14052 ( .A(n12564), .B(n12563), .ZN(n12767) );
  NAND2_X1 U14053 ( .A1(n12767), .A2(n16849), .ZN(n12569) );
  INV_X1 U14054 ( .A(n12565), .ZN(n12567) );
  INV_X1 U14055 ( .A(n12566), .ZN(n12581) );
  NAND2_X1 U14056 ( .A1(n12567), .A2(n12581), .ZN(n12568) );
  NAND2_X1 U14057 ( .A1(n12583), .A2(n12568), .ZN(n15947) );
  NAND2_X1 U14058 ( .A1(n12569), .A2(n15947), .ZN(n15065) );
  INV_X1 U14059 ( .A(n12758), .ZN(n12572) );
  NAND2_X1 U14060 ( .A1(n11741), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12570) );
  NAND2_X1 U14061 ( .A1(n12571), .A2(n12570), .ZN(n12741) );
  INV_X1 U14062 ( .A(n12741), .ZN(n14105) );
  MUX2_X1 U14063 ( .A(n12572), .B(n14105), .S(n11893), .Z(n12573) );
  MUX2_X1 U14064 ( .A(n12573), .B(P2_EBX_REG_0__SCAN_IN), .S(n12574), .Z(
        n14284) );
  INV_X1 U14065 ( .A(n14284), .ZN(n18634) );
  INV_X1 U14066 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18993) );
  NOR2_X1 U14067 ( .A1(n18634), .A2(n18993), .ZN(n12576) );
  NAND3_X1 U14068 ( .A1(n12574), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12575) );
  AND2_X1 U14069 ( .A1(n12578), .A2(n12575), .ZN(n18647) );
  NOR2_X1 U14070 ( .A1(n12576), .A2(n18647), .ZN(n14244) );
  AND2_X1 U14071 ( .A1(n12576), .A2(n18647), .ZN(n14243) );
  NOR2_X1 U14072 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14243), .ZN(
        n14242) );
  NOR2_X1 U14073 ( .A1(n14244), .A2(n14242), .ZN(n14341) );
  INV_X1 U14074 ( .A(n12577), .ZN(n12579) );
  NAND2_X1 U14075 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  NAND2_X1 U14076 ( .A1(n12581), .A2(n12580), .ZN(n15542) );
  XNOR2_X1 U14077 ( .A(n15542), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14340) );
  INV_X1 U14078 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14379) );
  NOR2_X1 U14079 ( .A1(n15542), .A2(n14379), .ZN(n12582) );
  AOI21_X1 U14080 ( .B1(n14341), .B2(n14340), .A(n12582), .ZN(n15086) );
  OR2_X1 U14081 ( .A1(n12584), .A2(n11578), .ZN(n12585) );
  NAND2_X1 U14082 ( .A1(n11281), .A2(n12585), .ZN(n18658) );
  INV_X1 U14083 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15643) );
  AND2_X1 U14084 ( .A1(n18658), .A2(n15643), .ZN(n12587) );
  AOI21_X1 U14085 ( .B1(n15086), .B2(n19030), .A(n12587), .ZN(n12586) );
  NAND2_X1 U14086 ( .A1(n15065), .A2(n12586), .ZN(n12592) );
  INV_X1 U14087 ( .A(n15086), .ZN(n15066) );
  INV_X1 U14088 ( .A(n12587), .ZN(n12588) );
  AND2_X1 U14089 ( .A1(n12588), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12590) );
  INV_X1 U14090 ( .A(n18658), .ZN(n12589) );
  AOI22_X1 U14091 ( .A1(n15066), .A2(n12590), .B1(n12589), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U14092 ( .A1(n12592), .A2(n12591), .ZN(n15640) );
  NAND2_X1 U14093 ( .A1(n12593), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12594) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12532), .B1(
        n12544), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U14095 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12545), .B1(
        n12533), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U14096 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12547), .B1(
        n12538), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U14097 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12546), .B1(
        n12539), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U14098 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12607) );
  AOI22_X1 U14099 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19615), .B1(
        n19678), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U14100 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12531), .B1(
        n12549), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12604) );
  OAI22_X1 U14101 ( .A1(n12599), .A2(n12550), .B1(n12551), .B2(n13899), .ZN(
        n12600) );
  INV_X1 U14102 ( .A(n12600), .ZN(n12603) );
  INV_X1 U14103 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13902) );
  OAI22_X1 U14104 ( .A1(n15670), .A2(n12534), .B1(n12535), .B2(n13902), .ZN(
        n12601) );
  INV_X1 U14105 ( .A(n12601), .ZN(n12602) );
  NAND4_X1 U14106 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        n12606) );
  INV_X1 U14107 ( .A(n12608), .ZN(n12610) );
  NAND2_X1 U14108 ( .A1(n12610), .A2(n12609), .ZN(n12611) );
  NAND2_X1 U14109 ( .A1(n12616), .A2(n11579), .ZN(n12617) );
  INV_X1 U14110 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15787) );
  NAND2_X1 U14111 ( .A1(n12618), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12619) );
  XNOR2_X1 U14112 ( .A(n12621), .B(n12620), .ZN(n18702) );
  AND2_X1 U14113 ( .A1(n18702), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15778) );
  INV_X1 U14114 ( .A(n18702), .ZN(n12622) );
  NAND2_X1 U14115 ( .A1(n12622), .A2(n15788), .ZN(n15779) );
  INV_X1 U14116 ( .A(n12623), .ZN(n16005) );
  INV_X1 U14117 ( .A(n12624), .ZN(n12625) );
  NAND2_X1 U14118 ( .A1(n16005), .A2(n12625), .ZN(n12626) );
  AND2_X1 U14119 ( .A1(n12631), .A2(n12626), .ZN(n18710) );
  NAND2_X1 U14120 ( .A1(n18710), .A2(n11468), .ZN(n12629) );
  INV_X1 U14121 ( .A(n12629), .ZN(n12627) );
  NAND2_X1 U14122 ( .A1(n12627), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17437) );
  AND2_X1 U14123 ( .A1(n12629), .A2(n12628), .ZN(n17438) );
  XNOR2_X1 U14124 ( .A(n12631), .B(n12630), .ZN(n18724) );
  NAND2_X1 U14125 ( .A1(n18724), .A2(n11468), .ZN(n12632) );
  NAND2_X1 U14126 ( .A1(n12632), .A2(n16884), .ZN(n17150) );
  XNOR2_X1 U14127 ( .A(n12634), .B(n12633), .ZN(n18733) );
  NAND2_X1 U14128 ( .A1(n18733), .A2(n11468), .ZN(n12642) );
  INV_X1 U14129 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17140) );
  INV_X1 U14130 ( .A(n12635), .ZN(n12638) );
  INV_X1 U14131 ( .A(n12636), .ZN(n12637) );
  NAND2_X1 U14132 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  NAND2_X1 U14133 ( .A1(n12645), .A2(n12639), .ZN(n18748) );
  NOR2_X1 U14134 ( .A1(n18748), .A2(n16849), .ZN(n12641) );
  INV_X1 U14135 ( .A(n12641), .ZN(n12640) );
  INV_X1 U14136 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17123) );
  NAND2_X1 U14137 ( .A1(n12641), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16879) );
  OR2_X1 U14138 ( .A1(n12642), .A2(n17140), .ZN(n17135) );
  AND2_X1 U14139 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12643) );
  NAND2_X1 U14140 ( .A1(n18724), .A2(n12643), .ZN(n17149) );
  AND2_X1 U14141 ( .A1(n17135), .A2(n17149), .ZN(n16878) );
  XNOR2_X1 U14142 ( .A(n12645), .B(n12644), .ZN(n18761) );
  NAND2_X1 U14143 ( .A1(n18761), .A2(n11468), .ZN(n17109) );
  INV_X1 U14144 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17464) );
  NOR2_X1 U14145 ( .A1(n17109), .A2(n17464), .ZN(n12685) );
  INV_X1 U14146 ( .A(n12646), .ZN(n12654) );
  INV_X1 U14147 ( .A(n12647), .ZN(n12648) );
  NAND2_X1 U14148 ( .A1(n12654), .A2(n12648), .ZN(n12649) );
  NAND2_X1 U14149 ( .A1(n12696), .A2(n12649), .ZN(n18845) );
  INV_X1 U14150 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17024) );
  NAND2_X1 U14151 ( .A1(n12691), .A2(n17024), .ZN(n16806) );
  INV_X1 U14152 ( .A(n12650), .ZN(n12665) );
  INV_X1 U14153 ( .A(n12651), .ZN(n12652) );
  NAND2_X1 U14154 ( .A1(n12665), .A2(n12652), .ZN(n12653) );
  NAND2_X1 U14155 ( .A1(n12654), .A2(n12653), .ZN(n12687) );
  INV_X1 U14156 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17018) );
  OAI21_X1 U14157 ( .B1(n12687), .B2(n16849), .A(n17018), .ZN(n16821) );
  NAND2_X1 U14158 ( .A1(n16806), .A2(n16821), .ZN(n16779) );
  INV_X1 U14159 ( .A(n12655), .ZN(n12663) );
  NAND2_X1 U14160 ( .A1(n12669), .A2(n12656), .ZN(n12657) );
  NAND2_X1 U14161 ( .A1(n12663), .A2(n12657), .ZN(n18806) );
  OAI21_X1 U14162 ( .B1(n18806), .B2(n16849), .A(n12658), .ZN(n12660) );
  NAND2_X1 U14163 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12659) );
  INV_X1 U14164 ( .A(n12661), .ZN(n12662) );
  NAND2_X1 U14165 ( .A1(n12663), .A2(n12662), .ZN(n12664) );
  NAND2_X1 U14166 ( .A1(n12665), .A2(n12664), .ZN(n18823) );
  OR2_X1 U14167 ( .A1(n18823), .A2(n16849), .ZN(n12666) );
  INV_X1 U14168 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17055) );
  NAND2_X1 U14169 ( .A1(n12666), .A2(n17055), .ZN(n16829) );
  NAND2_X1 U14170 ( .A1(n12672), .A2(n12667), .ZN(n12668) );
  AND2_X1 U14171 ( .A1(n12669), .A2(n12668), .ZN(n18792) );
  AOI21_X1 U14172 ( .B1(n18792), .B2(n11468), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16845) );
  INV_X1 U14173 ( .A(n17109), .ZN(n16771) );
  NAND2_X1 U14174 ( .A1(n12675), .A2(n12670), .ZN(n12671) );
  NAND2_X1 U14175 ( .A1(n12672), .A2(n12671), .ZN(n18785) );
  OR2_X1 U14176 ( .A1(n18785), .A2(n16849), .ZN(n12673) );
  INV_X1 U14177 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17084) );
  NAND2_X1 U14178 ( .A1(n12673), .A2(n17084), .ZN(n16852) );
  NAND2_X1 U14179 ( .A1(n11268), .A2(n11308), .ZN(n12674) );
  NAND2_X1 U14180 ( .A1(n12675), .A2(n12674), .ZN(n18770) );
  OR2_X1 U14181 ( .A1(n18770), .A2(n16849), .ZN(n12676) );
  NAND2_X1 U14182 ( .A1(n12676), .A2(n17099), .ZN(n16868) );
  OAI211_X1 U14183 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16771), .A(
        n16852), .B(n16868), .ZN(n12677) );
  NOR2_X1 U14184 ( .A1(n16845), .A2(n12677), .ZN(n12678) );
  NAND3_X1 U14185 ( .A1(n16836), .A2(n16829), .A3(n12678), .ZN(n12679) );
  NOR2_X1 U14186 ( .A1(n16779), .A2(n12679), .ZN(n12683) );
  XNOR2_X1 U14187 ( .A(n12681), .B(n12680), .ZN(n18863) );
  NAND2_X1 U14188 ( .A1(n18863), .A2(n11468), .ZN(n12682) );
  INV_X1 U14189 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U14190 ( .A1(n12682), .A2(n12792), .ZN(n16786) );
  INV_X1 U14191 ( .A(n12695), .ZN(n12694) );
  AND2_X1 U14192 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12686) );
  NAND2_X1 U14193 ( .A1(n18863), .A2(n12686), .ZN(n16785) );
  INV_X1 U14194 ( .A(n12687), .ZN(n18834) );
  AND2_X1 U14195 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U14196 ( .A1(n18834), .A2(n12688), .ZN(n16820) );
  NAND2_X1 U14197 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12689) );
  NAND2_X1 U14198 ( .A1(n18792), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16846) );
  OR2_X1 U14199 ( .A1(n18770), .A2(n17099), .ZN(n16848) );
  OR2_X1 U14200 ( .A1(n18785), .A2(n17084), .ZN(n16850) );
  NAND3_X1 U14201 ( .A1(n16846), .A2(n16848), .A3(n16850), .ZN(n12690) );
  NAND2_X1 U14202 ( .A1(n12690), .A2(n11468), .ZN(n16775) );
  AND4_X1 U14203 ( .A1(n16820), .A2(n16776), .A3(n16828), .A4(n16775), .ZN(
        n12693) );
  INV_X1 U14204 ( .A(n12691), .ZN(n12692) );
  NAND2_X1 U14205 ( .A1(n12692), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16807) );
  XNOR2_X1 U14206 ( .A(n12696), .B(n11320), .ZN(n18854) );
  NAND2_X1 U14207 ( .A1(n18854), .A2(n11468), .ZN(n16780) );
  INV_X1 U14208 ( .A(n16780), .ZN(n12697) );
  NAND2_X1 U14209 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  XNOR2_X1 U14210 ( .A(n12702), .B(n12701), .ZN(n18873) );
  INV_X1 U14211 ( .A(n12703), .ZN(n12706) );
  INV_X1 U14212 ( .A(n12704), .ZN(n12705) );
  NAND2_X1 U14213 ( .A1(n12706), .A2(n12705), .ZN(n12707) );
  NAND2_X1 U14214 ( .A1(n12711), .A2(n12707), .ZN(n18886) );
  OR2_X1 U14215 ( .A1(n18886), .A2(n16849), .ZN(n12708) );
  NAND2_X1 U14216 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12709) );
  NAND2_X1 U14217 ( .A1(n16745), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12712) );
  XNOR2_X1 U14218 ( .A(n12711), .B(n12710), .ZN(n18896) );
  INV_X1 U14219 ( .A(n16745), .ZN(n12713) );
  XNOR2_X1 U14220 ( .A(n12715), .B(n12714), .ZN(n18919) );
  NAND2_X1 U14221 ( .A1(n18919), .A2(n11468), .ZN(n12716) );
  XNOR2_X1 U14222 ( .A(n12716), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16726) );
  XNOR2_X1 U14223 ( .A(n11256), .B(n12717), .ZN(n18909) );
  NAND2_X1 U14224 ( .A1(n18909), .A2(n11468), .ZN(n12718) );
  INV_X1 U14225 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16929) );
  NAND2_X1 U14226 ( .A1(n12718), .A2(n16929), .ZN(n16727) );
  INV_X1 U14227 ( .A(n12719), .ZN(n12722) );
  INV_X1 U14228 ( .A(n12720), .ZN(n12721) );
  NAND2_X1 U14229 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  NAND2_X1 U14230 ( .A1(n12726), .A2(n12723), .ZN(n18933) );
  NAND2_X1 U14231 ( .A1(n11279), .A2(n16893), .ZN(n12724) );
  NAND2_X1 U14232 ( .A1(n12726), .A2(n12725), .ZN(n12727) );
  NAND2_X1 U14233 ( .A1(n12728), .A2(n12727), .ZN(n18944) );
  INV_X1 U14234 ( .A(n16704), .ZN(n12731) );
  INV_X1 U14235 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16907) );
  NAND2_X1 U14236 ( .A1(n11191), .A2(n12732), .ZN(n12735) );
  NAND3_X1 U14237 ( .A1(n18919), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11468), .ZN(n12734) );
  AND2_X1 U14238 ( .A1(n11468), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12733) );
  NAND2_X1 U14239 ( .A1(n18909), .A2(n12733), .ZN(n16725) );
  XOR2_X1 U14240 ( .A(n12737), .B(n12736), .Z(n18953) );
  NAND2_X1 U14241 ( .A1(n18953), .A2(n11468), .ZN(n12739) );
  INV_X1 U14242 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12738) );
  NAND2_X1 U14243 ( .A1(n12739), .A2(n12738), .ZN(n15962) );
  INV_X1 U14244 ( .A(n12739), .ZN(n12740) );
  NAND2_X1 U14245 ( .A1(n12740), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15999) );
  NOR3_X1 U14246 ( .A1(n14109), .A2(n14108), .A3(n12741), .ZN(n12742) );
  NAND2_X1 U14247 ( .A1(n14096), .A2(n12742), .ZN(n12743) );
  NAND2_X1 U14248 ( .A1(n12743), .A2(n14913), .ZN(n12744) );
  OR2_X1 U14249 ( .A1(n14759), .A2(n12744), .ZN(n12749) );
  CLKBUF_X1 U14250 ( .A(n12745), .Z(n14745) );
  NAND2_X1 U14251 ( .A1(n14745), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12746) );
  NAND2_X1 U14252 ( .A1(n12746), .A2(n18987), .ZN(n14775) );
  INV_X1 U14253 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12747) );
  OAI21_X1 U14254 ( .B1(n13928), .B2(n14775), .A(n12747), .ZN(n12748) );
  NAND2_X1 U14255 ( .A1(n12748), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17476) );
  AND2_X1 U14256 ( .A1(n14314), .A2(n14102), .ZN(n14765) );
  INV_X1 U14257 ( .A(n14765), .ZN(n12757) );
  NAND2_X1 U14258 ( .A1(n12752), .A2(n12751), .ZN(n14113) );
  INV_X1 U14259 ( .A(n14108), .ZN(n14099) );
  NAND2_X1 U14260 ( .A1(n11893), .A2(n14099), .ZN(n14098) );
  NAND2_X1 U14261 ( .A1(n14105), .A2(n12753), .ZN(n14101) );
  AND2_X1 U14262 ( .A1(n14098), .A2(n14101), .ZN(n12754) );
  NOR2_X1 U14263 ( .A1(n14113), .A2(n12754), .ZN(n12755) );
  OR2_X1 U14264 ( .A1(n12755), .A2(n14118), .ZN(n14761) );
  INV_X1 U14265 ( .A(n14761), .ZN(n12756) );
  AND2_X1 U14266 ( .A1(n14314), .A2(n14327), .ZN(n14760) );
  NAND2_X1 U14267 ( .A1(n12756), .A2(n14760), .ZN(n14332) );
  OAI21_X1 U14268 ( .B1(n19043), .B2(n12757), .A(n14332), .ZN(n14777) );
  NAND2_X1 U14269 ( .A1(n14777), .A2(n18631), .ZN(n19057) );
  OR2_X1 U14270 ( .A1(n19057), .A2(n12609), .ZN(n17445) );
  XOR2_X1 U14271 ( .A(n12759), .B(n12758), .Z(n12761) );
  OR2_X1 U14272 ( .A1(n14285), .A2(n18993), .ZN(n14287) );
  INV_X1 U14273 ( .A(n14287), .ZN(n12760) );
  NAND2_X1 U14274 ( .A1(n12761), .A2(n12760), .ZN(n12762) );
  XOR2_X1 U14275 ( .A(n12761), .B(n12760), .Z(n14246) );
  NAND2_X1 U14276 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14246), .ZN(
        n14245) );
  NAND2_X1 U14277 ( .A1(n12762), .A2(n14245), .ZN(n12765) );
  XOR2_X1 U14278 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12765), .Z(
        n14371) );
  XOR2_X1 U14279 ( .A(n12764), .B(n12763), .Z(n14370) );
  NAND2_X1 U14280 ( .A1(n14371), .A2(n14370), .ZN(n14369) );
  NAND2_X1 U14281 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12765), .ZN(
        n12766) );
  NAND2_X1 U14282 ( .A1(n14369), .A2(n12766), .ZN(n12768) );
  XNOR2_X1 U14283 ( .A(n12768), .B(n19030), .ZN(n15085) );
  NAND2_X1 U14284 ( .A1(n12768), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12769) );
  INV_X1 U14285 ( .A(n12776), .ZN(n12772) );
  AND2_X1 U14286 ( .A1(n12776), .A2(n15642), .ZN(n12774) );
  NAND3_X1 U14287 ( .A1(n12772), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n12777), .ZN(n12778) );
  INV_X1 U14288 ( .A(n12785), .ZN(n12786) );
  AND2_X1 U14289 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17124) );
  NAND2_X1 U14290 ( .A1(n17124), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16798) );
  NAND3_X1 U14291 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12790) );
  NOR2_X1 U14292 ( .A1(n16798), .A2(n12790), .ZN(n17005) );
  NAND3_X1 U14293 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17004) );
  NAND3_X1 U14294 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16960) );
  NOR2_X1 U14295 ( .A1(n17004), .A2(n16960), .ZN(n12791) );
  NAND2_X1 U14296 ( .A1(n17005), .A2(n12791), .ZN(n15975) );
  INV_X1 U14297 ( .A(n15975), .ZN(n16961) );
  INV_X1 U14298 ( .A(n16768), .ZN(n12793) );
  INV_X1 U14299 ( .A(n16719), .ZN(n12794) );
  AOI21_X1 U14300 ( .B1(n12794), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12795) );
  NAND2_X1 U14301 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15974) );
  NOR2_X1 U14302 ( .A1(n12795), .A2(n16019), .ZN(n16899) );
  OR2_X1 U14303 ( .A1(n19057), .A2(n12069), .ZN(n17446) );
  INV_X1 U14304 ( .A(n17446), .ZN(n17467) );
  NAND2_X1 U14305 ( .A1(n16899), .A2(n17467), .ZN(n12804) );
  AND2_X1 U14306 ( .A1(n16544), .A2(n12796), .ZN(n12797) );
  NAND2_X1 U14307 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n14914) );
  NAND2_X1 U14308 ( .A1(n19593), .A2(n14914), .ZN(n18630) );
  OR2_X1 U14309 ( .A1(n18630), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12798) );
  AND2_X1 U14310 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17340) );
  NAND2_X1 U14311 ( .A1(n11739), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U14312 ( .A1(n22141), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U14313 ( .A1(n14805), .A2(n12799), .ZN(n14290) );
  NAND2_X1 U14314 ( .A1(n17443), .A2(n18960), .ZN(n12800) );
  NAND2_X1 U14315 ( .A1(n11167), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16890) );
  OAI211_X1 U14316 ( .C1(n17452), .C2(n12801), .A(n12800), .B(n16890), .ZN(
        n12802) );
  AOI21_X1 U14317 ( .B1(n18958), .B2(n17457), .A(n12802), .ZN(n12803) );
  AND2_X2 U14318 ( .A1(n17369), .A2(n12810), .ZN(n13544) );
  AOI22_X1 U14319 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U14320 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13390), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U14321 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12950), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12806) );
  AND2_X2 U14322 ( .A1(n12811), .A2(n14597), .ZN(n12895) );
  BUF_X4 U14323 ( .A(n12895), .Z(n13719) );
  AOI22_X1 U14324 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14325 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12815) );
  AND2_X2 U14326 ( .A1(n12811), .A2(n12809), .ZN(n13088) );
  AOI22_X1 U14327 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12814) );
  AND2_X2 U14328 ( .A1(n14598), .A2(n14597), .ZN(n13422) );
  AOI22_X1 U14329 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12813) );
  AND2_X2 U14330 ( .A1(n14597), .A2(n17368), .ZN(n13358) );
  AOI22_X1 U14331 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U14332 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12950), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U14333 ( .A1(n12896), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U14334 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U14335 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12825) );
  AOI22_X1 U14336 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U14337 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13544), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U14338 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U14339 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13390), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U14340 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12824) );
  AOI22_X1 U14341 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U14342 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U14343 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U14344 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12826) );
  NAND4_X1 U14345 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        n12835) );
  AOI22_X1 U14346 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13390), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U14347 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12950), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U14348 ( .A1(n12896), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12831) );
  AOI22_X1 U14349 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12830) );
  NAND4_X1 U14350 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n12834) );
  NAND2_X1 U14351 ( .A1(n14588), .A2(n14636), .ZN(n13244) );
  AOI22_X1 U14352 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U14353 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13390), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U14354 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12950), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12837) );
  BUF_X2 U14355 ( .A(n12895), .Z(n13692) );
  AOI22_X1 U14356 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12836) );
  NAND4_X1 U14357 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        n12845) );
  AOI22_X1 U14358 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U14359 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U14360 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U14361 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12840) );
  NAND4_X1 U14362 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12844) );
  NAND2_X1 U14363 ( .A1(n12869), .A2(n14637), .ZN(n12932) );
  INV_X1 U14364 ( .A(n14637), .ZN(n14455) );
  NAND2_X2 U14365 ( .A1(n14455), .A2(n12846), .ZN(n16505) );
  NAND2_X1 U14366 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U14367 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12850) );
  NAND2_X1 U14368 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12849) );
  NAND2_X1 U14369 ( .A1(n12874), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12848) );
  NAND2_X1 U14370 ( .A1(n13544), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12856) );
  NAND2_X1 U14371 ( .A1(n12852), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12855) );
  NAND2_X1 U14372 ( .A1(n12896), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12854) );
  NAND2_X1 U14373 ( .A1(n13390), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12853) );
  NAND2_X1 U14374 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U14375 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12859) );
  NAND2_X1 U14376 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12858) );
  NAND2_X1 U14377 ( .A1(n13363), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12857) );
  NAND2_X1 U14378 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12864) );
  NAND2_X1 U14379 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12863) );
  NAND2_X1 U14380 ( .A1(n13422), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12862) );
  NAND2_X1 U14381 ( .A1(n13358), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12861) );
  INV_X4 U14382 ( .A(n14268), .ZN(n14467) );
  NAND3_X1 U14383 ( .A1(n12932), .A2(n16505), .A3(n14467), .ZN(n12924) );
  INV_X1 U14384 ( .A(n12869), .ZN(n12890) );
  NAND2_X1 U14385 ( .A1(n13544), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12873) );
  NAND2_X1 U14386 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12872) );
  NAND2_X1 U14387 ( .A1(n12896), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U14388 ( .A1(n13390), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U14389 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12878) );
  NAND2_X1 U14390 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U14391 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12876) );
  NAND2_X1 U14392 ( .A1(n12874), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12875) );
  NAND2_X1 U14393 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12882) );
  NAND2_X1 U14394 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12881) );
  NAND2_X1 U14395 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12880) );
  NAND2_X1 U14396 ( .A1(n11160), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U14397 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12886) );
  NAND2_X1 U14398 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12885) );
  NAND2_X1 U14399 ( .A1(n13422), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12884) );
  NAND2_X1 U14400 ( .A1(n13358), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12883) );
  AND2_X2 U14401 ( .A1(n22386), .A2(n15821), .ZN(n17412) );
  NAND2_X1 U14402 ( .A1(n12890), .A2(n17412), .ZN(n12933) );
  AOI22_X1 U14403 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U14404 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U14405 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U14406 ( .A1(n13390), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12891) );
  NAND4_X1 U14407 ( .A1(n12894), .A2(n12893), .A3(n12892), .A4(n12891), .ZN(
        n12902) );
  AOI22_X1 U14408 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13544), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U14409 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U14410 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U14411 ( .A1(n12950), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12897) );
  NAND4_X1 U14412 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12901) );
  AOI22_X1 U14413 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U14414 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12874), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U14415 ( .A1(n12945), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U14416 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12904) );
  NAND4_X1 U14417 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12913) );
  AOI22_X1 U14418 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U14419 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13390), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U14420 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12950), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U14421 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12908) );
  NAND4_X1 U14422 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12912) );
  AND2_X1 U14423 ( .A1(n15821), .A2(n14459), .ZN(n12935) );
  AOI21_X1 U14424 ( .B1(n17364), .B2(n13247), .A(n12935), .ZN(n15900) );
  NOR2_X1 U14425 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n22116) );
  INV_X1 U14426 ( .A(n22116), .ZN(n16529) );
  NOR2_X1 U14427 ( .A1(n16529), .A2(n22122), .ZN(n12914) );
  NAND2_X1 U14428 ( .A1(n22236), .A2(n14467), .ZN(n14886) );
  AND4_X1 U14429 ( .A1(n12933), .A2(n15900), .A3(n12914), .A4(n14886), .ZN(
        n12923) );
  NAND2_X1 U14430 ( .A1(n14637), .A2(n12977), .ZN(n12915) );
  NOR2_X2 U14431 ( .A1(n15821), .A2(n14467), .ZN(n14307) );
  INV_X2 U14432 ( .A(n14307), .ZN(n14881) );
  AOI21_X1 U14433 ( .B1(n12915), .B2(n14881), .A(n16057), .ZN(n12916) );
  INV_X1 U14434 ( .A(n14270), .ZN(n12918) );
  NAND2_X1 U14435 ( .A1(n15825), .A2(n14477), .ZN(n12917) );
  NAND4_X1 U14436 ( .A1(n12918), .A2(n22457), .A3(n12917), .A4(n14636), .ZN(
        n14256) );
  NAND2_X1 U14437 ( .A1(n14256), .A2(n16505), .ZN(n12921) );
  NAND2_X1 U14438 ( .A1(n12919), .A2(n14459), .ZN(n12920) );
  NAND2_X1 U14439 ( .A1(n12921), .A2(n12920), .ZN(n12931) );
  NAND2_X1 U14440 ( .A1(n12931), .A2(n14307), .ZN(n14473) );
  NAND4_X1 U14441 ( .A1(n12924), .A2(n12923), .A3(n12922), .A4(n14473), .ZN(
        n12944) );
  AND2_X2 U14442 ( .A1(n12925), .A2(n15821), .ZN(n15895) );
  INV_X1 U14443 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20212) );
  NAND2_X1 U14444 ( .A1(n20212), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22164) );
  INV_X1 U14445 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U14446 ( .A1(n12926), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n12927) );
  AND2_X1 U14447 ( .A1(n22164), .A2(n12927), .ZN(n14265) );
  NAND2_X1 U14448 ( .A1(n22386), .A2(n14265), .ZN(n12930) );
  NAND2_X1 U14449 ( .A1(n14471), .A2(n14307), .ZN(n12928) );
  NAND2_X1 U14450 ( .A1(n14636), .A2(n15524), .ZN(n15820) );
  INV_X1 U14451 ( .A(n15820), .ZN(n13248) );
  NAND4_X1 U14452 ( .A1(n17364), .A2(n14307), .A3(n22528), .A4(n13248), .ZN(
        n15893) );
  NAND2_X1 U14453 ( .A1(n14476), .A2(n15893), .ZN(n12929) );
  OAI21_X1 U14454 ( .B1(n12931), .B2(n17364), .A(n22236), .ZN(n12940) );
  NAND2_X1 U14455 ( .A1(n12932), .A2(n16505), .ZN(n12934) );
  AOI21_X1 U14456 ( .B1(n14471), .B2(n16057), .A(n12935), .ZN(n12938) );
  INV_X1 U14457 ( .A(n14271), .ZN(n14587) );
  NAND2_X1 U14458 ( .A1(n15897), .A2(n14587), .ZN(n12937) );
  NAND2_X1 U14459 ( .A1(n22116), .A2(n22122), .ZN(n13752) );
  INV_X1 U14460 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n22121) );
  AND2_X1 U14461 ( .A1(n22121), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13242) );
  MUX2_X1 U14462 ( .A(n13752), .B(n13242), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n12942) );
  OAI21_X2 U14463 ( .B1(n13018), .B2(n14483), .A(n12942), .ZN(n12943) );
  OAI21_X2 U14464 ( .B1(n12944), .B2(n12943), .A(n12988), .ZN(n14894) );
  AOI22_X1 U14465 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U14466 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U14467 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U14468 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12946) );
  NAND4_X1 U14469 ( .A1(n12949), .A2(n12948), .A3(n12947), .A4(n12946), .ZN(
        n12956) );
  AOI22_X1 U14470 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U14471 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U14472 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U14473 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12951) );
  NAND4_X1 U14474 ( .A1(n12954), .A2(n12953), .A3(n12952), .A4(n12951), .ZN(
        n12955) );
  INV_X1 U14475 ( .A(n13165), .ZN(n12967) );
  AOI22_X1 U14476 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U14477 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U14478 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U14479 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12957) );
  NAND4_X1 U14480 ( .A1(n12960), .A2(n12959), .A3(n12958), .A4(n12957), .ZN(
        n12966) );
  AOI22_X1 U14481 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U14482 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U14483 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U14484 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12961) );
  NAND4_X1 U14485 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12965) );
  OR2_X1 U14486 ( .A1(n12966), .A2(n12965), .ZN(n13050) );
  XNOR2_X1 U14487 ( .A(n12967), .B(n13050), .ZN(n12968) );
  INV_X1 U14488 ( .A(n13038), .ZN(n13160) );
  NAND2_X1 U14489 ( .A1(n12968), .A2(n13160), .ZN(n12974) );
  INV_X1 U14490 ( .A(n12969), .ZN(n13043) );
  INV_X1 U14491 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12972) );
  AOI21_X1 U14492 ( .B1(n15837), .B2(n13165), .A(n22122), .ZN(n12971) );
  NAND2_X1 U14493 ( .A1(n22236), .A2(n13050), .ZN(n12970) );
  OAI211_X1 U14494 ( .C1(n13232), .C2(n12972), .A(n12971), .B(n12970), .ZN(
        n12973) );
  NAND2_X1 U14495 ( .A1(n13043), .A2(n12973), .ZN(n12976) );
  OR2_X1 U14496 ( .A1(n12974), .A2(n12973), .ZN(n12975) );
  NAND2_X1 U14497 ( .A1(n14843), .A2(n13190), .ZN(n12980) );
  INV_X1 U14498 ( .A(n13050), .ZN(n12978) );
  AND2_X1 U14499 ( .A1(n22236), .A2(n12977), .ZN(n13053) );
  AOI21_X1 U14500 ( .B1(n12978), .B2(n17412), .A(n13053), .ZN(n12979) );
  NAND2_X1 U14501 ( .A1(n12980), .A2(n12979), .ZN(n14488) );
  NAND2_X1 U14502 ( .A1(n14488), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14489) );
  NAND2_X1 U14503 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13016) );
  OAI21_X1 U14504 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n13016), .ZN(n22323) );
  INV_X1 U14505 ( .A(n13242), .ZN(n17417) );
  NAND2_X1 U14506 ( .A1(n17417), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13010) );
  OAI21_X1 U14507 ( .B1(n13752), .B2(n22323), .A(n13010), .ZN(n12982) );
  INV_X1 U14508 ( .A(n12982), .ZN(n12983) );
  INV_X1 U14509 ( .A(n12984), .ZN(n12985) );
  INV_X1 U14510 ( .A(n14847), .ZN(n12987) );
  INV_X1 U14511 ( .A(n12988), .ZN(n12989) );
  AOI22_X1 U14512 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U14513 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U14514 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U14515 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12990) );
  NAND4_X1 U14516 ( .A1(n12993), .A2(n12992), .A3(n12991), .A4(n12990), .ZN(
        n12999) );
  AOI22_X1 U14517 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U14518 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14519 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U14520 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12994) );
  NAND4_X1 U14521 ( .A1(n12997), .A2(n12996), .A3(n12995), .A4(n12994), .ZN(
        n12998) );
  OR2_X1 U14522 ( .A1(n12999), .A2(n12998), .ZN(n13049) );
  NAND2_X1 U14523 ( .A1(n13160), .A2(n13049), .ZN(n13000) );
  INV_X1 U14524 ( .A(n13049), .ZN(n13001) );
  XNOR2_X1 U14525 ( .A(n13001), .B(n13050), .ZN(n13002) );
  NAND2_X1 U14526 ( .A1(n13002), .A2(n17412), .ZN(n13003) );
  AND3_X1 U14527 ( .A1(n13003), .A2(n14271), .A3(n14477), .ZN(n13004) );
  XNOR2_X1 U14528 ( .A(n14489), .B(n13006), .ZN(n14649) );
  NAND2_X1 U14529 ( .A1(n14649), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14650) );
  INV_X1 U14530 ( .A(n13006), .ZN(n13007) );
  OR2_X1 U14531 ( .A1(n13007), .A2(n14489), .ZN(n13008) );
  INV_X1 U14532 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21748) );
  XNOR2_X1 U14533 ( .A(n13056), .B(n21748), .ZN(n14673) );
  INV_X1 U14534 ( .A(n13009), .ZN(n13012) );
  NAND2_X1 U14535 ( .A1(n13010), .A2(n12981), .ZN(n13011) );
  NAND2_X1 U14536 ( .A1(n13012), .A2(n13011), .ZN(n13013) );
  INV_X1 U14537 ( .A(n13016), .ZN(n13015) );
  NAND2_X1 U14538 ( .A1(n13015), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15023) );
  NAND2_X1 U14539 ( .A1(n13016), .A2(n22237), .ZN(n13017) );
  NAND2_X1 U14540 ( .A1(n15023), .A2(n13017), .ZN(n15528) );
  NAND2_X1 U14541 ( .A1(n17417), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13020) );
  NAND2_X2 U14542 ( .A1(n17321), .A2(n13024), .ZN(n16514) );
  NAND2_X1 U14543 ( .A1(n22236), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14544 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U14545 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U14546 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U14547 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13025) );
  NAND4_X1 U14548 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13034) );
  AOI22_X1 U14549 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U14550 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14551 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13030) );
  AOI22_X1 U14552 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13029) );
  NAND4_X1 U14553 ( .A1(n13032), .A2(n13031), .A3(n13030), .A4(n13029), .ZN(
        n13033) );
  OR2_X1 U14554 ( .A1(n13034), .A2(n13033), .ZN(n13048) );
  AOI22_X1 U14555 ( .A1(n13239), .A2(n13048), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13220), .ZN(n13035) );
  INV_X1 U14556 ( .A(n13046), .ZN(n13044) );
  INV_X1 U14557 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13040) );
  INV_X1 U14558 ( .A(n13036), .ZN(n13037) );
  NAND2_X1 U14559 ( .A1(n13037), .A2(n13049), .ZN(n13039) );
  OAI211_X1 U14560 ( .C1(n13232), .C2(n13040), .A(n13039), .B(n13038), .ZN(
        n13041) );
  INV_X1 U14561 ( .A(n13041), .ZN(n13042) );
  NAND2_X1 U14562 ( .A1(n13044), .A2(n13265), .ZN(n13047) );
  NAND2_X1 U14563 ( .A1(n13047), .A2(n13076), .ZN(n13253) );
  INV_X1 U14564 ( .A(n13190), .ZN(n13206) );
  INV_X1 U14565 ( .A(n13048), .ZN(n13052) );
  NAND2_X1 U14566 ( .A1(n13050), .A2(n13049), .ZN(n13051) );
  NAND2_X1 U14567 ( .A1(n13051), .A2(n13052), .ZN(n13080) );
  OAI21_X1 U14568 ( .B1(n13052), .B2(n13051), .A(n13080), .ZN(n13054) );
  AOI21_X1 U14569 ( .B1(n13054), .B2(n17412), .A(n13053), .ZN(n13055) );
  OAI21_X1 U14570 ( .B1(n13253), .B2(n13206), .A(n13055), .ZN(n14672) );
  NAND2_X1 U14571 ( .A1(n14673), .A2(n14672), .ZN(n14671) );
  NAND2_X1 U14572 ( .A1(n13056), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13057) );
  INV_X1 U14573 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15909) );
  OR2_X1 U14574 ( .A1(n13059), .A2(n13058), .ZN(n13064) );
  INV_X1 U14575 ( .A(n15023), .ZN(n13060) );
  INV_X1 U14576 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13197) );
  NAND2_X1 U14577 ( .A1(n13060), .A2(n13197), .ZN(n22589) );
  NAND2_X1 U14578 ( .A1(n15023), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13061) );
  NAND2_X1 U14579 ( .A1(n22589), .A2(n13061), .ZN(n22309) );
  INV_X1 U14580 ( .A(n13752), .ZN(n13062) );
  AOI22_X1 U14581 ( .A1(n22309), .A2(n13062), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17417), .ZN(n13063) );
  XNOR2_X2 U14582 ( .A(n17321), .B(n14988), .ZN(n17360) );
  AOI22_X1 U14583 ( .A1(n13088), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U14584 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U14585 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U14586 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13065) );
  NAND4_X1 U14587 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13065), .ZN(
        n13074) );
  AOI22_X1 U14588 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13719), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U14589 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U14590 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U14591 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13069) );
  NAND4_X1 U14592 ( .A1(n13072), .A2(n13071), .A3(n13070), .A4(n13069), .ZN(
        n13073) );
  OR2_X1 U14593 ( .A1(n13074), .A2(n13073), .ZN(n13079) );
  AOI22_X1 U14594 ( .A1(n13239), .A2(n13079), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13220), .ZN(n13075) );
  NAND2_X1 U14595 ( .A1(n14641), .A2(n13076), .ZN(n13078) );
  AND2_X1 U14596 ( .A1(n13080), .A2(n13079), .ZN(n13123) );
  OAI21_X1 U14597 ( .B1(n13080), .B2(n13079), .A(n17412), .ZN(n13081) );
  OAI22_X1 U14598 ( .A1(n15517), .A2(n13206), .B1(n13123), .B2(n13081), .ZN(
        n14825) );
  NAND2_X1 U14599 ( .A1(n14826), .A2(n14825), .ZN(n14824) );
  NAND2_X1 U14600 ( .A1(n13082), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13083) );
  NAND2_X1 U14601 ( .A1(n14824), .A2(n13083), .ZN(n20329) );
  AOI22_X1 U14602 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U14603 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13693), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U14604 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13708), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14605 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n13692), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U14606 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13095) );
  AOI22_X1 U14607 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13720), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U14608 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U14609 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U14610 ( .A1(n13089), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13090) );
  NAND4_X1 U14611 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        n13094) );
  OR2_X1 U14612 ( .A1(n13095), .A2(n13094), .ZN(n13122) );
  NAND2_X1 U14613 ( .A1(n13239), .A2(n13122), .ZN(n13097) );
  NAND2_X1 U14614 ( .A1(n13220), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13096) );
  NAND2_X1 U14615 ( .A1(n13097), .A2(n13096), .ZN(n13118) );
  XNOR2_X1 U14616 ( .A(n13115), .B(n13118), .ZN(n13286) );
  NAND2_X1 U14617 ( .A1(n13286), .A2(n13190), .ZN(n13101) );
  INV_X1 U14618 ( .A(n13122), .ZN(n13098) );
  XNOR2_X1 U14619 ( .A(n13123), .B(n13098), .ZN(n13099) );
  NAND2_X1 U14620 ( .A1(n13099), .A2(n17412), .ZN(n13100) );
  NAND2_X1 U14621 ( .A1(n13101), .A2(n13100), .ZN(n13102) );
  INV_X1 U14622 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15910) );
  XNOR2_X1 U14623 ( .A(n13102), .B(n15910), .ZN(n20328) );
  NAND2_X1 U14624 ( .A1(n20329), .A2(n20328), .ZN(n20327) );
  NAND2_X1 U14625 ( .A1(n13102), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13103) );
  INV_X1 U14626 ( .A(n13118), .ZN(n13114) );
  AOI22_X1 U14627 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U14628 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U14629 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U14630 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13104) );
  NAND4_X1 U14631 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13113) );
  AOI22_X1 U14632 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U14633 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U14634 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U14635 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13108) );
  NAND4_X1 U14636 ( .A1(n13111), .A2(n13110), .A3(n13109), .A4(n13108), .ZN(
        n13112) );
  OR2_X1 U14637 ( .A1(n13113), .A2(n13112), .ZN(n13141) );
  AOI22_X1 U14638 ( .A1(n13239), .A2(n13141), .B1(n13220), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U14639 ( .B1(n13115), .B2(n13114), .A(n13116), .ZN(n13121) );
  INV_X1 U14640 ( .A(n13116), .ZN(n13117) );
  NAND2_X1 U14641 ( .A1(n13121), .A2(n13140), .ZN(n13293) );
  OR2_X1 U14642 ( .A1(n13293), .A2(n13206), .ZN(n13126) );
  NAND2_X1 U14643 ( .A1(n13123), .A2(n13122), .ZN(n13142) );
  XNOR2_X1 U14644 ( .A(n13141), .B(n13142), .ZN(n13124) );
  NAND2_X1 U14645 ( .A1(n17412), .A2(n13124), .ZN(n13125) );
  NAND2_X1 U14646 ( .A1(n13126), .A2(n13125), .ZN(n13127) );
  INV_X1 U14647 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21777) );
  XNOR2_X1 U14648 ( .A(n13127), .B(n21777), .ZN(n20334) );
  NAND2_X1 U14649 ( .A1(n20335), .A2(n20334), .ZN(n20333) );
  NAND2_X1 U14650 ( .A1(n13127), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U14651 ( .A1(n20333), .A2(n13128), .ZN(n20340) );
  AOI22_X1 U14652 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U14653 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U14654 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U14655 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13129) );
  NAND4_X1 U14656 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13138) );
  AOI22_X1 U14657 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U14658 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U14659 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U14660 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13133) );
  NAND4_X1 U14661 ( .A1(n13136), .A2(n13135), .A3(n13134), .A4(n13133), .ZN(
        n13137) );
  OR2_X1 U14662 ( .A1(n13138), .A2(n13137), .ZN(n13153) );
  AOI22_X1 U14663 ( .A1(n13239), .A2(n13153), .B1(n13220), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13139) );
  NAND2_X1 U14664 ( .A1(n13140), .A2(n13139), .ZN(n13298) );
  NAND3_X1 U14665 ( .A1(n13162), .A2(n13190), .A3(n13298), .ZN(n13147) );
  INV_X1 U14666 ( .A(n13141), .ZN(n13143) );
  NOR2_X1 U14667 ( .A1(n13143), .A2(n13142), .ZN(n13154) );
  INV_X1 U14668 ( .A(n13154), .ZN(n13144) );
  XNOR2_X1 U14669 ( .A(n13153), .B(n13144), .ZN(n13145) );
  NAND2_X1 U14670 ( .A1(n17412), .A2(n13145), .ZN(n13146) );
  NAND2_X1 U14671 ( .A1(n13147), .A2(n13146), .ZN(n13148) );
  INV_X1 U14672 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21762) );
  XNOR2_X1 U14673 ( .A(n13148), .B(n21762), .ZN(n20339) );
  NAND2_X1 U14674 ( .A1(n20340), .A2(n20339), .ZN(n20342) );
  NAND2_X1 U14675 ( .A1(n13148), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13149) );
  NAND2_X1 U14676 ( .A1(n13239), .A2(n13165), .ZN(n13151) );
  NAND2_X1 U14677 ( .A1(n13220), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13150) );
  NAND2_X1 U14678 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U14679 ( .A1(n13305), .A2(n13190), .ZN(n13157) );
  NAND2_X1 U14680 ( .A1(n13154), .A2(n13153), .ZN(n13163) );
  XNOR2_X1 U14681 ( .A(n13165), .B(n13163), .ZN(n13155) );
  NAND2_X1 U14682 ( .A1(n17412), .A2(n13155), .ZN(n13156) );
  NAND2_X1 U14683 ( .A1(n13157), .A2(n13156), .ZN(n13158) );
  INV_X1 U14684 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21789) );
  XNOR2_X1 U14685 ( .A(n13158), .B(n21789), .ZN(n20347) );
  NAND2_X1 U14686 ( .A1(n13158), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13159) );
  AND3_X1 U14687 ( .A1(n13190), .A2(n13160), .A3(n13165), .ZN(n13161) );
  INV_X1 U14688 ( .A(n13163), .ZN(n13164) );
  NAND3_X1 U14689 ( .A1(n17412), .A2(n13165), .A3(n13164), .ZN(n13166) );
  NAND2_X1 U14690 ( .A1(n13169), .A2(n13166), .ZN(n13167) );
  INV_X1 U14691 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21798) );
  XNOR2_X1 U14692 ( .A(n13167), .B(n21798), .ZN(n15696) );
  XNOR2_X1 U14693 ( .A(n13169), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15730) );
  INV_X1 U14694 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21811) );
  NAND2_X2 U14695 ( .A1(n15729), .A2(n13168), .ZN(n16388) );
  AOI21_X1 U14696 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n20353), .ZN(n16400) );
  NOR2_X1 U14697 ( .A1(n20353), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16403) );
  INV_X1 U14698 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21729) );
  NOR3_X1 U14699 ( .A1(n16400), .A2(n16403), .A3(n16404), .ZN(n16391) );
  INV_X1 U14700 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21730) );
  NAND2_X1 U14701 ( .A1(n13169), .A2(n21730), .ZN(n13170) );
  NAND2_X1 U14702 ( .A1(n16391), .A2(n13170), .ZN(n20373) );
  NAND2_X1 U14703 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21870) );
  INV_X1 U14704 ( .A(n21870), .ZN(n13172) );
  AND2_X1 U14705 ( .A1(n13169), .A2(n13172), .ZN(n20376) );
  NOR2_X1 U14706 ( .A1(n13169), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20377) );
  AOI21_X1 U14707 ( .B1(n20376), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n20377), .ZN(n13178) );
  OR2_X1 U14708 ( .A1(n13169), .A2(n21730), .ZN(n13173) );
  INV_X1 U14709 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15685) );
  INV_X1 U14710 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20354) );
  INV_X1 U14711 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21822) );
  AND3_X1 U14712 ( .A1(n15685), .A2(n20354), .A3(n21822), .ZN(n13174) );
  NOR2_X1 U14713 ( .A1(n13169), .A2(n13174), .ZN(n16390) );
  INV_X1 U14714 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21865) );
  INV_X1 U14715 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21842) );
  NAND2_X1 U14716 ( .A1(n21865), .A2(n21842), .ZN(n21869) );
  NOR2_X1 U14717 ( .A1(n21869), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13175) );
  NOR2_X1 U14718 ( .A1(n13169), .A2(n13175), .ZN(n13176) );
  NOR2_X1 U14719 ( .A1(n16377), .A2(n13176), .ZN(n13177) );
  AND2_X1 U14720 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16485) );
  NAND2_X1 U14721 ( .A1(n16485), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21888) );
  INV_X1 U14722 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16357) );
  NOR2_X1 U14723 ( .A1(n21888), .A2(n16357), .ZN(n13179) );
  INV_X1 U14724 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21874) );
  INV_X1 U14725 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16359) );
  INV_X1 U14726 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16490) );
  NAND4_X1 U14727 ( .A1(n21874), .A2(n16359), .A3(n16357), .A4(n16490), .ZN(
        n13180) );
  OAI21_X1 U14728 ( .B1(n16356), .B2(n13180), .A(n20353), .ZN(n16349) );
  NAND2_X1 U14729 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15926) );
  INV_X1 U14730 ( .A(n15926), .ZN(n15904) );
  NAND2_X1 U14731 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16301) );
  NAND2_X1 U14732 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16433) );
  INV_X1 U14733 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21912) );
  INV_X1 U14734 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16461) );
  INV_X1 U14735 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20389) );
  NAND3_X1 U14736 ( .A1(n21912), .A2(n16461), .A3(n20389), .ZN(n16302) );
  OAI21_X1 U14737 ( .B1(n16300), .B2(n16302), .A(n20353), .ZN(n16324) );
  NOR2_X1 U14738 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16442) );
  NAND3_X1 U14739 ( .A1(n16324), .A2(n13181), .A3(n16442), .ZN(n16283) );
  INV_X1 U14740 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16432) );
  INV_X1 U14741 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16508) );
  XNOR2_X1 U14742 ( .A(n13169), .B(n16508), .ZN(n13187) );
  INV_X1 U14743 ( .A(n13187), .ZN(n13183) );
  NOR2_X1 U14744 ( .A1(n20353), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13185) );
  INV_X1 U14745 ( .A(n13185), .ZN(n13182) );
  NAND2_X1 U14746 ( .A1(n13183), .A2(n13182), .ZN(n13189) );
  OAI21_X1 U14747 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n20353), .ZN(n13186) );
  INV_X1 U14748 ( .A(n13186), .ZN(n13184) );
  OAI21_X1 U14749 ( .B1(n13185), .B2(n13184), .A(n16508), .ZN(n13188) );
  NAND2_X1 U14750 ( .A1(n22238), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13192) );
  NAND2_X1 U14751 ( .A1(n12981), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13191) );
  NAND2_X1 U14752 ( .A1(n13192), .A2(n13191), .ZN(n13203) );
  NAND2_X1 U14753 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n22251), .ZN(
        n13207) );
  NAND2_X1 U14754 ( .A1(n13193), .A2(n13192), .ZN(n13218) );
  OR2_X1 U14755 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n22237), .ZN(
        n13194) );
  NAND2_X1 U14756 ( .A1(n13218), .A2(n13194), .ZN(n13196) );
  NAND2_X1 U14757 ( .A1(n22237), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13195) );
  NAND2_X1 U14758 ( .A1(n13196), .A2(n13195), .ZN(n13231) );
  NAND2_X1 U14759 ( .A1(n13197), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13227) );
  NAND2_X1 U14760 ( .A1(n13058), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13198) );
  AND2_X1 U14761 ( .A1(n13227), .A2(n13198), .ZN(n13230) );
  NAND2_X1 U14762 ( .A1(n13231), .A2(n13230), .ZN(n13200) );
  INV_X1 U14763 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17424) );
  NAND2_X1 U14764 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17424), .ZN(
        n13199) );
  NAND3_X1 U14765 ( .A1(n13200), .A2(n13227), .A3(n13199), .ZN(n13201) );
  INV_X1 U14766 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17326) );
  NAND2_X1 U14767 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17326), .ZN(
        n13228) );
  INV_X1 U14768 ( .A(n13207), .ZN(n13202) );
  XNOR2_X1 U14769 ( .A(n13203), .B(n13202), .ZN(n14260) );
  OAI22_X1 U14770 ( .A1(n13232), .A2(n14260), .B1(n22122), .B2(n14477), .ZN(
        n13208) );
  INV_X1 U14771 ( .A(n13208), .ZN(n13204) );
  OAI21_X1 U14772 ( .B1(n13219), .B2(n22386), .A(n13204), .ZN(n13216) );
  INV_X1 U14773 ( .A(n14260), .ZN(n13205) );
  OAI21_X1 U14774 ( .B1(n13206), .B2(n13239), .A(n13205), .ZN(n13215) );
  OAI21_X1 U14775 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n22251), .A(
        n13207), .ZN(n13209) );
  AOI211_X1 U14776 ( .C1(n14471), .C2(n15821), .A(n13209), .B(n13221), .ZN(
        n13213) );
  NOR3_X1 U14777 ( .A1(n13208), .A2(n14467), .A3(n14260), .ZN(n13212) );
  INV_X1 U14778 ( .A(n13209), .ZN(n13210) );
  AOI21_X1 U14779 ( .B1(n13239), .B2(n13210), .A(n13238), .ZN(n13211) );
  NOR3_X1 U14780 ( .A1(n13213), .A2(n13212), .A3(n13211), .ZN(n13214) );
  AOI21_X1 U14781 ( .B1(n13216), .B2(n13215), .A(n13214), .ZN(n13226) );
  XNOR2_X1 U14782 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13217) );
  XNOR2_X1 U14783 ( .A(n13218), .B(n13217), .ZN(n14257) );
  AOI211_X1 U14784 ( .C1(n13220), .C2(n14257), .A(n13221), .B(n13222), .ZN(
        n13225) );
  INV_X1 U14785 ( .A(n13221), .ZN(n13224) );
  INV_X1 U14786 ( .A(n13222), .ZN(n13223) );
  OAI22_X1 U14787 ( .A1(n13226), .A2(n13225), .B1(n13224), .B2(n13223), .ZN(
        n13234) );
  INV_X1 U14788 ( .A(n13227), .ZN(n13229) );
  OAI22_X1 U14789 ( .A1(n13231), .A2(n13230), .B1(n13229), .B2(n13228), .ZN(
        n14258) );
  NAND2_X1 U14790 ( .A1(n13232), .A2(n14258), .ZN(n13233) );
  AOI22_X1 U14791 ( .A1(n13234), .A2(n13233), .B1(n13238), .B2(n14258), .ZN(
        n13235) );
  INV_X1 U14792 ( .A(n13235), .ZN(n13236) );
  NAND2_X1 U14793 ( .A1(n13242), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22135) );
  NOR2_X2 U14794 ( .A1(n15830), .A2(n22135), .ZN(n14305) );
  NAND2_X1 U14795 ( .A1(n16505), .A2(n22236), .ZN(n13243) );
  NAND2_X1 U14796 ( .A1(n13243), .A2(n14271), .ZN(n13246) );
  NOR2_X1 U14797 ( .A1(n14637), .A2(n15892), .ZN(n13245) );
  OR2_X1 U14798 ( .A1(n13245), .A2(n13244), .ZN(n14466) );
  NOR2_X1 U14799 ( .A1(n13246), .A2(n14466), .ZN(n14458) );
  AND2_X1 U14800 ( .A1(n14458), .A2(n14471), .ZN(n17399) );
  NAND2_X1 U14801 ( .A1(n13247), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13398) );
  AND2_X1 U14802 ( .A1(n13248), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13280) );
  INV_X1 U14803 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13250) );
  INV_X1 U14804 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22282) );
  NAND2_X1 U14805 ( .A1(n22253), .A2(n22282), .ZN(n14876) );
  INV_X1 U14806 ( .A(n14876), .ZN(n13736) );
  XNOR2_X1 U14807 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14904) );
  AND2_X1 U14808 ( .A1(n22253), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13740) );
  AOI21_X1 U14809 ( .B1(n13736), .B2(n14904), .A(n13740), .ZN(n13249) );
  OAI21_X1 U14810 ( .B1(n13734), .B2(n13250), .A(n13249), .ZN(n13251) );
  AOI21_X1 U14811 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13280), .A(
        n13251), .ZN(n13252) );
  NAND2_X1 U14812 ( .A1(n13740), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13272) );
  NAND2_X1 U14813 ( .A1(n13254), .A2(n13272), .ZN(n14677) );
  INV_X1 U14814 ( .A(n14677), .ZN(n13271) );
  OAI21_X1 U14815 ( .B1(n14843), .B2(n15524), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n14485) );
  OR2_X1 U14816 ( .A1(n14894), .A2(n13398), .ZN(n13259) );
  INV_X1 U14817 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U14818 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n22253), .ZN(
        n13255) );
  OAI21_X1 U14819 ( .B1(n13734), .B2(n13256), .A(n13255), .ZN(n13257) );
  AOI21_X1 U14820 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13280), .A(
        n13257), .ZN(n13258) );
  OR2_X1 U14821 ( .A1(n14485), .A2(n14484), .ZN(n14487) );
  NAND2_X1 U14822 ( .A1(n14484), .A2(n13736), .ZN(n13260) );
  NAND2_X1 U14823 ( .A1(n14487), .A2(n13260), .ZN(n14586) );
  INV_X1 U14824 ( .A(n13261), .ZN(n13264) );
  INV_X1 U14825 ( .A(n13262), .ZN(n13263) );
  NAND2_X1 U14826 ( .A1(n13264), .A2(n13263), .ZN(n13266) );
  INV_X1 U14827 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n13267) );
  INV_X1 U14828 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14646) );
  OAI22_X1 U14829 ( .A1(n13734), .A2(n13267), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14646), .ZN(n13268) );
  AOI21_X1 U14830 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13280), .A(
        n13268), .ZN(n13269) );
  NAND2_X1 U14831 ( .A1(n14586), .A2(n14585), .ZN(n14676) );
  NAND2_X1 U14832 ( .A1(n13271), .A2(n13270), .ZN(n14674) );
  INV_X1 U14833 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n14822) );
  NAND3_X1 U14834 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13289) );
  INV_X1 U14835 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U14836 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U14837 ( .A1(n13274), .A2(n13273), .ZN(n13275) );
  NAND2_X1 U14838 ( .A1(n13289), .A2(n13275), .ZN(n15052) );
  AOI22_X1 U14839 ( .A1(n13736), .A2(n15052), .B1(n13740), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13276) );
  OAI21_X1 U14840 ( .B1(n13734), .B2(n14822), .A(n13276), .ZN(n13277) );
  AOI21_X1 U14841 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13280), .A(
        n13277), .ZN(n13278) );
  OAI21_X1 U14842 ( .B1(n15517), .B2(n13398), .A(n13278), .ZN(n14813) );
  NAND2_X1 U14843 ( .A1(n14814), .A2(n14813), .ZN(n14717) );
  INV_X1 U14844 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13279) );
  XNOR2_X1 U14845 ( .A(n13289), .B(n13279), .ZN(n21948) );
  INV_X1 U14846 ( .A(n13280), .ZN(n13283) );
  NAND2_X1 U14847 ( .A1(n22253), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13282) );
  NAND2_X1 U14848 ( .A1(n13741), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13281) );
  OAI211_X1 U14849 ( .C1(n13283), .C2(n17326), .A(n13282), .B(n13281), .ZN(
        n13284) );
  MUX2_X1 U14850 ( .A(n21948), .B(n13284), .S(n14876), .Z(n13285) );
  INV_X1 U14851 ( .A(n13289), .ZN(n13287) );
  AOI21_X1 U14852 ( .B1(n13287), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U14853 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13288) );
  OR2_X1 U14854 ( .A1(n13290), .A2(n13294), .ZN(n21960) );
  AOI22_X1 U14855 ( .A1(n21960), .A2(n13736), .B1(n13740), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U14856 ( .A1(n13741), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n13291) );
  OAI211_X1 U14857 ( .C1(n13293), .C2(n13398), .A(n13292), .B(n13291), .ZN(
        n14857) );
  NAND2_X1 U14858 ( .A1(n14718), .A2(n14857), .ZN(n14856) );
  INV_X1 U14859 ( .A(n14856), .ZN(n13300) );
  INV_X1 U14860 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n15092) );
  NOR2_X1 U14861 ( .A1(n13294), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13295) );
  OR2_X1 U14862 ( .A1(n13301), .A2(n13295), .ZN(n21975) );
  AOI22_X1 U14863 ( .A1(n21975), .A2(n13736), .B1(n13740), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13296) );
  OAI21_X1 U14864 ( .B1(n13734), .B2(n15092), .A(n13296), .ZN(n13297) );
  INV_X1 U14865 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15117) );
  NAND2_X1 U14866 ( .A1(n13301), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13322) );
  OR2_X1 U14867 ( .A1(n13301), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13302) );
  NAND2_X1 U14868 ( .A1(n13322), .A2(n13302), .ZN(n21986) );
  AOI22_X1 U14869 ( .A1(n21986), .A2(n13736), .B1(n13740), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13303) );
  OAI21_X1 U14870 ( .B1(n13734), .B2(n15117), .A(n13303), .ZN(n13304) );
  INV_X1 U14871 ( .A(n15108), .ZN(n13306) );
  AOI22_X1 U14872 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U14873 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13719), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U14874 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U14875 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13307) );
  NAND4_X1 U14876 ( .A1(n13310), .A2(n13309), .A3(n13308), .A4(n13307), .ZN(
        n13316) );
  AOI22_X1 U14877 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14878 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U14879 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U14880 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13311) );
  NAND4_X1 U14881 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n13311), .ZN(
        n13315) );
  OAI21_X1 U14882 ( .B1(n13316), .B2(n13315), .A(n13463), .ZN(n13321) );
  NAND2_X1 U14883 ( .A1(n13741), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13320) );
  INV_X1 U14884 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13317) );
  XNOR2_X1 U14885 ( .A(n13322), .B(n13317), .ZN(n15699) );
  NAND2_X1 U14886 ( .A1(n15699), .A2(n13736), .ZN(n13319) );
  NAND2_X1 U14887 ( .A1(n13740), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13318) );
  AND4_X1 U14888 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n15120) );
  XOR2_X1 U14889 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13346), .Z(n15732) );
  AOI22_X1 U14890 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13326) );
  AOI22_X1 U14891 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U14892 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U14893 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13323) );
  NAND4_X1 U14894 ( .A1(n13326), .A2(n13325), .A3(n13324), .A4(n13323), .ZN(
        n13332) );
  AOI22_X1 U14895 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13330) );
  AOI22_X1 U14896 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U14897 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14898 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13327) );
  NAND4_X1 U14899 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        n13331) );
  OR2_X1 U14900 ( .A1(n13332), .A2(n13331), .ZN(n13333) );
  AOI22_X1 U14901 ( .A1(n13463), .A2(n13333), .B1(n13740), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U14902 ( .A1(n13741), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13334) );
  OAI211_X1 U14903 ( .C1(n15732), .C2(n14876), .A(n13335), .B(n13334), .ZN(
        n15572) );
  AOI22_X1 U14904 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U14905 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U14906 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U14907 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13358), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13336) );
  NAND4_X1 U14908 ( .A1(n13339), .A2(n13338), .A3(n13337), .A4(n13336), .ZN(
        n13345) );
  AOI22_X1 U14909 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U14910 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14911 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U14912 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13340) );
  NAND4_X1 U14913 ( .A1(n13343), .A2(n13342), .A3(n13341), .A4(n13340), .ZN(
        n13344) );
  NOR2_X1 U14914 ( .A1(n13345), .A2(n13344), .ZN(n13350) );
  NAND2_X1 U14915 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13351) );
  INV_X1 U14916 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13347) );
  XNOR2_X1 U14917 ( .A(n13351), .B(n13347), .ZN(n16416) );
  NAND2_X1 U14918 ( .A1(n16416), .A2(n13736), .ZN(n13349) );
  AOI22_X1 U14919 ( .A1(n13741), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13740), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13348) );
  OAI211_X1 U14920 ( .C1(n13350), .C2(n13398), .A(n13349), .B(n13348), .ZN(
        n15679) );
  OR2_X1 U14921 ( .A1(n13352), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13353) );
  NAND2_X1 U14922 ( .A1(n13352), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13399) );
  NAND2_X1 U14923 ( .A1(n13353), .A2(n13399), .ZN(n21995) );
  NAND2_X1 U14924 ( .A1(n21995), .A2(n13736), .ZN(n13357) );
  INV_X1 U14925 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15765) );
  INV_X1 U14926 ( .A(n13740), .ZN(n13481) );
  INV_X1 U14927 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13354) );
  OAI22_X1 U14928 ( .A1(n13734), .A2(n15765), .B1(n13481), .B2(n13354), .ZN(
        n13355) );
  INV_X1 U14929 ( .A(n13355), .ZN(n13356) );
  NAND2_X1 U14930 ( .A1(n13357), .A2(n13356), .ZN(n15763) );
  AOI22_X1 U14931 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U14932 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U14933 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13360) );
  AOI22_X1 U14934 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13359) );
  NAND4_X1 U14935 ( .A1(n13362), .A2(n13361), .A3(n13360), .A4(n13359), .ZN(
        n13369) );
  AOI22_X1 U14936 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U14937 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U14938 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U14939 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13364) );
  NAND4_X1 U14940 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n13364), .ZN(
        n13368) );
  OR2_X1 U14941 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  AND2_X1 U14942 ( .A1(n13463), .A2(n13370), .ZN(n16144) );
  INV_X1 U14943 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13371) );
  XOR2_X1 U14944 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13403), .Z(
        n16409) );
  AOI22_X1 U14945 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13717), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U14946 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U14947 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U14948 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13372) );
  NAND4_X1 U14949 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13381) );
  AOI22_X1 U14950 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U14951 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U14952 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U14953 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13376) );
  NAND4_X1 U14954 ( .A1(n13379), .A2(n13378), .A3(n13377), .A4(n13376), .ZN(
        n13380) );
  OAI21_X1 U14955 ( .B1(n13381), .B2(n13380), .A(n13463), .ZN(n13384) );
  NAND2_X1 U14956 ( .A1(n13741), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13383) );
  NAND2_X1 U14957 ( .A1(n13740), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13382) );
  AND3_X1 U14958 ( .A1(n13384), .A2(n13383), .A3(n13382), .ZN(n13385) );
  OAI21_X1 U14959 ( .B1(n16409), .B2(n14876), .A(n13385), .ZN(n16148) );
  INV_X1 U14960 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n16280) );
  AOI22_X1 U14961 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13720), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U14962 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U14963 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n13692), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13387) );
  AOI22_X1 U14964 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13386) );
  NAND4_X1 U14965 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13396) );
  AOI22_X1 U14966 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13708), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U14967 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13422), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U14968 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13693), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13392) );
  AOI22_X1 U14969 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13391) );
  NAND4_X1 U14970 ( .A1(n13394), .A2(n13393), .A3(n13392), .A4(n13391), .ZN(
        n13395) );
  NOR2_X1 U14971 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  OR2_X1 U14972 ( .A1(n13398), .A2(n13397), .ZN(n13402) );
  XNOR2_X1 U14973 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n13399), .ZN(
        n22000) );
  OAI22_X1 U14974 ( .A1(n22000), .A2(n14876), .B1(n13481), .B2(n13371), .ZN(
        n13400) );
  INV_X1 U14975 ( .A(n13400), .ZN(n13401) );
  OAI211_X1 U14976 ( .C1(n13734), .C2(n16280), .A(n13402), .B(n13401), .ZN(
        n16210) );
  AND2_X1 U14977 ( .A1(n16148), .A2(n16210), .ZN(n15800) );
  NAND2_X1 U14978 ( .A1(n13469), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13487) );
  XNOR2_X1 U14979 ( .A(n13487), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n22030) );
  NAND2_X1 U14980 ( .A1(n22030), .A2(n13736), .ZN(n13420) );
  AOI22_X1 U14981 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U14982 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U14983 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U14984 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13404) );
  NAND4_X1 U14985 ( .A1(n13407), .A2(n13406), .A3(n13405), .A4(n13404), .ZN(
        n13416) );
  AOI22_X1 U14986 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U14987 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13412) );
  NAND2_X1 U14988 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13409) );
  NAND2_X1 U14989 ( .A1(n13709), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13408) );
  AND3_X1 U14990 ( .A1(n13409), .A2(n13408), .A3(n14876), .ZN(n13411) );
  AOI22_X1 U14991 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13410) );
  NAND4_X1 U14992 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13415) );
  INV_X1 U14993 ( .A(n16505), .ZN(n13414) );
  NAND2_X1 U14994 ( .A1(n13414), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13702) );
  NAND2_X1 U14995 ( .A1(n13702), .A2(n14876), .ZN(n13551) );
  OAI21_X1 U14996 ( .B1(n13416), .B2(n13415), .A(n13551), .ZN(n13418) );
  AOI22_X1 U14997 ( .A1(n13741), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22253), .ZN(n13417) );
  NAND2_X1 U14998 ( .A1(n13418), .A2(n13417), .ZN(n13419) );
  NAND2_X1 U14999 ( .A1(n13420), .A2(n13419), .ZN(n16192) );
  INV_X1 U15000 ( .A(n16192), .ZN(n13486) );
  INV_X1 U15001 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16384) );
  XNOR2_X1 U15002 ( .A(n13421), .B(n16384), .ZN(n22019) );
  NAND2_X1 U15003 ( .A1(n22019), .A2(n13736), .ZN(n13438) );
  AOI22_X1 U15004 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U15005 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15006 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U15008 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13423) );
  NAND4_X1 U15009 ( .A1(n13426), .A2(n13425), .A3(n13424), .A4(n13423), .ZN(
        n13434) );
  NAND2_X1 U15010 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13428) );
  NAND2_X1 U15011 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13427) );
  AND3_X1 U15012 ( .A1(n13428), .A2(n13427), .A3(n14876), .ZN(n13432) );
  AOI22_X1 U15013 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U15014 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15015 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13429) );
  NAND4_X1 U15016 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n13429), .ZN(
        n13433) );
  OAI21_X1 U15017 ( .B1(n13434), .B2(n13433), .A(n13551), .ZN(n13436) );
  AOI22_X1 U15018 ( .A1(n13741), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n22253), .ZN(n13435) );
  NAND2_X1 U15019 ( .A1(n13436), .A2(n13435), .ZN(n13437) );
  NAND2_X1 U15020 ( .A1(n13438), .A2(n13437), .ZN(n16195) );
  INV_X1 U15021 ( .A(n16195), .ZN(n13468) );
  XOR2_X1 U15022 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n13439), .Z(
        n20366) );
  INV_X1 U15023 ( .A(n20366), .ZN(n16140) );
  AOI22_X1 U15024 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U15025 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U15026 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U15027 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13440) );
  NAND4_X1 U15028 ( .A1(n13443), .A2(n13442), .A3(n13441), .A4(n13440), .ZN(
        n13449) );
  AOI22_X1 U15029 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13447) );
  AOI22_X1 U15030 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13693), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U15031 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U15032 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13444) );
  NAND4_X1 U15033 ( .A1(n13447), .A2(n13446), .A3(n13445), .A4(n13444), .ZN(
        n13448) );
  OAI21_X1 U15034 ( .B1(n13449), .B2(n13448), .A(n13463), .ZN(n13452) );
  NAND2_X1 U15035 ( .A1(n13741), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U15036 ( .A1(n13740), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13450) );
  NAND3_X1 U15037 ( .A1(n13452), .A2(n13451), .A3(n13450), .ZN(n13453) );
  AOI21_X1 U15038 ( .B1(n16140), .B2(n13736), .A(n13453), .ZN(n16133) );
  INV_X1 U15039 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16395) );
  XNOR2_X1 U15040 ( .A(n13454), .B(n16395), .ZN(n22010) );
  AOI22_X1 U15041 ( .A1(n13741), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13740), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15042 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U15043 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15044 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U15045 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13455) );
  NAND4_X1 U15046 ( .A1(n13458), .A2(n13457), .A3(n13456), .A4(n13455), .ZN(
        n13465) );
  AOI22_X1 U15047 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U15048 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13722), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U15049 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U15050 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13459) );
  NAND4_X1 U15051 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13459), .ZN(
        n13464) );
  OAI21_X1 U15052 ( .B1(n13465), .B2(n13464), .A(n13463), .ZN(n13466) );
  OAI211_X1 U15053 ( .C1(n22010), .C2(n14876), .A(n13467), .B(n13466), .ZN(
        n15802) );
  INV_X1 U15054 ( .A(n15802), .ZN(n15801) );
  NOR2_X1 U15055 ( .A1(n16133), .A2(n15801), .ZN(n16130) );
  AND2_X1 U15056 ( .A1(n13468), .A2(n16130), .ZN(n16118) );
  XOR2_X1 U15057 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13469), .Z(
        n20380) );
  INV_X1 U15058 ( .A(n13702), .ZN(n13731) );
  AOI22_X1 U15059 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U15060 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15061 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U15062 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13470) );
  NAND4_X1 U15063 ( .A1(n13473), .A2(n13472), .A3(n13471), .A4(n13470), .ZN(
        n13479) );
  AOI22_X1 U15064 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U15065 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U15066 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U15067 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13474) );
  NAND4_X1 U15068 ( .A1(n13477), .A2(n13476), .A3(n13475), .A4(n13474), .ZN(
        n13478) );
  OR2_X1 U15069 ( .A1(n13479), .A2(n13478), .ZN(n13484) );
  INV_X1 U15070 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13482) );
  INV_X1 U15071 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13480) );
  OAI22_X1 U15072 ( .A1(n13734), .A2(n13482), .B1(n13481), .B2(n13480), .ZN(
        n13483) );
  AOI21_X1 U15073 ( .B1(n13731), .B2(n13484), .A(n13483), .ZN(n13485) );
  OAI21_X1 U15074 ( .B1(n20380), .B2(n14876), .A(n13485), .ZN(n16119) );
  AND2_X1 U15075 ( .A1(n16118), .A2(n16119), .ZN(n16120) );
  AND2_X1 U15076 ( .A1(n13486), .A2(n16120), .ZN(n16189) );
  INV_X1 U15077 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n22027) );
  OR2_X1 U15078 ( .A1(n13488), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13489) );
  NAND2_X1 U15079 ( .A1(n13488), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13535) );
  NAND2_X1 U15080 ( .A1(n13489), .A2(n13535), .ZN(n22041) );
  AOI22_X1 U15081 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13493) );
  AOI22_X1 U15082 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13492) );
  AOI22_X1 U15083 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U15084 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13490) );
  NAND4_X1 U15085 ( .A1(n13493), .A2(n13492), .A3(n13491), .A4(n13490), .ZN(
        n13499) );
  AOI22_X1 U15086 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U15087 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13496) );
  AOI22_X1 U15088 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U15089 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13494) );
  NAND4_X1 U15090 ( .A1(n13497), .A2(n13496), .A3(n13495), .A4(n13494), .ZN(
        n13498) );
  OAI21_X1 U15091 ( .B1(n13499), .B2(n13498), .A(n13731), .ZN(n13502) );
  NAND2_X1 U15092 ( .A1(n13741), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U15093 ( .A1(n22253), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13500) );
  NAND4_X1 U15094 ( .A1(n13502), .A2(n14876), .A3(n13501), .A4(n13500), .ZN(
        n13503) );
  OAI21_X1 U15095 ( .B1(n22041), .B2(n14876), .A(n13503), .ZN(n20305) );
  INV_X1 U15096 ( .A(n20305), .ZN(n13504) );
  AND2_X1 U15097 ( .A1(n16189), .A2(n13504), .ZN(n13505) );
  AOI22_X1 U15098 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U15099 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U15100 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13507) );
  AOI22_X1 U15101 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13506) );
  NAND4_X1 U15102 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        n13515) );
  AOI22_X1 U15103 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13693), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U15104 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13708), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U15105 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13511) );
  AOI22_X1 U15106 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13510) );
  NAND4_X1 U15107 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        n13514) );
  NOR2_X1 U15108 ( .A1(n13515), .A2(n13514), .ZN(n13518) );
  INV_X1 U15109 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16366) );
  AOI21_X1 U15110 ( .B1(n16366), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13516) );
  AOI21_X1 U15111 ( .B1(n13741), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13516), .ZN(
        n13517) );
  OAI21_X1 U15112 ( .B1(n13702), .B2(n13518), .A(n13517), .ZN(n13520) );
  XNOR2_X1 U15113 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n13535), .ZN(
        n22049) );
  NAND2_X1 U15114 ( .A1(n13736), .A2(n22049), .ZN(n13519) );
  AND2_X1 U15115 ( .A1(n13520), .A2(n13519), .ZN(n16186) );
  AOI22_X1 U15116 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13719), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U15117 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U15118 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U15119 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13521) );
  NAND4_X1 U15120 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n13521), .ZN(
        n13530) );
  AOI22_X1 U15121 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U15122 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U15123 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U15124 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13525) );
  NAND4_X1 U15125 ( .A1(n13528), .A2(n13527), .A3(n13526), .A4(n13525), .ZN(
        n13529) );
  NOR2_X1 U15126 ( .A1(n13530), .A2(n13529), .ZN(n13534) );
  INV_X1 U15127 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15598) );
  NAND2_X1 U15128 ( .A1(n22253), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13531) );
  OAI211_X1 U15129 ( .C1(n13734), .C2(n15598), .A(n14876), .B(n13531), .ZN(
        n13532) );
  INV_X1 U15130 ( .A(n13532), .ZN(n13533) );
  OAI21_X1 U15131 ( .B1(n13702), .B2(n13534), .A(n13533), .ZN(n13539) );
  INV_X1 U15132 ( .A(n13535), .ZN(n13536) );
  NAND2_X1 U15133 ( .A1(n13537), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13583) );
  OAI21_X1 U15134 ( .B1(n13537), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n13583), .ZN(n22068) );
  OR2_X1 U15135 ( .A1(n22068), .A2(n14876), .ZN(n13538) );
  AND2_X1 U15136 ( .A1(n13539), .A2(n13538), .ZN(n16355) );
  AOI22_X1 U15137 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13708), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U15138 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13719), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U15139 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15140 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13540) );
  NAND4_X1 U15141 ( .A1(n13543), .A2(n13542), .A3(n13541), .A4(n13540), .ZN(
        n13553) );
  AOI22_X1 U15142 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13544), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U15143 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13546) );
  NAND2_X1 U15144 ( .A1(n13707), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13545) );
  AND3_X1 U15145 ( .A1(n13546), .A2(n13545), .A3(n14876), .ZN(n13549) );
  AOI22_X1 U15146 ( .A1(n13710), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U15147 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13547) );
  NAND4_X1 U15148 ( .A1(n13550), .A2(n13549), .A3(n13548), .A4(n13547), .ZN(
        n13552) );
  OAI21_X1 U15149 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(n13556) );
  NAND2_X1 U15150 ( .A1(n13741), .A2(P1_EAX_REG_22__SCAN_IN), .ZN(n13555) );
  NAND2_X1 U15151 ( .A1(n22253), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13554) );
  NAND3_X1 U15152 ( .A1(n13556), .A2(n13555), .A3(n13554), .ZN(n13558) );
  XNOR2_X1 U15153 ( .A(n13583), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n22080) );
  NAND2_X1 U15154 ( .A1(n22080), .A2(n13736), .ZN(n13557) );
  NAND2_X1 U15155 ( .A1(n13558), .A2(n13557), .ZN(n16173) );
  AOI22_X1 U15156 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U15157 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13561) );
  AOI22_X1 U15158 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13560) );
  AOI22_X1 U15159 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13559) );
  NAND4_X1 U15160 ( .A1(n13562), .A2(n13561), .A3(n13560), .A4(n13559), .ZN(
        n13568) );
  AOI22_X1 U15161 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U15162 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U15163 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U15164 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13563) );
  NAND4_X1 U15165 ( .A1(n13566), .A2(n13565), .A3(n13564), .A4(n13563), .ZN(
        n13567) );
  NOR2_X1 U15166 ( .A1(n13568), .A2(n13567), .ZN(n13598) );
  AOI22_X1 U15167 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13572) );
  AOI22_X1 U15168 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U15169 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U15170 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13569) );
  NAND4_X1 U15171 ( .A1(n13572), .A2(n13571), .A3(n13570), .A4(n13569), .ZN(
        n13578) );
  AOI22_X1 U15172 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13576) );
  AOI22_X1 U15173 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13575) );
  AOI22_X1 U15174 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13574) );
  AOI22_X1 U15175 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13573) );
  NAND4_X1 U15176 ( .A1(n13576), .A2(n13575), .A3(n13574), .A4(n13573), .ZN(
        n13577) );
  NOR2_X1 U15177 ( .A1(n13578), .A2(n13577), .ZN(n13599) );
  XNOR2_X1 U15178 ( .A(n13598), .B(n13599), .ZN(n13582) );
  INV_X1 U15179 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n15583) );
  NAND2_X1 U15180 ( .A1(n22253), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13579) );
  OAI211_X1 U15181 ( .C1(n13734), .C2(n15583), .A(n14876), .B(n13579), .ZN(
        n13580) );
  INV_X1 U15182 ( .A(n13580), .ZN(n13581) );
  OAI21_X1 U15183 ( .B1(n13702), .B2(n13582), .A(n13581), .ZN(n13587) );
  INV_X1 U15184 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n22074) );
  NOR2_X1 U15185 ( .A1(n13583), .A2(n22074), .ZN(n13584) );
  OR2_X1 U15186 ( .A1(n13584), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13585) );
  NAND2_X1 U15187 ( .A1(n13584), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13604) );
  NAND2_X1 U15188 ( .A1(n13585), .A2(n13604), .ZN(n22097) );
  OR2_X1 U15189 ( .A1(n22097), .A2(n14876), .ZN(n13586) );
  NAND2_X1 U15190 ( .A1(n13587), .A2(n13586), .ZN(n20295) );
  XNOR2_X1 U15191 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n13604), .ZN(
        n22106) );
  AOI22_X1 U15192 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13591) );
  AOI22_X1 U15193 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13590) );
  AOI22_X1 U15194 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U15195 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13588) );
  NAND4_X1 U15196 ( .A1(n13591), .A2(n13590), .A3(n13589), .A4(n13588), .ZN(
        n13597) );
  AOI22_X1 U15197 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U15198 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U15199 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U15200 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13592) );
  NAND4_X1 U15201 ( .A1(n13595), .A2(n13594), .A3(n13593), .A4(n13592), .ZN(
        n13596) );
  OR2_X1 U15202 ( .A1(n13597), .A2(n13596), .ZN(n13617) );
  NOR2_X1 U15203 ( .A1(n13599), .A2(n13598), .ZN(n13618) );
  XOR2_X1 U15204 ( .A(n13617), .B(n13618), .Z(n13602) );
  INV_X1 U15205 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15592) );
  OAI21_X1 U15206 ( .B1(n22282), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n22253), .ZN(n13600) );
  OAI21_X1 U15207 ( .B1(n13734), .B2(n15592), .A(n13600), .ZN(n13601) );
  AOI21_X1 U15208 ( .B1(n13602), .B2(n13731), .A(n13601), .ZN(n13603) );
  AOI21_X1 U15209 ( .B1(n13736), .B2(n22106), .A(n13603), .ZN(n16169) );
  INV_X1 U15210 ( .A(n13604), .ZN(n13605) );
  NAND2_X1 U15211 ( .A1(n13606), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13639) );
  OAI21_X1 U15212 ( .B1(n13606), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n13639), .ZN(n16334) );
  AOI22_X1 U15213 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U15214 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U15215 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15216 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13607) );
  NAND4_X1 U15217 ( .A1(n13610), .A2(n13609), .A3(n13608), .A4(n13607), .ZN(
        n13616) );
  AOI22_X1 U15218 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U15219 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U15220 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15221 ( .A1(n13718), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13611) );
  NAND4_X1 U15222 ( .A1(n13614), .A2(n13613), .A3(n13612), .A4(n13611), .ZN(
        n13615) );
  NOR2_X1 U15223 ( .A1(n13616), .A2(n13615), .ZN(n13634) );
  NAND2_X1 U15224 ( .A1(n13618), .A2(n13617), .ZN(n13633) );
  XNOR2_X1 U15225 ( .A(n13634), .B(n13633), .ZN(n13621) );
  OAI21_X1 U15226 ( .B1(n22282), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n22253), .ZN(n13620) );
  NAND2_X1 U15227 ( .A1(n13741), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n13619) );
  OAI211_X1 U15228 ( .C1(n13621), .C2(n13702), .A(n13620), .B(n13619), .ZN(
        n13622) );
  OAI21_X1 U15229 ( .B1(n14876), .B2(n16334), .A(n13622), .ZN(n16107) );
  XNOR2_X1 U15230 ( .A(n13639), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16322) );
  AOI22_X1 U15231 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U15232 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13625) );
  AOI22_X1 U15233 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U15234 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13623) );
  NAND4_X1 U15235 ( .A1(n13626), .A2(n13625), .A3(n13624), .A4(n13623), .ZN(
        n13632) );
  AOI22_X1 U15236 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U15237 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13629) );
  AOI22_X1 U15238 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U15239 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13627) );
  NAND4_X1 U15240 ( .A1(n13630), .A2(n13629), .A3(n13628), .A4(n13627), .ZN(
        n13631) );
  OR2_X1 U15241 ( .A1(n13632), .A2(n13631), .ZN(n13644) );
  NOR2_X1 U15242 ( .A1(n13634), .A2(n13633), .ZN(n13645) );
  XOR2_X1 U15243 ( .A(n13644), .B(n13645), .Z(n13637) );
  INV_X1 U15244 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n15600) );
  OAI21_X1 U15245 ( .B1(n22282), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n22253), .ZN(n13635) );
  OAI21_X1 U15246 ( .B1(n13734), .B2(n15600), .A(n13635), .ZN(n13636) );
  AOI21_X1 U15247 ( .B1(n13637), .B2(n13731), .A(n13636), .ZN(n13638) );
  AOI21_X1 U15248 ( .B1(n13736), .B2(n16322), .A(n13638), .ZN(n16095) );
  INV_X1 U15249 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16320) );
  NOR2_X1 U15250 ( .A1(n13639), .A2(n16320), .ZN(n13640) );
  NAND2_X1 U15251 ( .A1(n13640), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13678) );
  INV_X1 U15252 ( .A(n13640), .ZN(n13642) );
  INV_X1 U15253 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U15254 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  NAND2_X1 U15255 ( .A1(n13678), .A2(n13643), .ZN(n16316) );
  NAND2_X1 U15256 ( .A1(n13645), .A2(n13644), .ZN(n13672) );
  AOI22_X1 U15257 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U15258 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13693), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13650) );
  AOI22_X1 U15259 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13722), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U15260 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13712), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13648) );
  NAND4_X1 U15261 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13657) );
  AOI22_X1 U15262 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U15263 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13708), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U15264 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U15265 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13652) );
  NAND4_X1 U15266 ( .A1(n13655), .A2(n13654), .A3(n13653), .A4(n13652), .ZN(
        n13656) );
  NOR2_X1 U15267 ( .A1(n13657), .A2(n13656), .ZN(n13673) );
  XNOR2_X1 U15268 ( .A(n13672), .B(n13673), .ZN(n13660) );
  AOI21_X1 U15269 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n22253), .A(
        n13736), .ZN(n13659) );
  NAND2_X1 U15270 ( .A1(n13741), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n13658) );
  OAI211_X1 U15271 ( .C1(n13660), .C2(n13702), .A(n13659), .B(n13658), .ZN(
        n13661) );
  OAI21_X1 U15272 ( .B1(n14876), .B2(n16316), .A(n13661), .ZN(n16087) );
  XNOR2_X1 U15273 ( .A(n13678), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16311) );
  AOI22_X1 U15274 ( .A1(n13646), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U15275 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13664) );
  AOI22_X1 U15276 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U15277 ( .A1(n13691), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13662) );
  NAND4_X1 U15278 ( .A1(n13665), .A2(n13664), .A3(n13663), .A4(n13662), .ZN(
        n13671) );
  AOI22_X1 U15279 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U15280 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U15281 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13667) );
  AOI22_X1 U15282 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13666) );
  NAND4_X1 U15283 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n13670) );
  OR2_X1 U15284 ( .A1(n13671), .A2(n13670), .ZN(n13684) );
  NOR2_X1 U15285 ( .A1(n13673), .A2(n13672), .ZN(n13685) );
  XOR2_X1 U15286 ( .A(n13684), .B(n13685), .Z(n13676) );
  INV_X1 U15287 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15604) );
  OAI21_X1 U15288 ( .B1(n22282), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n22253), .ZN(n13674) );
  OAI21_X1 U15289 ( .B1(n13734), .B2(n15604), .A(n13674), .ZN(n13675) );
  AOI21_X1 U15290 ( .B1(n13676), .B2(n13731), .A(n13675), .ZN(n13677) );
  AOI21_X1 U15291 ( .B1(n13736), .B2(n16311), .A(n13677), .ZN(n16074) );
  INV_X1 U15292 ( .A(n13678), .ZN(n13679) );
  NAND2_X1 U15293 ( .A1(n13680), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13749) );
  INV_X1 U15294 ( .A(n13680), .ZN(n13682) );
  INV_X1 U15295 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13681) );
  NAND2_X1 U15296 ( .A1(n13682), .A2(n13681), .ZN(n13683) );
  NAND2_X1 U15297 ( .A1(n13749), .A2(n13683), .ZN(n16296) );
  NAND2_X1 U15298 ( .A1(n13685), .A2(n13684), .ZN(n13705) );
  AOI22_X1 U15299 ( .A1(n13686), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13647), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13690) );
  AOI22_X1 U15300 ( .A1(n12903), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13689) );
  AOI22_X1 U15301 ( .A1(n13721), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11160), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U15302 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13687) );
  NAND4_X1 U15303 ( .A1(n13690), .A2(n13689), .A3(n13688), .A4(n13687), .ZN(
        n13699) );
  AOI22_X1 U15304 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13710), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U15305 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13696) );
  AOI22_X1 U15306 ( .A1(n13692), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13691), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13695) );
  AOI22_X1 U15307 ( .A1(n13693), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13694) );
  NAND4_X1 U15308 ( .A1(n13697), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        n13698) );
  NOR2_X1 U15309 ( .A1(n13699), .A2(n13698), .ZN(n13706) );
  XNOR2_X1 U15310 ( .A(n13705), .B(n13706), .ZN(n13703) );
  AOI21_X1 U15311 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22253), .A(
        n13736), .ZN(n13701) );
  NAND2_X1 U15312 ( .A1(n13741), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13700) );
  OAI211_X1 U15313 ( .C1(n13703), .C2(n13702), .A(n13701), .B(n13700), .ZN(
        n13704) );
  OAI21_X1 U15314 ( .B1(n14876), .B2(n16296), .A(n13704), .ZN(n16066) );
  NOR2_X1 U15315 ( .A1(n13706), .A2(n13705), .ZN(n13730) );
  AOI22_X1 U15316 ( .A1(n13708), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13707), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U15317 ( .A1(n13710), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13709), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U15318 ( .A1(n13647), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13363), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U15319 ( .A1(n13712), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13711), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13713) );
  NAND4_X1 U15320 ( .A1(n13716), .A2(n13715), .A3(n13714), .A4(n13713), .ZN(
        n13728) );
  AOI22_X1 U15321 ( .A1(n13717), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13646), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U15322 ( .A1(n13719), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13718), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U15323 ( .A1(n13720), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12903), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13724) );
  AOI22_X1 U15324 ( .A1(n13722), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13721), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13723) );
  NAND4_X1 U15325 ( .A1(n13726), .A2(n13725), .A3(n13724), .A4(n13723), .ZN(
        n13727) );
  NOR2_X1 U15326 ( .A1(n13728), .A2(n13727), .ZN(n13729) );
  XNOR2_X1 U15327 ( .A(n13730), .B(n13729), .ZN(n13732) );
  NAND2_X1 U15328 ( .A1(n13732), .A2(n13731), .ZN(n13739) );
  INV_X1 U15329 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15606) );
  OAI21_X1 U15330 ( .B1(n22282), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n22253), .ZN(n13733) );
  OAI21_X1 U15331 ( .B1(n13734), .B2(n15606), .A(n13733), .ZN(n13735) );
  INV_X1 U15332 ( .A(n13735), .ZN(n13738) );
  XNOR2_X1 U15333 ( .A(n13749), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16287) );
  AND2_X1 U15334 ( .A1(n16287), .A2(n13736), .ZN(n13737) );
  AOI21_X1 U15335 ( .B1(n13739), .B2(n13738), .A(n13737), .ZN(n16053) );
  NAND2_X1 U15336 ( .A1(n16065), .A2(n16053), .ZN(n13744) );
  AOI22_X1 U15337 ( .A1(n13741), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13740), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13742) );
  INV_X1 U15338 ( .A(n13742), .ZN(n13743) );
  AND3_X1 U15339 ( .A1(n22122), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13745) );
  NOR2_X2 U15340 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22292) );
  INV_X1 U15341 ( .A(n20385), .ZN(n16413) );
  INV_X1 U15342 ( .A(n22292), .ZN(n22358) );
  NAND2_X1 U15343 ( .A1(n22358), .A2(n13752), .ZN(n21695) );
  AND2_X1 U15344 ( .A1(n21695), .A2(n22122), .ZN(n13746) );
  NAND2_X1 U15345 ( .A1(n22122), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17411) );
  NAND2_X1 U15346 ( .A1(n22282), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13747) );
  AND2_X1 U15347 ( .A1(n17411), .A2(n13747), .ZN(n14491) );
  INV_X1 U15348 ( .A(n14491), .ZN(n13748) );
  INV_X1 U15349 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16289) );
  INV_X1 U15350 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13750) );
  XNOR2_X1 U15351 ( .A(n13751), .B(n13750), .ZN(n14896) );
  OR2_X1 U15352 ( .A1(n13752), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21915) );
  INV_X1 U15353 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20257) );
  NOR2_X1 U15354 ( .A1(n21915), .A2(n20257), .ZN(n15923) );
  AOI21_X1 U15355 ( .B1(n20388), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15923), .ZN(n13753) );
  OAI21_X1 U15356 ( .B1(n20395), .B2(n14896), .A(n13753), .ZN(n13754) );
  OAI21_X1 U15357 ( .B1(n15934), .B2(n22113), .A(n13755), .ZN(P1_U2968) );
  INV_X1 U15358 ( .A(n14805), .ZN(n13781) );
  NAND2_X1 U15359 ( .A1(n11881), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U15360 ( .A1(n13788), .A2(n19593), .ZN(n13778) );
  AND2_X1 U15361 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13767) );
  NAND2_X1 U15362 ( .A1(n13767), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13769) );
  NAND2_X1 U15363 ( .A1(n19594), .A2(n19593), .ZN(n19694) );
  AOI21_X1 U15364 ( .B1(n13769), .B2(n19563), .A(n19694), .ZN(n13758) );
  INV_X1 U15365 ( .A(n13769), .ZN(n13757) );
  NAND2_X1 U15366 ( .A1(n13757), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19714) );
  AND2_X1 U15367 ( .A1(n13758), .A2(n19714), .ZN(n19555) );
  AOI21_X1 U15368 ( .B1(n13778), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19555), .ZN(n13759) );
  NAND2_X1 U15369 ( .A1(n13760), .A2(n13759), .ZN(n13765) );
  NAND2_X1 U15370 ( .A1(n13762), .A2(n13761), .ZN(n13793) );
  NOR2_X1 U15371 ( .A1(n13793), .A2(n13763), .ZN(n13764) );
  OAI21_X1 U15372 ( .B1(n13765), .B2(n13764), .A(n13787), .ZN(n13766) );
  INV_X1 U15373 ( .A(n13767), .ZN(n19659) );
  NAND2_X1 U15374 ( .A1(n19659), .A2(n19592), .ZN(n13768) );
  NAND2_X1 U15375 ( .A1(n13769), .A2(n13768), .ZN(n19556) );
  NOR2_X1 U15376 ( .A1(n19556), .A2(n19694), .ZN(n13770) );
  AOI21_X1 U15377 ( .B1(n13778), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13770), .ZN(n13771) );
  INV_X1 U15378 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13772) );
  NOR2_X1 U15379 ( .A1(n13793), .A2(n13772), .ZN(n13773) );
  NAND2_X1 U15380 ( .A1(n13774), .A2(n13773), .ZN(n13785) );
  NAND2_X1 U15381 ( .A1(n18637), .A2(n13781), .ZN(n13777) );
  AOI22_X1 U15382 ( .A1(n13778), .A2(n11196), .B1(n19708), .B2(n19612), .ZN(
        n13776) );
  INV_X1 U15383 ( .A(n13793), .ZN(n14035) );
  NAND2_X1 U15384 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13782) );
  NAND2_X1 U15385 ( .A1(n13778), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13779) );
  OAI21_X1 U15386 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19659), .ZN(n19614) );
  OR2_X1 U15387 ( .A1(n19614), .A2(n19694), .ZN(n19672) );
  NAND2_X1 U15388 ( .A1(n13779), .A2(n19672), .ZN(n13780) );
  INV_X1 U15389 ( .A(n13782), .ZN(n13783) );
  NOR2_X1 U15390 ( .A1(n15632), .A2(n13783), .ZN(n13784) );
  NAND2_X1 U15391 ( .A1(n14415), .A2(n14416), .ZN(n13786) );
  INV_X1 U15392 ( .A(n13788), .ZN(n13789) );
  NAND2_X1 U15393 ( .A1(n13789), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13790) );
  NOR2_X1 U15394 ( .A1(n13793), .A2(n13792), .ZN(n14531) );
  NAND2_X1 U15395 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U15396 ( .A1(n15098), .A2(n15552), .ZN(n15551) );
  AOI22_X1 U15397 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U15398 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13798) );
  NAND2_X1 U15399 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13797) );
  AND2_X1 U15400 ( .A1(n13798), .A2(n13797), .ZN(n13801) );
  AOI22_X1 U15401 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U15402 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13799) );
  NAND4_X1 U15403 ( .A1(n13802), .A2(n13801), .A3(n13800), .A4(n13799), .ZN(
        n13811) );
  INV_X1 U15404 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13804) );
  INV_X1 U15405 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13803) );
  OAI22_X1 U15406 ( .A1(n13926), .A2(n13804), .B1(n13924), .B2(n13803), .ZN(
        n13805) );
  INV_X1 U15407 ( .A(n13805), .ZN(n13809) );
  AOI22_X1 U15408 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U15409 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13807) );
  NAND2_X1 U15410 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13806) );
  NAND4_X1 U15411 ( .A1(n13809), .A2(n13808), .A3(n13807), .A4(n13806), .ZN(
        n13810) );
  NOR2_X1 U15412 ( .A1(n13811), .A2(n13810), .ZN(n15576) );
  AOI22_X1 U15413 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U15414 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U15415 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13813) );
  AND2_X1 U15416 ( .A1(n13814), .A2(n13813), .ZN(n13817) );
  AOI22_X1 U15417 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U15418 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13815) );
  NAND4_X1 U15419 ( .A1(n13818), .A2(n13817), .A3(n13816), .A4(n13815), .ZN(
        n13827) );
  INV_X1 U15420 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13820) );
  INV_X1 U15421 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13819) );
  OAI22_X1 U15422 ( .A1(n13926), .A2(n13820), .B1(n13924), .B2(n13819), .ZN(
        n13821) );
  INV_X1 U15423 ( .A(n13821), .ZN(n13825) );
  AOI22_X1 U15424 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13824) );
  AOI22_X1 U15425 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13823) );
  NAND2_X1 U15426 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13822) );
  NAND4_X1 U15427 ( .A1(n13825), .A2(n13824), .A3(n13823), .A4(n13822), .ZN(
        n13826) );
  NOR2_X1 U15428 ( .A1(n13827), .A2(n13826), .ZN(n15716) );
  AOI22_X1 U15429 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U15430 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U15431 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13828) );
  AND2_X1 U15432 ( .A1(n13829), .A2(n13828), .ZN(n13832) );
  AOI22_X1 U15433 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U15434 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13830) );
  NAND4_X1 U15435 ( .A1(n13833), .A2(n13832), .A3(n13831), .A4(n13830), .ZN(
        n13842) );
  INV_X1 U15436 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13835) );
  INV_X1 U15437 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13834) );
  OAI22_X1 U15438 ( .A1(n13926), .A2(n13835), .B1(n13924), .B2(n13834), .ZN(
        n13836) );
  INV_X1 U15439 ( .A(n13836), .ZN(n13840) );
  AOI22_X1 U15440 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U15441 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U15442 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13837) );
  NAND4_X1 U15443 ( .A1(n13840), .A2(n13839), .A3(n13838), .A4(n13837), .ZN(
        n13841) );
  OR2_X1 U15444 ( .A1(n13842), .A2(n13841), .ZN(n15768) );
  AOI22_X1 U15445 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U15446 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U15447 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13843) );
  AND2_X1 U15448 ( .A1(n13844), .A2(n13843), .ZN(n13847) );
  AOI22_X1 U15449 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U15450 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13845) );
  NAND4_X1 U15451 ( .A1(n13848), .A2(n13847), .A3(n13846), .A4(n13845), .ZN(
        n13857) );
  INV_X1 U15452 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13849) );
  OAI22_X1 U15453 ( .A1(n13926), .A2(n13850), .B1(n13924), .B2(n13849), .ZN(
        n13851) );
  INV_X1 U15454 ( .A(n13851), .ZN(n13855) );
  AOI22_X1 U15455 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U15456 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U15457 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n13852) );
  NAND4_X1 U15458 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  OR2_X1 U15459 ( .A1(n13857), .A2(n13856), .ZN(n16599) );
  AOI22_X1 U15460 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U15461 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U15462 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13858) );
  AND2_X1 U15463 ( .A1(n13859), .A2(n13858), .ZN(n13862) );
  AOI22_X1 U15464 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U15465 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13860) );
  NAND4_X1 U15466 ( .A1(n13863), .A2(n13862), .A3(n13861), .A4(n13860), .ZN(
        n13872) );
  INV_X1 U15467 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13864) );
  OAI22_X1 U15468 ( .A1(n13926), .A2(n13865), .B1(n13924), .B2(n13864), .ZN(
        n13866) );
  INV_X1 U15469 ( .A(n13866), .ZN(n13870) );
  AOI22_X1 U15470 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13869) );
  AOI22_X1 U15471 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U15472 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13867) );
  NAND4_X1 U15473 ( .A1(n13870), .A2(n13869), .A3(n13868), .A4(n13867), .ZN(
        n13871) );
  NOR2_X1 U15474 ( .A1(n13872), .A2(n13871), .ZN(n15808) );
  INV_X1 U15475 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U15476 ( .A1(n13912), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U15477 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13913), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13874) );
  OAI211_X1 U15478 ( .C1(n13877), .C2(n13876), .A(n13875), .B(n13874), .ZN(
        n13888) );
  INV_X1 U15479 ( .A(n13930), .ZN(n13903) );
  AOI22_X1 U15480 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U15481 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13878) );
  OAI211_X1 U15482 ( .C1(n13903), .C2(n13880), .A(n13879), .B(n13878), .ZN(
        n13887) );
  AOI22_X1 U15483 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U15484 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13881) );
  NAND2_X1 U15485 ( .A1(n13882), .A2(n13881), .ZN(n13886) );
  INV_X1 U15486 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13883) );
  OAI22_X1 U15487 ( .A1(n13926), .A2(n13884), .B1(n13924), .B2(n13883), .ZN(
        n13885) );
  NOR4_X1 U15488 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n16595) );
  INV_X1 U15489 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13891) );
  INV_X1 U15490 ( .A(n13913), .ZN(n13890) );
  INV_X1 U15491 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13889) );
  OAI22_X1 U15492 ( .A1(n13892), .A2(n13891), .B1(n13890), .B2(n13889), .ZN(
        n13898) );
  INV_X1 U15493 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13895) );
  INV_X1 U15494 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13893) );
  OAI22_X1 U15495 ( .A1(n13896), .A2(n13895), .B1(n13894), .B2(n13893), .ZN(
        n13897) );
  AOI211_X1 U15496 ( .C1(n13914), .C2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n13898), .B(n13897), .ZN(n13910) );
  NOR2_X1 U15497 ( .A1(n13926), .A2(n13899), .ZN(n13905) );
  AOI22_X1 U15498 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15499 ( .A1(n12101), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13900) );
  OAI211_X1 U15500 ( .C1(n13903), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        n13904) );
  AOI211_X1 U15501 ( .C1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .C2(n13906), .A(
        n13905), .B(n13904), .ZN(n13909) );
  AOI22_X1 U15502 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U15503 ( .A1(n12144), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13918), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13907) );
  NAND4_X1 U15504 ( .A1(n13910), .A2(n13909), .A3(n13908), .A4(n13907), .ZN(
        n16587) );
  AOI22_X1 U15505 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n13912), .B1(
        n13911), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U15506 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13913), .B1(
        n12096), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U15507 ( .A1(n13914), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13915) );
  AND2_X1 U15508 ( .A1(n13916), .A2(n13915), .ZN(n13921) );
  AOI22_X1 U15509 ( .A1(n13917), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12241), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13918), .B1(
        n12144), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13919) );
  NAND4_X1 U15511 ( .A1(n13922), .A2(n13921), .A3(n13920), .A4(n13919), .ZN(
        n13936) );
  INV_X1 U15512 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13925) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13923) );
  OAI22_X1 U15514 ( .A1(n13926), .A2(n13925), .B1(n13924), .B2(n13923), .ZN(
        n13927) );
  INV_X1 U15515 ( .A(n13927), .ZN(n13934) );
  AOI22_X1 U15516 ( .A1(n12176), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13928), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U15517 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12101), .B1(
        n13929), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13932) );
  NAND2_X1 U15518 ( .A1(n13930), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13931) );
  NAND4_X1 U15519 ( .A1(n13934), .A2(n13933), .A3(n13932), .A4(n13931), .ZN(
        n13935) );
  NOR2_X1 U15520 ( .A1(n13936), .A2(n13935), .ZN(n13957) );
  AOI22_X1 U15521 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13948) );
  AND2_X1 U15522 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13939) );
  OR2_X1 U15523 ( .A1(n13939), .A2(n13938), .ZN(n14087) );
  INV_X1 U15524 ( .A(n14087), .ZN(n14041) );
  NAND2_X1 U15525 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13942) );
  NAND2_X1 U15526 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13941) );
  AND3_X1 U15527 ( .A1(n14041), .A2(n13942), .A3(n13941), .ZN(n13947) );
  AOI22_X1 U15528 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U15529 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13945) );
  NAND4_X1 U15530 ( .A1(n13948), .A2(n13947), .A3(n13946), .A4(n13945), .ZN(
        n13956) );
  AOI22_X1 U15531 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U15532 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U15533 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13952) );
  NAND2_X1 U15534 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13950) );
  NAND2_X1 U15535 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13949) );
  AND3_X1 U15536 ( .A1(n13950), .A2(n14087), .A3(n13949), .ZN(n13951) );
  NAND4_X1 U15537 ( .A1(n13954), .A2(n13953), .A3(n13952), .A4(n13951), .ZN(
        n13955) );
  NAND2_X1 U15538 ( .A1(n13956), .A2(n13955), .ZN(n13958) );
  XNOR2_X1 U15539 ( .A(n13957), .B(n13958), .ZN(n16583) );
  INV_X1 U15540 ( .A(n13957), .ZN(n13960) );
  INV_X1 U15541 ( .A(n13958), .ZN(n13959) );
  NAND2_X1 U15542 ( .A1(n13960), .A2(n13959), .ZN(n13976) );
  AOI22_X1 U15543 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U15544 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13962) );
  NAND2_X1 U15545 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13961) );
  AND3_X1 U15546 ( .A1(n14041), .A2(n13962), .A3(n13961), .ZN(n13965) );
  AOI22_X1 U15547 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U15548 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13963) );
  NAND4_X1 U15549 ( .A1(n13966), .A2(n13965), .A3(n13964), .A4(n13963), .ZN(
        n13974) );
  AOI22_X1 U15550 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U15551 ( .A1(n11163), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13971) );
  AOI22_X1 U15552 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U15553 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13968) );
  NAND2_X1 U15554 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13967) );
  AND3_X1 U15555 ( .A1(n13968), .A2(n14087), .A3(n13967), .ZN(n13969) );
  NAND4_X1 U15556 ( .A1(n13972), .A2(n13971), .A3(n13970), .A4(n13969), .ZN(
        n13973) );
  NAND2_X1 U15557 ( .A1(n13974), .A2(n13973), .ZN(n13978) );
  INV_X1 U15558 ( .A(n13976), .ZN(n13975) );
  NAND2_X1 U15559 ( .A1(n14035), .A2(n13975), .ZN(n13977) );
  NOR2_X1 U15560 ( .A1(n13976), .A2(n13978), .ZN(n13993) );
  AOI22_X1 U15561 ( .A1(n13978), .A2(n13977), .B1(n13993), .B2(n12069), .ZN(
        n16575) );
  NAND2_X1 U15562 ( .A1(n16574), .A2(n16575), .ZN(n13997) );
  AOI22_X1 U15563 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13984) );
  NAND2_X1 U15564 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13980) );
  NAND2_X1 U15565 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13979) );
  AND3_X1 U15566 ( .A1(n14041), .A2(n13980), .A3(n13979), .ZN(n13983) );
  AOI22_X1 U15567 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U15568 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13981) );
  NAND4_X1 U15569 ( .A1(n13984), .A2(n13983), .A3(n13982), .A4(n13981), .ZN(
        n13992) );
  AOI22_X1 U15570 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U15571 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U15572 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13988) );
  NAND2_X1 U15573 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13986) );
  NAND2_X1 U15574 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13985) );
  AND3_X1 U15575 ( .A1(n13986), .A2(n14087), .A3(n13985), .ZN(n13987) );
  NAND4_X1 U15576 ( .A1(n13990), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13991) );
  AND2_X1 U15577 ( .A1(n13992), .A2(n13991), .ZN(n13995) );
  NAND2_X1 U15578 ( .A1(n13993), .A2(n13995), .ZN(n14033) );
  OAI211_X1 U15579 ( .C1(n13993), .C2(n13995), .A(n14033), .B(n14035), .ZN(
        n13998) );
  INV_X1 U15580 ( .A(n13998), .ZN(n13994) );
  INV_X1 U15581 ( .A(n13995), .ZN(n13996) );
  NOR2_X1 U15582 ( .A1(n12069), .A2(n13996), .ZN(n16565) );
  AOI22_X1 U15583 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14004) );
  NAND2_X1 U15584 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14000) );
  NAND2_X1 U15585 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13999) );
  AND3_X1 U15586 ( .A1(n14041), .A2(n14000), .A3(n13999), .ZN(n14003) );
  AOI22_X1 U15587 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U15588 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14001) );
  NAND4_X1 U15589 ( .A1(n14004), .A2(n14003), .A3(n14002), .A4(n14001), .ZN(
        n14012) );
  AOI22_X1 U15590 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U15591 ( .A1(n11162), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14084), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U15592 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12083), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14008) );
  NAND2_X1 U15593 ( .A1(n11204), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14006) );
  NAND2_X1 U15594 ( .A1(n14080), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14005) );
  AND3_X1 U15595 ( .A1(n14006), .A2(n14005), .A3(n14087), .ZN(n14007) );
  NAND4_X1 U15596 ( .A1(n14010), .A2(n14009), .A3(n14008), .A4(n14007), .ZN(
        n14011) );
  AND2_X1 U15597 ( .A1(n14012), .A2(n14011), .ZN(n14031) );
  XNOR2_X1 U15598 ( .A(n14033), .B(n14031), .ZN(n14013) );
  AND2_X1 U15599 ( .A1(n14013), .A2(n14035), .ZN(n14014) );
  NAND2_X1 U15600 ( .A1(n12609), .A2(n14031), .ZN(n16560) );
  AOI22_X1 U15601 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14022) );
  AOI22_X1 U15602 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U15603 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14020) );
  NAND2_X1 U15604 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14018) );
  NAND2_X1 U15605 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14017) );
  AND3_X1 U15606 ( .A1(n14018), .A2(n14087), .A3(n14017), .ZN(n14019) );
  NAND4_X1 U15607 ( .A1(n14022), .A2(n14021), .A3(n14020), .A4(n14019), .ZN(
        n14030) );
  AOI22_X1 U15608 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U15609 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14024) );
  NAND2_X1 U15610 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14023) );
  AND3_X1 U15611 ( .A1(n14041), .A2(n14024), .A3(n14023), .ZN(n14027) );
  AOI22_X1 U15612 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U15613 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14025) );
  NAND4_X1 U15614 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        n14029) );
  NAND2_X1 U15615 ( .A1(n14030), .A2(n14029), .ZN(n14038) );
  INV_X1 U15616 ( .A(n14038), .ZN(n14037) );
  INV_X1 U15617 ( .A(n14031), .ZN(n14032) );
  OR2_X1 U15618 ( .A1(n14033), .A2(n14032), .ZN(n14034) );
  INV_X1 U15619 ( .A(n14034), .ZN(n14036) );
  OR2_X1 U15620 ( .A1(n14034), .A2(n14038), .ZN(n16540) );
  OAI211_X1 U15621 ( .C1(n14037), .C2(n14036), .A(n16540), .B(n14035), .ZN(
        n14054) );
  NOR2_X1 U15622 ( .A1(n12069), .A2(n14038), .ZN(n16552) );
  AOI22_X1 U15623 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14045) );
  NAND2_X1 U15624 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14040) );
  NAND2_X1 U15625 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n14039) );
  AND3_X1 U15626 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(n14044) );
  AOI22_X1 U15627 ( .A1(n11163), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U15628 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14042) );
  NAND4_X1 U15629 ( .A1(n14045), .A2(n14044), .A3(n14043), .A4(n14042), .ZN(
        n14053) );
  AOI22_X1 U15630 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U15631 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14084), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U15632 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14049) );
  NAND2_X1 U15633 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14047) );
  NAND2_X1 U15634 ( .A1(n14080), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14046) );
  AND3_X1 U15635 ( .A1(n14047), .A2(n14046), .A3(n14087), .ZN(n14048) );
  NAND4_X1 U15636 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14052) );
  AND2_X1 U15637 ( .A1(n14053), .A2(n14052), .ZN(n16541) );
  NAND2_X1 U15638 ( .A1(n14055), .A2(n14054), .ZN(n16549) );
  AOI22_X1 U15639 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11162), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U15640 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U15641 ( .A1(n14057), .A2(n14056), .ZN(n14069) );
  AOI21_X1 U15642 ( .B1(n14084), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n14087), .ZN(n14059) );
  AOI22_X1 U15643 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14058) );
  OAI211_X1 U15644 ( .C1(n11201), .C2(n15670), .A(n14059), .B(n14058), .ZN(
        n14068) );
  AOI22_X1 U15645 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11163), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U15646 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14061) );
  NAND2_X1 U15647 ( .A1(n14062), .A2(n14061), .ZN(n14067) );
  AOI22_X1 U15648 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14065) );
  NAND2_X1 U15649 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14064) );
  NAND2_X1 U15650 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14063) );
  NAND4_X1 U15651 ( .A1(n14065), .A2(n14064), .A3(n14063), .A4(n14087), .ZN(
        n14066) );
  OAI22_X1 U15652 ( .A1(n14069), .A2(n14068), .B1(n14067), .B2(n14066), .ZN(
        n14070) );
  NAND2_X1 U15653 ( .A1(n12069), .A2(n16541), .ZN(n14072) );
  NOR2_X1 U15654 ( .A1(n16540), .A2(n14072), .ZN(n16534) );
  NAND2_X1 U15655 ( .A1(n11250), .A2(n14073), .ZN(n14095) );
  AOI22_X1 U15656 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11162), .B1(
        n14079), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U15657 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14074) );
  NAND2_X1 U15658 ( .A1(n14075), .A2(n14074), .ZN(n14092) );
  INV_X1 U15659 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19532) );
  AOI21_X1 U15660 ( .B1(n14084), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n14087), .ZN(n14077) );
  AOI22_X1 U15661 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14076) );
  OAI211_X1 U15662 ( .C1(n13944), .C2(n19532), .A(n14077), .B(n14076), .ZN(
        n14091) );
  AOI22_X1 U15663 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U15664 ( .A1(n11163), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14080), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U15665 ( .A1(n14082), .A2(n14081), .ZN(n14090) );
  AOI22_X1 U15666 ( .A1(n14083), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11204), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U15667 ( .A1(n12083), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14086) );
  NAND2_X1 U15668 ( .A1(n14084), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14085) );
  NAND4_X1 U15669 ( .A1(n14088), .A2(n14087), .A3(n14086), .A4(n14085), .ZN(
        n14089) );
  OAI22_X1 U15670 ( .A1(n14092), .A2(n14091), .B1(n14090), .B2(n14089), .ZN(
        n14093) );
  INV_X1 U15671 ( .A(n14093), .ZN(n14094) );
  NOR2_X1 U15672 ( .A1(n14096), .A2(n11893), .ZN(n14097) );
  OR2_X1 U15673 ( .A1(n14118), .A2(n14097), .ZN(n14115) );
  AND2_X1 U15674 ( .A1(n14117), .A2(n12069), .ZN(n14100) );
  OAI21_X1 U15675 ( .B1(n14100), .B2(n14099), .A(n14098), .ZN(n14111) );
  NAND2_X1 U15676 ( .A1(n14102), .A2(n14101), .ZN(n14107) );
  INV_X1 U15677 ( .A(n14103), .ZN(n14104) );
  OAI211_X1 U15678 ( .C1(n12069), .C2(n14105), .A(n11861), .B(n14104), .ZN(
        n14106) );
  OAI211_X1 U15679 ( .C1(n11855), .C2(n14108), .A(n14107), .B(n14106), .ZN(
        n14110) );
  AOI21_X1 U15680 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14112) );
  AOI21_X1 U15681 ( .B1(n14113), .B2(n11893), .A(n14112), .ZN(n14114) );
  NOR2_X1 U15682 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  MUX2_X1 U15683 ( .A(n18987), .B(n14116), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14311) );
  INV_X1 U15684 ( .A(n14117), .ZN(n14300) );
  AND2_X1 U15685 ( .A1(n14118), .A2(n14300), .ZN(n14119) );
  INV_X1 U15686 ( .A(n14912), .ZN(n14121) );
  NAND2_X1 U15687 ( .A1(n14120), .A2(n11656), .ZN(n14363) );
  INV_X1 U15688 ( .A(n14363), .ZN(n14766) );
  NAND2_X1 U15689 ( .A1(n14121), .A2(n14766), .ZN(n14738) );
  NAND2_X1 U15690 ( .A1(n14738), .A2(n11240), .ZN(n14122) );
  NAND2_X1 U15691 ( .A1(n16571), .A2(n15617), .ZN(n16606) );
  OAI21_X1 U15692 ( .B1(n15961), .B2(n16606), .A(n14123), .ZN(P2_U2857) );
  NOR4_X1 U15693 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14127) );
  NOR4_X1 U15694 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14126) );
  NOR4_X1 U15695 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14125) );
  NOR4_X1 U15696 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14124) );
  AND4_X1 U15697 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14132) );
  NOR4_X1 U15698 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n14130) );
  NOR4_X1 U15699 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14129) );
  NOR4_X1 U15700 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14128) );
  INV_X1 U15701 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20213) );
  AND4_X1 U15702 ( .A1(n14130), .A2(n14129), .A3(n14128), .A4(n20213), .ZN(
        n14131) );
  NAND2_X1 U15703 ( .A1(n14132), .A2(n14131), .ZN(n14133) );
  AND2_X2 U15704 ( .A1(n14133), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15813)
         );
  INV_X1 U15705 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20458) );
  INV_X1 U15706 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22750) );
  NOR4_X1 U15707 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20458), .A4(n22750), .ZN(n14135) );
  NOR4_X1 U15708 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14134) );
  NAND3_X1 U15709 ( .A1(n15813), .A2(n14135), .A3(n14134), .ZN(U214) );
  NOR4_X1 U15710 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14139) );
  NOR4_X1 U15711 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14138) );
  NOR4_X1 U15712 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14137) );
  NOR4_X1 U15713 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14136) );
  NAND4_X1 U15714 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14144) );
  NOR4_X1 U15715 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14142) );
  NOR4_X1 U15716 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14141) );
  NOR4_X1 U15717 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14140) );
  INV_X1 U15718 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20120) );
  NAND4_X1 U15719 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n20120), .ZN(
        n14143) );
  OAI21_X1 U15720 ( .B1(n14144), .B2(n14143), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14211) );
  NOR2_X1 U15721 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14146) );
  NOR4_X1 U15722 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14145) );
  NAND4_X1 U15723 ( .A1(n14146), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14145), .ZN(n14147) );
  OR2_X1 U15724 ( .A1(n14211), .A2(n14147), .ZN(n20401) );
  OR2_X1 U15725 ( .A1(n20401), .A2(n20446), .ZN(U212) );
  NOR2_X1 U15726 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14147), .ZN(n19419)
         );
  INV_X1 U15727 ( .A(n18631), .ZN(n19054) );
  OR2_X1 U15728 ( .A1(n14148), .A2(n19054), .ZN(n14298) );
  NOR2_X1 U15729 ( .A1(n14759), .A2(n14298), .ZN(n18653) );
  INV_X1 U15730 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n17505) );
  INV_X1 U15731 ( .A(n14152), .ZN(n14150) );
  OAI211_X1 U15732 ( .C1(n18653), .C2(n17505), .A(n14150), .B(n14149), .ZN(
        P2_U2814) );
  OR3_X1 U15733 ( .A1(n14152), .A2(n17427), .A3(P2_READREQUEST_REG_SCAN_IN), 
        .ZN(n14153) );
  OAI22_X1 U15734 ( .A1(n14151), .A2(n18628), .B1(n14153), .B2(n18653), .ZN(
        n14154) );
  INV_X1 U15735 ( .A(n14154), .ZN(P2_U3612) );
  INV_X1 U15736 ( .A(n14221), .ZN(n14226) );
  INV_X1 U15737 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14156) );
  INV_X1 U15738 ( .A(n14297), .ZN(n14222) );
  INV_X1 U15739 ( .A(n14211), .ZN(n15619) );
  AOI22_X1 U15740 ( .A1(n15619), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15622), .ZN(n19527) );
  NOR2_X1 U15741 ( .A1(n14226), .A2(n19527), .ZN(n14189) );
  AOI21_X1 U15742 ( .B1(n14222), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14189), .ZN(
        n14155) );
  OAI21_X1 U15743 ( .B1(n14227), .B2(n14156), .A(n14155), .ZN(P2_U2959) );
  INV_X1 U15744 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14158) );
  OAI22_X1 U15745 ( .A1(n14211), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15619), .ZN(n19724) );
  NOR2_X1 U15746 ( .A1(n14226), .A2(n19724), .ZN(n14186) );
  AOI21_X1 U15747 ( .B1(n14222), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14186), .ZN(
        n14157) );
  OAI21_X1 U15748 ( .B1(n14227), .B2(n14158), .A(n14157), .ZN(P2_U2958) );
  INV_X1 U15749 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U15750 ( .A1(n15619), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15622), .ZN(n20006) );
  NOR2_X1 U15751 ( .A1(n14226), .A2(n20006), .ZN(n14163) );
  AOI21_X1 U15752 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n14222), .A(n14163), .ZN(
        n14159) );
  OAI21_X1 U15753 ( .B1(n14227), .B2(n14160), .A(n14159), .ZN(P2_U2967) );
  INV_X1 U15754 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14162) );
  OAI22_X1 U15755 ( .A1(n15622), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15619), .ZN(n19827) );
  NOR2_X1 U15756 ( .A1(n14226), .A2(n19827), .ZN(n14180) );
  AOI21_X1 U15757 ( .B1(n14222), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14180), .ZN(
        n14161) );
  OAI21_X1 U15758 ( .B1(n14227), .B2(n14162), .A(n14161), .ZN(P2_U2956) );
  INV_X1 U15759 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14165) );
  AOI21_X1 U15760 ( .B1(n14222), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14163), .ZN(
        n14164) );
  OAI21_X1 U15761 ( .B1(n14227), .B2(n14165), .A(n14164), .ZN(P2_U2952) );
  INV_X1 U15762 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U15763 ( .A1(n15619), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14211), .ZN(n16663) );
  NOR2_X1 U15764 ( .A1(n14226), .A2(n16663), .ZN(n14170) );
  AOI21_X1 U15765 ( .B1(P2_EAX_REG_8__SCAN_IN), .B2(n14222), .A(n14170), .ZN(
        n14166) );
  OAI21_X1 U15766 ( .B1(n14227), .B2(n14167), .A(n14166), .ZN(P2_U2975) );
  INV_X1 U15767 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U15768 ( .A1(n15619), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14211), .ZN(n19772) );
  NOR2_X1 U15769 ( .A1(n14226), .A2(n19772), .ZN(n14177) );
  AOI21_X1 U15770 ( .B1(n14222), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14177), .ZN(
        n14168) );
  OAI21_X1 U15771 ( .B1(n14227), .B2(n14169), .A(n14168), .ZN(P2_U2972) );
  INV_X1 U15772 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14172) );
  AOI21_X1 U15773 ( .B1(n14222), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14170), .ZN(
        n14171) );
  OAI21_X1 U15774 ( .B1(n14227), .B2(n14172), .A(n14171), .ZN(P2_U2960) );
  INV_X1 U15775 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U15776 ( .A1(n15619), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15622), .ZN(n16693) );
  NOR2_X1 U15777 ( .A1(n14226), .A2(n16693), .ZN(n14183) );
  AOI21_X1 U15778 ( .B1(n14222), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14183), .ZN(
        n14173) );
  OAI21_X1 U15779 ( .B1(n14227), .B2(n14174), .A(n14173), .ZN(P2_U2955) );
  INV_X1 U15780 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14176) );
  OAI22_X1 U15781 ( .A1(n14211), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15619), .ZN(n19918) );
  NOR2_X1 U15782 ( .A1(n14226), .A2(n19918), .ZN(n14192) );
  AOI21_X1 U15783 ( .B1(n14222), .B2(P2_EAX_REG_2__SCAN_IN), .A(n14192), .ZN(
        n14175) );
  OAI21_X1 U15784 ( .B1(n14227), .B2(n14176), .A(n14175), .ZN(P2_U2969) );
  INV_X1 U15785 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14179) );
  AOI21_X1 U15786 ( .B1(n14222), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14177), .ZN(
        n14178) );
  OAI21_X1 U15787 ( .B1(n14227), .B2(n14179), .A(n14178), .ZN(P2_U2957) );
  INV_X1 U15788 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14182) );
  AOI21_X1 U15789 ( .B1(n14222), .B2(P2_EAX_REG_4__SCAN_IN), .A(n14180), .ZN(
        n14181) );
  OAI21_X1 U15790 ( .B1(n14227), .B2(n14182), .A(n14181), .ZN(P2_U2971) );
  INV_X1 U15791 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14185) );
  AOI21_X1 U15792 ( .B1(n14222), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14183), .ZN(
        n14184) );
  OAI21_X1 U15793 ( .B1(n14227), .B2(n14185), .A(n14184), .ZN(P2_U2970) );
  INV_X1 U15794 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14188) );
  AOI21_X1 U15795 ( .B1(n14222), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14186), .ZN(
        n14187) );
  OAI21_X1 U15796 ( .B1(n14227), .B2(n14188), .A(n14187), .ZN(P2_U2973) );
  INV_X1 U15797 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14191) );
  AOI21_X1 U15798 ( .B1(n14222), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14189), .ZN(
        n14190) );
  OAI21_X1 U15799 ( .B1(n14227), .B2(n14191), .A(n14190), .ZN(P2_U2974) );
  INV_X1 U15800 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14194) );
  AOI21_X1 U15801 ( .B1(n14222), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14192), .ZN(
        n14193) );
  OAI21_X1 U15802 ( .B1(n14227), .B2(n14194), .A(n14193), .ZN(P2_U2954) );
  INV_X1 U15803 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U15804 ( .A1(n15619), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15622), .ZN(n19963) );
  NOR2_X1 U15805 ( .A1(n14226), .A2(n19963), .ZN(n14197) );
  AOI21_X1 U15806 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14222), .A(n14197), .ZN(
        n14195) );
  OAI21_X1 U15807 ( .B1(n14227), .B2(n14196), .A(n14195), .ZN(P2_U2968) );
  INV_X1 U15808 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14199) );
  AOI21_X1 U15809 ( .B1(n14222), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14197), .ZN(
        n14198) );
  OAI21_X1 U15810 ( .B1(n14227), .B2(n14199), .A(n14198), .ZN(P2_U2953) );
  INV_X1 U15811 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U15812 ( .A1(n15619), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n14211), .ZN(n16620) );
  INV_X1 U15813 ( .A(n16620), .ZN(n14200) );
  NAND2_X1 U15814 ( .A1(n14221), .A2(n14200), .ZN(n14228) );
  NAND2_X1 U15815 ( .A1(n14222), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n14201) );
  OAI211_X1 U15816 ( .C1(n14227), .C2(n14202), .A(n14228), .B(n14201), .ZN(
        P2_U2979) );
  INV_X1 U15817 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n14207) );
  INV_X1 U15818 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14203) );
  OR2_X1 U15819 ( .A1(n15622), .A2(n14203), .ZN(n14205) );
  NAND2_X1 U15820 ( .A1(n14211), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U15821 ( .A1(n14205), .A2(n14204), .ZN(n16642) );
  NAND2_X1 U15822 ( .A1(n14221), .A2(n16642), .ZN(n14230) );
  NAND2_X1 U15823 ( .A1(n14222), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n14206) );
  OAI211_X1 U15824 ( .C1(n14227), .C2(n14207), .A(n14230), .B(n14206), .ZN(
        P2_U2977) );
  INV_X1 U15825 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n14210) );
  AOI22_X1 U15826 ( .A1(n15619), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n15622), .ZN(n15955) );
  INV_X1 U15827 ( .A(n15955), .ZN(n14208) );
  NAND2_X1 U15828 ( .A1(n14221), .A2(n14208), .ZN(n14232) );
  NAND2_X1 U15829 ( .A1(n14222), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n14209) );
  OAI211_X1 U15830 ( .C1(n14227), .C2(n14210), .A(n14232), .B(n14209), .ZN(
        P2_U2981) );
  INV_X1 U15831 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14216) );
  INV_X1 U15832 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20421) );
  OR2_X1 U15833 ( .A1(n14211), .A2(n20421), .ZN(n14213) );
  NAND2_X1 U15834 ( .A1(n14211), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14212) );
  AND2_X1 U15835 ( .A1(n14213), .A2(n14212), .ZN(n16651) );
  INV_X1 U15836 ( .A(n16651), .ZN(n14214) );
  NAND2_X1 U15837 ( .A1(n14221), .A2(n14214), .ZN(n14236) );
  NAND2_X1 U15838 ( .A1(n14222), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n14215) );
  OAI211_X1 U15839 ( .C1(n14227), .C2(n14216), .A(n14236), .B(n14215), .ZN(
        P2_U2976) );
  INV_X1 U15840 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14219) );
  AOI22_X1 U15841 ( .A1(n15619), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15622), .ZN(n16631) );
  INV_X1 U15842 ( .A(n16631), .ZN(n14217) );
  NAND2_X1 U15843 ( .A1(n14221), .A2(n14217), .ZN(n14239) );
  NAND2_X1 U15844 ( .A1(n14222), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14218) );
  OAI211_X1 U15845 ( .C1(n14227), .C2(n14219), .A(n14239), .B(n14218), .ZN(
        P2_U2978) );
  INV_X1 U15846 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U15847 ( .A1(n15619), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15622), .ZN(n16612) );
  INV_X1 U15848 ( .A(n16612), .ZN(n14220) );
  NAND2_X1 U15849 ( .A1(n14221), .A2(n14220), .ZN(n14234) );
  NAND2_X1 U15850 ( .A1(n14222), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14223) );
  OAI211_X1 U15851 ( .C1(n14227), .C2(n14224), .A(n14234), .B(n14223), .ZN(
        P2_U2980) );
  AOI22_X1 U15852 ( .A1(n15619), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15622), .ZN(n15106) );
  INV_X1 U15853 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17545) );
  INV_X1 U15854 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14225) );
  OAI222_X1 U15855 ( .A1(n14226), .A2(n15106), .B1(n14297), .B2(n17545), .C1(
        n14227), .C2(n14225), .ZN(P2_U2982) );
  INV_X1 U15856 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n16619) );
  INV_X1 U15857 ( .A(n14227), .ZN(n14238) );
  NAND2_X1 U15858 ( .A1(n14238), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14229) );
  OAI211_X1 U15859 ( .C1(n14297), .C2(n16619), .A(n14229), .B(n14228), .ZN(
        P2_U2964) );
  INV_X1 U15860 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U15861 ( .A1(n14238), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14231) );
  OAI211_X1 U15862 ( .C1(n14297), .C2(n14512), .A(n14231), .B(n14230), .ZN(
        P2_U2962) );
  INV_X1 U15863 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n15954) );
  NAND2_X1 U15864 ( .A1(n14238), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14233) );
  OAI211_X1 U15865 ( .C1(n14297), .C2(n15954), .A(n14233), .B(n14232), .ZN(
        P2_U2966) );
  INV_X1 U15866 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16611) );
  NAND2_X1 U15867 ( .A1(n14238), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14235) );
  OAI211_X1 U15868 ( .C1(n14297), .C2(n16611), .A(n14235), .B(n14234), .ZN(
        P2_U2965) );
  INV_X1 U15869 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U15870 ( .A1(n14238), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14237) );
  OAI211_X1 U15871 ( .C1(n14297), .C2(n14504), .A(n14237), .B(n14236), .ZN(
        P2_U2961) );
  INV_X1 U15872 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n16630) );
  NAND2_X1 U15873 ( .A1(n14238), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14240) );
  OAI211_X1 U15874 ( .C1(n14297), .C2(n16630), .A(n14240), .B(n14239), .ZN(
        P2_U2963) );
  INV_X1 U15875 ( .A(n14244), .ZN(n14241) );
  AOI222_X1 U15876 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14244), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14243), .C1(n14242), .C2(
        n14241), .ZN(n17167) );
  INV_X1 U15877 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14249) );
  NOR2_X1 U15878 ( .A1(n17452), .A2(n14249), .ZN(n14248) );
  OAI21_X1 U15879 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14246), .A(
        n14245), .ZN(n17165) );
  NAND2_X1 U15880 ( .A1(n11167), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n17164) );
  OAI21_X1 U15881 ( .B1(n17446), .B2(n17165), .A(n17164), .ZN(n14247) );
  AOI211_X1 U15882 ( .C1(n17443), .C2(n14249), .A(n14248), .B(n14247), .ZN(
        n14251) );
  NAND2_X1 U15883 ( .A1(n17457), .A2(n18648), .ZN(n14250) );
  OAI211_X1 U15884 ( .C1(n17167), .C2(n17445), .A(n14251), .B(n14250), .ZN(
        P2_U3013) );
  NAND2_X1 U15885 ( .A1(n12069), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14252) );
  AND4_X1 U15886 ( .A1(n13761), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14252), 
        .A4(n19593), .ZN(n14253) );
  MUX2_X1 U15887 ( .A(n11912), .B(n18992), .S(n16571), .Z(n14254) );
  OAI21_X1 U15888 ( .B1(n16606), .B2(n17477), .A(n14254), .ZN(P2_U2887) );
  NAND2_X1 U15889 ( .A1(n14471), .A2(n22236), .ZN(n14255) );
  OR2_X1 U15890 ( .A1(n14256), .A2(n14255), .ZN(n14276) );
  NOR2_X1 U15891 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  AND2_X1 U15892 ( .A1(n14260), .A2(n14259), .ZN(n14261) );
  OR2_X1 U15893 ( .A1(n14262), .A2(n14261), .ZN(n15818) );
  NOR2_X1 U15894 ( .A1(n14276), .A2(n15818), .ZN(n16040) );
  NOR2_X1 U15895 ( .A1(n16040), .A2(n15895), .ZN(n14263) );
  AOI21_X1 U15896 ( .B1(n15830), .B2(n14881), .A(n14263), .ZN(n20396) );
  INV_X1 U15897 ( .A(n14886), .ZN(n14264) );
  NOR2_X1 U15898 ( .A1(n14264), .A2(n17412), .ZN(n16515) );
  INV_X1 U15899 ( .A(n16515), .ZN(n14266) );
  OR2_X1 U15900 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n14265), .ZN(n14882) );
  NAND2_X1 U15901 ( .A1(n14266), .A2(n14882), .ZN(n14267) );
  NAND2_X1 U15902 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21697) );
  NAND2_X1 U15903 ( .A1(n14267), .A2(n21697), .ZN(n21701) );
  NAND2_X1 U15904 ( .A1(n20396), .A2(n21701), .ZN(n17403) );
  INV_X1 U15905 ( .A(n22135), .ZN(n15833) );
  AND2_X1 U15906 ( .A1(n17403), .A2(n15833), .ZN(n22114) );
  INV_X1 U15907 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n14283) );
  NAND2_X1 U15908 ( .A1(n15841), .A2(n14271), .ZN(n14269) );
  NOR2_X1 U15909 ( .A1(n14269), .A2(n16505), .ZN(n15905) );
  INV_X1 U15910 ( .A(n15905), .ZN(n14279) );
  NAND2_X1 U15911 ( .A1(n14271), .A2(n15821), .ZN(n15898) );
  NAND2_X1 U15912 ( .A1(n14270), .A2(n22528), .ZN(n14274) );
  NAND2_X1 U15913 ( .A1(n14271), .A2(n14307), .ZN(n14272) );
  NOR2_X1 U15914 ( .A1(n14272), .A2(n16505), .ZN(n14452) );
  OR2_X1 U15915 ( .A1(n17399), .A2(n14452), .ZN(n15839) );
  INV_X1 U15916 ( .A(n15839), .ZN(n14273) );
  OAI21_X1 U15917 ( .B1(n15898), .B2(n14274), .A(n14273), .ZN(n14275) );
  NAND2_X1 U15918 ( .A1(n15830), .A2(n14275), .ZN(n14278) );
  INV_X1 U15919 ( .A(n14276), .ZN(n14457) );
  NAND2_X1 U15920 ( .A1(n14457), .A2(n15818), .ZN(n14277) );
  OAI211_X1 U15921 ( .C1(n15830), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n14280) );
  NAND2_X1 U15922 ( .A1(n14280), .A2(n14636), .ZN(n17400) );
  INV_X1 U15923 ( .A(n17400), .ZN(n14281) );
  NAND2_X1 U15924 ( .A1(n22114), .A2(n14281), .ZN(n14282) );
  OAI21_X1 U15925 ( .B1(n22114), .B2(n14283), .A(n14282), .ZN(P1_U3484) );
  INV_X1 U15926 ( .A(n17457), .ZN(n17471) );
  INV_X1 U15927 ( .A(n17445), .ZN(n17462) );
  XNOR2_X1 U15928 ( .A(n14284), .B(n18993), .ZN(n18990) );
  NAND2_X1 U15929 ( .A1(n11167), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18995) );
  INV_X1 U15930 ( .A(n18995), .ZN(n14289) );
  NAND2_X1 U15931 ( .A1(n14285), .A2(n18993), .ZN(n14286) );
  NAND2_X1 U15932 ( .A1(n14287), .A2(n14286), .ZN(n18996) );
  NOR2_X1 U15933 ( .A1(n17446), .A2(n18996), .ZN(n14288) );
  AOI211_X1 U15934 ( .C1(n17462), .C2(n18990), .A(n14289), .B(n14288), .ZN(
        n14292) );
  INV_X1 U15935 ( .A(n17452), .ZN(n17461) );
  OAI21_X1 U15936 ( .B1(n17461), .B2(n14290), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14291) );
  OAI211_X1 U15937 ( .C1(n17471), .C2(n18992), .A(n14292), .B(n14291), .ZN(
        P2_U3014) );
  INV_X1 U15938 ( .A(n19551), .ZN(n17488) );
  MUX2_X1 U15939 ( .A(n12430), .B(n14295), .S(n16571), .Z(n14296) );
  OAI21_X1 U15940 ( .B1(n17488), .B2(n16606), .A(n14296), .ZN(P2_U2886) );
  INV_X1 U15941 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15721) );
  NAND2_X1 U15942 ( .A1(n14912), .A2(n12069), .ZN(n14731) );
  OAI21_X1 U15943 ( .B1(n14731), .B2(n14298), .A(n14297), .ZN(n14299) );
  NAND2_X1 U15944 ( .A1(n17509), .A2(n14300), .ZN(n14518) );
  NOR2_X1 U15945 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14914), .ZN(n17530) );
  AOI22_X1 U15946 ( .A1(n17530), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14301) );
  OAI21_X1 U15947 ( .B1(n15721), .B2(n14518), .A(n14301), .ZN(P2_U2934) );
  INV_X1 U15948 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14303) );
  AOI22_X1 U15949 ( .A1(n17530), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14302) );
  OAI21_X1 U15950 ( .B1(n14303), .B2(n14518), .A(n14302), .ZN(P2_U2933) );
  NAND2_X1 U15951 ( .A1(n22292), .A2(n22121), .ZN(n20399) );
  INV_X1 U15952 ( .A(n20399), .ZN(n14304) );
  NOR2_X1 U15953 ( .A1(n14304), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14309)
         );
  NAND2_X1 U15954 ( .A1(n16040), .A2(n22386), .ZN(n14453) );
  NAND2_X1 U15955 ( .A1(n14457), .A2(n14467), .ZN(n17375) );
  NOR2_X1 U15956 ( .A1(n17375), .A2(n22135), .ZN(n14306) );
  NAND2_X1 U15957 ( .A1(n15824), .A2(n14306), .ZN(n14868) );
  OAI21_X1 U15958 ( .B1(n16057), .B2(n14307), .A(n21696), .ZN(n14308) );
  OAI21_X1 U15959 ( .B1(n14309), .B2(n21696), .A(n14308), .ZN(P1_U3487) );
  INV_X1 U15960 ( .A(n14310), .ZN(n14771) );
  INV_X1 U15961 ( .A(n11877), .ZN(n14343) );
  NAND2_X1 U15962 ( .A1(n14771), .A2(n14343), .ZN(n14338) );
  OAI21_X1 U15963 ( .B1(n14311), .B2(n11854), .A(n11888), .ZN(n14312) );
  INV_X1 U15964 ( .A(n14312), .ZN(n14313) );
  NAND2_X1 U15965 ( .A1(n14313), .A2(n14731), .ZN(n14337) );
  NAND2_X1 U15966 ( .A1(n14314), .A2(n12069), .ZN(n14315) );
  NOR2_X1 U15967 ( .A1(n19043), .A2(n14315), .ZN(n14335) );
  MUX2_X1 U15968 ( .A(n14316), .B(n11877), .S(n12609), .Z(n14317) );
  INV_X1 U15969 ( .A(n22174), .ZN(n19035) );
  OR2_X1 U15970 ( .A1(n14317), .A2(n19035), .ZN(n14333) );
  NAND2_X1 U15971 ( .A1(n14804), .A2(n14771), .ZN(n14319) );
  OR2_X1 U15972 ( .A1(n14759), .A2(n14319), .ZN(n14331) );
  NAND2_X1 U15973 ( .A1(n14320), .A2(n11877), .ZN(n14321) );
  NAND2_X1 U15974 ( .A1(n14148), .A2(n14321), .ZN(n14330) );
  NAND2_X1 U15975 ( .A1(n12609), .A2(n11888), .ZN(n14358) );
  AOI21_X1 U15976 ( .B1(n14358), .B2(n11861), .A(n19528), .ZN(n14323) );
  OAI211_X1 U15977 ( .C1(n14323), .C2(n14343), .A(n14322), .B(n11923), .ZN(
        n14324) );
  INV_X1 U15978 ( .A(n14324), .ZN(n14329) );
  INV_X1 U15979 ( .A(n14325), .ZN(n14326) );
  NAND2_X1 U15980 ( .A1(n14326), .A2(n15617), .ZN(n14328) );
  NAND2_X1 U15981 ( .A1(n14328), .A2(n14327), .ZN(n14351) );
  AND3_X1 U15982 ( .A1(n14330), .A2(n14329), .A3(n14351), .ZN(n14360) );
  AND2_X1 U15983 ( .A1(n14331), .A2(n14360), .ZN(n14735) );
  OAI211_X1 U15984 ( .C1(n14759), .C2(n14333), .A(n14735), .B(n14332), .ZN(
        n14334) );
  NOR2_X1 U15985 ( .A1(n14335), .A2(n14334), .ZN(n14336) );
  OAI211_X1 U15986 ( .C1(n14731), .C2(n14338), .A(n14337), .B(n14336), .ZN(
        n14339) );
  NAND2_X1 U15987 ( .A1(n14378), .A2(n14765), .ZN(n17166) );
  XNOR2_X1 U15988 ( .A(n14341), .B(n14340), .ZN(n14393) );
  MUX2_X1 U15989 ( .A(n14342), .B(n14343), .S(n11854), .Z(n14348) );
  INV_X1 U15990 ( .A(n14151), .ZN(n18624) );
  OAI21_X1 U15991 ( .B1(n11852), .B2(n11888), .A(n18624), .ZN(n14346) );
  NOR2_X1 U15992 ( .A1(n11923), .A2(n11855), .ZN(n14345) );
  NAND2_X1 U15993 ( .A1(n14345), .A2(n14344), .ZN(n14394) );
  NAND2_X1 U15994 ( .A1(n14346), .A2(n14394), .ZN(n14347) );
  NOR2_X1 U15995 ( .A1(n14348), .A2(n14347), .ZN(n14356) );
  NAND3_X1 U15996 ( .A1(n11910), .A2(n11852), .A3(n14349), .ZN(n14355) );
  NAND2_X1 U15997 ( .A1(n14350), .A2(n12069), .ZN(n14782) );
  NAND2_X1 U15998 ( .A1(n14782), .A2(n14351), .ZN(n14353) );
  NAND2_X1 U15999 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  AND3_X1 U16000 ( .A1(n14356), .A2(n14355), .A3(n14354), .ZN(n14741) );
  NAND2_X1 U16001 ( .A1(n14741), .A2(n11240), .ZN(n14357) );
  NAND2_X1 U16002 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17171) );
  NAND2_X1 U16003 ( .A1(n14379), .A2(n17171), .ZN(n19026) );
  NAND3_X1 U16004 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15751) );
  AND2_X1 U16005 ( .A1(n19026), .A2(n15751), .ZN(n14362) );
  AND2_X1 U16006 ( .A1(n11167), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14384) );
  INV_X1 U16007 ( .A(n14358), .ZN(n14359) );
  INV_X1 U16008 ( .A(n17047), .ZN(n15072) );
  NOR2_X1 U16009 ( .A1(n15072), .A2(n14362), .ZN(n14361) );
  AOI211_X1 U16010 ( .C1(n17048), .C2(n14362), .A(n14384), .B(n14361), .ZN(
        n14383) );
  NAND2_X1 U16011 ( .A1(n12422), .A2(n12069), .ZN(n14364) );
  NAND2_X1 U16012 ( .A1(n14364), .A2(n14363), .ZN(n14365) );
  INV_X1 U16013 ( .A(n19003), .ZN(n19020) );
  INV_X1 U16014 ( .A(n14366), .ZN(n14367) );
  XNOR2_X1 U16015 ( .A(n14368), .B(n14367), .ZN(n15541) );
  OAI21_X1 U16016 ( .B1(n14371), .B2(n14370), .A(n14369), .ZN(n14388) );
  OAI22_X1 U16017 ( .A1(n19020), .A2(n15541), .B1(n14388), .B2(n19015), .ZN(
        n14381) );
  INV_X1 U16018 ( .A(n14378), .ZN(n14372) );
  NAND2_X1 U16019 ( .A1(n14372), .A2(n18830), .ZN(n18994) );
  NAND2_X1 U16020 ( .A1(n14374), .A2(n12609), .ZN(n14376) );
  NAND2_X1 U16021 ( .A1(n14376), .A2(n11198), .ZN(n14377) );
  NAND2_X1 U16022 ( .A1(n14378), .A2(n14377), .ZN(n18991) );
  OAI22_X1 U16023 ( .A1(n18994), .A2(n14379), .B1(n14730), .B2(n18991), .ZN(
        n14380) );
  NOR2_X1 U16024 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  OAI211_X1 U16025 ( .C1(n17166), .C2(n14393), .A(n14383), .B(n14382), .ZN(
        P2_U3044) );
  INV_X1 U16026 ( .A(n15539), .ZN(n14391) );
  INV_X1 U16027 ( .A(n14384), .ZN(n14387) );
  INV_X1 U16028 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14385) );
  OR2_X1 U16029 ( .A1(n17452), .A2(n14385), .ZN(n14386) );
  OAI211_X1 U16030 ( .C1(n14388), .C2(n17446), .A(n14387), .B(n14386), .ZN(
        n14390) );
  NOR2_X1 U16031 ( .A1(n17471), .A2(n14730), .ZN(n14389) );
  AOI211_X1 U16032 ( .C1(n17443), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        n14392) );
  OAI21_X1 U16033 ( .B1(n17445), .B2(n14393), .A(n14392), .ZN(P2_U3012) );
  NAND2_X1 U16034 ( .A1(n14912), .A2(n14758), .ZN(n14736) );
  NAND2_X1 U16035 ( .A1(n14736), .A2(n14394), .ZN(n14395) );
  NAND2_X1 U16036 ( .A1(n14395), .A2(n18631), .ZN(n14397) );
  NAND2_X1 U16037 ( .A1(n14151), .A2(n22174), .ZN(n14770) );
  OR2_X1 U16038 ( .A1(n18628), .A2(n14770), .ZN(n14396) );
  NAND2_X1 U16039 ( .A1(n19770), .A2(n14398), .ZN(n19773) );
  NOR2_X2 U16040 ( .A1(n19905), .A2(n15617), .ZN(n19822) );
  XNOR2_X1 U16041 ( .A(n14400), .B(n14399), .ZN(n18635) );
  INV_X1 U16042 ( .A(n18635), .ZN(n18989) );
  AOI22_X1 U16043 ( .A1(n19822), .A2(n18989), .B1(n19905), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U16044 ( .A1(n19770), .A2(n14401), .ZN(n19911) );
  INV_X1 U16045 ( .A(n19911), .ZN(n19821) );
  XNOR2_X1 U16046 ( .A(n19550), .B(n18635), .ZN(n14402) );
  NAND2_X1 U16047 ( .A1(n19821), .A2(n14402), .ZN(n14403) );
  OAI211_X1 U16048 ( .C1(n20006), .C2(n19773), .A(n14404), .B(n14403), .ZN(
        P2_U2919) );
  OR2_X1 U16049 ( .A1(n14406), .A2(n14405), .ZN(n14408) );
  NAND2_X1 U16050 ( .A1(n14408), .A2(n14407), .ZN(n18646) );
  XNOR2_X1 U16051 ( .A(n19551), .B(n18646), .ZN(n14410) );
  NOR2_X1 U16052 ( .A1(n17477), .A2(n18635), .ZN(n14409) );
  NOR2_X1 U16053 ( .A1(n14410), .A2(n14409), .ZN(n14619) );
  AOI21_X1 U16054 ( .B1(n14410), .B2(n14409), .A(n14619), .ZN(n14414) );
  AOI22_X1 U16055 ( .A1(n19822), .A2(n18646), .B1(n19905), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14413) );
  INV_X1 U16056 ( .A(n19773), .ZN(n14705) );
  INV_X1 U16057 ( .A(n19963), .ZN(n14411) );
  NAND2_X1 U16058 ( .A1(n14705), .A2(n14411), .ZN(n14412) );
  OAI211_X1 U16059 ( .C1(n14414), .C2(n19911), .A(n14413), .B(n14412), .ZN(
        P2_U2918) );
  INV_X1 U16060 ( .A(n14416), .ZN(n14417) );
  MUX2_X1 U16061 ( .A(n12429), .B(n14730), .S(n16571), .Z(n14418) );
  OAI21_X1 U16062 ( .B1(n17481), .B2(n16606), .A(n14418), .ZN(P2_U2885) );
  INV_X1 U16063 ( .A(n21697), .ZN(n22165) );
  OR2_X1 U16064 ( .A1(n22386), .A2(n22165), .ZN(n14419) );
  OR2_X1 U16065 ( .A1(n16043), .A2(n14419), .ZN(n14580) );
  INV_X1 U16066 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20413) );
  INV_X1 U16067 ( .A(n15813), .ZN(n15812) );
  NOR2_X1 U16068 ( .A1(n15813), .A2(DATAI_5_), .ZN(n14420) );
  AOI21_X1 U16069 ( .B1(n15813), .B2(n20413), .A(n14420), .ZN(n22527) );
  NAND2_X1 U16070 ( .A1(n14521), .A2(n22527), .ZN(n14553) );
  NOR2_X1 U16071 ( .A1(n17412), .A2(n21697), .ZN(n14421) );
  NOR2_X1 U16072 ( .A1(n16043), .A2(n14421), .ZN(n14579) );
  INV_X2 U16073 ( .A(n14579), .ZN(n14566) );
  NAND2_X1 U16074 ( .A1(n14566), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14422) );
  OAI211_X1 U16075 ( .C1(n14519), .C2(n15598), .A(n14553), .B(n14422), .ZN(
        P1_U2942) );
  INV_X1 U16076 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15608) );
  MUX2_X1 U16077 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n15813), .Z(
        n22223) );
  NAND2_X1 U16078 ( .A1(n14521), .A2(n22223), .ZN(n14557) );
  NAND2_X1 U16079 ( .A1(n14566), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14423) );
  OAI211_X1 U16080 ( .C1(n14519), .C2(n15608), .A(n14557), .B(n14423), .ZN(
        P1_U2943) );
  INV_X1 U16081 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15610) );
  INV_X1 U16082 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20409) );
  NOR2_X1 U16083 ( .A1(n15813), .A2(DATAI_3_), .ZN(n14424) );
  AOI21_X1 U16084 ( .B1(n15813), .B2(n20409), .A(n14424), .ZN(n22456) );
  NAND2_X1 U16085 ( .A1(n14521), .A2(n22456), .ZN(n14559) );
  NAND2_X1 U16086 ( .A1(n14566), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14425) );
  OAI211_X1 U16087 ( .C1(n15610), .C2(n14519), .A(n14559), .B(n14425), .ZN(
        P1_U2940) );
  INV_X1 U16088 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20417) );
  NOR2_X1 U16089 ( .A1(n15813), .A2(DATAI_7_), .ZN(n14426) );
  AOI21_X1 U16090 ( .B1(n15813), .B2(n20417), .A(n14426), .ZN(n22631) );
  NAND2_X1 U16091 ( .A1(n14521), .A2(n22631), .ZN(n14549) );
  NAND2_X1 U16092 ( .A1(n14566), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14427) );
  OAI211_X1 U16093 ( .C1(n14519), .C2(n15583), .A(n14549), .B(n14427), .ZN(
        P1_U2944) );
  INV_X1 U16094 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15594) );
  NAND2_X1 U16095 ( .A1(n15812), .A2(DATAI_4_), .ZN(n14429) );
  NAND2_X1 U16096 ( .A1(n15813), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14428) );
  AND2_X1 U16097 ( .A1(n14429), .A2(n14428), .ZN(n14861) );
  INV_X1 U16098 ( .A(n14861), .ZN(n16255) );
  NAND2_X1 U16099 ( .A1(n14521), .A2(n16255), .ZN(n14555) );
  NAND2_X1 U16100 ( .A1(n14566), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14430) );
  OAI211_X1 U16101 ( .C1(n15594), .C2(n14519), .A(n14555), .B(n14430), .ZN(
        P1_U2941) );
  INV_X1 U16102 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20419) );
  NAND2_X1 U16103 ( .A1(n15813), .A2(n20419), .ZN(n14431) );
  OAI21_X1 U16104 ( .B1(n15813), .B2(DATAI_8_), .A(n14431), .ZN(n15550) );
  INV_X1 U16105 ( .A(n15550), .ZN(n22376) );
  NAND2_X1 U16106 ( .A1(n14521), .A2(n22376), .ZN(n14561) );
  NAND2_X1 U16107 ( .A1(n14566), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14432) );
  OAI211_X1 U16108 ( .C1(n14519), .C2(n15592), .A(n14561), .B(n14432), .ZN(
        P1_U2945) );
  INV_X1 U16109 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15596) );
  INV_X1 U16110 ( .A(DATAI_9_), .ZN(n14434) );
  NAND2_X1 U16111 ( .A1(n15813), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U16112 ( .B1(n15813), .B2(n14434), .A(n14433), .ZN(n16249) );
  NAND2_X1 U16113 ( .A1(n14521), .A2(n16249), .ZN(n14543) );
  NAND2_X1 U16114 ( .A1(n14566), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14435) );
  OAI211_X1 U16115 ( .C1(n14519), .C2(n15596), .A(n14543), .B(n14435), .ZN(
        P1_U2946) );
  MUX2_X1 U16116 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n15813), .Z(
        n16243) );
  NAND2_X1 U16117 ( .A1(n14521), .A2(n16243), .ZN(n14547) );
  NAND2_X1 U16118 ( .A1(n14566), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14436) );
  OAI211_X1 U16119 ( .C1(n14519), .C2(n15600), .A(n14547), .B(n14436), .ZN(
        P1_U2947) );
  INV_X1 U16120 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n15613) );
  INV_X1 U16121 ( .A(DATAI_11_), .ZN(n15350) );
  NAND2_X1 U16122 ( .A1(n15813), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14437) );
  OAI21_X1 U16123 ( .B1(n15813), .B2(n15350), .A(n14437), .ZN(n16237) );
  NAND2_X1 U16124 ( .A1(n14521), .A2(n16237), .ZN(n14563) );
  NAND2_X1 U16125 ( .A1(n14566), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14438) );
  OAI211_X1 U16126 ( .C1(n14519), .C2(n15613), .A(n14563), .B(n14438), .ZN(
        P1_U2948) );
  INV_X1 U16127 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15570) );
  INV_X1 U16128 ( .A(DATAI_0_), .ZN(n14440) );
  NAND2_X1 U16129 ( .A1(n15813), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U16130 ( .B1(n15813), .B2(n14440), .A(n14439), .ZN(n22235) );
  NAND2_X1 U16131 ( .A1(n14521), .A2(n22235), .ZN(n14551) );
  NAND2_X1 U16132 ( .A1(n14566), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14441) );
  OAI211_X1 U16133 ( .C1(n15570), .C2(n14519), .A(n14551), .B(n14441), .ZN(
        P1_U2937) );
  MUX2_X1 U16134 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n15813), .Z(
        n22385) );
  NAND2_X1 U16135 ( .A1(n14521), .A2(n22385), .ZN(n14568) );
  NAND2_X1 U16136 ( .A1(n14566), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14442) );
  OAI211_X1 U16137 ( .C1(n13482), .C2(n14519), .A(n14568), .B(n14442), .ZN(
        P1_U2938) );
  INV_X1 U16138 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14873) );
  INV_X1 U16139 ( .A(DATAI_2_), .ZN(n15365) );
  NAND2_X1 U16140 ( .A1(n15812), .A2(n15365), .ZN(n14444) );
  INV_X1 U16141 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20407) );
  NAND2_X1 U16142 ( .A1(n15813), .A2(n20407), .ZN(n14443) );
  AND2_X1 U16143 ( .A1(n14444), .A2(n14443), .ZN(n16261) );
  NAND2_X1 U16144 ( .A1(n14521), .A2(n16261), .ZN(n14545) );
  NAND2_X1 U16145 ( .A1(n14566), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14445) );
  OAI211_X1 U16146 ( .C1(n14873), .C2(n14519), .A(n14545), .B(n14445), .ZN(
        P1_U2939) );
  INV_X1 U16147 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20205) );
  INV_X1 U16148 ( .A(DATAI_13_), .ZN(n14447) );
  NAND2_X1 U16149 ( .A1(n15813), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14446) );
  OAI21_X1 U16150 ( .B1(n15813), .B2(n14447), .A(n14446), .ZN(n16273) );
  NAND2_X1 U16151 ( .A1(n14521), .A2(n16273), .ZN(n14565) );
  NAND2_X1 U16152 ( .A1(n14566), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14448) );
  OAI211_X1 U16153 ( .C1(n20205), .C2(n14519), .A(n14565), .B(n14448), .ZN(
        P1_U2965) );
  INV_X1 U16154 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20207) );
  INV_X1 U16155 ( .A(DATAI_14_), .ZN(n15344) );
  NAND2_X1 U16156 ( .A1(n15813), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14449) );
  OAI21_X1 U16157 ( .B1(n15813), .B2(n15344), .A(n14449), .ZN(n16220) );
  NAND2_X1 U16158 ( .A1(n14521), .A2(n16220), .ZN(n14524) );
  NAND2_X1 U16159 ( .A1(n14566), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14450) );
  OAI211_X1 U16160 ( .C1(n20207), .C2(n14519), .A(n14524), .B(n14450), .ZN(
        P1_U2966) );
  NOR2_X1 U16161 ( .A1(n14882), .A2(n22165), .ZN(n14451) );
  NAND2_X1 U16162 ( .A1(n15824), .A2(n14451), .ZN(n17414) );
  AND2_X1 U16163 ( .A1(n17375), .A2(n17413), .ZN(n14464) );
  NOR2_X1 U16164 ( .A1(n17413), .A2(n11159), .ZN(n15835) );
  AOI21_X1 U16165 ( .B1(n15835), .B2(n21697), .A(n14452), .ZN(n14454) );
  OAI22_X1 U16166 ( .A1(n15830), .A2(n14454), .B1(n22165), .B2(n14453), .ZN(
        n14634) );
  INV_X1 U16167 ( .A(n14634), .ZN(n14463) );
  AOI21_X1 U16168 ( .B1(n14455), .B2(n14467), .A(n22236), .ZN(n14456) );
  NAND2_X1 U16169 ( .A1(n12932), .A2(n14456), .ZN(n14475) );
  AOI21_X1 U16170 ( .B1(n14475), .B2(n14458), .A(n14457), .ZN(n15828) );
  NOR2_X1 U16171 ( .A1(n14886), .A2(n14459), .ZN(n14460) );
  OR2_X1 U16172 ( .A1(n15828), .A2(n14460), .ZN(n14461) );
  AOI21_X1 U16173 ( .B1(n15830), .B2(n15905), .A(n14461), .ZN(n14462) );
  OAI211_X1 U16174 ( .C1(n17414), .C2(n14464), .A(n14463), .B(n14462), .ZN(
        n17383) );
  INV_X1 U16175 ( .A(n17383), .ZN(n17405) );
  NAND2_X1 U16176 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n17421) );
  NOR2_X1 U16177 ( .A1(n22122), .A2(n17421), .ZN(n14601) );
  NAND2_X1 U16178 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n14601), .ZN(n14465) );
  NAND2_X1 U16179 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22122), .ZN(n22126) );
  OAI211_X1 U16180 ( .C1(n17405), .C2(n22135), .A(n14465), .B(n22126), .ZN(
        n22119) );
  NAND2_X1 U16181 ( .A1(n14466), .A2(n16057), .ZN(n14470) );
  OAI21_X1 U16182 ( .B1(n15825), .B2(n15524), .A(n14636), .ZN(n14468) );
  OAI21_X1 U16183 ( .B1(n14468), .B2(n17364), .A(n14467), .ZN(n14469) );
  OAI211_X1 U16184 ( .C1(n14471), .C2(n14886), .A(n14470), .B(n14469), .ZN(
        n14472) );
  INV_X1 U16185 ( .A(n14472), .ZN(n14474) );
  NAND3_X1 U16186 ( .A1(n14475), .A2(n14474), .A3(n14473), .ZN(n15902) );
  OR2_X1 U16187 ( .A1(n15902), .A2(n14478), .ZN(n17359) );
  INV_X1 U16188 ( .A(n17359), .ZN(n17378) );
  OAI22_X1 U16189 ( .A1(n14894), .A2(n17378), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16505), .ZN(n17386) );
  INV_X1 U16190 ( .A(n17386), .ZN(n14480) );
  INV_X1 U16191 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21743) );
  AOI22_X1 U16192 ( .A1(n14483), .A2(n22129), .B1(n21743), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14479) );
  OAI21_X1 U16193 ( .B1(n14480), .B2(n16529), .A(n14479), .ZN(n14481) );
  NOR2_X1 U16194 ( .A1(n17375), .A2(n14483), .ZN(n17385) );
  AOI22_X1 U16195 ( .A1(n22119), .A2(n14481), .B1(n22116), .B2(n17385), .ZN(
        n14482) );
  OAI21_X1 U16196 ( .B1(n14483), .B2(n22119), .A(n14482), .ZN(P1_U3474) );
  NAND2_X1 U16197 ( .A1(n14485), .A2(n14484), .ZN(n14486) );
  NAND2_X1 U16198 ( .A1(n14487), .A2(n14486), .ZN(n14900) );
  OR2_X1 U16199 ( .A1(n14488), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14490) );
  AND2_X1 U16200 ( .A1(n14490), .A2(n14489), .ZN(n16492) );
  NAND2_X1 U16201 ( .A1(n20392), .A2(n16492), .ZN(n14495) );
  NAND2_X1 U16202 ( .A1(n14491), .A2(n16407), .ZN(n14493) );
  INV_X2 U16203 ( .A(n21915), .ZN(n21923) );
  NAND2_X1 U16204 ( .A1(n21923), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n16496) );
  INV_X1 U16205 ( .A(n16496), .ZN(n14492) );
  AOI21_X1 U16206 ( .B1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n14493), .A(
        n14492), .ZN(n14494) );
  OAI211_X1 U16207 ( .C1(n14900), .C2(n16413), .A(n14495), .B(n14494), .ZN(
        P1_U2999) );
  OAI21_X1 U16208 ( .B1(n14497), .B2(n14496), .A(n14582), .ZN(n18705) );
  OAI222_X1 U16209 ( .A1(n19773), .A2(n19527), .B1(n18705), .B2(n19781), .C1(
        n19770), .C2(n17524), .ZN(P2_U2912) );
  XOR2_X1 U16210 ( .A(n14499), .B(n14498), .Z(n18694) );
  INV_X1 U16211 ( .A(n18694), .ZN(n14500) );
  INV_X1 U16212 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17522) );
  OAI222_X1 U16213 ( .A1(n19773), .A2(n19724), .B1(n14500), .B2(n19781), .C1(
        n19770), .C2(n17522), .ZN(P2_U2913) );
  INV_X1 U16214 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U16215 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17541), .B1(n17542), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14501) );
  OAI21_X1 U16216 ( .B1(n15620), .B2(n14518), .A(n14501), .ZN(P2_U2935) );
  INV_X1 U16217 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U16218 ( .A1(n17542), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14502) );
  OAI21_X1 U16219 ( .B1(n16674), .B2(n14518), .A(n14502), .ZN(P2_U2928) );
  AOI22_X1 U16220 ( .A1(n17542), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14503) );
  OAI21_X1 U16221 ( .B1(n14504), .B2(n14518), .A(n14503), .ZN(P2_U2926) );
  INV_X1 U16222 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16223 ( .A1(n17542), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14505) );
  OAI21_X1 U16224 ( .B1(n14506), .B2(n14518), .A(n14505), .ZN(P2_U2929) );
  INV_X1 U16225 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16662) );
  AOI22_X1 U16226 ( .A1(n17542), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14507) );
  OAI21_X1 U16227 ( .B1(n16662), .B2(n14518), .A(n14507), .ZN(P2_U2927) );
  AOI22_X1 U16228 ( .A1(n17542), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14508) );
  OAI21_X1 U16229 ( .B1(n16611), .B2(n14518), .A(n14508), .ZN(P2_U2922) );
  AOI22_X1 U16230 ( .A1(n17542), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14509) );
  OAI21_X1 U16231 ( .B1(n16619), .B2(n14518), .A(n14509), .ZN(P2_U2923) );
  AOI22_X1 U16232 ( .A1(n17542), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14510) );
  OAI21_X1 U16233 ( .B1(n16630), .B2(n14518), .A(n14510), .ZN(P2_U2924) );
  AOI22_X1 U16234 ( .A1(n17542), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14511) );
  OAI21_X1 U16235 ( .B1(n14512), .B2(n14518), .A(n14511), .ZN(P2_U2925) );
  INV_X1 U16236 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n16683) );
  AOI22_X1 U16237 ( .A1(n17542), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14513) );
  OAI21_X1 U16238 ( .B1(n16683), .B2(n14518), .A(n14513), .ZN(P2_U2930) );
  INV_X1 U16239 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U16240 ( .A1(n17542), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14514) );
  OAI21_X1 U16241 ( .B1(n14515), .B2(n14518), .A(n14514), .ZN(P2_U2931) );
  INV_X1 U16242 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U16243 ( .A1(n17530), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14516) );
  OAI21_X1 U16244 ( .B1(n16692), .B2(n14518), .A(n14516), .ZN(P2_U2932) );
  AOI22_X1 U16245 ( .A1(n17530), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14517) );
  OAI21_X1 U16246 ( .B1(n15954), .B2(n14518), .A(n14517), .ZN(P2_U2921) );
  INV_X1 U16247 ( .A(DATAI_12_), .ZN(n15349) );
  NAND2_X1 U16248 ( .A1(n15813), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14520) );
  OAI21_X1 U16249 ( .B1(n15813), .B2(n15349), .A(n14520), .ZN(n16276) );
  NAND2_X1 U16250 ( .A1(n14521), .A2(n16276), .ZN(n14541) );
  NAND2_X1 U16251 ( .A1(n14566), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14522) );
  OAI211_X1 U16252 ( .C1(n14869), .C2(n15604), .A(n14541), .B(n14522), .ZN(
        P1_U2949) );
  NAND2_X1 U16253 ( .A1(n14566), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14523) );
  OAI211_X1 U16254 ( .C1(n14869), .C2(n15606), .A(n14524), .B(n14523), .ZN(
        P1_U2951) );
  XOR2_X1 U16255 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14525), .Z(n14530)
         );
  NAND2_X1 U16256 ( .A1(n14526), .A2(n14536), .ZN(n14528) );
  INV_X1 U16257 ( .A(n14572), .ZN(n14527) );
  AND2_X1 U16258 ( .A1(n14528), .A2(n14527), .ZN(n18683) );
  INV_X1 U16259 ( .A(n18683), .ZN(n15649) );
  MUX2_X1 U16260 ( .A(n12435), .B(n15649), .S(n16571), .Z(n14529) );
  OAI21_X1 U16261 ( .B1(n14530), .B2(n16606), .A(n14529), .ZN(P2_U2882) );
  OR2_X1 U16262 ( .A1(n14532), .A2(n14531), .ZN(n14533) );
  NAND2_X1 U16263 ( .A1(n14525), .A2(n14533), .ZN(n19775) );
  OR2_X1 U16264 ( .A1(n14535), .A2(n14534), .ZN(n14537) );
  NAND2_X1 U16265 ( .A1(n14537), .A2(n14536), .ZN(n18675) );
  NOR2_X1 U16266 ( .A1(n18675), .A2(n16604), .ZN(n14538) );
  AOI21_X1 U16267 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16604), .A(n14538), .ZN(
        n14539) );
  OAI21_X1 U16268 ( .B1(n19775), .B2(n16606), .A(n14539), .ZN(P2_U2883) );
  NAND2_X1 U16269 ( .A1(n14566), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14540) );
  OAI211_X1 U16270 ( .C1(n16280), .C2(n14869), .A(n14541), .B(n14540), .ZN(
        P1_U2964) );
  INV_X1 U16271 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20198) );
  NAND2_X1 U16272 ( .A1(n14566), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14542) );
  OAI211_X1 U16273 ( .C1(n20198), .C2(n14869), .A(n14543), .B(n14542), .ZN(
        P1_U2961) );
  NAND2_X1 U16274 ( .A1(n14566), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14544) );
  OAI211_X1 U16275 ( .C1(n13250), .C2(n14869), .A(n14545), .B(n14544), .ZN(
        P1_U2954) );
  INV_X1 U16276 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20201) );
  NAND2_X1 U16277 ( .A1(n14566), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14546) );
  OAI211_X1 U16278 ( .C1(n20201), .C2(n14869), .A(n14547), .B(n14546), .ZN(
        P1_U2962) );
  NAND2_X1 U16279 ( .A1(n14566), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14548) );
  OAI211_X1 U16280 ( .C1(n15117), .C2(n14869), .A(n14549), .B(n14548), .ZN(
        P1_U2959) );
  NAND2_X1 U16281 ( .A1(n14566), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14550) );
  OAI211_X1 U16282 ( .C1(n13256), .C2(n14869), .A(n14551), .B(n14550), .ZN(
        P1_U2952) );
  INV_X1 U16283 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20191) );
  NAND2_X1 U16284 ( .A1(n14566), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14552) );
  OAI211_X1 U16285 ( .C1(n20191), .C2(n14869), .A(n14553), .B(n14552), .ZN(
        P1_U2957) );
  INV_X1 U16286 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20189) );
  NAND2_X1 U16287 ( .A1(n14566), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14554) );
  OAI211_X1 U16288 ( .C1(n20189), .C2(n14869), .A(n14555), .B(n14554), .ZN(
        P1_U2956) );
  NAND2_X1 U16289 ( .A1(n14566), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14556) );
  OAI211_X1 U16290 ( .C1(n15092), .C2(n14869), .A(n14557), .B(n14556), .ZN(
        P1_U2958) );
  NAND2_X1 U16291 ( .A1(n14566), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14558) );
  OAI211_X1 U16292 ( .C1(n14822), .C2(n14869), .A(n14559), .B(n14558), .ZN(
        P1_U2955) );
  INV_X1 U16293 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20196) );
  NAND2_X1 U16294 ( .A1(n14566), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14560) );
  OAI211_X1 U16295 ( .C1(n20196), .C2(n14869), .A(n14561), .B(n14560), .ZN(
        P1_U2960) );
  NAND2_X1 U16296 ( .A1(n14566), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14562) );
  OAI211_X1 U16297 ( .C1(n15765), .C2(n14869), .A(n14563), .B(n14562), .ZN(
        P1_U2963) );
  INV_X1 U16298 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n15602) );
  NAND2_X1 U16299 ( .A1(n14566), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14564) );
  OAI211_X1 U16300 ( .C1(n15602), .C2(n14869), .A(n14565), .B(n14564), .ZN(
        P1_U2950) );
  NAND2_X1 U16301 ( .A1(n14566), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14567) );
  OAI211_X1 U16302 ( .C1(n13267), .C2(n14869), .A(n14568), .B(n14567), .ZN(
        P1_U2953) );
  NOR2_X1 U16303 ( .A1(n14525), .A2(n14569), .ZN(n14571) );
  OR2_X1 U16304 ( .A1(n14525), .A2(n14570), .ZN(n14612) );
  OAI211_X1 U16305 ( .C1(n14571), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16596), .B(n14612), .ZN(n14576) );
  OR2_X1 U16306 ( .A1(n14573), .A2(n14572), .ZN(n14574) );
  NAND2_X1 U16307 ( .A1(n14614), .A2(n14574), .ZN(n18698) );
  INV_X1 U16308 ( .A(n18698), .ZN(n15742) );
  NAND2_X1 U16309 ( .A1(n16571), .A2(n15742), .ZN(n14575) );
  OAI211_X1 U16310 ( .C1(n16571), .C2(n18687), .A(n14576), .B(n14575), .ZN(
        P2_U2881) );
  INV_X1 U16311 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20211) );
  INV_X1 U16312 ( .A(DATAI_15_), .ZN(n15343) );
  NOR2_X1 U16313 ( .A1(n15813), .A2(n15343), .ZN(n14577) );
  AOI21_X1 U16314 ( .B1(n15813), .B2(BUF1_REG_15__SCAN_IN), .A(n14577), .ZN(
        n16271) );
  INV_X1 U16315 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14578) );
  OAI222_X1 U16316 ( .A1(n14869), .A2(n20211), .B1(n14580), .B2(n16271), .C1(
        n14579), .C2(n14578), .ZN(P1_U2967) );
  AOI21_X1 U16317 ( .B1(n14583), .B2(n14582), .A(n14581), .ZN(n19002) );
  INV_X1 U16318 ( .A(n19002), .ZN(n14584) );
  INV_X1 U16319 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17526) );
  OAI222_X1 U16320 ( .A1(n19773), .A2(n16663), .B1(n14584), .B2(n19781), .C1(
        n19770), .C2(n17526), .ZN(P2_U2911) );
  OAI21_X1 U16321 ( .B1(n14586), .B2(n14585), .A(n14676), .ZN(n15567) );
  NOR2_X1 U16322 ( .A1(n14587), .A2(n16505), .ZN(n16516) );
  NAND2_X1 U16323 ( .A1(n15830), .A2(n16516), .ZN(n14590) );
  INV_X1 U16324 ( .A(n14588), .ZN(n14589) );
  INV_X1 U16325 ( .A(n14636), .ZN(n22633) );
  NAND4_X1 U16326 ( .A1(n14589), .A2(n17364), .A3(n15837), .A4(n22633), .ZN(
        n14632) );
  NAND2_X1 U16327 ( .A1(n14590), .A2(n14632), .ZN(n14592) );
  NOR2_X1 U16328 ( .A1(n11159), .A2(n22135), .ZN(n14591) );
  AND2_X2 U16329 ( .A1(n14592), .A2(n14591), .ZN(n20326) );
  NAND2_X1 U16330 ( .A1(n20326), .A2(n14636), .ZN(n16219) );
  INV_X1 U16331 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n15559) );
  INV_X1 U16332 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21936) );
  NAND2_X1 U16333 ( .A1(n15883), .A2(n21936), .ZN(n14593) );
  OAI211_X1 U16334 ( .C1(n11159), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14593), .B(
        n15889), .ZN(n14594) );
  INV_X1 U16335 ( .A(n15883), .ZN(n14595) );
  MUX2_X1 U16336 ( .A(n16057), .B(n14595), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14630) );
  XNOR2_X1 U16337 ( .A(n15558), .B(n11159), .ZN(n21924) );
  INV_X1 U16338 ( .A(n21924), .ZN(n14596) );
  OAI222_X1 U16339 ( .A1(n15567), .A2(n16219), .B1(n15559), .B2(n20326), .C1(
        n14596), .C2(n16217), .ZN(P1_U2871) );
  NOR2_X1 U16340 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22130) );
  INV_X1 U16341 ( .A(n22130), .ZN(n14875) );
  INV_X1 U16342 ( .A(n14597), .ZN(n14599) );
  OAI21_X1 U16343 ( .B1(n14599), .B2(n14598), .A(n17326), .ZN(n14600) );
  INV_X1 U16344 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n14602) );
  NAND2_X1 U16345 ( .A1(n14600), .A2(n14602), .ZN(n16498) );
  INV_X1 U16346 ( .A(n14601), .ZN(n22125) );
  AOI21_X1 U16347 ( .B1(n16498), .B2(n14602), .A(n22125), .ZN(n14603) );
  OR2_X1 U16348 ( .A1(n22632), .A2(n14603), .ZN(n17423) );
  INV_X1 U16349 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n22316) );
  NAND2_X1 U16350 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22316), .ZN(n16500) );
  NAND2_X1 U16351 ( .A1(n17423), .A2(n16500), .ZN(n14670) );
  NAND2_X1 U16352 ( .A1(n17423), .A2(n22292), .ZN(n14666) );
  OR2_X1 U16353 ( .A1(n14971), .A2(n22282), .ZN(n14844) );
  XNOR2_X1 U16354 ( .A(n13253), .B(n14844), .ZN(n14604) );
  OAI222_X1 U16355 ( .A1(n14670), .A2(n16514), .B1(n17423), .B2(n22237), .C1(
        n14666), .C2(n14604), .ZN(P1_U3476) );
  INV_X1 U16356 ( .A(n14657), .ZN(n14605) );
  OAI21_X1 U16357 ( .B1(n14615), .B2(n14606), .A(n14605), .ZN(n18720) );
  OAI211_X1 U16358 ( .C1(n14609), .C2(n14608), .A(n14607), .B(n16596), .ZN(
        n14611) );
  NAND2_X1 U16359 ( .A1(n16604), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14610) );
  OAI211_X1 U16360 ( .C1(n18720), .C2(n16604), .A(n14611), .B(n14610), .ZN(
        P2_U2879) );
  XOR2_X1 U16361 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14612), .Z(n14618)
         );
  AND2_X1 U16362 ( .A1(n14614), .A2(n14613), .ZN(n14616) );
  OR2_X1 U16363 ( .A1(n14616), .A2(n14615), .ZN(n18704) );
  MUX2_X1 U16364 ( .A(n12436), .B(n18704), .S(n16571), .Z(n14617) );
  OAI21_X1 U16365 ( .B1(n14618), .B2(n16606), .A(n14617), .ZN(P2_U2880) );
  INV_X1 U16366 ( .A(n18646), .ZN(n14620) );
  AOI21_X1 U16367 ( .B1(n14620), .B2(n17488), .A(n14619), .ZN(n14698) );
  XNOR2_X1 U16368 ( .A(n14698), .B(n15541), .ZN(n14693) );
  XNOR2_X1 U16369 ( .A(n14693), .B(n17481), .ZN(n14621) );
  NAND2_X1 U16370 ( .A1(n14621), .A2(n19821), .ZN(n14623) );
  INV_X1 U16371 ( .A(n15541), .ZN(n17484) );
  AOI22_X1 U16372 ( .A1(n19822), .A2(n17484), .B1(n19905), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14622) );
  OAI211_X1 U16373 ( .C1(n19918), .C2(n19773), .A(n14623), .B(n14622), .ZN(
        P2_U2917) );
  INV_X1 U16374 ( .A(n14624), .ZN(n14663) );
  INV_X1 U16375 ( .A(n14625), .ZN(n14627) );
  INV_X1 U16376 ( .A(n14581), .ZN(n14626) );
  NAND2_X1 U16377 ( .A1(n14627), .A2(n14626), .ZN(n14628) );
  NAND2_X1 U16378 ( .A1(n14663), .A2(n14628), .ZN(n18728) );
  INV_X1 U16379 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17528) );
  OAI222_X1 U16380 ( .A1(n18728), .A2(n19781), .B1(n19773), .B2(n16651), .C1(
        n19770), .C2(n17528), .ZN(P2_U2910) );
  NOR2_X1 U16381 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14629) );
  NOR2_X1 U16382 ( .A1(n14630), .A2(n14629), .ZN(n16494) );
  INV_X1 U16383 ( .A(n20326), .ZN(n16167) );
  AOI22_X1 U16384 ( .A1(n20322), .A2(n16494), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n16167), .ZN(n14631) );
  OAI21_X1 U16385 ( .B1(n16219), .B2(n14900), .A(n14631), .ZN(P1_U2872) );
  NOR2_X1 U16386 ( .A1(n14632), .A2(n14881), .ZN(n14633) );
  NAND2_X1 U16387 ( .A1(n14637), .A2(n14636), .ZN(n14638) );
  NOR2_X1 U16388 ( .A1(n22375), .A2(n14638), .ZN(n16274) );
  INV_X1 U16389 ( .A(n22235), .ZN(n14639) );
  OAI222_X1 U16390 ( .A1(n16281), .A2(n14900), .B1(n16279), .B2(n13256), .C1(
        n16278), .C2(n14639), .ZN(P1_U2904) );
  INV_X1 U16391 ( .A(n22385), .ZN(n14640) );
  OAI222_X1 U16392 ( .A1(n16281), .A2(n15567), .B1(n16279), .B2(n13267), .C1(
        n16278), .C2(n14640), .ZN(P1_U2903) );
  INV_X1 U16393 ( .A(n17360), .ZN(n14645) );
  INV_X1 U16394 ( .A(n15517), .ZN(n14643) );
  NAND2_X1 U16395 ( .A1(n15028), .A2(n22265), .ZN(n15024) );
  INV_X1 U16396 ( .A(n13253), .ZN(n14842) );
  NAND2_X1 U16397 ( .A1(n15016), .A2(n22265), .ZN(n15012) );
  INV_X1 U16398 ( .A(n15012), .ZN(n14642) );
  AOI21_X1 U16399 ( .B1(n14643), .B2(n15024), .A(n14642), .ZN(n14644) );
  OAI222_X1 U16400 ( .A1(n14670), .A2(n14645), .B1(n17423), .B2(n13197), .C1(
        n14666), .C2(n14644), .ZN(P1_U3475) );
  INV_X1 U16401 ( .A(n15567), .ZN(n14648) );
  INV_X1 U16402 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20275) );
  OAI22_X1 U16403 ( .A1(n16407), .A2(n14646), .B1(n21915), .B2(n20275), .ZN(
        n14647) );
  AOI21_X1 U16404 ( .B1(n20385), .B2(n14648), .A(n14647), .ZN(n14652) );
  OR2_X1 U16405 ( .A1(n14649), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21926) );
  NAND3_X1 U16406 ( .A1(n21926), .A2(n20392), .A3(n21927), .ZN(n14651) );
  OAI211_X1 U16407 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20395), .A(
        n14652), .B(n14651), .ZN(P1_U2998) );
  INV_X1 U16408 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n18726) );
  INV_X1 U16409 ( .A(n14607), .ZN(n14655) );
  OAI211_X1 U16410 ( .C1(n14655), .C2(n13795), .A(n16596), .B(n14654), .ZN(
        n14660) );
  OR2_X1 U16411 ( .A1(n14657), .A2(n14656), .ZN(n14658) );
  AND2_X1 U16412 ( .A1(n14709), .A2(n14658), .ZN(n17449) );
  NAND2_X1 U16413 ( .A1(n16571), .A2(n17449), .ZN(n14659) );
  OAI211_X1 U16414 ( .C1(n16571), .C2(n18726), .A(n14660), .B(n14659), .ZN(
        P2_U2878) );
  INV_X1 U16415 ( .A(n14661), .ZN(n14664) );
  AOI21_X1 U16416 ( .B1(n14664), .B2(n14663), .A(n14662), .ZN(n18741) );
  INV_X1 U16417 ( .A(n18741), .ZN(n17142) );
  INV_X1 U16418 ( .A(n16642), .ZN(n14665) );
  INV_X1 U16419 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17532) );
  OAI222_X1 U16420 ( .A1(n17142), .A2(n19781), .B1(n19773), .B2(n14665), .C1(
        n19770), .C2(n17532), .ZN(P2_U2909) );
  INV_X1 U16421 ( .A(n17423), .ZN(n14668) );
  AOI211_X1 U16422 ( .C1(n22282), .C2(n14971), .A(n22265), .B(n14666), .ZN(
        n14667) );
  AOI21_X1 U16423 ( .B1(n14668), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n14667), .ZN(n14669) );
  OAI21_X1 U16424 ( .B1(n22339), .B2(n14670), .A(n14669), .ZN(P1_U3477) );
  OAI21_X1 U16425 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n21737) );
  INV_X1 U16426 ( .A(n14674), .ZN(n14675) );
  AOI21_X1 U16427 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(n14903) );
  NAND2_X1 U16428 ( .A1(n21923), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n21739) );
  NAND2_X1 U16429 ( .A1(n20388), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14678) );
  OAI211_X1 U16430 ( .C1(n20395), .C2(n14904), .A(n21739), .B(n14678), .ZN(
        n14679) );
  AOI21_X1 U16431 ( .B1(n14903), .B2(n20385), .A(n14679), .ZN(n14680) );
  OAI21_X1 U16432 ( .B1(n22113), .B2(n21737), .A(n14680), .ZN(P1_U2997) );
  INV_X1 U16433 ( .A(n14903), .ZN(n14688) );
  INV_X1 U16434 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15490) );
  NAND2_X1 U16435 ( .A1(n15886), .A2(n15490), .ZN(n14683) );
  OAI21_X1 U16436 ( .B1(n16057), .B2(n21748), .A(n15883), .ZN(n14681) );
  OAI21_X1 U16437 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n11159), .A(n14681), .ZN(
        n14682) );
  AOI21_X1 U16438 ( .B1(n14686), .B2(n14685), .A(n14817), .ZN(n14905) );
  INV_X1 U16439 ( .A(n14905), .ZN(n21740) );
  OAI222_X1 U16440 ( .A1(n14688), .A2(n16219), .B1(n15490), .B2(n20326), .C1(
        n21740), .C2(n16217), .ZN(P1_U2870) );
  INV_X1 U16441 ( .A(n16261), .ZN(n14687) );
  OAI222_X1 U16442 ( .A1(n14688), .A2(n16281), .B1(n16279), .B2(n13250), .C1(
        n16278), .C2(n14687), .ZN(P1_U2902) );
  OR2_X1 U16443 ( .A1(n14690), .A2(n14689), .ZN(n14692) );
  NAND2_X1 U16444 ( .A1(n14692), .A2(n14691), .ZN(n19021) );
  NAND2_X1 U16445 ( .A1(n14693), .A2(n19642), .ZN(n14701) );
  XNOR2_X1 U16446 ( .A(n19660), .B(n19021), .ZN(n14699) );
  NAND2_X1 U16447 ( .A1(n14698), .A2(n17484), .ZN(n14700) );
  NAND3_X1 U16448 ( .A1(n14701), .A2(n14699), .A3(n14700), .ZN(n14830) );
  INV_X1 U16449 ( .A(n14830), .ZN(n14703) );
  AOI21_X1 U16450 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14702) );
  OAI21_X1 U16451 ( .B1(n14703), .B2(n14702), .A(n19821), .ZN(n14707) );
  INV_X1 U16452 ( .A(n16693), .ZN(n14704) );
  AOI22_X1 U16453 ( .A1(n14705), .A2(n14704), .B1(n19905), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n14706) );
  OAI211_X1 U16454 ( .C1(n19021), .C2(n19912), .A(n14707), .B(n14706), .ZN(
        P2_U2916) );
  OAI21_X1 U16455 ( .B1(n14662), .B2(n14708), .A(n14721), .ZN(n18746) );
  INV_X1 U16456 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17534) );
  OAI222_X1 U16457 ( .A1(n19773), .A2(n16631), .B1(n18746), .B2(n19781), .C1(
        n19770), .C2(n17534), .ZN(P2_U2908) );
  OAI21_X1 U16458 ( .B1(n11976), .B2(n11684), .A(n14710), .ZN(n18744) );
  INV_X1 U16459 ( .A(n14711), .ZN(n14713) );
  OAI211_X1 U16460 ( .C1(n13796), .C2(n14713), .A(n16596), .B(n14712), .ZN(
        n14715) );
  NAND2_X1 U16461 ( .A1(n16604), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14714) );
  OAI211_X1 U16462 ( .C1(n18744), .C2(n16604), .A(n14715), .B(n14714), .ZN(
        P2_U2877) );
  AND2_X1 U16463 ( .A1(n14717), .A2(n14716), .ZN(n14719) );
  OR2_X1 U16464 ( .A1(n14719), .A2(n14718), .ZN(n20320) );
  OAI222_X1 U16465 ( .A1(n16281), .A2(n20320), .B1(n16279), .B2(n20189), .C1(
        n16278), .C2(n14861), .ZN(P1_U2900) );
  INV_X1 U16466 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17536) );
  XNOR2_X1 U16467 ( .A(n14721), .B(n14720), .ZN(n18763) );
  OAI222_X1 U16468 ( .A1(n19773), .A2(n16620), .B1(n19770), .B2(n17536), .C1(
        n18763), .C2(n19781), .ZN(P2_U2907) );
  OR2_X1 U16469 ( .A1(n14758), .A2(n14766), .ZN(n14744) );
  INV_X1 U16470 ( .A(n12085), .ZN(n14723) );
  NAND2_X1 U16471 ( .A1(n14723), .A2(n14722), .ZN(n14747) );
  NAND2_X1 U16472 ( .A1(n11178), .A2(n14747), .ZN(n14728) );
  AND2_X1 U16473 ( .A1(n11198), .A2(n11240), .ZN(n14749) );
  NOR2_X1 U16474 ( .A1(n14724), .A2(n14745), .ZN(n14725) );
  NAND2_X1 U16475 ( .A1(n14374), .A2(n14725), .ZN(n14726) );
  OAI21_X1 U16476 ( .B1(n14749), .B2(n14728), .A(n14726), .ZN(n14727) );
  AOI21_X1 U16477 ( .B1(n14744), .B2(n14728), .A(n14727), .ZN(n14729) );
  OAI21_X1 U16478 ( .B1(n14730), .B2(n14741), .A(n14729), .ZN(n15675) );
  INV_X1 U16479 ( .A(n14731), .ZN(n14733) );
  INV_X1 U16480 ( .A(n14148), .ZN(n14732) );
  NAND3_X1 U16481 ( .A1(n14733), .A2(n14732), .A3(n14771), .ZN(n14740) );
  INV_X1 U16482 ( .A(n14734), .ZN(n14773) );
  OAI211_X1 U16483 ( .C1(n14773), .C2(n14770), .A(n14736), .B(n14735), .ZN(
        n14737) );
  INV_X1 U16484 ( .A(n14737), .ZN(n14739) );
  MUX2_X1 U16485 ( .A(n15675), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15630), .Z(n14802) );
  INV_X1 U16486 ( .A(n14741), .ZN(n14784) );
  NAND2_X1 U16487 ( .A1(n13756), .A2(n14784), .ZN(n14754) );
  NAND2_X1 U16488 ( .A1(n14374), .A2(n14745), .ZN(n14742) );
  NAND2_X1 U16489 ( .A1(n14742), .A2(n11178), .ZN(n14743) );
  AOI21_X1 U16490 ( .B1(n14744), .B2(n14747), .A(n14743), .ZN(n14752) );
  INV_X1 U16491 ( .A(n14745), .ZN(n14746) );
  NAND2_X1 U16492 ( .A1(n14374), .A2(n14746), .ZN(n14748) );
  OAI211_X1 U16493 ( .C1(n14749), .C2(n11204), .A(n14748), .B(n14747), .ZN(
        n14750) );
  INV_X1 U16494 ( .A(n14750), .ZN(n14751) );
  MUX2_X1 U16495 ( .A(n14752), .B(n14751), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14753) );
  NAND2_X1 U16496 ( .A1(n14754), .A2(n14753), .ZN(n15935) );
  OR2_X1 U16497 ( .A1(n15935), .A2(n15630), .ZN(n14757) );
  NAND2_X1 U16498 ( .A1(n15630), .A2(n14755), .ZN(n14756) );
  NAND2_X1 U16499 ( .A1(n14757), .A2(n14756), .ZN(n14796) );
  INV_X1 U16500 ( .A(n14796), .ZN(n14801) );
  INV_X1 U16501 ( .A(n15630), .ZN(n14793) );
  INV_X1 U16502 ( .A(n14758), .ZN(n14769) );
  NAND2_X1 U16503 ( .A1(n14759), .A2(n12422), .ZN(n14763) );
  NAND2_X1 U16504 ( .A1(n14761), .A2(n14760), .ZN(n14762) );
  NAND2_X1 U16505 ( .A1(n14763), .A2(n14762), .ZN(n14764) );
  AOI21_X1 U16506 ( .B1(n19043), .B2(n14765), .A(n14764), .ZN(n14768) );
  NAND2_X1 U16507 ( .A1(n14912), .A2(n14766), .ZN(n14767) );
  OAI211_X1 U16508 ( .C1(n14912), .C2(n14769), .A(n14768), .B(n14767), .ZN(
        n19056) );
  INV_X1 U16509 ( .A(n19056), .ZN(n14781) );
  INV_X1 U16510 ( .A(n14770), .ZN(n14772) );
  NOR3_X1 U16511 ( .A1(n14773), .A2(n14772), .A3(n14771), .ZN(n19055) );
  OR2_X1 U16512 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14779) );
  NAND2_X1 U16513 ( .A1(n14774), .A2(n14775), .ZN(n18984) );
  NOR3_X1 U16514 ( .A1(n18984), .A2(n14776), .A3(n11855), .ZN(n14778) );
  AOI211_X1 U16515 ( .C1(n19055), .C2(n14779), .A(n14778), .B(n14777), .ZN(
        n14780) );
  OAI211_X1 U16516 ( .C1(n14793), .C2(n18987), .A(n14781), .B(n14780), .ZN(
        n14800) );
  NOR2_X1 U16517 ( .A1(n14802), .A2(n19592), .ZN(n14795) );
  NAND2_X1 U16518 ( .A1(n14782), .A2(n11921), .ZN(n14786) );
  MUX2_X1 U16519 ( .A(n14374), .B(n14786), .S(n11741), .Z(n14783) );
  AOI21_X1 U16520 ( .B1(n18637), .B2(n14784), .A(n14783), .ZN(n15631) );
  AND2_X1 U16521 ( .A1(n15631), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14790) );
  NAND2_X1 U16522 ( .A1(n18648), .A2(n14784), .ZN(n14789) );
  NOR2_X1 U16523 ( .A1(n14785), .A2(n12085), .ZN(n14787) );
  AOI22_X1 U16524 ( .A1(n14374), .A2(n12073), .B1(n14787), .B2(n14786), .ZN(
        n14788) );
  AND2_X1 U16525 ( .A1(n14789), .A2(n14788), .ZN(n17176) );
  AND2_X1 U16526 ( .A1(n14790), .A2(n17176), .ZN(n14791) );
  OAI22_X1 U16527 ( .A1(n14791), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17176), .B2(n14790), .ZN(n14792) );
  AOI22_X1 U16528 ( .A1(n14802), .A2(n19592), .B1(n14793), .B2(n14792), .ZN(
        n14794) );
  AOI211_X1 U16529 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n14796), .A(
        n14795), .B(n14794), .ZN(n14797) );
  AOI21_X1 U16530 ( .B1(n14801), .B2(n19563), .A(n14797), .ZN(n14798) );
  NOR2_X1 U16531 ( .A1(n14798), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n14799) );
  AOI211_X1 U16532 ( .C1(n14802), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        n19053) );
  NAND3_X1 U16533 ( .A1(n19053), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n14913), 
        .ZN(n14806) );
  AOI22_X1 U16534 ( .A1(n14806), .A2(n14805), .B1(n14804), .B2(n14803), .ZN(
        n19046) );
  OAI21_X1 U16535 ( .B1(n19046), .B2(n11739), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14807) );
  NOR2_X1 U16536 ( .A1(n11739), .A2(n14914), .ZN(n17342) );
  INV_X1 U16537 ( .A(n17342), .ZN(n19042) );
  NAND2_X1 U16538 ( .A1(n14807), .A2(n19042), .ZN(P2_U3593) );
  XNOR2_X1 U16539 ( .A(n14712), .B(n14808), .ZN(n14812) );
  NAND2_X1 U16540 ( .A1(n14710), .A2(n14809), .ZN(n14810) );
  NAND2_X1 U16541 ( .A1(n14933), .A2(n14810), .ZN(n18758) );
  MUX2_X1 U16542 ( .A(n18758), .B(n11977), .S(n16604), .Z(n14811) );
  OAI21_X1 U16543 ( .B1(n14812), .B2(n16606), .A(n14811), .ZN(P2_U2876) );
  XOR2_X1 U16544 ( .A(n14814), .B(n14813), .Z(n15059) );
  INV_X1 U16545 ( .A(n15059), .ZN(n14823) );
  NOR2_X1 U16546 ( .A1(n11159), .A2(n16057), .ZN(n15868) );
  MUX2_X1 U16547 ( .A(n15868), .B(n16057), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n14816) );
  NOR2_X1 U16548 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14815) );
  NOR2_X1 U16549 ( .A1(n14816), .A2(n14815), .ZN(n14818) );
  OR2_X1 U16550 ( .A1(n14817), .A2(n14818), .ZN(n14819) );
  AND2_X1 U16551 ( .A1(n14947), .A2(n14819), .ZN(n21754) );
  AOI22_X1 U16552 ( .A1(n20322), .A2(n21754), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n16167), .ZN(n14820) );
  OAI21_X1 U16553 ( .B1(n14823), .B2(n16219), .A(n14820), .ZN(P1_U2869) );
  INV_X1 U16554 ( .A(n22456), .ZN(n14821) );
  OAI222_X1 U16555 ( .A1(n14823), .A2(n16281), .B1(n14822), .B2(n16279), .C1(
        n16278), .C2(n14821), .ZN(P1_U2901) );
  OAI21_X1 U16556 ( .B1(n14826), .B2(n14825), .A(n14824), .ZN(n21755) );
  AOI22_X1 U16557 ( .A1(n20388), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21923), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14827) );
  OAI21_X1 U16558 ( .B1(n20395), .B2(n15052), .A(n14827), .ZN(n14828) );
  AOI21_X1 U16559 ( .B1(n15059), .B2(n20385), .A(n14828), .ZN(n14829) );
  OAI21_X1 U16560 ( .B1(n21755), .B2(n22113), .A(n14829), .ZN(P1_U2996) );
  INV_X1 U16561 ( .A(n19021), .ZN(n17491) );
  OAI21_X1 U16562 ( .B1(n17491), .B2(n19660), .A(n14830), .ZN(n14835) );
  NAND2_X1 U16563 ( .A1(n14831), .A2(n14691), .ZN(n14834) );
  INV_X1 U16564 ( .A(n14832), .ZN(n14833) );
  NAND2_X1 U16565 ( .A1(n14834), .A2(n14833), .ZN(n18659) );
  NAND2_X1 U16566 ( .A1(n14835), .A2(n18659), .ZN(n19777) );
  XNOR2_X1 U16567 ( .A(n19777), .B(n19775), .ZN(n14836) );
  NAND2_X1 U16568 ( .A1(n14836), .A2(n19821), .ZN(n14839) );
  INV_X1 U16569 ( .A(n18659), .ZN(n14837) );
  AOI22_X1 U16570 ( .A1(n19822), .A2(n14837), .B1(n19905), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14838) );
  OAI211_X1 U16571 ( .C1(n19827), .C2(n19773), .A(n14839), .B(n14838), .ZN(
        P2_U2915) );
  NOR2_X1 U16572 ( .A1(n15813), .A2(n16413), .ZN(n22636) );
  NAND2_X1 U16573 ( .A1(n22636), .A2(DATAI_26_), .ZN(n14841) );
  AND2_X1 U16574 ( .A1(n15813), .A2(n20385), .ZN(n22635) );
  NAND2_X1 U16575 ( .A1(n22635), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14840) );
  AND2_X1 U16576 ( .A1(n14841), .A2(n14840), .ZN(n15043) );
  NAND3_X1 U16577 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n22237), .ZN(n22327) );
  INV_X1 U16578 ( .A(n22327), .ZN(n14850) );
  NOR3_X1 U16579 ( .A1(n14972), .A2(n22358), .A3(n14844), .ZN(n14845) );
  OAI21_X1 U16580 ( .B1(n14850), .B2(n14845), .A(n22268), .ZN(n22712) );
  NAND2_X1 U16581 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14855) );
  NOR2_X2 U16582 ( .A1(n14972), .A2(n22274), .ZN(n22718) );
  AOI22_X1 U16583 ( .A1(DATAI_18_), .A2(n22636), .B1(n22635), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n22455) );
  INV_X1 U16584 ( .A(n22455), .ZN(n22446) );
  INV_X1 U16585 ( .A(n22451), .ZN(n15036) );
  NOR2_X1 U16586 ( .A1(n22251), .A2(n22327), .ZN(n22711) );
  INV_X1 U16587 ( .A(n22711), .ZN(n22603) );
  NAND2_X1 U16588 ( .A1(n22632), .A2(n16261), .ZN(n22449) );
  NAND2_X1 U16589 ( .A1(n17360), .A2(n16514), .ZN(n22322) );
  INV_X1 U16590 ( .A(n14894), .ZN(n16501) );
  AND2_X1 U16591 ( .A1(n14847), .A2(n16501), .ZN(n22263) );
  INV_X1 U16592 ( .A(n22263), .ZN(n14848) );
  OAI21_X1 U16593 ( .B1(n22322), .B2(n14848), .A(n22603), .ZN(n14849) );
  NAND2_X1 U16594 ( .A1(n14849), .A2(n22292), .ZN(n14852) );
  NAND2_X1 U16595 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14850), .ZN(n14851) );
  AND2_X1 U16596 ( .A1(n14852), .A2(n14851), .ZN(n22602) );
  OAI22_X1 U16597 ( .A1(n15036), .A2(n22603), .B1(n22449), .B2(n22602), .ZN(
        n14853) );
  AOI21_X1 U16598 ( .B1(n22718), .B2(n22446), .A(n14853), .ZN(n14854) );
  OAI211_X1 U16599 ( .C1(n15043), .C2(n22715), .A(n14855), .B(n14854), .ZN(
        P1_U3123) );
  OR2_X1 U16600 ( .A1(n14718), .A2(n14857), .ZN(n14858) );
  AND2_X1 U16601 ( .A1(n14856), .A2(n14858), .ZN(n21958) );
  INV_X1 U16602 ( .A(n21958), .ZN(n14860) );
  AOI22_X1 U16603 ( .A1(n16274), .A2(n22527), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n22375), .ZN(n14859) );
  OAI21_X1 U16604 ( .B1(n14860), .B2(n16281), .A(n14859), .ZN(P1_U2899) );
  NOR2_X1 U16605 ( .A1(n22285), .A2(n14861), .ZN(n22522) );
  NAND2_X1 U16606 ( .A1(n22712), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14867) );
  NAND2_X1 U16607 ( .A1(n22636), .A2(DATAI_28_), .ZN(n14863) );
  NAND2_X1 U16608 ( .A1(n22635), .A2(BUF1_REG_28__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U16609 ( .A1(n14863), .A2(n14862), .ZN(n22523) );
  INV_X1 U16610 ( .A(n22718), .ZN(n14864) );
  INV_X1 U16611 ( .A(DATAI_20_), .ZN(n16258) );
  INV_X1 U16612 ( .A(n22636), .ZN(n22640) );
  INV_X1 U16613 ( .A(n22635), .ZN(n22639) );
  INV_X1 U16614 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20439) );
  OAI22_X1 U16615 ( .A1(n16258), .A2(n22640), .B1(n22639), .B2(n20439), .ZN(
        n22517) );
  INV_X1 U16616 ( .A(n22517), .ZN(n22526) );
  INV_X1 U16617 ( .A(n22634), .ZN(n15525) );
  NAND2_X1 U16618 ( .A1(n15525), .A2(n15892), .ZN(n14984) );
  OAI22_X1 U16619 ( .A1(n14864), .A2(n22526), .B1(n14984), .B2(n22603), .ZN(
        n14865) );
  AOI21_X1 U16620 ( .B1(n22704), .B2(n22523), .A(n14865), .ZN(n14866) );
  OAI211_X1 U16621 ( .C1(n22602), .C2(n22520), .A(n14867), .B(n14866), .ZN(
        P1_U3125) );
  NAND2_X1 U16622 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  INV_X1 U16623 ( .A(n14882), .ZN(n22161) );
  NAND2_X1 U16624 ( .A1(n20183), .A2(n15821), .ZN(n15612) );
  NOR2_X1 U16625 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17421), .ZN(n20194) );
  AOI22_X1 U16626 ( .A1(n20194), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14871) );
  OAI21_X1 U16627 ( .B1(n13482), .B2(n15612), .A(n14871), .ZN(P1_U2919) );
  AOI22_X1 U16628 ( .A1(n21698), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14872) );
  OAI21_X1 U16629 ( .B1(n14873), .B2(n15612), .A(n14872), .ZN(P1_U2918) );
  INV_X1 U16630 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17538) );
  OAI21_X1 U16631 ( .B1(n11314), .B2(n14874), .A(n15062), .ZN(n18780) );
  OAI222_X1 U16632 ( .A1(n19773), .A2(n16612), .B1(n19770), .B2(n17538), .C1(
        n18780), .C2(n19781), .ZN(P2_U2906) );
  OAI21_X1 U16633 ( .B1(n22316), .B2(n14875), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n17358) );
  OAI21_X1 U16634 ( .B1(n22121), .B2(n14876), .A(n22122), .ZN(n14877) );
  NAND2_X1 U16635 ( .A1(n17358), .A2(n14877), .ZN(n14878) );
  NAND2_X1 U16636 ( .A1(n14878), .A2(n21915), .ZN(n14879) );
  OR2_X2 U16637 ( .A1(n21696), .A2(n14879), .ZN(n22050) );
  INV_X1 U16638 ( .A(n14889), .ZN(n14885) );
  NOR2_X1 U16639 ( .A1(n14896), .A2(n22121), .ZN(n14880) );
  OAI21_X1 U16640 ( .B1(n14881), .B2(n14885), .A(n22052), .ZN(n21957) );
  INV_X1 U16641 ( .A(n21957), .ZN(n15568) );
  NAND2_X1 U16642 ( .A1(n22386), .A2(n14882), .ZN(n14883) );
  NAND2_X1 U16643 ( .A1(n14883), .A2(n21697), .ZN(n15822) );
  NAND2_X1 U16644 ( .A1(n22282), .A2(n14889), .ZN(n14884) );
  OR3_X2 U16645 ( .A1(n15822), .A2(n22236), .A3(n14884), .ZN(n22069) );
  NAND2_X1 U16646 ( .A1(n22050), .A2(n22069), .ZN(n22040) );
  OR2_X1 U16647 ( .A1(n14886), .A2(n14885), .ZN(n21940) );
  NAND2_X1 U16648 ( .A1(n21697), .A2(n22282), .ZN(n14887) );
  NAND3_X1 U16649 ( .A1(n14887), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n14889), 
        .ZN(n14888) );
  NOR2_X2 U16650 ( .A1(n11159), .A2(n14888), .ZN(n22093) );
  INV_X1 U16651 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16159) );
  OAI211_X1 U16652 ( .C1(n22386), .C2(n16159), .A(n15821), .B(n14889), .ZN(
        n14890) );
  INV_X1 U16653 ( .A(n14890), .ZN(n14892) );
  OR2_X1 U16654 ( .A1(n15822), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14891) );
  AOI22_X1 U16655 ( .A1(n16494), .A2(n22093), .B1(n22079), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n14893) );
  OAI21_X1 U16656 ( .B1(n14894), .B2(n21940), .A(n14893), .ZN(n14895) );
  AOI21_X1 U16657 ( .B1(n22040), .B2(P1_REIP_REG_0__SCAN_IN), .A(n14895), .ZN(
        n14899) );
  AND2_X1 U16658 ( .A1(n14896), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14897) );
  OAI21_X1 U16659 ( .B1(n22061), .B2(n22107), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14898) );
  OAI211_X1 U16660 ( .C1(n15568), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        P1_U2840) );
  INV_X1 U16661 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14911) );
  NOR2_X1 U16662 ( .A1(n20275), .A2(n22069), .ZN(n15048) );
  NAND2_X1 U16663 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n15048), .ZN(n15046) );
  INV_X1 U16664 ( .A(n22040), .ZN(n22085) );
  INV_X1 U16665 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20214) );
  INV_X1 U16666 ( .A(n15048), .ZN(n14901) );
  OAI21_X1 U16667 ( .B1(n22085), .B2(n20214), .A(n14901), .ZN(n14902) );
  AOI22_X1 U16668 ( .A1(n14903), .A2(n21957), .B1(n15046), .B2(n14902), .ZN(
        n14910) );
  INV_X1 U16669 ( .A(n14904), .ZN(n14908) );
  AOI22_X1 U16670 ( .A1(n14905), .A2(n22093), .B1(n22079), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14906) );
  OAI21_X1 U16671 ( .B1(n16514), .B2(n21940), .A(n14906), .ZN(n14907) );
  AOI21_X1 U16672 ( .B1(n22107), .B2(n14908), .A(n14907), .ZN(n14909) );
  OAI211_X1 U16673 ( .C1(n14911), .C2(n22098), .A(n14910), .B(n14909), .ZN(
        P1_U2838) );
  NAND2_X1 U16674 ( .A1(n19551), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19605) );
  NAND3_X1 U16675 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19534) );
  OAI21_X1 U16676 ( .B1(n19552), .B2(n19605), .A(n19534), .ZN(n14919) );
  AOI21_X1 U16677 ( .B1(n14913), .B2(n19594), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19049) );
  AND2_X1 U16678 ( .A1(n14914), .A2(n19049), .ZN(n14916) );
  INV_X1 U16679 ( .A(n14916), .ZN(n14915) );
  NAND2_X1 U16680 ( .A1(n19593), .A2(n14916), .ZN(n19699) );
  INV_X1 U16681 ( .A(n19699), .ZN(n19712) );
  NAND2_X1 U16682 ( .A1(n12533), .A2(n19712), .ZN(n14917) );
  OAI211_X1 U16683 ( .C1(n20005), .C2(n19714), .A(n14917), .B(n19648), .ZN(
        n14918) );
  NAND2_X1 U16684 ( .A1(n14919), .A2(n14918), .ZN(n20012) );
  INV_X1 U16685 ( .A(n20012), .ZN(n19533) );
  INV_X1 U16686 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14926) );
  INV_X1 U16687 ( .A(n19714), .ZN(n20008) );
  OAI21_X1 U16688 ( .B1(n12533), .B2(n20008), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14920) );
  OAI21_X1 U16689 ( .B1(n19534), .B2(n19694), .A(n14920), .ZN(n20009) );
  NOR2_X2 U16690 ( .A1(n16693), .A2(n20005), .ZN(n19901) );
  NOR2_X2 U16691 ( .A1(n14921), .A2(n20007), .ZN(n19898) );
  INV_X1 U16692 ( .A(n19898), .ZN(n14923) );
  NAND2_X1 U16693 ( .A1(n19551), .A2(n19550), .ZN(n19643) );
  AOI22_X1 U16694 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20010), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20011), .ZN(n19895) );
  NAND2_X1 U16695 ( .A1(n19551), .A2(n17477), .ZN(n19657) );
  AOI22_X1 U16696 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20010), .ZN(n19904) );
  INV_X1 U16697 ( .A(n19904), .ZN(n19892) );
  AOI22_X1 U16698 ( .A1(n20109), .A2(n19900), .B1(n19966), .B2(n19892), .ZN(
        n14922) );
  OAI21_X1 U16699 ( .B1(n14923), .B2(n19714), .A(n14922), .ZN(n14924) );
  AOI21_X1 U16700 ( .B1(n20009), .B2(n19901), .A(n14924), .ZN(n14925) );
  OAI21_X1 U16701 ( .B1(n19533), .B2(n14926), .A(n14925), .ZN(P2_U3171) );
  INV_X1 U16702 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14931) );
  NOR2_X2 U16703 ( .A1(n19772), .A2(n20005), .ZN(n19815) );
  NOR2_X2 U16704 ( .A1(n12574), .A2(n20007), .ZN(n19813) );
  INV_X1 U16705 ( .A(n19813), .ZN(n14928) );
  INV_X1 U16706 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21028) );
  INV_X1 U16707 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n22531) );
  OAI22_X1 U16708 ( .A1(n21028), .A2(n19961), .B1(n22531), .B2(n19960), .ZN(
        n19814) );
  AOI22_X1 U16709 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20010), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20011), .ZN(n19818) );
  AOI22_X1 U16710 ( .A1(n20109), .A2(n19814), .B1(n19966), .B2(n19808), .ZN(
        n14927) );
  OAI21_X1 U16711 ( .B1(n14928), .B2(n19714), .A(n14927), .ZN(n14929) );
  AOI21_X1 U16712 ( .B1(n20009), .B2(n19815), .A(n14929), .ZN(n14930) );
  OAI21_X1 U16713 ( .B1(n19533), .B2(n14931), .A(n14930), .ZN(P2_U3173) );
  AND2_X1 U16714 ( .A1(n14933), .A2(n14932), .ZN(n14934) );
  OR2_X1 U16715 ( .A1(n14934), .A2(n14941), .ZN(n18764) );
  OAI211_X1 U16716 ( .C1(n11315), .C2(n14936), .A(n14935), .B(n16596), .ZN(
        n14938) );
  NAND2_X1 U16717 ( .A1(n16604), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14937) );
  OAI211_X1 U16718 ( .C1(n18764), .C2(n16604), .A(n14938), .B(n14937), .ZN(
        P2_U2875) );
  XOR2_X1 U16719 ( .A(n15100), .B(n14939), .Z(n14945) );
  OR2_X1 U16720 ( .A1(n14941), .A2(n14940), .ZN(n14942) );
  AND2_X1 U16721 ( .A1(n15096), .A2(n14942), .ZN(n18777) );
  INV_X1 U16722 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18769) );
  NOR2_X1 U16723 ( .A1(n16571), .A2(n18769), .ZN(n14943) );
  AOI21_X1 U16724 ( .B1(n18777), .B2(n16571), .A(n14943), .ZN(n14944) );
  OAI21_X1 U16725 ( .B1(n14945), .B2(n16606), .A(n14944), .ZN(P2_U2874) );
  XNOR2_X1 U16726 ( .A(n14856), .B(n13299), .ZN(n21968) );
  INV_X1 U16727 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20319) );
  NAND2_X1 U16728 ( .A1(n15868), .A2(n20319), .ZN(n14950) );
  NAND2_X1 U16729 ( .A1(n15889), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14948) );
  OAI211_X1 U16730 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n11159), .A(n14948), .B(
        n15883), .ZN(n14949) );
  AND2_X1 U16731 ( .A1(n14950), .A2(n14949), .ZN(n20313) );
  NAND2_X1 U16732 ( .A1(n15883), .A2(n15910), .ZN(n14951) );
  OAI211_X1 U16733 ( .C1(n11159), .C2(P1_EBX_REG_4__SCAN_IN), .A(n14951), .B(
        n15889), .ZN(n14952) );
  OAI21_X1 U16734 ( .B1(n15878), .B2(P1_EBX_REG_4__SCAN_IN), .A(n14952), .ZN(
        n20321) );
  INV_X1 U16735 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n14959) );
  NAND2_X1 U16736 ( .A1(n15886), .A2(n14959), .ZN(n14956) );
  NAND2_X1 U16737 ( .A1(n15883), .A2(n21762), .ZN(n14954) );
  OAI211_X1 U16738 ( .C1(n11159), .C2(P1_EBX_REG_6__SCAN_IN), .A(n14954), .B(
        n15889), .ZN(n14955) );
  AND2_X1 U16739 ( .A1(n20316), .A2(n14957), .ZN(n14958) );
  OR2_X1 U16740 ( .A1(n14958), .A2(n15113), .ZN(n21966) );
  OAI22_X1 U16741 ( .A1(n16217), .A2(n21966), .B1(n14959), .B2(n20326), .ZN(
        n14960) );
  AOI21_X1 U16742 ( .B1(n21968), .B2(n20323), .A(n14960), .ZN(n14961) );
  INV_X1 U16743 ( .A(n14961), .ZN(P1_U2866) );
  OR2_X1 U16744 ( .A1(n22322), .A2(n14979), .ZN(n14962) );
  NAND3_X1 U16745 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n22238), .A3(
        n22237), .ZN(n22307) );
  NOR2_X1 U16746 ( .A1(n22251), .A2(n22307), .ZN(n22698) );
  INV_X1 U16747 ( .A(n22698), .ZN(n14973) );
  NAND2_X1 U16748 ( .A1(n14962), .A2(n14973), .ZN(n14965) );
  NAND2_X1 U16749 ( .A1(n14965), .A2(n22292), .ZN(n14964) );
  INV_X1 U16750 ( .A(n22307), .ZN(n14968) );
  NAND2_X1 U16751 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14968), .ZN(n14963) );
  NAND2_X1 U16752 ( .A1(n14964), .A2(n14963), .ZN(n22697) );
  INV_X1 U16753 ( .A(n22697), .ZN(n14978) );
  INV_X1 U16754 ( .A(n14965), .ZN(n14966) );
  OAI21_X1 U16755 ( .B1(n14972), .B2(n22282), .A(n14966), .ZN(n14967) );
  OAI221_X1 U16756 ( .B1(n22292), .B2(n14968), .C1(n22358), .C2(n14967), .A(
        n22268), .ZN(n22699) );
  NAND2_X1 U16757 ( .A1(n22699), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14977) );
  INV_X1 U16758 ( .A(n22702), .ZN(n22311) );
  NAND2_X1 U16759 ( .A1(n14971), .A2(n14970), .ZN(n15518) );
  NOR2_X2 U16760 ( .A1(n14972), .A2(n15518), .ZN(n22705) );
  INV_X1 U16761 ( .A(n22705), .ZN(n14974) );
  OAI22_X1 U16762 ( .A1(n14974), .A2(n22526), .B1(n14973), .B2(n14984), .ZN(
        n14975) );
  AOI21_X1 U16763 ( .B1(n22311), .B2(n22523), .A(n14975), .ZN(n14976) );
  OAI211_X1 U16764 ( .C1(n14978), .C2(n22520), .A(n14977), .B(n14976), .ZN(
        P1_U3109) );
  NOR2_X1 U16765 ( .A1(n16514), .A2(n14988), .ZN(n22295) );
  INV_X1 U16766 ( .A(n14979), .ZN(n22252) );
  NAND3_X1 U16767 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n22238), .A3(
        n13197), .ZN(n22278) );
  NOR2_X1 U16768 ( .A1(n22251), .A2(n22278), .ZN(n22673) );
  AOI21_X1 U16769 ( .B1(n22295), .B2(n22252), .A(n22673), .ZN(n14980) );
  OAI22_X1 U16770 ( .A1(n14980), .A2(n22358), .B1(n22278), .B2(n22253), .ZN(
        n22672) );
  INV_X1 U16771 ( .A(n22672), .ZN(n15001) );
  INV_X1 U16772 ( .A(n22278), .ZN(n14983) );
  INV_X1 U16773 ( .A(n15016), .ZN(n14981) );
  OAI21_X1 U16774 ( .B1(n14981), .B2(n22282), .A(n14980), .ZN(n14982) );
  OAI221_X1 U16775 ( .B1(n22292), .B2(n14983), .C1(n22358), .C2(n14982), .A(
        n22268), .ZN(n22675) );
  NAND2_X1 U16776 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14987) );
  INV_X1 U16777 ( .A(n22523), .ZN(n15037) );
  INV_X1 U16778 ( .A(n15518), .ZN(n14997) );
  OAI22_X1 U16779 ( .A1(n15037), .A2(n22671), .B1(n22683), .B2(n22526), .ZN(
        n14985) );
  AOI21_X1 U16780 ( .B1(n22521), .B2(n22673), .A(n14985), .ZN(n14986) );
  OAI211_X1 U16781 ( .C1(n15001), .C2(n22520), .A(n14987), .B(n14986), .ZN(
        P1_U3077) );
  INV_X1 U16782 ( .A(n14988), .ZN(n17320) );
  NOR2_X1 U16783 ( .A1(n16514), .A2(n17320), .ZN(n22355) );
  NAND2_X1 U16784 ( .A1(n22355), .A2(n22252), .ZN(n14989) );
  NAND3_X1 U16785 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(n22238), .ZN(n22343) );
  NOR2_X1 U16786 ( .A1(n22251), .A2(n22343), .ZN(n22725) );
  INV_X1 U16787 ( .A(n22725), .ZN(n22612) );
  NAND2_X1 U16788 ( .A1(n14989), .A2(n22612), .ZN(n14992) );
  NAND2_X1 U16789 ( .A1(n14992), .A2(n22292), .ZN(n14991) );
  INV_X1 U16790 ( .A(n22343), .ZN(n14996) );
  NAND2_X1 U16791 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14996), .ZN(n14990) );
  AND2_X1 U16792 ( .A1(n14991), .A2(n14990), .ZN(n22611) );
  INV_X1 U16793 ( .A(n15028), .ZN(n14994) );
  INV_X1 U16794 ( .A(n14992), .ZN(n14993) );
  OAI21_X1 U16795 ( .B1(n14994), .B2(n22282), .A(n14993), .ZN(n14995) );
  OAI221_X1 U16796 ( .B1(n22292), .B2(n14996), .C1(n22358), .C2(n14995), .A(
        n22268), .ZN(n22726) );
  NAND2_X1 U16797 ( .A1(n22726), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n15000) );
  INV_X1 U16798 ( .A(n22733), .ZN(n15006) );
  NAND2_X1 U16799 ( .A1(n15028), .A2(n22230), .ZN(n22729) );
  OAI22_X1 U16800 ( .A1(n15006), .A2(n22526), .B1(n15037), .B2(n22729), .ZN(
        n14998) );
  AOI21_X1 U16801 ( .B1(n22521), .B2(n22725), .A(n14998), .ZN(n14999) );
  OAI211_X1 U16802 ( .C1(n22611), .C2(n22520), .A(n15000), .B(n14999), .ZN(
        P1_U3141) );
  INV_X1 U16803 ( .A(n22673), .ZN(n15005) );
  NAND2_X1 U16804 ( .A1(n22675), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n15004) );
  INV_X1 U16805 ( .A(n15043), .ZN(n22452) );
  OAI22_X1 U16806 ( .A1(n22683), .A2(n22455), .B1(n22449), .B2(n15001), .ZN(
        n15002) );
  AOI21_X1 U16807 ( .B1(n22674), .B2(n22452), .A(n15002), .ZN(n15003) );
  OAI211_X1 U16808 ( .C1(n15036), .C2(n15005), .A(n15004), .B(n15003), .ZN(
        P1_U3075) );
  NAND2_X1 U16809 ( .A1(n22726), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n15009) );
  OAI22_X1 U16810 ( .A1(n15006), .A2(n22455), .B1(n22449), .B2(n22611), .ZN(
        n15007) );
  AOI21_X1 U16811 ( .B1(n22717), .B2(n22452), .A(n15007), .ZN(n15008) );
  OAI211_X1 U16812 ( .C1(n15036), .C2(n22612), .A(n15009), .B(n15008), .ZN(
        P1_U3139) );
  INV_X1 U16813 ( .A(n22589), .ZN(n22685) );
  AOI21_X1 U16814 ( .B1(n22295), .B2(n22263), .A(n22685), .ZN(n15013) );
  OR2_X1 U16815 ( .A1(n15013), .A2(n22358), .ZN(n15011) );
  NAND3_X1 U16816 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(n13197), .ZN(n22291) );
  INV_X1 U16817 ( .A(n22291), .ZN(n15015) );
  NAND2_X1 U16818 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15015), .ZN(n15010) );
  AND2_X1 U16819 ( .A1(n15011), .A2(n15010), .ZN(n22588) );
  NAND2_X1 U16820 ( .A1(n15013), .A2(n15012), .ZN(n15014) );
  OAI221_X1 U16821 ( .B1(n22292), .B2(n15015), .C1(n22358), .C2(n15014), .A(
        n22268), .ZN(n22687) );
  NAND2_X1 U16822 ( .A1(n22687), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n15019) );
  INV_X1 U16823 ( .A(n22693), .ZN(n22690) );
  OAI22_X1 U16824 ( .A1(n15037), .A2(n22593), .B1(n22690), .B2(n22526), .ZN(
        n15017) );
  AOI21_X1 U16825 ( .B1(n22685), .B2(n22521), .A(n15017), .ZN(n15018) );
  OAI211_X1 U16826 ( .C1(n22588), .C2(n22520), .A(n15019), .B(n15018), .ZN(
        P1_U3093) );
  NAND2_X1 U16827 ( .A1(n22687), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n15022) );
  OAI22_X1 U16828 ( .A1(n22690), .A2(n22455), .B1(n22449), .B2(n22588), .ZN(
        n15020) );
  AOI21_X1 U16829 ( .B1(n22686), .B2(n22452), .A(n15020), .ZN(n15021) );
  OAI211_X1 U16830 ( .C1(n15036), .C2(n22589), .A(n15022), .B(n15021), .ZN(
        P1_U3091) );
  NOR2_X1 U16831 ( .A1(n15023), .A2(n13197), .ZN(n22741) );
  INV_X1 U16832 ( .A(n22741), .ZN(n22624) );
  NAND3_X1 U16833 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22353) );
  INV_X1 U16834 ( .A(n22353), .ZN(n15030) );
  AOI21_X1 U16835 ( .B1(n22355), .B2(n22263), .A(n22741), .ZN(n15029) );
  NAND2_X1 U16836 ( .A1(n15024), .A2(n15029), .ZN(n15025) );
  OAI221_X1 U16837 ( .B1(n22292), .B2(n15030), .C1(n22358), .C2(n15025), .A(
        n22268), .ZN(n22744) );
  NAND2_X1 U16838 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n15035) );
  INV_X1 U16839 ( .A(n22747), .ZN(n22359) );
  OR2_X1 U16840 ( .A1(n15029), .A2(n22358), .ZN(n15032) );
  NAND2_X1 U16841 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15030), .ZN(n15031) );
  AND2_X1 U16842 ( .A1(n15032), .A2(n15031), .ZN(n22622) );
  OAI22_X1 U16843 ( .A1(n22232), .A2(n22455), .B1(n22449), .B2(n22622), .ZN(
        n15033) );
  AOI21_X1 U16844 ( .B1(n22359), .B2(n22452), .A(n15033), .ZN(n15034) );
  OAI211_X1 U16845 ( .C1(n15036), .C2(n22624), .A(n15035), .B(n15034), .ZN(
        P1_U3155) );
  NAND2_X1 U16846 ( .A1(n22744), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n15040) );
  OAI22_X1 U16847 ( .A1(n22232), .A2(n22526), .B1(n15037), .B2(n22747), .ZN(
        n15038) );
  AOI21_X1 U16848 ( .B1(n22521), .B2(n22741), .A(n15038), .ZN(n15039) );
  OAI211_X1 U16849 ( .C1(n22622), .C2(n22520), .A(n15040), .B(n15039), .ZN(
        P1_U3157) );
  INV_X1 U16850 ( .A(n22449), .ZN(n22450) );
  AOI22_X1 U16851 ( .A1(n22451), .A2(n22698), .B1(n22450), .B2(n22697), .ZN(
        n15042) );
  NAND2_X1 U16852 ( .A1(n22705), .A2(n22446), .ZN(n15041) );
  OAI211_X1 U16853 ( .C1(n15043), .C2(n22702), .A(n15042), .B(n15041), .ZN(
        n15044) );
  AOI21_X1 U16854 ( .B1(n22699), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n15044), .ZN(n15045) );
  INV_X1 U16855 ( .A(n15045), .ZN(P1_U3107) );
  INV_X1 U16856 ( .A(n15046), .ZN(n15047) );
  AOI21_X1 U16857 ( .B1(n22040), .B2(P1_REIP_REG_3__SCAN_IN), .A(n15047), .ZN(
        n15057) );
  NAND3_X1 U16858 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(n15048), .ZN(n21942) );
  INV_X1 U16859 ( .A(n21942), .ZN(n15056) );
  INV_X1 U16860 ( .A(n21940), .ZN(n15562) );
  NAND2_X1 U16861 ( .A1(n17360), .A2(n15562), .ZN(n15050) );
  AOI22_X1 U16862 ( .A1(n21754), .A2(n22093), .B1(n22079), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n15049) );
  NAND2_X1 U16863 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  AOI21_X1 U16864 ( .B1(n22061), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15051), .ZN(n15055) );
  INV_X1 U16865 ( .A(n15052), .ZN(n15053) );
  NAND2_X1 U16866 ( .A1(n22107), .A2(n15053), .ZN(n15054) );
  OAI211_X1 U16867 ( .C1(n15057), .C2(n15056), .A(n15055), .B(n15054), .ZN(
        n15058) );
  AOI21_X1 U16868 ( .B1(n15059), .B2(n21957), .A(n15058), .ZN(n15060) );
  INV_X1 U16869 ( .A(n15060), .ZN(P1_U2837) );
  AOI21_X1 U16870 ( .B1(n15063), .B2(n15062), .A(n15061), .ZN(n18787) );
  INV_X1 U16871 ( .A(n18787), .ZN(n15064) );
  INV_X1 U16872 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17540) );
  OAI222_X1 U16873 ( .A1(n19773), .A2(n15955), .B1(n15064), .B2(n19781), .C1(
        n19770), .C2(n17540), .ZN(P2_U2905) );
  XNOR2_X1 U16874 ( .A(n15065), .B(n19030), .ZN(n15087) );
  AOI22_X1 U16875 ( .A1(n15087), .A2(n15066), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15065), .ZN(n15068) );
  XNOR2_X1 U16876 ( .A(n18658), .B(n15643), .ZN(n15067) );
  XNOR2_X1 U16877 ( .A(n15068), .B(n15067), .ZN(n15084) );
  OAI21_X1 U16878 ( .B1(n15070), .B2(n15643), .A(n11185), .ZN(n15082) );
  INV_X1 U16879 ( .A(n19015), .ZN(n19007) );
  AND2_X1 U16880 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19026), .ZN(
        n15749) );
  INV_X1 U16881 ( .A(n17048), .ZN(n15071) );
  OAI21_X1 U16882 ( .B1(n15071), .B2(n15751), .A(n15072), .ZN(n19027) );
  NAND2_X1 U16883 ( .A1(n15749), .A2(n19027), .ZN(n15641) );
  NOR2_X1 U16884 ( .A1(n17047), .A2(n17048), .ZN(n19001) );
  INV_X1 U16885 ( .A(n18994), .ZN(n17170) );
  NOR2_X1 U16886 ( .A1(n15072), .A2(n19026), .ZN(n15073) );
  AOI211_X1 U16887 ( .C1(n17048), .C2(n15751), .A(n17170), .B(n15073), .ZN(
        n19031) );
  OAI21_X1 U16888 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19001), .A(
        n19031), .ZN(n15646) );
  INV_X1 U16889 ( .A(n15646), .ZN(n15075) );
  NAND2_X1 U16890 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n11167), .ZN(n15074) );
  OAI221_X1 U16891 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15641), .C1(
        n15643), .C2(n15075), .A(n15074), .ZN(n15077) );
  OAI22_X1 U16892 ( .A1(n18675), .A2(n18991), .B1(n19020), .B2(n18659), .ZN(
        n15076) );
  AOI211_X1 U16893 ( .C1(n15082), .C2(n19007), .A(n15077), .B(n15076), .ZN(
        n15078) );
  OAI21_X1 U16894 ( .B1(n15084), .B2(n17166), .A(n15078), .ZN(P2_U3042) );
  OAI22_X1 U16895 ( .A1(n11952), .A2(n18830), .B1(n17475), .B2(n18668), .ZN(
        n15079) );
  AOI21_X1 U16896 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17461), .A(
        n15079), .ZN(n15080) );
  OAI21_X1 U16897 ( .B1(n17471), .B2(n18675), .A(n15080), .ZN(n15081) );
  AOI21_X1 U16898 ( .B1(n15082), .B2(n17467), .A(n15081), .ZN(n15083) );
  OAI21_X1 U16899 ( .B1(n15084), .B2(n17445), .A(n15083), .ZN(P2_U3010) );
  XNOR2_X1 U16900 ( .A(n12767), .B(n15085), .ZN(n19016) );
  XNOR2_X1 U16901 ( .A(n15087), .B(n15086), .ZN(n19025) );
  NAND2_X1 U16902 ( .A1(n19025), .A2(n17462), .ZN(n15091) );
  NAND2_X1 U16903 ( .A1(n17443), .A2(n15944), .ZN(n15088) );
  NAND2_X1 U16904 ( .A1(n11167), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n19019) );
  OAI211_X1 U16905 ( .C1(n15946), .C2(n17452), .A(n15088), .B(n19019), .ZN(
        n15089) );
  AOI21_X1 U16906 ( .B1(n17457), .B2(n13756), .A(n15089), .ZN(n15090) );
  OAI211_X1 U16907 ( .C1(n19016), .C2(n17446), .A(n15091), .B(n15090), .ZN(
        P2_U3011) );
  INV_X1 U16908 ( .A(n22223), .ZN(n15094) );
  INV_X1 U16909 ( .A(n21968), .ZN(n15093) );
  OAI222_X1 U16910 ( .A1(n16278), .A2(n15094), .B1(n16281), .B2(n15093), .C1(
        n15092), .C2(n16279), .ZN(P1_U2898) );
  AOI21_X1 U16911 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n18788) );
  INV_X1 U16912 ( .A(n18788), .ZN(n17089) );
  INV_X1 U16913 ( .A(n15098), .ZN(n15102) );
  OAI21_X1 U16914 ( .B1(n14935), .B2(n15100), .A(n15099), .ZN(n15101) );
  NAND3_X1 U16915 ( .A1(n15102), .A2(n15101), .A3(n16596), .ZN(n15104) );
  NAND2_X1 U16916 ( .A1(n16604), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15103) );
  OAI211_X1 U16917 ( .C1(n17089), .C2(n16604), .A(n15104), .B(n15103), .ZN(
        P2_U2873) );
  XNOR2_X1 U16918 ( .A(n15061), .B(n15105), .ZN(n18804) );
  OAI222_X1 U16919 ( .A1(n19773), .A2(n15106), .B1(n19770), .B2(n17545), .C1(
        n19781), .C2(n18804), .ZN(P2_U2904) );
  NAND2_X1 U16920 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  AND2_X1 U16921 ( .A1(n15107), .A2(n15110), .ZN(n21983) );
  INV_X1 U16922 ( .A(n21983), .ZN(n15116) );
  INV_X1 U16923 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21980) );
  MUX2_X1 U16924 ( .A(n15868), .B(n16057), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n15112) );
  NOR2_X1 U16925 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15111) );
  NOR2_X1 U16926 ( .A1(n15112), .A2(n15111), .ZN(n15114) );
  NOR2_X1 U16927 ( .A1(n15113), .A2(n15114), .ZN(n15115) );
  OR2_X1 U16928 ( .A1(n15125), .A2(n15115), .ZN(n21976) );
  OAI222_X1 U16929 ( .A1(n15116), .A2(n16219), .B1(n20326), .B2(n21980), .C1(
        n21976), .C2(n16217), .ZN(P1_U2865) );
  INV_X1 U16930 ( .A(n22631), .ZN(n15118) );
  OAI222_X1 U16931 ( .A1(n15118), .A2(n16278), .B1(n15117), .B2(n16279), .C1(
        n15116), .C2(n16281), .ZN(P1_U2897) );
  AOI21_X1 U16932 ( .B1(n15120), .B2(n15107), .A(n15119), .ZN(n15701) );
  INV_X1 U16933 ( .A(n15701), .ZN(n15549) );
  INV_X1 U16934 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21977) );
  INV_X1 U16935 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20223) );
  INV_X1 U16936 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21955) );
  NAND4_X1 U16937 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n21950)
         );
  NOR2_X1 U16938 ( .A1(n21955), .A2(n21950), .ZN(n21963) );
  NAND2_X1 U16939 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21963), .ZN(n21965) );
  NOR3_X1 U16940 ( .A1(n21977), .A2(n20223), .A3(n21965), .ZN(n15703) );
  OAI21_X1 U16941 ( .B1(n15703), .B2(n22069), .A(n22050), .ZN(n15585) );
  INV_X1 U16942 ( .A(n21965), .ZN(n21961) );
  INV_X2 U16943 ( .A(n22069), .ZN(n22073) );
  NAND2_X1 U16944 ( .A1(n21961), .A2(n22073), .ZN(n21981) );
  OAI21_X1 U16945 ( .B1(n21977), .B2(n21981), .A(n20223), .ZN(n15129) );
  NOR2_X1 U16946 ( .A1(n21964), .A2(n20399), .ZN(n22044) );
  AOI21_X1 U16947 ( .B1(n22079), .B2(P1_EBX_REG_8__SCAN_IN), .A(n22044), .ZN(
        n15121) );
  OAI21_X1 U16948 ( .B1(n22096), .B2(n15699), .A(n15121), .ZN(n15128) );
  NAND2_X1 U16949 ( .A1(n15883), .A2(n21798), .ZN(n15122) );
  OAI211_X1 U16950 ( .C1(n11159), .C2(P1_EBX_REG_8__SCAN_IN), .A(n15122), .B(
        n15889), .ZN(n15123) );
  OAI21_X1 U16951 ( .B1(n15878), .B2(P1_EBX_REG_8__SCAN_IN), .A(n15123), .ZN(
        n15124) );
  OR2_X1 U16952 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  NAND2_X1 U16953 ( .A1(n15684), .A2(n15126), .ZN(n21792) );
  OAI22_X1 U16954 ( .A1(n13317), .A2(n22098), .B1(n22111), .B2(n21792), .ZN(
        n15127) );
  AOI211_X1 U16955 ( .C1(n15585), .C2(n15129), .A(n15128), .B(n15127), .ZN(
        n15130) );
  OAI21_X1 U16956 ( .B1(n15549), .B2(n22052), .A(n15130), .ZN(P1_U2832) );
  INV_X1 U16957 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15131) );
  OAI222_X1 U16958 ( .A1(n15549), .A2(n16219), .B1(n15131), .B2(n20326), .C1(
        n21792), .C2(n16217), .ZN(P1_U2864) );
  XOR2_X1 U16959 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_128), .Z(n15134) );
  INV_X1 U16960 ( .A(DATAI_31_), .ZN(n15817) );
  XNOR2_X1 U16961 ( .A(n15817), .B(keyinput_129), .ZN(n15133) );
  INV_X1 U16962 ( .A(DATAI_30_), .ZN(n16223) );
  XNOR2_X1 U16963 ( .A(n16223), .B(keyinput_130), .ZN(n15132) );
  AOI21_X1 U16964 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(n15138) );
  XOR2_X1 U16965 ( .A(DATAI_28_), .B(keyinput_132), .Z(n15137) );
  XOR2_X1 U16966 ( .A(DATAI_29_), .B(keyinput_131), .Z(n15136) );
  XNOR2_X1 U16967 ( .A(DATAI_27_), .B(keyinput_133), .ZN(n15135) );
  NOR4_X1 U16968 ( .A1(n15138), .A2(n15137), .A3(n15136), .A4(n15135), .ZN(
        n15141) );
  XNOR2_X1 U16969 ( .A(DATAI_26_), .B(keyinput_134), .ZN(n15140) );
  XNOR2_X1 U16970 ( .A(DATAI_25_), .B(keyinput_135), .ZN(n15139) );
  OAI21_X1 U16971 ( .B1(n15141), .B2(n15140), .A(n15139), .ZN(n15147) );
  XOR2_X1 U16972 ( .A(DATAI_24_), .B(keyinput_136), .Z(n15146) );
  XNOR2_X1 U16973 ( .A(DATAI_22_), .B(keyinput_138), .ZN(n15144) );
  XNOR2_X1 U16974 ( .A(DATAI_21_), .B(keyinput_139), .ZN(n15143) );
  XNOR2_X1 U16975 ( .A(DATAI_23_), .B(keyinput_137), .ZN(n15142) );
  NAND3_X1 U16976 ( .A1(n15144), .A2(n15143), .A3(n15142), .ZN(n15145) );
  AOI21_X1 U16977 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15151) );
  XOR2_X1 U16978 ( .A(DATAI_19_), .B(keyinput_141), .Z(n15150) );
  XOR2_X1 U16979 ( .A(DATAI_20_), .B(keyinput_140), .Z(n15149) );
  XNOR2_X1 U16980 ( .A(DATAI_18_), .B(keyinput_142), .ZN(n15148) );
  NOR4_X1 U16981 ( .A1(n15151), .A2(n15150), .A3(n15149), .A4(n15148), .ZN(
        n15154) );
  XOR2_X1 U16982 ( .A(DATAI_17_), .B(keyinput_143), .Z(n15153) );
  XOR2_X1 U16983 ( .A(DATAI_16_), .B(keyinput_144), .Z(n15152) );
  OAI21_X1 U16984 ( .B1(n15154), .B2(n15153), .A(n15152), .ZN(n15158) );
  XNOR2_X1 U16985 ( .A(n15343), .B(keyinput_145), .ZN(n15157) );
  XNOR2_X1 U16986 ( .A(n15344), .B(keyinput_146), .ZN(n15156) );
  XNOR2_X1 U16987 ( .A(DATAI_13_), .B(keyinput_147), .ZN(n15155) );
  AOI211_X1 U16988 ( .C1(n15158), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        n15161) );
  XNOR2_X1 U16989 ( .A(n15349), .B(keyinput_148), .ZN(n15160) );
  XNOR2_X1 U16990 ( .A(n15350), .B(keyinput_149), .ZN(n15159) );
  OAI21_X1 U16991 ( .B1(n15161), .B2(n15160), .A(n15159), .ZN(n15165) );
  XOR2_X1 U16992 ( .A(DATAI_8_), .B(keyinput_152), .Z(n15164) );
  XNOR2_X1 U16993 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n15163) );
  XNOR2_X1 U16994 ( .A(DATAI_9_), .B(keyinput_151), .ZN(n15162) );
  NAND4_X1 U16995 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15168) );
  XOR2_X1 U16996 ( .A(DATAI_7_), .B(keyinput_153), .Z(n15167) );
  XOR2_X1 U16997 ( .A(DATAI_6_), .B(keyinput_154), .Z(n15166) );
  AOI21_X1 U16998 ( .B1(n15168), .B2(n15167), .A(n15166), .ZN(n15172) );
  XNOR2_X1 U16999 ( .A(DATAI_5_), .B(keyinput_155), .ZN(n15171) );
  XOR2_X1 U17000 ( .A(DATAI_4_), .B(keyinput_156), .Z(n15170) );
  XOR2_X1 U17001 ( .A(DATAI_3_), .B(keyinput_157), .Z(n15169) );
  OAI211_X1 U17002 ( .C1(n15172), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        n15175) );
  XNOR2_X1 U17003 ( .A(DATAI_2_), .B(keyinput_158), .ZN(n15174) );
  XOR2_X1 U17004 ( .A(DATAI_1_), .B(keyinput_159), .Z(n15173) );
  AOI21_X1 U17005 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15188) );
  INV_X1 U17006 ( .A(READY1), .ZN(n15177) );
  INV_X1 U17007 ( .A(NA), .ZN(n22175) );
  OAI22_X1 U17008 ( .A1(n15177), .A2(keyinput_164), .B1(n22175), .B2(
        keyinput_162), .ZN(n15176) );
  AOI221_X1 U17009 ( .B1(n15177), .B2(keyinput_164), .C1(keyinput_162), .C2(
        n22175), .A(n15176), .ZN(n15178) );
  INV_X1 U17010 ( .A(n15178), .ZN(n15187) );
  OAI22_X1 U17011 ( .A1(READY2), .A2(keyinput_165), .B1(DATAI_0_), .B2(
        keyinput_160), .ZN(n15179) );
  AOI221_X1 U17012 ( .B1(READY2), .B2(keyinput_165), .C1(keyinput_160), .C2(
        DATAI_0_), .A(n15179), .ZN(n15185) );
  INV_X1 U17013 ( .A(keyinput_161), .ZN(n15180) );
  XNOR2_X1 U17014 ( .A(n15180), .B(HOLD), .ZN(n15184) );
  INV_X1 U17015 ( .A(keyinput_166), .ZN(n15181) );
  XNOR2_X1 U17016 ( .A(n15181), .B(P1_READREQUEST_REG_SCAN_IN), .ZN(n15183) );
  XNOR2_X1 U17017 ( .A(BS16), .B(keyinput_163), .ZN(n15182) );
  NAND4_X1 U17018 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15186) );
  NOR3_X1 U17019 ( .A1(n15188), .A2(n15187), .A3(n15186), .ZN(n15195) );
  XNOR2_X1 U17020 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_167), .ZN(n15194) );
  XOR2_X1 U17021 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_168), .Z(n15192)
         );
  XOR2_X1 U17022 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_169), .Z(n15191) );
  INV_X1 U17023 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20400) );
  XNOR2_X1 U17024 ( .A(n20400), .B(keyinput_170), .ZN(n15190) );
  XNOR2_X1 U17025 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_171), .ZN(
        n15189) );
  NOR4_X1 U17026 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15193) );
  OAI21_X1 U17027 ( .B1(n15195), .B2(n15194), .A(n15193), .ZN(n15199) );
  XNOR2_X1 U17028 ( .A(n22282), .B(keyinput_172), .ZN(n15198) );
  XNOR2_X1 U17029 ( .A(P1_MORE_REG_SCAN_IN), .B(keyinput_173), .ZN(n15197) );
  XNOR2_X1 U17030 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_174), .ZN(n15196) );
  AOI211_X1 U17031 ( .C1(n15199), .C2(n15198), .A(n15197), .B(n15196), .ZN(
        n15202) );
  XNOR2_X1 U17032 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_175), .ZN(n15201) );
  XNOR2_X1 U17033 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_176), .ZN(
        n15200) );
  NOR3_X1 U17034 ( .A1(n15202), .A2(n15201), .A3(n15200), .ZN(n15224) );
  XOR2_X1 U17035 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_180), .Z(n15223)
         );
  XOR2_X1 U17036 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_177), .Z(
        n15222) );
  INV_X1 U17037 ( .A(keyinput_179), .ZN(n15203) );
  NAND2_X1 U17038 ( .A1(n15203), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n15209) );
  AOI22_X1 U17039 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_187), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_184), .ZN(n15207) );
  INV_X1 U17040 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20278) );
  AOI22_X1 U17041 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_186), .B1(
        n20278), .B2(keyinput_178), .ZN(n15206) );
  INV_X1 U17042 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20252) );
  INV_X1 U17043 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20248) );
  AOI22_X1 U17044 ( .A1(n20252), .A2(keyinput_183), .B1(keyinput_185), .B2(
        n20248), .ZN(n15205) );
  INV_X1 U17045 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20262) );
  INV_X1 U17046 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20255) );
  AOI22_X1 U17047 ( .A1(n20262), .A2(keyinput_179), .B1(keyinput_182), .B2(
        n20255), .ZN(n15204) );
  AND4_X1 U17048 ( .A1(n15207), .A2(n15206), .A3(n15205), .A4(n15204), .ZN(
        n15208) );
  OAI211_X1 U17049 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(keyinput_186), .A(
        n15209), .B(n15208), .ZN(n15211) );
  OAI22_X1 U17050 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(keyinput_187), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_184), .ZN(n15210) );
  NOR2_X1 U17051 ( .A1(n15211), .A2(n15210), .ZN(n15220) );
  INV_X1 U17052 ( .A(keyinput_181), .ZN(n15212) );
  XNOR2_X1 U17053 ( .A(n15212), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n15219) );
  INV_X1 U17054 ( .A(keyinput_183), .ZN(n15214) );
  INV_X1 U17055 ( .A(keyinput_178), .ZN(n15213) );
  AOI22_X1 U17056 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n15214), .B1(n15213), 
        .B2(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n15218) );
  INV_X1 U17057 ( .A(keyinput_182), .ZN(n15216) );
  INV_X1 U17058 ( .A(keyinput_185), .ZN(n15215) );
  AOI22_X1 U17059 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n15216), .B1(n15215), 
        .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n15217) );
  NAND4_X1 U17060 ( .A1(n15220), .A2(n15219), .A3(n15218), .A4(n15217), .ZN(
        n15221) );
  NOR4_X1 U17061 ( .A1(n15224), .A2(n15223), .A3(n15222), .A4(n15221), .ZN(
        n15227) );
  XOR2_X1 U17062 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .Z(n15226)
         );
  XNOR2_X1 U17063 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .ZN(n15225)
         );
  OAI21_X1 U17064 ( .B1(n15227), .B2(n15226), .A(n15225), .ZN(n15229) );
  XNOR2_X1 U17065 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n15228)
         );
  NAND2_X1 U17066 ( .A1(n15229), .A2(n15228), .ZN(n15233) );
  XNOR2_X1 U17067 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_193), .ZN(n15232)
         );
  XNOR2_X1 U17068 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .ZN(n15231)
         );
  XNOR2_X1 U17069 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .ZN(n15230)
         );
  NAND4_X1 U17070 ( .A1(n15233), .A2(n15232), .A3(n15231), .A4(n15230), .ZN(
        n15236) );
  XNOR2_X1 U17071 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n15235)
         );
  XOR2_X1 U17072 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_195), .Z(n15234)
         );
  AOI21_X1 U17073 ( .B1(n15236), .B2(n15235), .A(n15234), .ZN(n15242) );
  INV_X1 U17074 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20231) );
  INV_X1 U17075 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21711) );
  AOI22_X1 U17076 ( .A1(n20231), .A2(keyinput_196), .B1(keyinput_198), .B2(
        n21711), .ZN(n15237) );
  OAI221_X1 U17077 ( .B1(n20231), .B2(keyinput_196), .C1(n21711), .C2(
        keyinput_198), .A(n15237), .ZN(n15241) );
  INV_X1 U17078 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21828) );
  AOI22_X1 U17079 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_200), .B1(
        n21828), .B2(keyinput_199), .ZN(n15238) );
  OAI221_X1 U17080 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_200), .C1(
        n21828), .C2(keyinput_199), .A(n15238), .ZN(n15240) );
  XNOR2_X1 U17081 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n15239)
         );
  NOR4_X1 U17082 ( .A1(n15242), .A2(n15241), .A3(n15240), .A4(n15239), .ZN(
        n15245) );
  XOR2_X1 U17083 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .Z(n15244)
         );
  XNOR2_X1 U17084 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .ZN(n15243)
         );
  OAI21_X1 U17085 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(n15251) );
  XOR2_X1 U17086 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .Z(n15247) );
  XOR2_X1 U17087 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_204), .Z(n15246) );
  NOR2_X1 U17088 ( .A1(n15247), .A2(n15246), .ZN(n15250) );
  XNOR2_X1 U17089 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .ZN(n15249)
         );
  XNOR2_X1 U17090 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_206), .ZN(n15248)
         );
  AOI211_X1 U17091 ( .C1(n15251), .C2(n15250), .A(n15249), .B(n15248), .ZN(
        n15255) );
  XNOR2_X1 U17092 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_207), .ZN(n15254)
         );
  XNOR2_X1 U17093 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_209), .ZN(n15253)
         );
  XNOR2_X1 U17094 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_208), .ZN(n15252)
         );
  OAI211_X1 U17095 ( .C1(n15255), .C2(n15254), .A(n15253), .B(n15252), .ZN(
        n15258) );
  XNOR2_X1 U17096 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_210), .ZN(n15257)
         );
  XNOR2_X1 U17097 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_211), .ZN(n15256)
         );
  NAND3_X1 U17098 ( .A1(n15258), .A2(n15257), .A3(n15256), .ZN(n15261) );
  XOR2_X1 U17099 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .Z(n15260) );
  INV_X1 U17100 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16162) );
  XNOR2_X1 U17101 ( .A(n16162), .B(keyinput_213), .ZN(n15259) );
  NAND3_X1 U17102 ( .A1(n15261), .A2(n15260), .A3(n15259), .ZN(n15267) );
  XOR2_X1 U17103 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_214), .Z(n15266) );
  INV_X1 U17104 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15885) );
  XNOR2_X1 U17105 ( .A(n15885), .B(keyinput_215), .ZN(n15264) );
  XNOR2_X1 U17106 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_217), .ZN(n15263)
         );
  XNOR2_X1 U17107 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_216), .ZN(n15262)
         );
  NAND3_X1 U17108 ( .A1(n15264), .A2(n15263), .A3(n15262), .ZN(n15265) );
  AOI21_X1 U17109 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15270) );
  INV_X1 U17110 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n22101) );
  XNOR2_X1 U17111 ( .A(n22101), .B(keyinput_219), .ZN(n15269) );
  XNOR2_X1 U17112 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .ZN(n15268)
         );
  NOR3_X1 U17113 ( .A1(n15270), .A2(n15269), .A3(n15268), .ZN(n15273) );
  INV_X1 U17114 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n22089) );
  XNOR2_X1 U17115 ( .A(n22089), .B(keyinput_220), .ZN(n15272) );
  XNOR2_X1 U17116 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_221), .ZN(n15271)
         );
  NOR3_X1 U17117 ( .A1(n15273), .A2(n15272), .A3(n15271), .ZN(n15280) );
  XOR2_X1 U17118 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_222), .Z(n15279) );
  XOR2_X1 U17119 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .Z(n15277) );
  XOR2_X1 U17120 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_225), .Z(n15276) );
  INV_X1 U17121 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n22058) );
  XNOR2_X1 U17122 ( .A(n22058), .B(keyinput_223), .ZN(n15275) );
  XNOR2_X1 U17123 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .ZN(n15274)
         );
  NOR4_X1 U17124 ( .A1(n15277), .A2(n15276), .A3(n15275), .A4(n15274), .ZN(
        n15278) );
  OAI21_X1 U17125 ( .B1(n15280), .B2(n15279), .A(n15278), .ZN(n15283) );
  XOR2_X1 U17126 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_227), .Z(n15282) );
  XNOR2_X1 U17127 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_228), .ZN(n15281)
         );
  NAND3_X1 U17128 ( .A1(n15283), .A2(n15282), .A3(n15281), .ZN(n15286) );
  INV_X1 U17129 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n16206) );
  XNOR2_X1 U17130 ( .A(n16206), .B(keyinput_229), .ZN(n15285) );
  XNOR2_X1 U17131 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_230), .ZN(n15284)
         );
  NAND3_X1 U17132 ( .A1(n15286), .A2(n15285), .A3(n15284), .ZN(n15293) );
  XOR2_X1 U17133 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .Z(n15290) );
  INV_X1 U17134 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16218) );
  XNOR2_X1 U17135 ( .A(n16218), .B(keyinput_231), .ZN(n15289) );
  XNOR2_X1 U17136 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_233), .ZN(n15288)
         );
  XNOR2_X1 U17137 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n15287)
         );
  NOR4_X1 U17138 ( .A1(n15290), .A2(n15289), .A3(n15288), .A4(n15287), .ZN(
        n15292) );
  XOR2_X1 U17139 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .Z(n15291) );
  AOI21_X1 U17140 ( .B1(n15293), .B2(n15292), .A(n15291), .ZN(n15300) );
  XNOR2_X1 U17141 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .ZN(n15299)
         );
  XNOR2_X1 U17142 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n15297)
         );
  XNOR2_X1 U17143 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n15296)
         );
  XNOR2_X1 U17144 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_237), .ZN(n15295)
         );
  XNOR2_X1 U17145 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n15294)
         );
  NOR4_X1 U17146 ( .A1(n15297), .A2(n15296), .A3(n15295), .A4(n15294), .ZN(
        n15298) );
  OAI21_X1 U17147 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15303) );
  XNOR2_X1 U17148 ( .A(n15490), .B(keyinput_241), .ZN(n15302) );
  XNOR2_X1 U17149 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .ZN(n15301)
         );
  AOI21_X1 U17150 ( .B1(n15303), .B2(n15302), .A(n15301), .ZN(n15306) );
  XOR2_X1 U17151 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .Z(n15305) );
  XNOR2_X1 U17152 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .ZN(n15304)
         );
  NOR3_X1 U17153 ( .A1(n15306), .A2(n15305), .A3(n15304), .ZN(n15313) );
  XOR2_X1 U17154 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .Z(n15310) );
  XOR2_X1 U17155 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .Z(n15309) );
  XNOR2_X1 U17156 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .ZN(n15308)
         );
  XNOR2_X1 U17157 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n15307)
         );
  NAND4_X1 U17158 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15312) );
  XNOR2_X1 U17159 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n15311)
         );
  OAI21_X1 U17160 ( .B1(n15313), .B2(n15312), .A(n15311), .ZN(n15319) );
  XOR2_X1 U17161 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .Z(n15318) );
  XOR2_X1 U17162 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .Z(n15316) );
  XNOR2_X1 U17163 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .ZN(n15315)
         );
  XNOR2_X1 U17164 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .ZN(n15314)
         );
  NAND3_X1 U17165 ( .A1(n15316), .A2(n15315), .A3(n15314), .ZN(n15317) );
  AOI21_X1 U17166 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(n15516) );
  XOR2_X1 U17167 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .Z(n15515) );
  XNOR2_X1 U17168 ( .A(n15817), .B(keyinput_1), .ZN(n15322) );
  XOR2_X1 U17169 ( .A(keyinput_0), .B(P1_MEMORYFETCH_REG_SCAN_IN), .Z(n15321)
         );
  XNOR2_X1 U17170 ( .A(n16223), .B(keyinput_2), .ZN(n15320) );
  AOI21_X1 U17171 ( .B1(n15322), .B2(n15321), .A(n15320), .ZN(n15326) );
  XOR2_X1 U17172 ( .A(DATAI_28_), .B(keyinput_4), .Z(n15325) );
  XNOR2_X1 U17173 ( .A(DATAI_29_), .B(keyinput_3), .ZN(n15324) );
  XNOR2_X1 U17174 ( .A(DATAI_27_), .B(keyinput_5), .ZN(n15323) );
  NOR4_X1 U17175 ( .A1(n15326), .A2(n15325), .A3(n15324), .A4(n15323), .ZN(
        n15329) );
  XNOR2_X1 U17176 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n15328) );
  XOR2_X1 U17177 ( .A(DATAI_25_), .B(keyinput_7), .Z(n15327) );
  OAI21_X1 U17178 ( .B1(n15329), .B2(n15328), .A(n15327), .ZN(n15335) );
  XOR2_X1 U17179 ( .A(keyinput_8), .B(DATAI_24_), .Z(n15334) );
  XOR2_X1 U17180 ( .A(keyinput_9), .B(DATAI_23_), .Z(n15332) );
  XOR2_X1 U17181 ( .A(keyinput_11), .B(DATAI_21_), .Z(n15331) );
  INV_X1 U17182 ( .A(DATAI_22_), .ZN(n22227) );
  XNOR2_X1 U17183 ( .A(n22227), .B(keyinput_10), .ZN(n15330) );
  NAND3_X1 U17184 ( .A1(n15332), .A2(n15331), .A3(n15330), .ZN(n15333) );
  AOI21_X1 U17185 ( .B1(n15335), .B2(n15334), .A(n15333), .ZN(n15339) );
  XOR2_X1 U17186 ( .A(keyinput_13), .B(DATAI_19_), .Z(n15338) );
  XOR2_X1 U17187 ( .A(DATAI_20_), .B(keyinput_12), .Z(n15337) );
  XNOR2_X1 U17188 ( .A(keyinput_14), .B(DATAI_18_), .ZN(n15336) );
  NOR4_X1 U17189 ( .A1(n15339), .A2(n15338), .A3(n15337), .A4(n15336), .ZN(
        n15342) );
  XNOR2_X1 U17190 ( .A(keyinput_15), .B(DATAI_17_), .ZN(n15341) );
  XNOR2_X1 U17191 ( .A(keyinput_16), .B(DATAI_16_), .ZN(n15340) );
  OAI21_X1 U17192 ( .B1(n15342), .B2(n15341), .A(n15340), .ZN(n15348) );
  XNOR2_X1 U17193 ( .A(n15343), .B(keyinput_17), .ZN(n15347) );
  XNOR2_X1 U17194 ( .A(n15344), .B(keyinput_18), .ZN(n15346) );
  XNOR2_X1 U17195 ( .A(DATAI_13_), .B(keyinput_19), .ZN(n15345) );
  AOI211_X1 U17196 ( .C1(n15348), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15353) );
  XNOR2_X1 U17197 ( .A(n15349), .B(keyinput_20), .ZN(n15352) );
  XNOR2_X1 U17198 ( .A(n15350), .B(keyinput_21), .ZN(n15351) );
  OAI21_X1 U17199 ( .B1(n15353), .B2(n15352), .A(n15351), .ZN(n15357) );
  XNOR2_X1 U17200 ( .A(DATAI_9_), .B(keyinput_23), .ZN(n15356) );
  XNOR2_X1 U17201 ( .A(DATAI_10_), .B(keyinput_22), .ZN(n15355) );
  XNOR2_X1 U17202 ( .A(keyinput_24), .B(DATAI_8_), .ZN(n15354) );
  NAND4_X1 U17203 ( .A1(n15357), .A2(n15356), .A3(n15355), .A4(n15354), .ZN(
        n15360) );
  XOR2_X1 U17204 ( .A(keyinput_25), .B(DATAI_7_), .Z(n15359) );
  XNOR2_X1 U17205 ( .A(keyinput_26), .B(DATAI_6_), .ZN(n15358) );
  AOI21_X1 U17206 ( .B1(n15360), .B2(n15359), .A(n15358), .ZN(n15364) );
  XOR2_X1 U17207 ( .A(keyinput_27), .B(DATAI_5_), .Z(n15363) );
  XOR2_X1 U17208 ( .A(DATAI_4_), .B(keyinput_28), .Z(n15362) );
  XNOR2_X1 U17209 ( .A(keyinput_29), .B(DATAI_3_), .ZN(n15361) );
  OAI211_X1 U17210 ( .C1(n15364), .C2(n15363), .A(n15362), .B(n15361), .ZN(
        n15368) );
  XNOR2_X1 U17211 ( .A(n15365), .B(keyinput_30), .ZN(n15367) );
  XNOR2_X1 U17212 ( .A(keyinput_31), .B(DATAI_1_), .ZN(n15366) );
  AOI21_X1 U17213 ( .B1(n15368), .B2(n15367), .A(n15366), .ZN(n15379) );
  AOI22_X1 U17214 ( .A1(keyinput_32), .A2(DATAI_0_), .B1(n22175), .B2(
        keyinput_34), .ZN(n15369) );
  OAI221_X1 U17215 ( .B1(keyinput_32), .B2(DATAI_0_), .C1(n22175), .C2(
        keyinput_34), .A(n15369), .ZN(n15378) );
  INV_X1 U17216 ( .A(READY2), .ZN(n15372) );
  INV_X1 U17217 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n15371) );
  AOI22_X1 U17218 ( .A1(n15372), .A2(keyinput_37), .B1(keyinput_38), .B2(
        n15371), .ZN(n15370) );
  OAI221_X1 U17219 ( .B1(n15372), .B2(keyinput_37), .C1(n15371), .C2(
        keyinput_38), .A(n15370), .ZN(n15377) );
  XOR2_X1 U17220 ( .A(keyinput_35), .B(BS16), .Z(n15375) );
  XOR2_X1 U17221 ( .A(HOLD), .B(keyinput_33), .Z(n15374) );
  XOR2_X1 U17222 ( .A(READY1), .B(keyinput_36), .Z(n15373) );
  NAND3_X1 U17223 ( .A1(n15375), .A2(n15374), .A3(n15373), .ZN(n15376) );
  NOR4_X1 U17224 ( .A1(n15379), .A2(n15378), .A3(n15377), .A4(n15376), .ZN(
        n15386) );
  XOR2_X1 U17225 ( .A(P1_ADS_N_REG_SCAN_IN), .B(keyinput_39), .Z(n15385) );
  XOR2_X1 U17226 ( .A(keyinput_41), .B(P1_M_IO_N_REG_SCAN_IN), .Z(n15383) );
  XOR2_X1 U17227 ( .A(keyinput_43), .B(P1_REQUESTPENDING_REG_SCAN_IN), .Z(
        n15382) );
  XNOR2_X1 U17228 ( .A(n20400), .B(keyinput_42), .ZN(n15381) );
  XNOR2_X1 U17229 ( .A(keyinput_40), .B(P1_CODEFETCH_REG_SCAN_IN), .ZN(n15380)
         );
  NOR4_X1 U17230 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15384) );
  OAI21_X1 U17231 ( .B1(n15386), .B2(n15385), .A(n15384), .ZN(n15390) );
  XNOR2_X1 U17232 ( .A(P1_STATEBS16_REG_SCAN_IN), .B(keyinput_44), .ZN(n15389)
         );
  XNOR2_X1 U17233 ( .A(keyinput_46), .B(P1_FLUSH_REG_SCAN_IN), .ZN(n15388) );
  XNOR2_X1 U17234 ( .A(keyinput_45), .B(P1_MORE_REG_SCAN_IN), .ZN(n15387) );
  AOI211_X1 U17235 ( .C1(n15390), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15393) );
  XOR2_X1 U17236 ( .A(keyinput_47), .B(P1_W_R_N_REG_SCAN_IN), .Z(n15392) );
  XNOR2_X1 U17237 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .ZN(
        n15391) );
  NOR3_X1 U17238 ( .A1(n15393), .A2(n15392), .A3(n15391), .ZN(n15415) );
  INV_X1 U17239 ( .A(keyinput_50), .ZN(n15395) );
  INV_X1 U17240 ( .A(keyinput_51), .ZN(n15394) );
  OAI22_X1 U17241 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(n15395), .B1(n15394), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n15409) );
  INV_X1 U17242 ( .A(keyinput_59), .ZN(n15403) );
  AOI22_X1 U17243 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_57), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .ZN(n15402) );
  INV_X1 U17244 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20259) );
  OAI22_X1 U17245 ( .A1(n20259), .A2(keyinput_53), .B1(n20278), .B2(
        keyinput_50), .ZN(n15399) );
  OAI22_X1 U17246 ( .A1(n20262), .A2(keyinput_51), .B1(n20255), .B2(
        keyinput_54), .ZN(n15398) );
  OAI22_X1 U17247 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_57), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .ZN(n15397) );
  INV_X1 U17248 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n22103) );
  OAI22_X1 U17249 ( .A1(n22103), .A2(keyinput_59), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_49), .ZN(n15396) );
  OR4_X1 U17250 ( .A1(n15399), .A2(n15398), .A3(n15397), .A4(n15396), .ZN(
        n15400) );
  AOI21_X1 U17251 ( .B1(keyinput_49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), .A(
        n15400), .ZN(n15401) );
  OAI211_X1 U17252 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n15403), .A(n15402), 
        .B(n15401), .ZN(n15408) );
  INV_X1 U17253 ( .A(keyinput_54), .ZN(n15405) );
  INV_X1 U17254 ( .A(keyinput_53), .ZN(n15404) );
  OAI22_X1 U17255 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n15405), .B1(n15404), 
        .B2(P1_REIP_REG_30__SCAN_IN), .ZN(n15407) );
  XNOR2_X1 U17256 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .ZN(n15406)
         );
  NOR4_X1 U17257 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15412) );
  XOR2_X1 U17258 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .Z(n15411) );
  XNOR2_X1 U17259 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .ZN(n15410)
         );
  NAND3_X1 U17260 ( .A1(n15412), .A2(n15411), .A3(n15410), .ZN(n15414) );
  XNOR2_X1 U17261 ( .A(keyinput_60), .B(P1_REIP_REG_23__SCAN_IN), .ZN(n15413)
         );
  OAI21_X1 U17262 ( .B1(n15415), .B2(n15414), .A(n15413), .ZN(n15418) );
  XOR2_X1 U17263 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_61), .Z(n15417) );
  XNOR2_X1 U17264 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .ZN(n15416)
         );
  AOI21_X1 U17265 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15422) );
  XOR2_X1 U17266 ( .A(keyinput_64), .B(P1_REIP_REG_19__SCAN_IN), .Z(n15421) );
  XOR2_X1 U17267 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_65), .Z(n15420) );
  XNOR2_X1 U17268 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .ZN(n15419)
         );
  NOR4_X1 U17269 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15425) );
  XNOR2_X1 U17270 ( .A(keyinput_66), .B(P1_REIP_REG_17__SCAN_IN), .ZN(n15424)
         );
  XNOR2_X1 U17271 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .ZN(n15423)
         );
  OAI21_X1 U17272 ( .B1(n15425), .B2(n15424), .A(n15423), .ZN(n15431) );
  OAI22_X1 U17273 ( .A1(n21711), .A2(keyinput_70), .B1(P1_REIP_REG_12__SCAN_IN), .B2(keyinput_71), .ZN(n15426) );
  AOI221_X1 U17274 ( .B1(n21711), .B2(keyinput_70), .C1(keyinput_71), .C2(
        P1_REIP_REG_12__SCAN_IN), .A(n15426), .ZN(n15430) );
  XOR2_X1 U17275 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_68), .Z(n15429) );
  INV_X1 U17276 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21721) );
  OAI22_X1 U17277 ( .A1(n21721), .A2(keyinput_69), .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_72), .ZN(n15427) );
  AOI221_X1 U17278 ( .B1(n21721), .B2(keyinput_69), .C1(keyinput_72), .C2(
        P1_REIP_REG_11__SCAN_IN), .A(n15427), .ZN(n15428) );
  NAND4_X1 U17279 ( .A1(n15431), .A2(n15430), .A3(n15429), .A4(n15428), .ZN(
        n15434) );
  XNOR2_X1 U17280 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .ZN(n15433)
         );
  XNOR2_X1 U17281 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .ZN(n15432)
         );
  AOI21_X1 U17282 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15437) );
  XOR2_X1 U17283 ( .A(keyinput_76), .B(P1_REIP_REG_7__SCAN_IN), .Z(n15436) );
  XOR2_X1 U17284 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .Z(n15435) );
  NOR3_X1 U17285 ( .A1(n15437), .A2(n15436), .A3(n15435), .ZN(n15440) );
  XOR2_X1 U17286 ( .A(keyinput_77), .B(P1_REIP_REG_6__SCAN_IN), .Z(n15439) );
  XOR2_X1 U17287 ( .A(keyinput_78), .B(P1_REIP_REG_5__SCAN_IN), .Z(n15438) );
  NOR3_X1 U17288 ( .A1(n15440), .A2(n15439), .A3(n15438), .ZN(n15444) );
  XOR2_X1 U17289 ( .A(keyinput_79), .B(P1_REIP_REG_4__SCAN_IN), .Z(n15443) );
  XOR2_X1 U17290 ( .A(keyinput_80), .B(P1_REIP_REG_3__SCAN_IN), .Z(n15442) );
  XOR2_X1 U17291 ( .A(keyinput_81), .B(P1_REIP_REG_2__SCAN_IN), .Z(n15441) );
  OAI211_X1 U17292 ( .C1(n15444), .C2(n15443), .A(n15442), .B(n15441), .ZN(
        n15447) );
  XOR2_X1 U17293 ( .A(keyinput_82), .B(P1_REIP_REG_1__SCAN_IN), .Z(n15446) );
  XNOR2_X1 U17294 ( .A(keyinput_83), .B(P1_REIP_REG_0__SCAN_IN), .ZN(n15445)
         );
  NAND3_X1 U17295 ( .A1(n15447), .A2(n15446), .A3(n15445), .ZN(n15450) );
  XOR2_X1 U17296 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .Z(n15449) );
  XNOR2_X1 U17297 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .ZN(n15448)
         );
  NAND3_X1 U17298 ( .A1(n15450), .A2(n15449), .A3(n15448), .ZN(n15456) );
  XOR2_X1 U17299 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .Z(n15455) );
  XOR2_X1 U17300 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_88), .Z(n15453) );
  XNOR2_X1 U17301 ( .A(n15885), .B(keyinput_87), .ZN(n15452) );
  XNOR2_X1 U17302 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .ZN(n15451)
         );
  NAND3_X1 U17303 ( .A1(n15453), .A2(n15452), .A3(n15451), .ZN(n15454) );
  AOI21_X1 U17304 ( .B1(n15456), .B2(n15455), .A(n15454), .ZN(n15459) );
  XOR2_X1 U17305 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n15458) );
  XNOR2_X1 U17306 ( .A(n22101), .B(keyinput_91), .ZN(n15457) );
  NOR3_X1 U17307 ( .A1(n15459), .A2(n15458), .A3(n15457), .ZN(n15462) );
  XNOR2_X1 U17308 ( .A(n22089), .B(keyinput_92), .ZN(n15461) );
  XNOR2_X1 U17309 ( .A(P1_EBX_REG_22__SCAN_IN), .B(keyinput_93), .ZN(n15460)
         );
  NOR3_X1 U17310 ( .A1(n15462), .A2(n15461), .A3(n15460), .ZN(n15469) );
  XOR2_X1 U17311 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .Z(n15468) );
  XOR2_X1 U17312 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .Z(n15466) );
  XNOR2_X1 U17313 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .ZN(n15465)
         );
  XNOR2_X1 U17314 ( .A(P1_EBX_REG_18__SCAN_IN), .B(keyinput_97), .ZN(n15464)
         );
  XNOR2_X1 U17315 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_96), .ZN(n15463)
         );
  NOR4_X1 U17316 ( .A1(n15466), .A2(n15465), .A3(n15464), .A4(n15463), .ZN(
        n15467) );
  OAI21_X1 U17317 ( .B1(n15469), .B2(n15468), .A(n15467), .ZN(n15472) );
  XOR2_X1 U17318 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .Z(n15471) );
  XNOR2_X1 U17319 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_100), .ZN(n15470)
         );
  NAND3_X1 U17320 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n15475) );
  XOR2_X1 U17321 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .Z(n15474) );
  XNOR2_X1 U17322 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n15473)
         );
  NAND3_X1 U17323 ( .A1(n15475), .A2(n15474), .A3(n15473), .ZN(n15482) );
  XNOR2_X1 U17324 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n15479)
         );
  XNOR2_X1 U17325 ( .A(keyinput_105), .B(P1_EBX_REG_10__SCAN_IN), .ZN(n15478)
         );
  XNOR2_X1 U17326 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .ZN(n15477)
         );
  XNOR2_X1 U17327 ( .A(P1_EBX_REG_12__SCAN_IN), .B(keyinput_103), .ZN(n15476)
         );
  NOR4_X1 U17328 ( .A1(n15479), .A2(n15478), .A3(n15477), .A4(n15476), .ZN(
        n15481) );
  XOR2_X1 U17329 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .Z(n15480) );
  AOI21_X1 U17330 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15489) );
  XNOR2_X1 U17331 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .ZN(n15488)
         );
  INV_X1 U17332 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20325) );
  XNOR2_X1 U17333 ( .A(n20325), .B(keyinput_111), .ZN(n15486) );
  XNOR2_X1 U17334 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .ZN(n15485)
         );
  XNOR2_X1 U17335 ( .A(n20319), .B(keyinput_110), .ZN(n15484) );
  XNOR2_X1 U17336 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .ZN(n15483)
         );
  NOR4_X1 U17337 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        n15487) );
  OAI21_X1 U17338 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15493) );
  XNOR2_X1 U17339 ( .A(n15490), .B(keyinput_113), .ZN(n15492) );
  XNOR2_X1 U17340 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .ZN(n15491)
         );
  AOI21_X1 U17341 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n15496) );
  XOR2_X1 U17342 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .Z(n15495) );
  XOR2_X1 U17343 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .Z(n15494) );
  NOR3_X1 U17344 ( .A1(n15496), .A2(n15495), .A3(n15494), .ZN(n15503) );
  XOR2_X1 U17345 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .Z(n15500) );
  XOR2_X1 U17346 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_120), .Z(n15499) );
  XNOR2_X1 U17347 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .ZN(n15498)
         );
  XNOR2_X1 U17348 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n15497)
         );
  NAND4_X1 U17349 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15502) );
  XOR2_X1 U17350 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_121), .Z(n15501) );
  OAI21_X1 U17351 ( .B1(n15503), .B2(n15502), .A(n15501), .ZN(n15509) );
  XNOR2_X1 U17352 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_122), .ZN(n15508)
         );
  XOR2_X1 U17353 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_123), .Z(n15506) );
  XNOR2_X1 U17354 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .ZN(n15505)
         );
  XNOR2_X1 U17355 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .ZN(n15504)
         );
  NAND3_X1 U17356 ( .A1(n15506), .A2(n15505), .A3(n15504), .ZN(n15507) );
  AOI21_X1 U17357 ( .B1(n15509), .B2(n15508), .A(n15507), .ZN(n15512) );
  XNOR2_X1 U17358 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n15511)
         );
  XNOR2_X1 U17359 ( .A(keyinput_255), .B(keyinput_127), .ZN(n15510) );
  OAI21_X1 U17360 ( .B1(n15512), .B2(n15511), .A(n15510), .ZN(n15514) );
  XNOR2_X1 U17361 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n15513)
         );
  OAI211_X1 U17362 ( .C1(n15516), .C2(n15515), .A(n15514), .B(n15513), .ZN(
        n15537) );
  NAND2_X1 U17363 ( .A1(n15517), .A2(n13253), .ZN(n22275) );
  OR2_X1 U17364 ( .A1(n22275), .A2(n15519), .ZN(n15526) );
  NOR3_X1 U17365 ( .A1(n22654), .A2(n22660), .A3(n22358), .ZN(n15520) );
  NOR2_X1 U17366 ( .A1(n22358), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22337) );
  NOR2_X1 U17367 ( .A1(n15520), .A2(n22337), .ZN(n15533) );
  INV_X1 U17368 ( .A(n15533), .ZN(n15523) );
  INV_X1 U17369 ( .A(n16514), .ZN(n15521) );
  OR2_X1 U17370 ( .A1(n17360), .A2(n15521), .ZN(n22250) );
  NOR2_X1 U17371 ( .A1(n22250), .A2(n22339), .ZN(n15532) );
  AND2_X1 U17372 ( .A1(n15528), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22325) );
  OR2_X1 U17373 ( .A1(n22323), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22300) );
  INV_X1 U17374 ( .A(n22300), .ZN(n15522) );
  AOI22_X1 U17375 ( .A1(n15523), .A2(n15532), .B1(n22325), .B2(n15522), .ZN(
        n22658) );
  NAND2_X1 U17376 ( .A1(n22632), .A2(n22223), .ZN(n22623) );
  AOI22_X1 U17377 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n22635), .B1(DATAI_30_), 
        .B2(n22636), .ZN(n22630) );
  INV_X1 U17378 ( .A(n22630), .ZN(n22618) );
  AOI22_X1 U17379 ( .A1(DATAI_22_), .A2(n22636), .B1(n22635), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n22621) );
  NAND2_X1 U17380 ( .A1(n15525), .A2(n15524), .ZN(n22625) );
  NOR3_X1 U17381 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(n22238), .ZN(n22273) );
  NAND2_X1 U17382 ( .A1(n22273), .A2(n22251), .ZN(n22260) );
  OAI22_X1 U17383 ( .A1(n22621), .A2(n15526), .B1(n22625), .B2(n22260), .ZN(
        n15527) );
  AOI21_X1 U17384 ( .B1(n22654), .B2(n22618), .A(n15527), .ZN(n15535) );
  NAND2_X1 U17385 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22300), .ZN(n22297) );
  INV_X1 U17386 ( .A(n22297), .ZN(n15530) );
  INV_X1 U17387 ( .A(n15528), .ZN(n15529) );
  NAND2_X1 U17388 ( .A1(n15529), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22356) );
  INV_X1 U17389 ( .A(n22314), .ZN(n22329) );
  AOI211_X1 U17390 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22260), .A(n15530), 
        .B(n22329), .ZN(n15531) );
  OAI21_X1 U17391 ( .B1(n15533), .B2(n15532), .A(n15531), .ZN(n22655) );
  NAND2_X1 U17392 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n15534) );
  OAI211_X1 U17393 ( .C1(n22658), .C2(n22623), .A(n15535), .B(n15534), .ZN(
        n15536) );
  XNOR2_X1 U17394 ( .A(n15537), .B(n15536), .ZN(P1_U3055) );
  INV_X1 U17395 ( .A(n18653), .ZN(n18666) );
  NOR2_X1 U17396 ( .A1(n18809), .A2(n15538), .ZN(n15671) );
  XNOR2_X1 U17397 ( .A(n15671), .B(n15539), .ZN(n15540) );
  NAND2_X1 U17398 ( .A1(n15540), .A2(n18980), .ZN(n15548) );
  INV_X1 U17399 ( .A(n18951), .ZN(n18884) );
  INV_X1 U17400 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17549) );
  INV_X1 U17401 ( .A(n18954), .ZN(n18968) );
  OAI22_X1 U17402 ( .A1(n15541), .A2(n18922), .B1(n17549), .B2(n18968), .ZN(
        n15544) );
  NOR2_X1 U17403 ( .A1(n18969), .A2(n15542), .ZN(n15543) );
  AOI211_X1 U17404 ( .C1(n18955), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15544), .B(n15543), .ZN(n15545) );
  OAI21_X1 U17405 ( .B1(n18884), .B2(n12429), .A(n15545), .ZN(n15546) );
  AOI21_X1 U17406 ( .B1(n18957), .B2(n12484), .A(n15546), .ZN(n15547) );
  OAI211_X1 U17407 ( .C1(n17481), .C2(n18666), .A(n15548), .B(n15547), .ZN(
        P2_U2853) );
  OAI222_X1 U17408 ( .A1(n15550), .A2(n16278), .B1(n20196), .B2(n16279), .C1(
        n15549), .C2(n16281), .ZN(P1_U2896) );
  OAI211_X1 U17409 ( .C1(n15098), .C2(n15552), .A(n15551), .B(n16596), .ZN(
        n15557) );
  AND2_X1 U17410 ( .A1(n15554), .A2(n15553), .ZN(n15555) );
  OR2_X1 U17411 ( .A1(n15555), .A2(n11252), .ZN(n16857) );
  INV_X1 U17412 ( .A(n16857), .ZN(n18801) );
  NAND2_X1 U17413 ( .A1(n18801), .A2(n16571), .ZN(n15556) );
  OAI211_X1 U17414 ( .C1(n16571), .C2(n12440), .A(n15557), .B(n15556), .ZN(
        P2_U2872) );
  INV_X1 U17415 ( .A(n22339), .ZN(n22354) );
  OAI22_X1 U17416 ( .A1(n15559), .A2(n22100), .B1(n15558), .B2(n22111), .ZN(
        n15561) );
  NOR2_X1 U17417 ( .A1(n22069), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15560) );
  AOI211_X1 U17418 ( .C1(n22354), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15563) );
  OAI21_X1 U17419 ( .B1(n22050), .B2(n20275), .A(n15563), .ZN(n15565) );
  NOR2_X1 U17420 ( .A1(n22096), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15564) );
  AOI211_X1 U17421 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15565), .B(n15564), .ZN(n15566) );
  OAI21_X1 U17422 ( .B1(n15568), .B2(n15567), .A(n15566), .ZN(P1_U2839) );
  AOI22_X1 U17423 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20208), .B1(n20194), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15569) );
  OAI21_X1 U17424 ( .B1(n15570), .B2(n15612), .A(n15569), .ZN(P1_U2920) );
  NOR2_X1 U17425 ( .A1(n15119), .A2(n15572), .ZN(n15573) );
  OR2_X1 U17426 ( .A1(n15571), .A2(n15573), .ZN(n15735) );
  AOI22_X1 U17427 ( .A1(n16274), .A2(n16249), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n22375), .ZN(n15574) );
  OAI21_X1 U17428 ( .B1(n15735), .B2(n16281), .A(n15574), .ZN(P1_U2895) );
  NAND2_X1 U17429 ( .A1(n15551), .A2(n15576), .ZN(n15577) );
  NAND2_X1 U17430 ( .A1(n15575), .A2(n15577), .ZN(n15628) );
  NAND2_X1 U17431 ( .A1(n16604), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15581) );
  OR2_X1 U17432 ( .A1(n11252), .A2(n15578), .ZN(n15579) );
  NAND2_X1 U17433 ( .A1(n15713), .A2(n15579), .ZN(n18813) );
  OR2_X1 U17434 ( .A1(n18813), .A2(n16604), .ZN(n15580) );
  OAI211_X1 U17435 ( .C1(n15628), .C2(n16606), .A(n15581), .B(n15580), .ZN(
        P2_U2871) );
  AOI22_X1 U17436 ( .A1(n20194), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15582) );
  OAI21_X1 U17437 ( .B1(n15583), .B2(n15612), .A(n15582), .ZN(P1_U2913) );
  INV_X1 U17438 ( .A(n15868), .ZN(n15879) );
  MUX2_X1 U17439 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n15584) );
  NAND2_X1 U17440 ( .A1(n15584), .A2(n11691), .ZN(n15683) );
  XNOR2_X1 U17441 ( .A(n15684), .B(n15683), .ZN(n21804) );
  AOI22_X1 U17442 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15585), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n22061), .ZN(n15586) );
  INV_X1 U17443 ( .A(n22044), .ZN(n22023) );
  OAI211_X1 U17444 ( .C1(n21804), .C2(n22111), .A(n15586), .B(n22023), .ZN(
        n15589) );
  INV_X1 U17445 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15637) );
  OR4_X1 U17446 ( .A1(n21977), .A2(n20223), .A3(n21981), .A4(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15587) );
  OAI21_X1 U17447 ( .B1(n22100), .B2(n15637), .A(n15587), .ZN(n15588) );
  AOI211_X1 U17448 ( .C1(n15732), .C2(n22107), .A(n15589), .B(n15588), .ZN(
        n15590) );
  OAI21_X1 U17449 ( .B1(n22052), .B2(n15735), .A(n15590), .ZN(P1_U2831) );
  AOI22_X1 U17450 ( .A1(n21698), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15591) );
  OAI21_X1 U17451 ( .B1(n15592), .B2(n15612), .A(n15591), .ZN(P1_U2912) );
  AOI22_X1 U17452 ( .A1(n21698), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15593) );
  OAI21_X1 U17453 ( .B1(n15594), .B2(n15612), .A(n15593), .ZN(P1_U2916) );
  AOI22_X1 U17454 ( .A1(n21698), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15595) );
  OAI21_X1 U17455 ( .B1(n15596), .B2(n15612), .A(n15595), .ZN(P1_U2911) );
  AOI22_X1 U17456 ( .A1(n21698), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15597) );
  OAI21_X1 U17457 ( .B1(n15598), .B2(n15612), .A(n15597), .ZN(P1_U2915) );
  AOI22_X1 U17458 ( .A1(n21698), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15599) );
  OAI21_X1 U17459 ( .B1(n15600), .B2(n15612), .A(n15599), .ZN(P1_U2910) );
  AOI22_X1 U17460 ( .A1(n21698), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15601) );
  OAI21_X1 U17461 ( .B1(n15602), .B2(n15612), .A(n15601), .ZN(P1_U2907) );
  AOI22_X1 U17462 ( .A1(n21698), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15603) );
  OAI21_X1 U17463 ( .B1(n15604), .B2(n15612), .A(n15603), .ZN(P1_U2908) );
  AOI22_X1 U17464 ( .A1(n21698), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15605) );
  OAI21_X1 U17465 ( .B1(n15606), .B2(n15612), .A(n15605), .ZN(P1_U2906) );
  AOI22_X1 U17466 ( .A1(n21698), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15607) );
  OAI21_X1 U17467 ( .B1(n15608), .B2(n15612), .A(n15607), .ZN(P1_U2914) );
  AOI22_X1 U17468 ( .A1(n21698), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15609) );
  OAI21_X1 U17469 ( .B1(n15610), .B2(n15612), .A(n15609), .ZN(P1_U2917) );
  AOI22_X1 U17470 ( .A1(n21698), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15611) );
  OAI21_X1 U17471 ( .B1(n15613), .B2(n15612), .A(n15611), .ZN(P1_U2909) );
  NAND2_X1 U17472 ( .A1(n15615), .A2(n15614), .ZN(n15616) );
  NAND2_X1 U17473 ( .A1(n15719), .A2(n15616), .ZN(n18812) );
  NAND2_X1 U17474 ( .A1(n11881), .A2(n15617), .ZN(n15618) );
  NOR2_X1 U17475 ( .A1(n19905), .A2(n15618), .ZN(n15623) );
  NAND2_X1 U17476 ( .A1(n19770), .A2(n11856), .ZN(n16694) );
  OAI22_X1 U17477 ( .A1(n16694), .A2(n20006), .B1(n15620), .B2(n19770), .ZN(
        n15621) );
  AOI21_X1 U17478 ( .B1(n19908), .B2(BUF1_REG_16__SCAN_IN), .A(n15621), .ZN(
        n15625) );
  AND2_X1 U17479 ( .A1(n15623), .A2(n15622), .ZN(n19909) );
  NAND2_X1 U17480 ( .A1(n19909), .A2(BUF2_REG_16__SCAN_IN), .ZN(n15624) );
  OAI211_X1 U17481 ( .C1(n18812), .C2(n19912), .A(n15625), .B(n15624), .ZN(
        n15626) );
  INV_X1 U17482 ( .A(n15626), .ZN(n15627) );
  OAI21_X1 U17483 ( .B1(n19911), .B2(n15628), .A(n15627), .ZN(P2_U2903) );
  AOI22_X1 U17484 ( .A1(n11739), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n17342), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n15629) );
  OAI21_X1 U17485 ( .B1(n15630), .B2(n19054), .A(n15629), .ZN(n18988) );
  INV_X1 U17486 ( .A(n18988), .ZN(n15938) );
  OAI21_X1 U17487 ( .B1(n15631), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n14913), 
        .ZN(n15634) );
  INV_X1 U17488 ( .A(n15673), .ZN(n18642) );
  OAI221_X1 U17489 ( .B1(n18809), .B2(n18642), .C1(n11165), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(P2_STATE2_REG_1__SCAN_IN), .ZN(
        n17178) );
  INV_X1 U17490 ( .A(n15632), .ZN(n15633) );
  INV_X1 U17491 ( .A(n17179), .ZN(n19047) );
  AOI22_X1 U17492 ( .A1(n15634), .A2(n17178), .B1(n15633), .B2(n19047), .ZN(
        n15636) );
  NAND2_X1 U17493 ( .A1(n15938), .A2(n11196), .ZN(n15635) );
  OAI21_X1 U17494 ( .B1(n15938), .B2(n15636), .A(n15635), .ZN(P2_U3601) );
  OAI222_X1 U17495 ( .A1(n15735), .A2(n16219), .B1(n20326), .B2(n15637), .C1(
        n21804), .C2(n16217), .ZN(P1_U2863) );
  XNOR2_X1 U17496 ( .A(n15638), .B(n15642), .ZN(n17430) );
  XNOR2_X1 U17497 ( .A(n15640), .B(n15639), .ZN(n17429) );
  AOI221_X1 U17498 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15643), .C2(n15642), .A(
        n15641), .ZN(n15645) );
  NOR2_X1 U17499 ( .A1(n11955), .A2(n18830), .ZN(n15644) );
  AOI211_X1 U17500 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15646), .A(
        n15645), .B(n15644), .ZN(n15652) );
  OAI21_X1 U17501 ( .B1(n14832), .B2(n15648), .A(n15647), .ZN(n19780) );
  OAI22_X1 U17502 ( .A1(n19780), .A2(n19020), .B1(n18991), .B2(n15649), .ZN(
        n15650) );
  INV_X1 U17503 ( .A(n15650), .ZN(n15651) );
  OAI211_X1 U17504 ( .C1(n17429), .C2(n17166), .A(n15652), .B(n15651), .ZN(
        n15653) );
  INV_X1 U17505 ( .A(n15653), .ZN(n15654) );
  OAI21_X1 U17506 ( .B1(n17430), .B2(n19015), .A(n15654), .ZN(P2_U3041) );
  NOR2_X2 U17507 ( .A1(n19581), .A2(n19657), .ZN(n20041) );
  INV_X1 U17508 ( .A(n20041), .ZN(n15655) );
  NAND3_X1 U17509 ( .A1(n15655), .A2(n19979), .A3(n19708), .ZN(n15656) );
  OR2_X1 U17510 ( .A1(n19694), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19709) );
  NAND3_X1 U17511 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19689), .A3(
        n19592), .ZN(n19590) );
  NOR2_X1 U17512 ( .A1(n19612), .A2(n19590), .ZN(n20047) );
  NAND3_X1 U17513 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19592), .ZN(n19572) );
  NOR2_X1 U17514 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19572), .ZN(
        n20040) );
  NOR2_X1 U17515 ( .A1(n20047), .A2(n20040), .ZN(n15666) );
  INV_X1 U17516 ( .A(n15666), .ZN(n15657) );
  OR2_X1 U17517 ( .A1(n15667), .A2(n15657), .ZN(n15660) );
  INV_X1 U17518 ( .A(n20040), .ZN(n15662) );
  OAI211_X1 U17519 ( .C1(n12534), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19694), 
        .B(n15662), .ZN(n15658) );
  AND2_X1 U17520 ( .A1(n15658), .A2(n19715), .ZN(n15659) );
  AOI22_X1 U17521 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20010), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20011), .ZN(n19761) );
  INV_X1 U17522 ( .A(n19761), .ZN(n19765) );
  AOI22_X1 U17523 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20010), .ZN(n19769) );
  INV_X1 U17524 ( .A(n20007), .ZN(n15661) );
  NAND2_X1 U17525 ( .A1(n11881), .A2(n15661), .ZN(n19732) );
  OAI22_X1 U17526 ( .A1(n19769), .A2(n19979), .B1(n19732), .B2(n15662), .ZN(
        n15663) );
  AOI21_X1 U17527 ( .B1(n19765), .B2(n20041), .A(n15663), .ZN(n15669) );
  INV_X1 U17528 ( .A(n12534), .ZN(n15664) );
  OAI21_X1 U17529 ( .B1(n15664), .B2(n20040), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15665) );
  NOR2_X2 U17530 ( .A1(n19724), .A2(n20005), .ZN(n19766) );
  NAND2_X1 U17531 ( .A1(n20042), .A2(n19766), .ZN(n15668) );
  OAI211_X1 U17532 ( .C1(n20046), .C2(n15670), .A(n15669), .B(n15668), .ZN(
        P2_U3134) );
  INV_X1 U17533 ( .A(n17178), .ZN(n15676) );
  OAI21_X1 U17534 ( .B1(n15673), .B2(n15672), .A(n15671), .ZN(n18656) );
  OAI21_X1 U17535 ( .B1(n11164), .B2(n15674), .A(n18656), .ZN(n17177) );
  AOI222_X1 U17536 ( .A1(n15676), .A2(n17177), .B1(n19047), .B2(n19642), .C1(
        n15675), .C2(n15936), .ZN(n15678) );
  NAND2_X1 U17537 ( .A1(n15938), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15677) );
  OAI21_X1 U17538 ( .B1(n15678), .B2(n15938), .A(n15677), .ZN(P2_U3599) );
  INV_X1 U17539 ( .A(n15679), .ZN(n15682) );
  INV_X1 U17540 ( .A(n15571), .ZN(n15681) );
  AOI21_X1 U17541 ( .B1(n15682), .B2(n15681), .A(n15680), .ZN(n16418) );
  INV_X1 U17542 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15692) );
  NAND2_X1 U17543 ( .A1(n15886), .A2(n15692), .ZN(n15688) );
  NAND2_X1 U17544 ( .A1(n15883), .A2(n15685), .ZN(n15686) );
  OAI211_X1 U17545 ( .C1(n11159), .C2(P1_EBX_REG_10__SCAN_IN), .A(n15686), .B(
        n15889), .ZN(n15687) );
  AND2_X1 U17546 ( .A1(n15688), .A2(n15687), .ZN(n15689) );
  OR2_X2 U17547 ( .A1(n15690), .A2(n15689), .ZN(n20288) );
  NAND2_X1 U17548 ( .A1(n15690), .A2(n15689), .ZN(n15691) );
  NAND2_X1 U17549 ( .A1(n20288), .A2(n15691), .ZN(n21812) );
  OAI22_X1 U17550 ( .A1(n16217), .A2(n21812), .B1(n15692), .B2(n20326), .ZN(
        n15693) );
  AOI21_X1 U17551 ( .B1(n16418), .B2(n20323), .A(n15693), .ZN(n15694) );
  INV_X1 U17552 ( .A(n15694), .ZN(P1_U2862) );
  OAI21_X1 U17553 ( .B1(n15697), .B2(n15696), .A(n15695), .ZN(n21787) );
  NOR2_X1 U17554 ( .A1(n21915), .A2(n20223), .ZN(n21790) );
  AOI21_X1 U17555 ( .B1(n20388), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21790), .ZN(n15698) );
  OAI21_X1 U17556 ( .B1(n20395), .B2(n15699), .A(n15698), .ZN(n15700) );
  AOI21_X1 U17557 ( .B1(n15701), .B2(n20385), .A(n15700), .ZN(n15702) );
  OAI21_X1 U17558 ( .B1(n21787), .B2(n22113), .A(n15702), .ZN(P1_U2991) );
  INV_X1 U17559 ( .A(n16418), .ZN(n15711) );
  INV_X1 U17560 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21813) );
  NAND2_X1 U17561 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15703), .ZN(n15704) );
  NOR2_X1 U17562 ( .A1(n21813), .A2(n15704), .ZN(n21987) );
  OAI21_X1 U17563 ( .B1(n21987), .B2(n22069), .A(n22050), .ZN(n22001) );
  OAI21_X1 U17564 ( .B1(n15704), .B2(n22069), .A(n21813), .ZN(n15708) );
  AOI21_X1 U17565 ( .B1(n22079), .B2(P1_EBX_REG_10__SCAN_IN), .A(n22044), .ZN(
        n15705) );
  OAI21_X1 U17566 ( .B1(n22096), .B2(n16416), .A(n15705), .ZN(n15707) );
  OAI22_X1 U17567 ( .A1(n13347), .A2(n22098), .B1(n22111), .B2(n21812), .ZN(
        n15706) );
  AOI211_X1 U17568 ( .C1(n22001), .C2(n15708), .A(n15707), .B(n15706), .ZN(
        n15709) );
  OAI21_X1 U17569 ( .B1(n15711), .B2(n22052), .A(n15709), .ZN(P1_U2830) );
  AOI22_X1 U17570 ( .A1(n16274), .A2(n16243), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n22375), .ZN(n15710) );
  OAI21_X1 U17571 ( .B1(n15711), .B2(n16281), .A(n15710), .ZN(P1_U2894) );
  AOI21_X1 U17572 ( .B1(n15714), .B2(n15713), .A(n15712), .ZN(n18826) );
  INV_X1 U17573 ( .A(n18826), .ZN(n17044) );
  AOI21_X1 U17574 ( .B1(n15716), .B2(n15575), .A(n15715), .ZN(n15726) );
  NAND2_X1 U17575 ( .A1(n15726), .A2(n16596), .ZN(n15718) );
  NAND2_X1 U17576 ( .A1(n16604), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15717) );
  OAI211_X1 U17577 ( .C1(n17044), .C2(n16604), .A(n15718), .B(n15717), .ZN(
        P2_U2870) );
  XOR2_X1 U17578 ( .A(n15720), .B(n15719), .Z(n18825) );
  INV_X1 U17579 ( .A(n18825), .ZN(n15728) );
  INV_X1 U17580 ( .A(n19909), .ZN(n16696) );
  INV_X1 U17581 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15724) );
  OAI22_X1 U17582 ( .A1(n16694), .A2(n19963), .B1(n15721), .B2(n19770), .ZN(
        n15722) );
  AOI21_X1 U17583 ( .B1(n19908), .B2(BUF1_REG_17__SCAN_IN), .A(n15722), .ZN(
        n15723) );
  OAI21_X1 U17584 ( .B1(n16696), .B2(n15724), .A(n15723), .ZN(n15725) );
  AOI21_X1 U17585 ( .B1(n15726), .B2(n19821), .A(n15725), .ZN(n15727) );
  OAI21_X1 U17586 ( .B1(n15728), .B2(n19912), .A(n15727), .ZN(P2_U2902) );
  OAI21_X1 U17587 ( .B1(n15731), .B2(n15730), .A(n15729), .ZN(n21805) );
  INV_X1 U17588 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20225) );
  NOR2_X1 U17589 ( .A1(n21915), .A2(n20225), .ZN(n21807) );
  AOI21_X1 U17590 ( .B1(n20388), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n21807), .ZN(n15734) );
  NAND2_X1 U17591 ( .A1(n20379), .A2(n15732), .ZN(n15733) );
  OAI211_X1 U17592 ( .C1(n15735), .C2(n16413), .A(n15734), .B(n15733), .ZN(
        n15736) );
  INV_X1 U17593 ( .A(n15736), .ZN(n15737) );
  OAI21_X1 U17594 ( .B1(n21805), .B2(n22113), .A(n15737), .ZN(P1_U2990) );
  XNOR2_X1 U17595 ( .A(n11192), .B(n15787), .ZN(n15748) );
  XNOR2_X1 U17596 ( .A(n15739), .B(n15741), .ZN(n15761) );
  AOI22_X1 U17597 ( .A1(n17457), .A2(n15742), .B1(n17461), .B2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15745) );
  OAI22_X1 U17598 ( .A1(n11961), .A2(n18830), .B1(n17475), .B2(n18692), .ZN(
        n15743) );
  INV_X1 U17599 ( .A(n15743), .ZN(n15744) );
  OAI211_X1 U17600 ( .C1(n15761), .C2(n17445), .A(n15745), .B(n15744), .ZN(
        n15746) );
  AOI21_X1 U17601 ( .B1(n15748), .B2(n17467), .A(n15746), .ZN(n15747) );
  INV_X1 U17602 ( .A(n15747), .ZN(P2_U3008) );
  NAND2_X1 U17603 ( .A1(n15748), .A2(n19007), .ZN(n15760) );
  NAND3_X1 U17604 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n15749), .ZN(n15754) );
  INV_X1 U17605 ( .A(n15754), .ZN(n15750) );
  NAND2_X1 U17606 ( .A1(n15750), .A2(n19027), .ZN(n15786) );
  NAND2_X1 U17607 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15750), .ZN(
        n15783) );
  NOR2_X1 U17608 ( .A1(n15783), .A2(n15751), .ZN(n15980) );
  INV_X1 U17609 ( .A(n15980), .ZN(n15752) );
  NAND2_X1 U17610 ( .A1(n17048), .A2(n15752), .ZN(n15753) );
  NAND2_X1 U17611 ( .A1(n15753), .A2(n18994), .ZN(n15782) );
  AOI21_X1 U17612 ( .B1(n17047), .B2(n15754), .A(n15782), .ZN(n15756) );
  NAND2_X1 U17613 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n11167), .ZN(n15755) );
  OAI221_X1 U17614 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15786), .C1(
        n15787), .C2(n15756), .A(n15755), .ZN(n15758) );
  NOR2_X1 U17615 ( .A1(n18991), .A2(n18698), .ZN(n15757) );
  AOI211_X1 U17616 ( .C1(n18694), .C2(n19003), .A(n15758), .B(n15757), .ZN(
        n15759) );
  OAI211_X1 U17617 ( .C1(n15761), .C2(n17166), .A(n15760), .B(n15759), .ZN(
        P2_U3040) );
  OAI21_X1 U17618 ( .B1(n15680), .B2(n15763), .A(n15762), .ZN(n16146) );
  XNOR2_X1 U17619 ( .A(n16146), .B(n16144), .ZN(n21992) );
  INV_X1 U17620 ( .A(n21992), .ZN(n15766) );
  INV_X1 U17621 ( .A(n16237), .ZN(n15764) );
  OAI222_X1 U17622 ( .A1(n15766), .A2(n16281), .B1(n15765), .B2(n16279), .C1(
        n16278), .C2(n15764), .ZN(P1_U2893) );
  NOR2_X1 U17623 ( .A1(n15715), .A2(n15768), .ZN(n15769) );
  OR2_X1 U17624 ( .A1(n15767), .A2(n15769), .ZN(n19910) );
  NAND2_X1 U17625 ( .A1(n15771), .A2(n15770), .ZN(n15772) );
  NAND2_X1 U17626 ( .A1(n16601), .A2(n15772), .ZN(n18843) );
  NOR2_X1 U17627 ( .A1(n18843), .A2(n16604), .ZN(n15773) );
  AOI21_X1 U17628 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n16604), .A(n15773), .ZN(
        n15774) );
  OAI21_X1 U17629 ( .B1(n19910), .B2(n16606), .A(n15774), .ZN(P2_U2869) );
  XNOR2_X1 U17630 ( .A(n15775), .B(n15776), .ZN(n15799) );
  INV_X1 U17631 ( .A(n15778), .ZN(n15780) );
  NAND2_X1 U17632 ( .A1(n15780), .A2(n15779), .ZN(n15781) );
  XNOR2_X1 U17633 ( .A(n15777), .B(n15781), .ZN(n15797) );
  INV_X1 U17634 ( .A(n15782), .ZN(n15784) );
  NAND2_X1 U17635 ( .A1(n17047), .A2(n15783), .ZN(n15983) );
  NAND2_X1 U17636 ( .A1(n15784), .A2(n15983), .ZN(n19004) );
  OAI22_X1 U17637 ( .A1(n18991), .A2(n18704), .B1(n17551), .B2(n18830), .ZN(
        n15785) );
  AOI21_X1 U17638 ( .B1(n19004), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15785), .ZN(n15790) );
  NOR2_X1 U17639 ( .A1(n15787), .A2(n15786), .ZN(n19010) );
  NAND2_X1 U17640 ( .A1(n19010), .A2(n15788), .ZN(n15789) );
  OAI211_X1 U17641 ( .C1(n18705), .C2(n19020), .A(n15790), .B(n15789), .ZN(
        n15791) );
  AOI21_X1 U17642 ( .B1(n15797), .B2(n19024), .A(n15791), .ZN(n15792) );
  OAI21_X1 U17643 ( .B1(n15799), .B2(n19015), .A(n15792), .ZN(P2_U3039) );
  OAI22_X1 U17644 ( .A1(n15793), .A2(n17452), .B1(n17551), .B2(n18830), .ZN(
        n15796) );
  INV_X1 U17645 ( .A(n18700), .ZN(n15794) );
  OAI22_X1 U17646 ( .A1(n17471), .A2(n18704), .B1(n17475), .B2(n15794), .ZN(
        n15795) );
  AOI211_X1 U17647 ( .C1(n15797), .C2(n17462), .A(n15796), .B(n15795), .ZN(
        n15798) );
  OAI21_X1 U17648 ( .B1(n15799), .B2(n17446), .A(n15798), .ZN(P2_U3007) );
  NAND2_X1 U17649 ( .A1(n11273), .A2(n15800), .ZN(n16147) );
  AOI22_X1 U17650 ( .A1(n16274), .A2(n16220), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n22375), .ZN(n15803) );
  OAI21_X1 U17651 ( .B1(n22008), .B2(n16281), .A(n15803), .ZN(P1_U2890) );
  OAI21_X1 U17652 ( .B1(n11285), .B2(n15805), .A(n15804), .ZN(n16801) );
  NAND2_X1 U17653 ( .A1(n15807), .A2(n15808), .ZN(n15809) );
  AND2_X1 U17654 ( .A1(n15806), .A2(n15809), .ZN(n19820) );
  NAND2_X1 U17655 ( .A1(n19820), .A2(n16596), .ZN(n15811) );
  NAND2_X1 U17656 ( .A1(n16604), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15810) );
  OAI211_X1 U17657 ( .C1(n16801), .C2(n16604), .A(n15811), .B(n15810), .ZN(
        P2_U2867) );
  NOR2_X1 U17658 ( .A1(n22375), .A2(n15820), .ZN(n15814) );
  NAND2_X1 U17659 ( .A1(n15814), .A2(n15812), .ZN(n22383) );
  NAND3_X1 U17660 ( .A1(n16044), .A2(n22633), .A3(n16279), .ZN(n15816) );
  AOI22_X1 U17661 ( .A1(n22378), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n22375), .ZN(n15815) );
  OAI211_X1 U17662 ( .C1(n22383), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        P1_U2873) );
  INV_X1 U17663 ( .A(n15818), .ZN(n15819) );
  OAI211_X1 U17664 ( .C1(n22386), .C2(n22161), .A(n15819), .B(n21697), .ZN(
        n15827) );
  OAI211_X1 U17665 ( .C1(n17413), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        n15823) );
  NAND2_X1 U17666 ( .A1(n15824), .A2(n15823), .ZN(n15826) );
  MUX2_X1 U17667 ( .A(n15827), .B(n15826), .S(n15825), .Z(n15832) );
  NOR2_X1 U17668 ( .A1(n16505), .A2(n22386), .ZN(n15829) );
  AOI21_X1 U17669 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(n15831) );
  NAND2_X1 U17670 ( .A1(n15832), .A2(n15831), .ZN(n15834) );
  INV_X1 U17671 ( .A(n15835), .ZN(n15836) );
  OAI211_X1 U17672 ( .C1(n15837), .C2(n15893), .A(n15836), .B(n17404), .ZN(
        n15838) );
  NOR2_X1 U17673 ( .A1(n15839), .A2(n15838), .ZN(n15840) );
  OAI22_X1 U17674 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n11159), .ZN(n15891) );
  OR2_X1 U17675 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15843) );
  NAND2_X1 U17676 ( .A1(n15841), .A2(n16162), .ZN(n15842) );
  NAND2_X1 U17677 ( .A1(n15843), .A2(n15842), .ZN(n16059) );
  MUX2_X1 U17678 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n15844) );
  NAND2_X1 U17679 ( .A1(n15844), .A2(n11678), .ZN(n20289) );
  NOR2_X2 U17680 ( .A1(n20288), .A2(n20289), .ZN(n20287) );
  OAI21_X1 U17681 ( .B1(n16057), .B2(n21822), .A(n15883), .ZN(n15845) );
  OAI21_X1 U17682 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(n11159), .A(n15845), .ZN(
        n15846) );
  OAI21_X1 U17683 ( .B1(n15878), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15846), .ZN(
        n16214) );
  MUX2_X1 U17684 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n15847) );
  NAND2_X1 U17685 ( .A1(n15847), .A2(n11690), .ZN(n16149) );
  NAND2_X1 U17686 ( .A1(n15886), .A2(n16206), .ZN(n15850) );
  NAND2_X1 U17687 ( .A1(n15883), .A2(n21730), .ZN(n15848) );
  OAI211_X1 U17688 ( .C1(n11159), .C2(P1_EBX_REG_14__SCAN_IN), .A(n15848), .B(
        n15889), .ZN(n15849) );
  AND2_X1 U17689 ( .A1(n15850), .A2(n15849), .ZN(n16204) );
  MUX2_X1 U17690 ( .A(n15868), .B(n16057), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n15852) );
  NOR2_X1 U17691 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15851) );
  NOR2_X1 U17692 ( .A1(n15852), .A2(n15851), .ZN(n16137) );
  NAND2_X1 U17693 ( .A1(n16136), .A2(n16137), .ZN(n16198) );
  INV_X1 U17694 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16200) );
  NAND2_X1 U17695 ( .A1(n15886), .A2(n16200), .ZN(n15855) );
  NAND2_X1 U17696 ( .A1(n15883), .A2(n21865), .ZN(n15853) );
  OAI211_X1 U17697 ( .C1(n11159), .C2(P1_EBX_REG_16__SCAN_IN), .A(n15853), .B(
        n15889), .ZN(n15854) );
  AND2_X1 U17698 ( .A1(n15855), .A2(n15854), .ZN(n16197) );
  MUX2_X1 U17699 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n15856) );
  NAND2_X1 U17700 ( .A1(n15856), .A2(n11689), .ZN(n16123) );
  NAND2_X1 U17701 ( .A1(n15883), .A2(n16357), .ZN(n15857) );
  OAI211_X1 U17702 ( .C1(n11159), .C2(P1_EBX_REG_18__SCAN_IN), .A(n15857), .B(
        n15889), .ZN(n15858) );
  OAI21_X1 U17703 ( .B1(n15878), .B2(P1_EBX_REG_18__SCAN_IN), .A(n15858), .ZN(
        n16187) );
  MUX2_X1 U17704 ( .A(n15868), .B(n16057), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n15860) );
  NOR2_X1 U17705 ( .A1(n15897), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15859) );
  NOR2_X1 U17706 ( .A1(n15860), .A2(n15859), .ZN(n20308) );
  NAND2_X1 U17707 ( .A1(n15886), .A2(n22058), .ZN(n15863) );
  NAND2_X1 U17708 ( .A1(n15883), .A2(n16359), .ZN(n15861) );
  OAI211_X1 U17709 ( .C1(n11159), .C2(P1_EBX_REG_20__SCAN_IN), .A(n15861), .B(
        n15889), .ZN(n15862) );
  AND2_X1 U17710 ( .A1(n15863), .A2(n15862), .ZN(n16181) );
  MUX2_X1 U17711 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n15864) );
  OAI21_X1 U17712 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15897), .A(
        n15864), .ZN(n16479) );
  INV_X1 U17713 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15865) );
  NAND2_X1 U17714 ( .A1(n15883), .A2(n15865), .ZN(n15866) );
  OAI211_X1 U17715 ( .C1(n11159), .C2(P1_EBX_REG_22__SCAN_IN), .A(n15866), .B(
        n15889), .ZN(n15867) );
  OAI21_X1 U17716 ( .B1(n15878), .B2(P1_EBX_REG_22__SCAN_IN), .A(n15867), .ZN(
        n16176) );
  NAND2_X1 U17717 ( .A1(n15868), .A2(n22089), .ZN(n15871) );
  NAND2_X1 U17718 ( .A1(n15889), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15869) );
  OAI211_X1 U17719 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n11159), .A(n15869), .B(
        n15883), .ZN(n15870) );
  AND2_X1 U17720 ( .A1(n15871), .A2(n15870), .ZN(n20300) );
  NAND2_X1 U17721 ( .A1(n15886), .A2(n22101), .ZN(n15874) );
  NAND2_X1 U17722 ( .A1(n15883), .A2(n16461), .ZN(n15872) );
  OAI211_X1 U17723 ( .C1(n11159), .C2(P1_EBX_REG_24__SCAN_IN), .A(n15872), .B(
        n15889), .ZN(n15873) );
  AND2_X1 U17724 ( .A1(n15874), .A2(n15873), .ZN(n16170) );
  MUX2_X1 U17725 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n15875) );
  NAND2_X1 U17726 ( .A1(n15875), .A2(n11687), .ZN(n16114) );
  INV_X1 U17727 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15927) );
  OAI21_X1 U17728 ( .B1(n16057), .B2(n15927), .A(n15883), .ZN(n15876) );
  OAI21_X1 U17729 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n11159), .A(n15876), .ZN(
        n15877) );
  OAI21_X1 U17730 ( .B1(n15878), .B2(P1_EBX_REG_26__SCAN_IN), .A(n15877), .ZN(
        n16099) );
  MUX2_X1 U17731 ( .A(n15879), .B(n15889), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n15880) );
  OAI21_X1 U17732 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15897), .A(
        n15880), .ZN(n16083) );
  INV_X1 U17733 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16445) );
  OAI21_X1 U17734 ( .B1(n11159), .B2(P1_EBX_REG_28__SCAN_IN), .A(n15889), .ZN(
        n15882) );
  AOI21_X1 U17735 ( .B1(n15883), .B2(n16445), .A(n15882), .ZN(n15884) );
  AOI21_X1 U17736 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n16076) );
  NOR2_X1 U17737 ( .A1(n11159), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n15888) );
  INV_X1 U17738 ( .A(n15897), .ZN(n15887) );
  AOI21_X1 U17739 ( .B1(n15887), .B2(n16432), .A(n15888), .ZN(n16056) );
  MUX2_X1 U17740 ( .A(n15888), .B(n16056), .S(n15889), .Z(n16064) );
  NAND2_X1 U17741 ( .A1(n16075), .A2(n16064), .ZN(n16058) );
  MUX2_X1 U17742 ( .A(n16059), .B(n15889), .S(n16058), .Z(n15890) );
  XOR2_X1 U17743 ( .A(n15891), .B(n15890), .Z(n16158) );
  NOR2_X1 U17744 ( .A1(n15893), .A2(n15892), .ZN(n15894) );
  AOI21_X1 U17745 ( .B1(n15895), .B2(n22386), .A(n15894), .ZN(n15896) );
  NOR2_X2 U17746 ( .A1(n15907), .A2(n15896), .ZN(n21925) );
  NAND2_X1 U17747 ( .A1(n15898), .A2(n15897), .ZN(n15899) );
  NAND2_X1 U17748 ( .A1(n15900), .A2(n15899), .ZN(n15901) );
  NOR2_X1 U17749 ( .A1(n15902), .A2(n15901), .ZN(n15903) );
  NOR2_X1 U17750 ( .A1(n15907), .A2(n15903), .ZN(n16491) );
  INV_X1 U17751 ( .A(n16491), .ZN(n21707) );
  INV_X1 U17752 ( .A(n15907), .ZN(n15906) );
  INV_X1 U17753 ( .A(n17375), .ZN(n16519) );
  NAND2_X1 U17754 ( .A1(n15906), .A2(n16519), .ZN(n21878) );
  OR2_X1 U17755 ( .A1(n21826), .A2(n15904), .ZN(n15921) );
  NAND2_X1 U17756 ( .A1(n15906), .A2(n15905), .ZN(n21705) );
  NAND2_X1 U17757 ( .A1(n16491), .A2(n21743), .ZN(n15908) );
  NAND2_X1 U17758 ( .A1(n21915), .A2(n15907), .ZN(n21935) );
  AND2_X1 U17759 ( .A1(n15908), .A2(n21935), .ZN(n21734) );
  NOR2_X1 U17760 ( .A1(n15910), .A2(n15909), .ZN(n21761) );
  NAND2_X1 U17761 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21761), .ZN(
        n21765) );
  NOR2_X1 U17762 ( .A1(n21762), .A2(n21765), .ZN(n21800) );
  NOR2_X1 U17763 ( .A1(n21798), .A2(n21789), .ZN(n21801) );
  NAND2_X1 U17764 ( .A1(n21800), .A2(n21801), .ZN(n21803) );
  NOR3_X1 U17765 ( .A1(n21811), .A2(n15685), .A3(n21803), .ZN(n21727) );
  OAI21_X1 U17766 ( .B1(n21743), .B2(n21936), .A(n21748), .ZN(n21779) );
  NAND3_X1 U17767 ( .A1(n21727), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n21779), .ZN(n21820) );
  NOR2_X1 U17768 ( .A1(n21822), .A2(n21820), .ZN(n21706) );
  NAND3_X1 U17769 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n21706), .ZN(n16471) );
  INV_X1 U17770 ( .A(n21888), .ZN(n15915) );
  INV_X1 U17771 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21855) );
  NOR2_X1 U17772 ( .A1(n21855), .A2(n21870), .ZN(n21850) );
  NAND2_X1 U17773 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21850), .ZN(
        n16474) );
  NOR2_X1 U17774 ( .A1(n15865), .A2(n16474), .ZN(n15911) );
  NAND2_X1 U17775 ( .A1(n15915), .A2(n15911), .ZN(n15912) );
  NOR2_X1 U17776 ( .A1(n16471), .A2(n15912), .ZN(n15924) );
  NAND2_X1 U17777 ( .A1(n15924), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15913) );
  NAND2_X1 U17778 ( .A1(n21821), .A2(n15913), .ZN(n15914) );
  AND2_X1 U17779 ( .A1(n21734), .A2(n15914), .ZN(n15918) );
  NAND3_X1 U17780 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21727), .ZN(n21823) );
  NAND2_X1 U17781 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21728) );
  NOR2_X1 U17782 ( .A1(n21823), .A2(n21728), .ZN(n21715) );
  NAND2_X1 U17783 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21715), .ZN(
        n21710) );
  NOR2_X1 U17784 ( .A1(n21730), .A2(n21710), .ZN(n16473) );
  INV_X1 U17785 ( .A(n16474), .ZN(n16482) );
  NAND2_X1 U17786 ( .A1(n16473), .A2(n16482), .ZN(n16483) );
  NAND2_X1 U17787 ( .A1(n15915), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15916) );
  NOR2_X1 U17788 ( .A1(n16483), .A2(n15916), .ZN(n15925) );
  OR2_X1 U17789 ( .A1(n21826), .A2(n15925), .ZN(n15917) );
  AND2_X1 U17790 ( .A1(n15918), .A2(n15917), .ZN(n16462) );
  OAI21_X1 U17791 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n21705), .A(
        n16462), .ZN(n15919) );
  INV_X1 U17792 ( .A(n15919), .ZN(n15920) );
  AND2_X1 U17793 ( .A1(n15921), .A2(n15920), .ZN(n21913) );
  NAND2_X1 U17794 ( .A1(n21913), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n21901) );
  OR2_X1 U17795 ( .A1(n21901), .A2(n21912), .ZN(n15922) );
  AND2_X1 U17796 ( .A1(n21826), .A2(n21705), .ZN(n21848) );
  NAND2_X1 U17797 ( .A1(n21848), .A2(n21734), .ZN(n21783) );
  NAND2_X1 U17798 ( .A1(n15922), .A2(n21783), .ZN(n16451) );
  NAND2_X1 U17799 ( .A1(n16451), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16422) );
  INV_X1 U17800 ( .A(n16433), .ZN(n16441) );
  NAND2_X1 U17801 ( .A1(n16441), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15928) );
  OAI211_X1 U17802 ( .C1(n16422), .C2(n15928), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n21783), .ZN(n15931) );
  INV_X1 U17803 ( .A(n15923), .ZN(n15930) );
  NAND2_X1 U17804 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16491), .ZN(
        n16480) );
  NAND2_X1 U17805 ( .A1(n21878), .A2(n16480), .ZN(n21725) );
  AOI22_X1 U17806 ( .A1(n15925), .A2(n21725), .B1(n21821), .B2(n15924), .ZN(
        n16466) );
  NOR2_X1 U17807 ( .A1(n16466), .A2(n15926), .ZN(n21900) );
  NAND2_X1 U17808 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21900), .ZN(
        n21899) );
  NOR2_X1 U17809 ( .A1(n21899), .A2(n15927), .ZN(n16455) );
  INV_X1 U17810 ( .A(n15928), .ZN(n16421) );
  NAND4_X1 U17811 ( .A1(n16455), .A2(n16421), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n16508), .ZN(n15929) );
  NAND3_X1 U17812 ( .A1(n15931), .A2(n15930), .A3(n15929), .ZN(n15932) );
  AOI21_X1 U17813 ( .B1(n16158), .B2(n21925), .A(n15932), .ZN(n15933) );
  OAI21_X1 U17814 ( .B1(n15934), .B2(n21862), .A(n15933), .ZN(P1_U3000) );
  AOI22_X1 U17815 ( .A1(n19660), .A2(n19047), .B1(n15936), .B2(n15935), .ZN(
        n15939) );
  NAND2_X1 U17816 ( .A1(n15938), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15937) );
  OAI21_X1 U17817 ( .B1(n15939), .B2(n15938), .A(n15937), .ZN(P2_U3596) );
  NOR2_X1 U17818 ( .A1(n16571), .A2(n12428), .ZN(n15940) );
  AOI21_X1 U17819 ( .B1(n16571), .B2(n13756), .A(n15940), .ZN(n15941) );
  OAI21_X1 U17820 ( .B1(n19573), .B2(n16606), .A(n15941), .ZN(P2_U2884) );
  NAND2_X1 U17821 ( .A1(n11164), .A2(n15942), .ZN(n15943) );
  XNOR2_X1 U17822 ( .A(n15944), .B(n15943), .ZN(n15945) );
  NAND2_X1 U17823 ( .A1(n15945), .A2(n18980), .ZN(n15953) );
  OAI22_X1 U17824 ( .A1(n15946), .A2(n18973), .B1(n18922), .B2(n19021), .ZN(
        n15949) );
  NOR2_X1 U17825 ( .A1(n18969), .A2(n15947), .ZN(n15948) );
  AOI211_X1 U17826 ( .C1(n18954), .C2(P2_REIP_REG_3__SCAN_IN), .A(n15949), .B(
        n15948), .ZN(n15950) );
  OAI21_X1 U17827 ( .B1(n18884), .B2(n12428), .A(n15950), .ZN(n15951) );
  AOI21_X1 U17828 ( .B1(n18957), .B2(n13756), .A(n15951), .ZN(n15952) );
  OAI211_X1 U17829 ( .C1(n18666), .C2(n19573), .A(n15953), .B(n15952), .ZN(
        P2_U2852) );
  INV_X1 U17830 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n15958) );
  OAI22_X1 U17831 ( .A1(n16694), .A2(n15955), .B1(n15954), .B2(n19770), .ZN(
        n15956) );
  AOI21_X1 U17832 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n19908), .A(n15956), .ZN(
        n15957) );
  OAI21_X1 U17833 ( .B1(n16696), .B2(n15958), .A(n15957), .ZN(n15959) );
  AOI21_X1 U17834 ( .B1(n15997), .B2(n19822), .A(n15959), .ZN(n15960) );
  OAI21_X1 U17835 ( .B1(n15961), .B2(n19911), .A(n15960), .ZN(P2_U2889) );
  INV_X1 U17836 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15965) );
  NOR2_X1 U17837 ( .A1(n16001), .A2(n11284), .ZN(n15967) );
  INV_X1 U17838 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15969) );
  NOR2_X1 U17839 ( .A1(n18830), .A2(n15969), .ZN(n15990) );
  AOI21_X1 U17840 ( .B1(n17461), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15990), .ZN(n15970) );
  OAI21_X1 U17841 ( .B1(n17475), .B2(n18978), .A(n15970), .ZN(n15972) );
  XNOR2_X1 U17842 ( .A(n16019), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15994) );
  NOR2_X1 U17843 ( .A1(n15994), .A2(n17446), .ZN(n15971) );
  AOI211_X1 U17844 ( .C1(n17457), .C2(n15977), .A(n15972), .B(n15971), .ZN(
        n15973) );
  OAI21_X1 U17845 ( .B1(n11184), .B2(n17445), .A(n15973), .ZN(P2_U2984) );
  NOR2_X1 U17846 ( .A1(n15974), .A2(n16893), .ZN(n15978) );
  NAND2_X1 U17847 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19009) );
  INV_X1 U17848 ( .A(n19009), .ZN(n15981) );
  NAND2_X1 U17849 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16963) );
  NOR3_X1 U17850 ( .A1(n15975), .A2(n16964), .A3(n16963), .ZN(n15979) );
  NAND2_X1 U17851 ( .A1(n17156), .A2(n15979), .ZN(n16953) );
  NAND2_X1 U17852 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15976) );
  OR2_X1 U17853 ( .A1(n16953), .A2(n15976), .ZN(n16925) );
  INV_X1 U17854 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16931) );
  NOR2_X1 U17855 ( .A1(n16925), .A2(n16931), .ZN(n16894) );
  NAND2_X1 U17856 ( .A1(n15978), .A2(n16894), .ZN(n15993) );
  INV_X1 U17857 ( .A(n18991), .ZN(n19017) );
  NAND2_X1 U17858 ( .A1(n15977), .A2(n19017), .ZN(n15992) );
  NAND2_X1 U17859 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15978), .ZN(
        n16028) );
  INV_X1 U17860 ( .A(n16028), .ZN(n15989) );
  OR2_X1 U17861 ( .A1(n19001), .A2(n15979), .ZN(n15986) );
  NAND2_X1 U17862 ( .A1(n17047), .A2(n19009), .ZN(n15985) );
  NAND2_X1 U17863 ( .A1(n15981), .A2(n15980), .ZN(n15982) );
  NAND2_X1 U17864 ( .A1(n17048), .A2(n15982), .ZN(n15984) );
  AND2_X1 U17865 ( .A1(n18994), .A2(n15983), .ZN(n15987) );
  AND3_X1 U17866 ( .A1(n15985), .A2(n15984), .A3(n15987), .ZN(n17121) );
  NAND3_X1 U17867 ( .A1(n15986), .A2(n17121), .A3(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16950) );
  NAND2_X1 U17868 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U17869 ( .A1(n19001), .A2(n15987), .ZN(n17122) );
  OAI21_X1 U17870 ( .B1(n16950), .B2(n15988), .A(n17122), .ZN(n16914) );
  OAI21_X1 U17871 ( .B1(n19001), .B2(n15989), .A(n16914), .ZN(n16032) );
  AOI21_X1 U17872 ( .B1(n16032), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15990), .ZN(n15991) );
  OAI211_X1 U17873 ( .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n15993), .A(
        n15992), .B(n15991), .ZN(n15996) );
  NOR2_X1 U17874 ( .A1(n15994), .A2(n19015), .ZN(n15995) );
  AOI211_X1 U17875 ( .C1(n19003), .C2(n15997), .A(n15996), .B(n15995), .ZN(
        n15998) );
  OAI21_X1 U17876 ( .B1(n11184), .B2(n17166), .A(n15998), .ZN(P2_U3016) );
  NOR2_X1 U17877 ( .A1(n16003), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n16006) );
  MUX2_X1 U17878 ( .A(n16006), .B(n16005), .S(n16004), .Z(n18966) );
  NAND2_X1 U17879 ( .A1(n18966), .A2(n11468), .ZN(n16007) );
  XNOR2_X1 U17880 ( .A(n16009), .B(n16008), .ZN(n16039) );
  INV_X1 U17881 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18967) );
  AOI22_X1 U17882 ( .A1(n16012), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n16013) );
  OAI21_X1 U17883 ( .B1(n16014), .B2(n18967), .A(n16013), .ZN(n16015) );
  AOI21_X1 U17884 ( .B1(n11865), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16015), .ZN(n16016) );
  AND2_X1 U17885 ( .A1(n11167), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n16031) );
  AOI21_X1 U17886 ( .B1(n17461), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16031), .ZN(n16017) );
  OAI21_X1 U17887 ( .B1(n17475), .B2(n16018), .A(n16017), .ZN(n16022) );
  NOR2_X1 U17888 ( .A1(n16035), .A2(n17446), .ZN(n16021) );
  OAI21_X1 U17889 ( .B1(n16039), .B2(n17445), .A(n16023), .ZN(P2_U2983) );
  AOI222_X1 U17890 ( .A1(n12093), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n16025), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11166), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16026) );
  XNOR2_X1 U17891 ( .A(n16027), .B(n16026), .ZN(n19524) );
  INV_X1 U17892 ( .A(n16894), .ZN(n16029) );
  NOR3_X1 U17893 ( .A1(n16029), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16028), .ZN(n16030) );
  AOI211_X1 U17894 ( .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16032), .A(
        n16031), .B(n16030), .ZN(n16033) );
  OAI21_X1 U17895 ( .B1(n16034), .B2(n18991), .A(n16033), .ZN(n16037) );
  NOR2_X1 U17896 ( .A1(n16035), .A2(n19015), .ZN(n16036) );
  OAI21_X1 U17897 ( .B1(n16039), .B2(n17166), .A(n16038), .ZN(P2_U3015) );
  INV_X1 U17898 ( .A(n16040), .ZN(n16041) );
  OAI21_X1 U17899 ( .B1(n16041), .B2(n22135), .A(P1_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n16042) );
  NAND3_X1 U17900 ( .A1(n16043), .A2(n20399), .A3(n16042), .ZN(P1_U2801) );
  INV_X1 U17901 ( .A(n16044), .ZN(n16052) );
  INV_X1 U17902 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n22086) );
  INV_X1 U17903 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n22075) );
  NAND2_X1 U17904 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21987), .ZN(n21997) );
  NOR2_X1 U17905 ( .A1(n21828), .A2(n21997), .ZN(n16152) );
  NAND2_X1 U17906 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16152), .ZN(n16151) );
  INV_X1 U17907 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20239) );
  INV_X1 U17908 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21864) );
  NOR4_X1 U17909 ( .A1(n20231), .A2(n20239), .A3(n21864), .A4(n21721), .ZN(
        n16045) );
  NAND4_X1 U17910 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_17__SCAN_IN), .A4(n16045), .ZN(n16046) );
  NOR2_X1 U17911 ( .A1(n16151), .A2(n16046), .ZN(n22060) );
  NAND2_X1 U17912 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22060), .ZN(n22070) );
  NOR2_X1 U17913 ( .A1(n22075), .A2(n22070), .ZN(n16108) );
  NAND2_X1 U17914 ( .A1(n16108), .A2(n22073), .ZN(n22087) );
  NOR2_X1 U17915 ( .A1(n22086), .A2(n22087), .ZN(n22104) );
  NAND2_X1 U17916 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n22104), .ZN(n16096) );
  INV_X1 U17917 ( .A(n16096), .ZN(n16112) );
  NAND3_X1 U17918 ( .A1(n16112), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_26__SCAN_IN), .ZN(n16104) );
  INV_X1 U17919 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20249) );
  NOR2_X1 U17920 ( .A1(n16104), .A2(n20249), .ZN(n16088) );
  NAND2_X1 U17921 ( .A1(n16088), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U17922 ( .A1(n16077), .A2(n20255), .ZN(n16067) );
  NAND2_X1 U17923 ( .A1(n16067), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16049) );
  NAND3_X1 U17924 ( .A1(n16049), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n22040), 
        .ZN(n16048) );
  AOI22_X1 U17925 ( .A1(n22061), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n22079), .ZN(n16047) );
  OAI211_X1 U17926 ( .C1(n16049), .C2(P1_REIP_REG_31__SCAN_IN), .A(n16048), 
        .B(n16047), .ZN(n16050) );
  AOI21_X1 U17927 ( .B1(n16158), .B2(n22093), .A(n16050), .ZN(n16051) );
  OAI21_X1 U17928 ( .B1(n16052), .B2(n22052), .A(n16051), .ZN(P1_U2809) );
  XOR2_X1 U17929 ( .A(n16053), .B(n16065), .Z(n16291) );
  INV_X1 U17930 ( .A(n16291), .ZN(n16226) );
  AOI22_X1 U17931 ( .A1(n22107), .A2(n16287), .B1(n22079), .B2(
        P1_EBX_REG_30__SCAN_IN), .ZN(n16054) );
  OAI21_X1 U17932 ( .B1(n22098), .B2(n16289), .A(n16054), .ZN(n16055) );
  INV_X1 U17933 ( .A(n16055), .ZN(n16061) );
  AOI22_X1 U17934 ( .A1(n16058), .A2(n16057), .B1(n16056), .B2(n16075), .ZN(
        n16060) );
  XNOR2_X1 U17935 ( .A(n16060), .B(n16059), .ZN(n16161) );
  INV_X1 U17936 ( .A(n16062), .ZN(n16063) );
  OAI21_X1 U17937 ( .B1(n16226), .B2(n22052), .A(n16063), .ZN(P1_U2810) );
  OAI21_X1 U17938 ( .B1(n16075), .B2(n16064), .A(n16058), .ZN(n16434) );
  AOI21_X1 U17939 ( .B1(n16066), .B2(n16073), .A(n16065), .ZN(n16298) );
  NAND2_X1 U17940 ( .A1(n16298), .A2(n22108), .ZN(n16072) );
  INV_X1 U17941 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16163) );
  OAI22_X1 U17942 ( .A1(n22096), .A2(n16296), .B1(n22100), .B2(n16163), .ZN(
        n16070) );
  NAND2_X1 U17943 ( .A1(n22040), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16068) );
  AOI21_X1 U17944 ( .B1(n16077), .B2(n16068), .A(n16067), .ZN(n16069) );
  AOI211_X1 U17945 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16070), .B(n16069), .ZN(n16071) );
  OAI211_X1 U17946 ( .C1(n22111), .C2(n16434), .A(n16072), .B(n16071), .ZN(
        P1_U2811) );
  OAI21_X1 U17947 ( .B1(n16086), .B2(n16074), .A(n16073), .ZN(n16308) );
  AOI21_X1 U17948 ( .B1(n16076), .B2(n11219), .A(n16075), .ZN(n16448) );
  INV_X1 U17949 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16307) );
  NOR2_X1 U17950 ( .A1(n22085), .A2(n20252), .ZN(n16078) );
  OAI21_X1 U17951 ( .B1(n16088), .B2(n16078), .A(n16077), .ZN(n16080) );
  AOI22_X1 U17952 ( .A1(n22107), .A2(n16311), .B1(n22079), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n16079) );
  OAI211_X1 U17953 ( .C1(n22098), .C2(n16307), .A(n16080), .B(n16079), .ZN(
        n16081) );
  AOI21_X1 U17954 ( .B1(n16448), .B2(n22093), .A(n16081), .ZN(n16082) );
  OAI21_X1 U17955 ( .B1(n16308), .B2(n22052), .A(n16082), .ZN(P1_U2812) );
  NAND2_X1 U17956 ( .A1(n11249), .A2(n16083), .ZN(n16084) );
  NAND2_X1 U17957 ( .A1(n11219), .A2(n16084), .ZN(n16456) );
  AOI21_X1 U17958 ( .B1(n16087), .B2(n16085), .A(n16086), .ZN(n16318) );
  NAND2_X1 U17959 ( .A1(n16318), .A2(n22108), .ZN(n16093) );
  INV_X1 U17960 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16165) );
  OAI22_X1 U17961 ( .A1(n22096), .A2(n16316), .B1(n22100), .B2(n16165), .ZN(
        n16091) );
  NAND2_X1 U17962 ( .A1(n22040), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16089) );
  AOI21_X1 U17963 ( .B1(n16104), .B2(n16089), .A(n16088), .ZN(n16090) );
  AOI211_X1 U17964 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16091), .B(n16090), .ZN(n16092) );
  OAI211_X1 U17965 ( .C1(n22111), .C2(n16456), .A(n16093), .B(n16092), .ZN(
        P1_U2813) );
  OAI21_X1 U17966 ( .B1(n16094), .B2(n16095), .A(n16085), .ZN(n16328) );
  INV_X1 U17967 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20246) );
  OAI22_X1 U17968 ( .A1(n16096), .A2(n20246), .B1(n22085), .B2(n20248), .ZN(
        n16103) );
  INV_X1 U17969 ( .A(n16322), .ZN(n16098) );
  AOI22_X1 U17970 ( .A1(n22061), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n22079), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n16097) );
  OAI21_X1 U17971 ( .B1(n22096), .B2(n16098), .A(n16097), .ZN(n16102) );
  OR2_X1 U17972 ( .A1(n16113), .A2(n16099), .ZN(n16100) );
  NAND2_X1 U17973 ( .A1(n11249), .A2(n16100), .ZN(n21905) );
  NOR2_X1 U17974 ( .A1(n21905), .A2(n22111), .ZN(n16101) );
  AOI211_X1 U17975 ( .C1(n16104), .C2(n16103), .A(n16102), .B(n16101), .ZN(
        n16105) );
  OAI21_X1 U17976 ( .B1(n16328), .B2(n22052), .A(n16105), .ZN(P1_U2814) );
  AOI21_X1 U17977 ( .B1(n16107), .B2(n16106), .A(n16094), .ZN(n16336) );
  INV_X1 U17978 ( .A(n16336), .ZN(n16254) );
  AND3_X1 U17979 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n16108), .A3(n22050), 
        .ZN(n22084) );
  AOI211_X1 U17980 ( .C1(n22084), .C2(P1_REIP_REG_24__SCAN_IN), .A(n22085), 
        .B(n20246), .ZN(n16111) );
  AOI22_X1 U17981 ( .A1(n22061), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n22079), .B2(P1_EBX_REG_25__SCAN_IN), .ZN(n16109) );
  OAI21_X1 U17982 ( .B1(n22096), .B2(n16334), .A(n16109), .ZN(n16110) );
  AOI211_X1 U17983 ( .C1(n16112), .C2(n20246), .A(n16111), .B(n16110), .ZN(
        n16116) );
  AOI21_X1 U17984 ( .B1(n16114), .B2(n16172), .A(n16113), .ZN(n21909) );
  NAND2_X1 U17985 ( .A1(n21909), .A2(n22093), .ZN(n16115) );
  OAI211_X1 U17986 ( .C1(n16254), .C2(n22052), .A(n16116), .B(n16115), .ZN(
        P1_U2815) );
  AND2_X1 U17987 ( .A1(n16117), .A2(n16118), .ZN(n16194) );
  NAND2_X1 U17988 ( .A1(n16117), .A2(n16120), .ZN(n16191) );
  INV_X1 U17989 ( .A(n22214), .ZN(n16129) );
  AND2_X1 U17990 ( .A1(n11247), .A2(n16123), .ZN(n16124) );
  NOR2_X1 U17991 ( .A1(n16122), .A2(n16124), .ZN(n21859) );
  INV_X1 U17992 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n20292) );
  AOI22_X1 U17993 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n22061), .B1(
        n20380), .B2(n22107), .ZN(n16125) );
  OAI211_X1 U17994 ( .C1(n22100), .C2(n20292), .A(n16125), .B(n22023), .ZN(
        n16127) );
  INV_X1 U17995 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20235) );
  NOR2_X1 U17996 ( .A1(n16151), .A2(n22069), .ZN(n22012) );
  NAND2_X1 U17997 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n22012), .ZN(n22011) );
  NAND2_X1 U17998 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22021), .ZN(n22020) );
  NOR2_X1 U17999 ( .A1(n20235), .A2(n22020), .ZN(n22026) );
  AOI211_X1 U18000 ( .C1(n20235), .C2(n22020), .A(n22026), .B(n22085), .ZN(
        n16126) );
  AOI211_X1 U18001 ( .C1(n21859), .C2(n22093), .A(n16127), .B(n16126), .ZN(
        n16128) );
  OAI21_X1 U18002 ( .B1(n16129), .B2(n22052), .A(n16128), .ZN(P1_U2823) );
  NAND2_X1 U18003 ( .A1(n16130), .A2(n16117), .ZN(n16196) );
  INV_X1 U18004 ( .A(n16196), .ZN(n16131) );
  INV_X1 U18005 ( .A(n22011), .ZN(n16134) );
  AOI21_X1 U18006 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n22040), .A(n16134), 
        .ZN(n16135) );
  INV_X1 U18007 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20294) );
  OAI22_X1 U18008 ( .A1(n22021), .A2(n16135), .B1(n20294), .B2(n22100), .ZN(
        n16142) );
  OAI21_X1 U18009 ( .B1(n16136), .B2(n16137), .A(n16198), .ZN(n16138) );
  INV_X1 U18010 ( .A(n16138), .ZN(n21843) );
  AOI22_X1 U18011 ( .A1(n21843), .A2(n22093), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n22061), .ZN(n16139) );
  OAI211_X1 U18012 ( .C1(n16140), .C2(n22096), .A(n16139), .B(n22023), .ZN(
        n16141) );
  AOI211_X1 U18013 ( .C1(n20367), .C2(n22108), .A(n16142), .B(n16141), .ZN(
        n16143) );
  INV_X1 U18014 ( .A(n16143), .ZN(P1_U2825) );
  INV_X1 U18015 ( .A(n16144), .ZN(n16145) );
  OAI21_X1 U18016 ( .B1(n16146), .B2(n16145), .A(n15762), .ZN(n16209) );
  AND2_X1 U18017 ( .A1(n16209), .A2(n16210), .ZN(n16211) );
  OAI21_X1 U18018 ( .B1(n16211), .B2(n16148), .A(n16147), .ZN(n16412) );
  NAND2_X1 U18019 ( .A1(n16215), .A2(n16149), .ZN(n16150) );
  AND2_X1 U18020 ( .A1(n16203), .A2(n16150), .ZN(n21717) );
  INV_X1 U18021 ( .A(n21717), .ZN(n16208) );
  INV_X1 U18022 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16406) );
  OAI22_X1 U18023 ( .A1(n16208), .A2(n22111), .B1(n16406), .B2(n22098), .ZN(
        n16156) );
  INV_X1 U18024 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16207) );
  AOI21_X1 U18025 ( .B1(n21964), .B2(P1_REIP_REG_13__SCAN_IN), .A(n22044), 
        .ZN(n16154) );
  OAI211_X1 U18026 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n16152), .A(n22073), 
        .B(n16151), .ZN(n16153) );
  OAI211_X1 U18027 ( .C1(n22100), .C2(n16207), .A(n16154), .B(n16153), .ZN(
        n16155) );
  AOI211_X1 U18028 ( .C1(n22107), .C2(n16409), .A(n16156), .B(n16155), .ZN(
        n16157) );
  OAI21_X1 U18029 ( .B1(n16412), .B2(n22052), .A(n16157), .ZN(P1_U2827) );
  INV_X1 U18030 ( .A(n16158), .ZN(n16160) );
  OAI22_X1 U18031 ( .A1(n16160), .A2(n16217), .B1(n20326), .B2(n16159), .ZN(
        P1_U2841) );
  OAI222_X1 U18032 ( .A1(n16226), .A2(n16219), .B1(n16162), .B2(n20326), .C1(
        n16217), .C2(n16161), .ZN(P1_U2842) );
  INV_X1 U18033 ( .A(n16298), .ZN(n16231) );
  OAI222_X1 U18034 ( .A1(n16219), .A2(n16231), .B1(n16163), .B2(n20326), .C1(
        n16434), .C2(n16217), .ZN(P1_U2843) );
  AOI22_X1 U18035 ( .A1(n16448), .A2(n20322), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n16167), .ZN(n16164) );
  OAI21_X1 U18036 ( .B1(n16308), .B2(n16219), .A(n16164), .ZN(P1_U2844) );
  INV_X1 U18037 ( .A(n16318), .ZN(n16242) );
  OAI222_X1 U18038 ( .A1(n16219), .A2(n16242), .B1(n16165), .B2(n20326), .C1(
        n16456), .C2(n16217), .ZN(P1_U2845) );
  INV_X1 U18039 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16166) );
  OAI222_X1 U18040 ( .A1(n21905), .A2(n16217), .B1(n16166), .B2(n20326), .C1(
        n16328), .C2(n16219), .ZN(P1_U2846) );
  AOI22_X1 U18041 ( .A1(n21909), .A2(n20322), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n16167), .ZN(n16168) );
  OAI21_X1 U18042 ( .B1(n16254), .B2(n16219), .A(n16168), .ZN(P1_U2847) );
  OAI21_X1 U18043 ( .B1(n20297), .B2(n16169), .A(n16106), .ZN(n16343) );
  NAND2_X1 U18044 ( .A1(n20299), .A2(n16170), .ZN(n16171) );
  NAND2_X1 U18045 ( .A1(n16172), .A2(n16171), .ZN(n22112) );
  OAI222_X1 U18046 ( .A1(n16219), .A2(n16343), .B1(n22101), .B2(n20326), .C1(
        n22112), .C2(n16217), .ZN(P1_U2848) );
  NAND2_X1 U18047 ( .A1(n16354), .A2(n16173), .ZN(n16174) );
  AND2_X1 U18048 ( .A1(n20296), .A2(n16174), .ZN(n22224) );
  NOR2_X1 U18049 ( .A1(n16477), .A2(n16176), .ZN(n16177) );
  OR2_X1 U18050 ( .A1(n16175), .A2(n16177), .ZN(n22083) );
  INV_X1 U18051 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16178) );
  OAI22_X1 U18052 ( .A1(n22083), .A2(n16217), .B1(n16178), .B2(n20326), .ZN(
        n16179) );
  AOI21_X1 U18053 ( .B1(n22224), .B2(n20323), .A(n16179), .ZN(n16180) );
  INV_X1 U18054 ( .A(n16180), .ZN(P1_U2850) );
  NAND2_X1 U18055 ( .A1(n20311), .A2(n16181), .ZN(n16182) );
  NAND2_X1 U18056 ( .A1(n16478), .A2(n16182), .ZN(n22051) );
  INV_X1 U18057 ( .A(n16184), .ZN(n16185) );
  OAI21_X1 U18058 ( .B1(n16183), .B2(n16186), .A(n16185), .ZN(n22053) );
  OAI222_X1 U18059 ( .A1(n22051), .A2(n16217), .B1(n22058), .B2(n20326), .C1(
        n22053), .C2(n16219), .ZN(P1_U2852) );
  NOR2_X1 U18060 ( .A1(n16122), .A2(n16187), .ZN(n16188) );
  OR2_X1 U18061 ( .A1(n20309), .A2(n16188), .ZN(n22031) );
  INV_X1 U18062 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n22028) );
  NAND2_X1 U18063 ( .A1(n16117), .A2(n16189), .ZN(n20306) );
  INV_X1 U18064 ( .A(n20306), .ZN(n16190) );
  AOI21_X1 U18065 ( .B1(n16192), .B2(n16191), .A(n16190), .ZN(n22033) );
  INV_X1 U18066 ( .A(n22033), .ZN(n16193) );
  OAI222_X1 U18067 ( .A1(n22031), .A2(n16217), .B1(n22028), .B2(n20326), .C1(
        n16193), .C2(n16219), .ZN(P1_U2854) );
  AOI21_X1 U18068 ( .B1(n16196), .B2(n16195), .A(n16194), .ZN(n16376) );
  NAND2_X1 U18069 ( .A1(n16198), .A2(n16197), .ZN(n16199) );
  NAND2_X1 U18070 ( .A1(n11247), .A2(n16199), .ZN(n22016) );
  OAI22_X1 U18071 ( .A1(n22016), .A2(n16217), .B1(n16200), .B2(n20326), .ZN(
        n16201) );
  AOI21_X1 U18072 ( .B1(n16376), .B2(n20323), .A(n16201), .ZN(n16202) );
  INV_X1 U18073 ( .A(n16202), .ZN(P1_U2856) );
  AOI21_X1 U18074 ( .B1(n16204), .B2(n16203), .A(n16136), .ZN(n16205) );
  INV_X1 U18075 ( .A(n16205), .ZN(n22007) );
  OAI222_X1 U18076 ( .A1(n22008), .A2(n16219), .B1(n16206), .B2(n20326), .C1(
        n16217), .C2(n22007), .ZN(P1_U2858) );
  OAI222_X1 U18077 ( .A1(n16208), .A2(n16217), .B1(n16207), .B2(n20326), .C1(
        n16412), .C2(n16219), .ZN(P1_U2859) );
  INV_X1 U18078 ( .A(n16209), .ZN(n16213) );
  INV_X1 U18079 ( .A(n16210), .ZN(n16212) );
  AOI21_X1 U18080 ( .B1(n16213), .B2(n16212), .A(n16211), .ZN(n21999) );
  INV_X1 U18081 ( .A(n21999), .ZN(n16282) );
  OR2_X1 U18082 ( .A1(n20287), .A2(n16214), .ZN(n16216) );
  AND2_X1 U18083 ( .A1(n16216), .A2(n16215), .ZN(n21996) );
  INV_X1 U18084 ( .A(n21996), .ZN(n21827) );
  OAI222_X1 U18085 ( .A1(n16282), .A2(n16219), .B1(n16218), .B2(n20326), .C1(
        n16217), .C2(n21827), .ZN(P1_U2860) );
  NAND2_X1 U18086 ( .A1(n22378), .A2(BUF1_REG_30__SCAN_IN), .ZN(n16222) );
  NOR2_X2 U18087 ( .A1(n22375), .A2(n11319), .ZN(n22377) );
  AOI22_X1 U18088 ( .A1(n22377), .A2(n16220), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n22375), .ZN(n16221) );
  OAI211_X1 U18089 ( .C1(n16223), .C2(n22383), .A(n16222), .B(n16221), .ZN(
        n16224) );
  INV_X1 U18090 ( .A(n16224), .ZN(n16225) );
  OAI21_X1 U18091 ( .B1(n16226), .B2(n16281), .A(n16225), .ZN(P1_U2874) );
  INV_X1 U18092 ( .A(DATAI_29_), .ZN(n22529) );
  NAND2_X1 U18093 ( .A1(n22378), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U18094 ( .A1(n22377), .A2(n16273), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n22375), .ZN(n16227) );
  OAI211_X1 U18095 ( .C1(n22529), .C2(n22383), .A(n16228), .B(n16227), .ZN(
        n16229) );
  INV_X1 U18096 ( .A(n16229), .ZN(n16230) );
  OAI21_X1 U18097 ( .B1(n16231), .B2(n16281), .A(n16230), .ZN(P1_U2875) );
  INV_X1 U18098 ( .A(DATAI_28_), .ZN(n16234) );
  NAND2_X1 U18099 ( .A1(n22378), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16233) );
  AOI22_X1 U18100 ( .A1(n22377), .A2(n16276), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n22375), .ZN(n16232) );
  OAI211_X1 U18101 ( .C1(n16234), .C2(n22383), .A(n16233), .B(n16232), .ZN(
        n16235) );
  INV_X1 U18102 ( .A(n16235), .ZN(n16236) );
  OAI21_X1 U18103 ( .B1(n16308), .B2(n16281), .A(n16236), .ZN(P1_U2876) );
  INV_X1 U18104 ( .A(DATAI_27_), .ZN(n22459) );
  NAND2_X1 U18105 ( .A1(n22378), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16239) );
  AOI22_X1 U18106 ( .A1(n22377), .A2(n16237), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n22375), .ZN(n16238) );
  OAI211_X1 U18107 ( .C1(n22459), .C2(n22383), .A(n16239), .B(n16238), .ZN(
        n16240) );
  INV_X1 U18108 ( .A(n16240), .ZN(n16241) );
  OAI21_X1 U18109 ( .B1(n16242), .B2(n16281), .A(n16241), .ZN(P1_U2877) );
  INV_X1 U18110 ( .A(DATAI_26_), .ZN(n16246) );
  NAND2_X1 U18111 ( .A1(n22378), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16245) );
  AOI22_X1 U18112 ( .A1(n22377), .A2(n16243), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n22375), .ZN(n16244) );
  OAI211_X1 U18113 ( .C1(n16246), .C2(n22383), .A(n16245), .B(n16244), .ZN(
        n16247) );
  INV_X1 U18114 ( .A(n16247), .ZN(n16248) );
  OAI21_X1 U18115 ( .B1(n16328), .B2(n16281), .A(n16248), .ZN(P1_U2878) );
  INV_X1 U18116 ( .A(DATAI_25_), .ZN(n22388) );
  NAND2_X1 U18117 ( .A1(n22378), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16251) );
  AOI22_X1 U18118 ( .A1(n22377), .A2(n16249), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n22375), .ZN(n16250) );
  OAI211_X1 U18119 ( .C1(n22388), .C2(n22383), .A(n16251), .B(n16250), .ZN(
        n16252) );
  INV_X1 U18120 ( .A(n16252), .ZN(n16253) );
  OAI21_X1 U18121 ( .B1(n16254), .B2(n16281), .A(n16253), .ZN(P1_U2879) );
  NAND2_X1 U18122 ( .A1(n22378), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16257) );
  AOI22_X1 U18123 ( .A1(n22377), .A2(n16255), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n22375), .ZN(n16256) );
  OAI211_X1 U18124 ( .C1(n16258), .C2(n22383), .A(n16257), .B(n16256), .ZN(
        n16259) );
  INV_X1 U18125 ( .A(n16259), .ZN(n16260) );
  OAI21_X1 U18126 ( .B1(n22053), .B2(n16281), .A(n16260), .ZN(P1_U2884) );
  INV_X1 U18127 ( .A(DATAI_18_), .ZN(n16264) );
  NAND2_X1 U18128 ( .A1(n22378), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16263) );
  AOI22_X1 U18129 ( .A1(n22377), .A2(n16261), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n22375), .ZN(n16262) );
  OAI211_X1 U18130 ( .C1(n16264), .C2(n22383), .A(n16263), .B(n16262), .ZN(
        n16265) );
  AOI21_X1 U18131 ( .B1(n22033), .B2(n22379), .A(n16265), .ZN(n16266) );
  INV_X1 U18132 ( .A(n16266), .ZN(P1_U2886) );
  INV_X1 U18133 ( .A(DATAI_16_), .ZN(n22247) );
  NAND2_X1 U18134 ( .A1(n22378), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16268) );
  AOI22_X1 U18135 ( .A1(n22377), .A2(n22235), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n22375), .ZN(n16267) );
  OAI211_X1 U18136 ( .C1(n22247), .C2(n22383), .A(n16268), .B(n16267), .ZN(
        n16269) );
  AOI21_X1 U18137 ( .B1(n16376), .B2(n22379), .A(n16269), .ZN(n16270) );
  INV_X1 U18138 ( .A(n16270), .ZN(P1_U2888) );
  INV_X1 U18139 ( .A(n20367), .ZN(n16272) );
  OAI222_X1 U18140 ( .A1(n16281), .A2(n16272), .B1(n16279), .B2(n20211), .C1(
        n16278), .C2(n16271), .ZN(P1_U2889) );
  AOI22_X1 U18141 ( .A1(n16274), .A2(n16273), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n22375), .ZN(n16275) );
  OAI21_X1 U18142 ( .B1(n16412), .B2(n16281), .A(n16275), .ZN(P1_U2891) );
  INV_X1 U18143 ( .A(n16276), .ZN(n16277) );
  OAI222_X1 U18144 ( .A1(n16282), .A2(n16281), .B1(n16280), .B2(n16279), .C1(
        n16278), .C2(n16277), .ZN(P1_U2892) );
  INV_X1 U18145 ( .A(n16283), .ZN(n16285) );
  XNOR2_X1 U18146 ( .A(n13169), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16293) );
  OAI211_X1 U18147 ( .C1(n16285), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16293), .B(n16284), .ZN(n16286) );
  XOR2_X1 U18148 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n16286), .Z(
        n16431) );
  NAND2_X1 U18149 ( .A1(n20379), .A2(n16287), .ZN(n16288) );
  NAND2_X1 U18150 ( .A1(n21923), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16425) );
  OAI211_X1 U18151 ( .C1(n16407), .C2(n16289), .A(n16288), .B(n16425), .ZN(
        n16290) );
  AOI21_X1 U18152 ( .B1(n16291), .B2(n20385), .A(n16290), .ZN(n16292) );
  OAI21_X1 U18153 ( .B1(n16431), .B2(n22113), .A(n16292), .ZN(P1_U2969) );
  XNOR2_X1 U18154 ( .A(n16294), .B(n16293), .ZN(n16440) );
  NOR2_X1 U18155 ( .A1(n21915), .A2(n20255), .ZN(n16436) );
  AOI21_X1 U18156 ( .B1(n20388), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16436), .ZN(n16295) );
  OAI21_X1 U18157 ( .B1(n20395), .B2(n16296), .A(n16295), .ZN(n16297) );
  AOI21_X1 U18158 ( .B1(n16298), .B2(n20385), .A(n16297), .ZN(n16299) );
  OAI21_X1 U18159 ( .B1(n22113), .B2(n16440), .A(n16299), .ZN(P1_U2970) );
  NAND2_X1 U18160 ( .A1(n13169), .A2(n16301), .ZN(n16323) );
  NAND2_X1 U18161 ( .A1(n20391), .A2(n16323), .ZN(n16305) );
  OAI21_X1 U18162 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16302), .A(
        n16305), .ZN(n16304) );
  INV_X1 U18163 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16454) );
  MUX2_X1 U18164 ( .A(n16454), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n13169), .Z(n16303) );
  OAI211_X1 U18165 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16305), .A(
        n16304), .B(n16303), .ZN(n16306) );
  XNOR2_X1 U18166 ( .A(n16306), .B(n16445), .ZN(n16450) );
  NAND2_X1 U18167 ( .A1(n21923), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16444) );
  OAI21_X1 U18168 ( .B1(n16407), .B2(n16307), .A(n16444), .ZN(n16310) );
  NOR2_X1 U18169 ( .A1(n16308), .A2(n16413), .ZN(n16309) );
  AOI211_X1 U18170 ( .C1(n20379), .C2(n16311), .A(n16310), .B(n16309), .ZN(
        n16312) );
  OAI21_X1 U18171 ( .B1(n22113), .B2(n16450), .A(n16312), .ZN(P1_U2971) );
  NAND2_X1 U18172 ( .A1(n16324), .A2(n13181), .ZN(n16314) );
  XNOR2_X1 U18173 ( .A(n13169), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16313) );
  XNOR2_X1 U18174 ( .A(n16314), .B(n16313), .ZN(n16460) );
  NOR2_X1 U18175 ( .A1(n21915), .A2(n20249), .ZN(n16453) );
  AOI21_X1 U18176 ( .B1(n20388), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16453), .ZN(n16315) );
  OAI21_X1 U18177 ( .B1(n20395), .B2(n16316), .A(n16315), .ZN(n16317) );
  AOI21_X1 U18178 ( .B1(n16318), .B2(n20385), .A(n16317), .ZN(n16319) );
  OAI21_X1 U18179 ( .B1(n16460), .B2(n22113), .A(n16319), .ZN(P1_U2972) );
  OAI22_X1 U18180 ( .A1(n16407), .A2(n16320), .B1(n21915), .B2(n20248), .ZN(
        n16321) );
  AOI21_X1 U18181 ( .B1(n16322), .B2(n20379), .A(n16321), .ZN(n16327) );
  NAND3_X1 U18182 ( .A1(n16324), .A2(n16330), .A3(n16323), .ZN(n16325) );
  XNOR2_X1 U18183 ( .A(n16325), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n21898) );
  NAND2_X1 U18184 ( .A1(n21898), .A2(n20392), .ZN(n16326) );
  OAI211_X1 U18185 ( .C1(n16328), .C2(n16413), .A(n16327), .B(n16326), .ZN(
        P1_U2973) );
  NAND2_X1 U18186 ( .A1(n20353), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16329) );
  OAI211_X1 U18187 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16461), .A(
        n16330), .B(n16329), .ZN(n16331) );
  AOI21_X1 U18188 ( .B1(n20391), .B2(n16461), .A(n16331), .ZN(n16332) );
  XNOR2_X1 U18189 ( .A(n16332), .B(n21912), .ZN(n21908) );
  INV_X1 U18190 ( .A(n21908), .ZN(n16338) );
  AOI22_X1 U18191 ( .A1(n20388), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n21923), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n16333) );
  OAI21_X1 U18192 ( .B1(n20395), .B2(n16334), .A(n16333), .ZN(n16335) );
  AOI21_X1 U18193 ( .B1(n16336), .B2(n20385), .A(n16335), .ZN(n16337) );
  OAI21_X1 U18194 ( .B1(n22113), .B2(n16338), .A(n16337), .ZN(P1_U2974) );
  INV_X1 U18195 ( .A(n20391), .ZN(n16339) );
  NAND2_X1 U18196 ( .A1(n16339), .A2(n20389), .ZN(n16341) );
  NAND2_X1 U18197 ( .A1(n20391), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16340) );
  MUX2_X1 U18198 ( .A(n16341), .B(n16340), .S(n13169), .Z(n16342) );
  XNOR2_X1 U18199 ( .A(n16342), .B(n16461), .ZN(n16470) );
  INV_X1 U18200 ( .A(n16343), .ZN(n22380) );
  INV_X1 U18201 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n22099) );
  NAND2_X1 U18202 ( .A1(n20379), .A2(n22106), .ZN(n16344) );
  NAND2_X1 U18203 ( .A1(n21923), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16463) );
  OAI211_X1 U18204 ( .C1(n16407), .C2(n22099), .A(n16344), .B(n16463), .ZN(
        n16345) );
  AOI21_X1 U18205 ( .B1(n22380), .B2(n20385), .A(n16345), .ZN(n16346) );
  OAI21_X1 U18206 ( .B1(n22113), .B2(n16470), .A(n16346), .ZN(P1_U2975) );
  INV_X1 U18207 ( .A(n22224), .ZN(n16353) );
  OAI22_X1 U18208 ( .A1(n16407), .A2(n22074), .B1(n21915), .B2(n22075), .ZN(
        n16347) );
  AOI21_X1 U18209 ( .B1(n22080), .B2(n20379), .A(n16347), .ZN(n16352) );
  NAND2_X1 U18210 ( .A1(n16349), .A2(n16348), .ZN(n16350) );
  XNOR2_X1 U18211 ( .A(n16350), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21892) );
  NAND2_X1 U18212 ( .A1(n21892), .A2(n20392), .ZN(n16351) );
  OAI211_X1 U18213 ( .C1(n16353), .C2(n16413), .A(n16352), .B(n16351), .ZN(
        P1_U2977) );
  OAI21_X1 U18214 ( .B1(n16184), .B2(n16355), .A(n16354), .ZN(n20303) );
  XNOR2_X1 U18215 ( .A(n13169), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16371) );
  NAND2_X1 U18216 ( .A1(n16356), .A2(n16371), .ZN(n16370) );
  OAI21_X1 U18217 ( .B1(n16357), .B2(n13169), .A(n16370), .ZN(n20384) );
  AOI22_X1 U18218 ( .A1(n20384), .A2(n21874), .B1(n13169), .B2(n16370), .ZN(
        n16364) );
  NAND2_X1 U18219 ( .A1(n16359), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16358) );
  OAI211_X1 U18220 ( .C1(n16359), .C2(n13169), .A(n16364), .B(n16358), .ZN(
        n16360) );
  XNOR2_X1 U18221 ( .A(n16360), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16476) );
  NAND2_X1 U18222 ( .A1(n16476), .A2(n20392), .ZN(n16363) );
  INV_X1 U18223 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22072) );
  NOR2_X1 U18224 ( .A1(n21915), .A2(n22072), .ZN(n16487) );
  NOR2_X1 U18225 ( .A1(n20395), .A2(n22068), .ZN(n16361) );
  AOI211_X1 U18226 ( .C1(n20388), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16487), .B(n16361), .ZN(n16362) );
  OAI211_X1 U18227 ( .C1(n16413), .C2(n20303), .A(n16363), .B(n16362), .ZN(
        P1_U2978) );
  OAI21_X1 U18228 ( .B1(n13169), .B2(n21874), .A(n16364), .ZN(n16365) );
  XNOR2_X1 U18229 ( .A(n16365), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n21879) );
  NAND2_X1 U18230 ( .A1(n21879), .A2(n20392), .ZN(n16369) );
  OAI22_X1 U18231 ( .A1(n16407), .A2(n16366), .B1(n21915), .B2(n20239), .ZN(
        n16367) );
  AOI21_X1 U18232 ( .B1(n20379), .B2(n22049), .A(n16367), .ZN(n16368) );
  OAI211_X1 U18233 ( .C1(n16413), .C2(n22053), .A(n16369), .B(n16368), .ZN(
        P1_U2979) );
  OAI21_X1 U18234 ( .B1(n16356), .B2(n16371), .A(n16370), .ZN(n21849) );
  INV_X1 U18235 ( .A(n22030), .ZN(n16373) );
  AOI22_X1 U18236 ( .A1(n20388), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n21923), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16372) );
  OAI21_X1 U18237 ( .B1(n20395), .B2(n16373), .A(n16372), .ZN(n16374) );
  AOI21_X1 U18238 ( .B1(n22033), .B2(n20385), .A(n16374), .ZN(n16375) );
  OAI21_X1 U18239 ( .B1(n22113), .B2(n21849), .A(n16375), .ZN(P1_U2981) );
  INV_X1 U18240 ( .A(n16376), .ZN(n22017) );
  AOI21_X1 U18241 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n13169), .A(
        n20377), .ZN(n16383) );
  INV_X1 U18242 ( .A(n16377), .ZN(n16378) );
  NAND2_X1 U18243 ( .A1(n16379), .A2(n16378), .ZN(n20364) );
  OR2_X1 U18244 ( .A1(n13169), .A2(n21842), .ZN(n20371) );
  NAND2_X1 U18245 ( .A1(n13169), .A2(n21842), .ZN(n16380) );
  NAND2_X1 U18246 ( .A1(n20371), .A2(n16380), .ZN(n20365) );
  NOR2_X1 U18247 ( .A1(n20364), .A2(n20365), .ZN(n16381) );
  AOI21_X1 U18248 ( .B1(n13169), .B2(n21842), .A(n16381), .ZN(n16382) );
  XNOR2_X1 U18249 ( .A(n16383), .B(n16382), .ZN(n21868) );
  NAND2_X1 U18250 ( .A1(n21868), .A2(n20392), .ZN(n16387) );
  OAI22_X1 U18251 ( .A1(n16407), .A2(n16384), .B1(n21915), .B2(n21864), .ZN(
        n16385) );
  AOI21_X1 U18252 ( .B1(n22019), .B2(n20379), .A(n16385), .ZN(n16386) );
  OAI211_X1 U18253 ( .C1(n16413), .C2(n22017), .A(n16387), .B(n16386), .ZN(
        P1_U2983) );
  NOR2_X1 U18254 ( .A1(n16389), .A2(n16390), .ZN(n20374) );
  INV_X1 U18255 ( .A(n16391), .ZN(n16392) );
  AOI22_X1 U18256 ( .A1(n20353), .A2(n21730), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n13169), .ZN(n16393) );
  XNOR2_X1 U18257 ( .A(n16394), .B(n16393), .ZN(n21731) );
  NAND2_X1 U18258 ( .A1(n21731), .A2(n20392), .ZN(n16398) );
  OAI22_X1 U18259 ( .A1(n16407), .A2(n16395), .B1(n21915), .B2(n21721), .ZN(
        n16396) );
  AOI21_X1 U18260 ( .B1(n22010), .B2(n20379), .A(n16396), .ZN(n16397) );
  OAI211_X1 U18261 ( .C1(n16413), .C2(n22008), .A(n16398), .B(n16397), .ZN(
        P1_U2985) );
  OAI21_X1 U18262 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n20353), .ZN(n16399) );
  OAI21_X1 U18263 ( .B1(n16401), .B2(n16400), .A(n16399), .ZN(n20361) );
  INV_X1 U18264 ( .A(n16403), .ZN(n16402) );
  OAI21_X1 U18265 ( .B1(n21822), .B2(n13169), .A(n16402), .ZN(n20360) );
  NOR2_X1 U18266 ( .A1(n20361), .A2(n20360), .ZN(n20359) );
  NOR2_X1 U18267 ( .A1(n16403), .A2(n20359), .ZN(n16405) );
  XNOR2_X1 U18268 ( .A(n16405), .B(n16404), .ZN(n21716) );
  NAND2_X1 U18269 ( .A1(n21716), .A2(n20392), .ZN(n16411) );
  OAI22_X1 U18270 ( .A1(n16407), .A2(n16406), .B1(n21915), .B2(n21711), .ZN(
        n16408) );
  AOI21_X1 U18271 ( .B1(n20379), .B2(n16409), .A(n16408), .ZN(n16410) );
  OAI211_X1 U18272 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        P1_U2986) );
  MUX2_X1 U18273 ( .A(n15729), .B(n16389), .S(n20353), .Z(n16414) );
  NOR2_X1 U18274 ( .A1(n16414), .A2(n15685), .ZN(n20352) );
  AOI21_X1 U18275 ( .B1(n15685), .B2(n16414), .A(n20352), .ZN(n21816) );
  INV_X1 U18276 ( .A(n21816), .ZN(n16420) );
  AOI22_X1 U18277 ( .A1(n20388), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n21923), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16415) );
  OAI21_X1 U18278 ( .B1(n20395), .B2(n16416), .A(n16415), .ZN(n16417) );
  AOI21_X1 U18279 ( .B1(n16418), .B2(n20385), .A(n16417), .ZN(n16419) );
  OAI21_X1 U18280 ( .B1(n16420), .B2(n22113), .A(n16419), .ZN(P1_U2989) );
  INV_X1 U18281 ( .A(n16161), .ZN(n16429) );
  NAND3_X1 U18282 ( .A1(n16455), .A2(n16422), .A3(n16421), .ZN(n16427) );
  OAI21_X1 U18283 ( .B1(n21848), .B2(n16441), .A(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16423) );
  INV_X1 U18284 ( .A(n16423), .ZN(n16424) );
  NAND2_X1 U18285 ( .A1(n16451), .A2(n16424), .ZN(n16438) );
  NAND3_X1 U18286 ( .A1(n16438), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n21783), .ZN(n16426) );
  NAND3_X1 U18287 ( .A1(n16427), .A2(n16426), .A3(n16425), .ZN(n16428) );
  AOI21_X1 U18288 ( .B1(n16429), .B2(n21925), .A(n16428), .ZN(n16430) );
  OAI21_X1 U18289 ( .B1(n16431), .B2(n21862), .A(n16430), .ZN(P1_U3001) );
  INV_X1 U18290 ( .A(n16455), .ZN(n16443) );
  OAI21_X1 U18291 ( .B1(n16443), .B2(n16433), .A(n16432), .ZN(n16437) );
  NOR2_X1 U18292 ( .A1(n16434), .A2(n21906), .ZN(n16435) );
  AOI211_X1 U18293 ( .C1(n16438), .C2(n16437), .A(n16436), .B(n16435), .ZN(
        n16439) );
  OAI21_X1 U18294 ( .B1(n16440), .B2(n21862), .A(n16439), .ZN(P1_U3002) );
  NOR3_X1 U18295 ( .A1(n16443), .A2(n16442), .A3(n16441), .ZN(n16447) );
  OAI21_X1 U18296 ( .B1(n16451), .B2(n16445), .A(n16444), .ZN(n16446) );
  AOI211_X1 U18297 ( .C1(n16448), .C2(n21925), .A(n16447), .B(n16446), .ZN(
        n16449) );
  OAI21_X1 U18298 ( .B1(n16450), .B2(n21862), .A(n16449), .ZN(P1_U3003) );
  NOR2_X1 U18299 ( .A1(n16451), .A2(n16454), .ZN(n16452) );
  AOI211_X1 U18300 ( .C1(n16455), .C2(n16454), .A(n16453), .B(n16452), .ZN(
        n16459) );
  INV_X1 U18301 ( .A(n16456), .ZN(n16457) );
  NAND2_X1 U18302 ( .A1(n16457), .A2(n21925), .ZN(n16458) );
  OAI211_X1 U18303 ( .C1(n16460), .C2(n21862), .A(n16459), .B(n16458), .ZN(
        P1_U3004) );
  INV_X1 U18304 ( .A(n22112), .ZN(n16468) );
  NAND2_X1 U18305 ( .A1(n16461), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16465) );
  NOR2_X1 U18306 ( .A1(n16466), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n21917) );
  INV_X1 U18307 ( .A(n16462), .ZN(n21918) );
  OAI21_X1 U18308 ( .B1(n21917), .B2(n21918), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16464) );
  OAI211_X1 U18309 ( .C1(n16466), .C2(n16465), .A(n16464), .B(n16463), .ZN(
        n16467) );
  AOI21_X1 U18310 ( .B1(n16468), .B2(n21925), .A(n16467), .ZN(n16469) );
  OAI21_X1 U18311 ( .B1(n16470), .B2(n21862), .A(n16469), .ZN(P1_U3007) );
  INV_X1 U18312 ( .A(n16485), .ZN(n16475) );
  AOI21_X1 U18313 ( .B1(n21821), .B2(n16471), .A(n21819), .ZN(n16472) );
  OAI21_X1 U18314 ( .B1(n21826), .B2(n16473), .A(n16472), .ZN(n21847) );
  OAI21_X1 U18315 ( .B1(n21847), .B2(n16474), .A(n21783), .ZN(n21876) );
  INV_X1 U18316 ( .A(n21876), .ZN(n21884) );
  AOI21_X1 U18317 ( .B1(n16475), .B2(n21783), .A(n21884), .ZN(n21893) );
  NAND2_X1 U18318 ( .A1(n16476), .A2(n11156), .ZN(n16489) );
  AOI21_X1 U18319 ( .B1(n16479), .B2(n16478), .A(n16477), .ZN(n22065) );
  NAND3_X1 U18320 ( .A1(n21727), .A2(n21821), .A3(n21779), .ZN(n16481) );
  AOI221_X1 U18321 ( .B1(n21823), .B2(n16481), .C1(n16480), .C2(n16481), .A(
        n21728), .ZN(n21712) );
  NAND4_X1 U18322 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n16482), .A4(n21712), .ZN(
        n21877) );
  OR2_X1 U18323 ( .A1(n21878), .A2(n16483), .ZN(n16484) );
  NAND2_X1 U18324 ( .A1(n21877), .A2(n16484), .ZN(n21883) );
  AND2_X1 U18325 ( .A1(n16485), .A2(n16490), .ZN(n16486) );
  AND2_X1 U18326 ( .A1(n21883), .A2(n16486), .ZN(n21895) );
  AOI211_X1 U18327 ( .C1(n22065), .C2(n21925), .A(n16487), .B(n21895), .ZN(
        n16488) );
  OAI211_X1 U18328 ( .C1(n21893), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        P1_U3010) );
  OAI21_X1 U18329 ( .B1(n21821), .B2(n16491), .A(n21743), .ZN(n21934) );
  NAND2_X1 U18330 ( .A1(n21878), .A2(n21935), .ZN(n16493) );
  AOI22_X1 U18331 ( .A1(n16493), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n11156), .B2(n16492), .ZN(n16497) );
  NAND2_X1 U18332 ( .A1(n21925), .A2(n16494), .ZN(n16495) );
  NAND4_X1 U18333 ( .A1(n21934), .A2(n16497), .A3(n16496), .A4(n16495), .ZN(
        P1_U3031) );
  INV_X1 U18334 ( .A(n16498), .ZN(n16499) );
  NOR2_X1 U18335 ( .A1(n16499), .A2(n17421), .ZN(n22133) );
  AOI21_X1 U18336 ( .B1(n16501), .B2(n16500), .A(n22133), .ZN(n16502) );
  OAI21_X1 U18337 ( .B1(n16503), .B2(n22358), .A(n16502), .ZN(n16504) );
  MUX2_X1 U18338 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16504), .S(
        n17423), .Z(P1_U3478) );
  NOR2_X1 U18339 ( .A1(n17375), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16507) );
  NOR3_X1 U18340 ( .A1(n16505), .A2(n14598), .A3(n17368), .ZN(n16506) );
  AOI211_X1 U18341 ( .C1(n22354), .C2(n17359), .A(n16507), .B(n16506), .ZN(
        n17388) );
  AOI22_X1 U18342 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n21936), .B2(n16508), .ZN(
        n16525) );
  INV_X1 U18343 ( .A(n16525), .ZN(n16511) );
  NOR2_X1 U18344 ( .A1(n22121), .A2(n21743), .ZN(n16526) );
  NOR3_X1 U18345 ( .A1(n14598), .A2(n17368), .A3(n16509), .ZN(n16510) );
  AOI21_X1 U18346 ( .B1(n16511), .B2(n16526), .A(n16510), .ZN(n16512) );
  OAI21_X1 U18347 ( .B1(n17388), .B2(n16529), .A(n16512), .ZN(n16513) );
  MUX2_X1 U18348 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16513), .S(
        n22119), .Z(P1_U3473) );
  OR2_X1 U18349 ( .A1(n16514), .A2(n17378), .ZN(n16524) );
  XNOR2_X1 U18350 ( .A(n17368), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16517) );
  INV_X1 U18351 ( .A(n16517), .ZN(n16527) );
  NAND2_X1 U18352 ( .A1(n17364), .A2(n16527), .ZN(n16521) );
  XNOR2_X1 U18353 ( .A(n12981), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16518) );
  AND2_X1 U18354 ( .A1(n16516), .A2(n16515), .ZN(n17367) );
  AOI22_X1 U18355 ( .A1(n16519), .A2(n16518), .B1(n17367), .B2(n16517), .ZN(
        n16520) );
  OAI21_X1 U18356 ( .B1(n17359), .B2(n16521), .A(n16520), .ZN(n16522) );
  INV_X1 U18357 ( .A(n16522), .ZN(n16523) );
  NAND2_X1 U18358 ( .A1(n16524), .A2(n16523), .ZN(n17384) );
  INV_X1 U18359 ( .A(n17384), .ZN(n16530) );
  AOI22_X1 U18360 ( .A1(n16527), .A2(n22129), .B1(n16526), .B2(n16525), .ZN(
        n16528) );
  OAI21_X1 U18361 ( .B1(n16530), .B2(n16529), .A(n16528), .ZN(n16531) );
  MUX2_X1 U18362 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16531), .S(
        n22119), .Z(P1_U3472) );
  NAND2_X1 U18363 ( .A1(n11600), .A2(n16571), .ZN(n16532) );
  OAI21_X1 U18364 ( .B1(n16571), .B2(n18972), .A(n16532), .ZN(P2_U2856) );
  XNOR2_X1 U18365 ( .A(n16535), .B(n16534), .ZN(n16618) );
  NOR2_X1 U18366 ( .A1(n16536), .A2(n16604), .ZN(n16537) );
  AOI21_X1 U18367 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16604), .A(n16537), .ZN(
        n16538) );
  OAI21_X1 U18368 ( .B1(n16618), .B2(n16606), .A(n16538), .ZN(P2_U2858) );
  INV_X1 U18369 ( .A(n16539), .ZN(n16550) );
  NAND2_X1 U18370 ( .A1(n16550), .A2(n16540), .ZN(n16542) );
  XNOR2_X1 U18371 ( .A(n16542), .B(n16541), .ZN(n16627) );
  NAND2_X1 U18372 ( .A1(n16604), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16548) );
  INV_X1 U18373 ( .A(n16544), .ZN(n16545) );
  AOI21_X1 U18374 ( .B1(n16546), .B2(n16543), .A(n16545), .ZN(n18948) );
  NAND2_X1 U18375 ( .A1(n18948), .A2(n16571), .ZN(n16547) );
  OAI211_X1 U18376 ( .C1(n16627), .C2(n16606), .A(n16548), .B(n16547), .ZN(
        P2_U2859) );
  NAND2_X1 U18377 ( .A1(n16550), .A2(n16549), .ZN(n16551) );
  XOR2_X1 U18378 ( .A(n16552), .B(n16551), .Z(n16637) );
  OAI21_X1 U18379 ( .B1(n16553), .B2(n16554), .A(n16543), .ZN(n16919) );
  NOR2_X1 U18380 ( .A1(n16919), .A2(n16604), .ZN(n16555) );
  AOI21_X1 U18381 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16604), .A(n16555), .ZN(
        n16556) );
  OAI21_X1 U18382 ( .B1(n16637), .B2(n16606), .A(n16556), .ZN(P2_U2860) );
  AND2_X1 U18383 ( .A1(n16568), .A2(n16557), .ZN(n16558) );
  AOI21_X1 U18384 ( .B1(n16561), .B2(n16560), .A(n16559), .ZN(n16641) );
  NAND2_X1 U18385 ( .A1(n16641), .A2(n16596), .ZN(n16563) );
  NAND2_X1 U18386 ( .A1(n16604), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16562) );
  OAI211_X1 U18387 ( .C1(n18924), .C2(n16604), .A(n16563), .B(n16562), .ZN(
        P2_U2861) );
  OAI21_X1 U18388 ( .B1(n16566), .B2(n16565), .A(n16564), .ZN(n16658) );
  NAND2_X1 U18389 ( .A1(n16604), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16573) );
  INV_X1 U18390 ( .A(n16568), .ZN(n16569) );
  AOI21_X1 U18391 ( .B1(n16570), .B2(n16567), .A(n16569), .ZN(n18914) );
  NAND2_X1 U18392 ( .A1(n18914), .A2(n16571), .ZN(n16572) );
  OAI211_X1 U18393 ( .C1(n16658), .C2(n16606), .A(n16573), .B(n16572), .ZN(
        P2_U2862) );
  OAI21_X1 U18394 ( .B1(n16574), .B2(n16575), .A(n13997), .ZN(n16670) );
  OAI21_X1 U18395 ( .B1(n16576), .B2(n16577), .A(n16567), .ZN(n18897) );
  NOR2_X1 U18396 ( .A1(n18897), .A2(n16604), .ZN(n16578) );
  AOI21_X1 U18397 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16604), .A(n16578), .ZN(
        n16579) );
  OAI21_X1 U18398 ( .B1(n16670), .B2(n16606), .A(n16579), .ZN(P2_U2863) );
  NOR2_X1 U18399 ( .A1(n16588), .A2(n16580), .ZN(n16581) );
  OR2_X1 U18400 ( .A1(n16576), .A2(n16581), .ZN(n16968) );
  XOR2_X1 U18401 ( .A(n16583), .B(n16582), .Z(n16679) );
  NAND2_X1 U18402 ( .A1(n16679), .A2(n16596), .ZN(n16585) );
  NAND2_X1 U18403 ( .A1(n16604), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16584) );
  OAI211_X1 U18404 ( .C1(n16968), .C2(n16604), .A(n16585), .B(n16584), .ZN(
        P2_U2864) );
  OAI21_X1 U18405 ( .B1(n16586), .B2(n16587), .A(n16582), .ZN(n19726) );
  AOI21_X1 U18406 ( .B1(n16589), .B2(n16592), .A(n16588), .ZN(n18874) );
  INV_X1 U18407 ( .A(n18874), .ZN(n16982) );
  NOR2_X1 U18408 ( .A1(n16982), .A2(n16604), .ZN(n16590) );
  AOI21_X1 U18409 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n16604), .A(n16590), .ZN(
        n16591) );
  OAI21_X1 U18410 ( .B1(n19726), .B2(n16606), .A(n16591), .ZN(P2_U2865) );
  INV_X1 U18411 ( .A(n16592), .ZN(n16593) );
  AOI21_X1 U18412 ( .B1(n16594), .B2(n15804), .A(n16593), .ZN(n18865) );
  INV_X1 U18413 ( .A(n18865), .ZN(n16993) );
  AOI21_X1 U18414 ( .B1(n16595), .B2(n15806), .A(n16586), .ZN(n16685) );
  NAND2_X1 U18415 ( .A1(n16685), .A2(n16596), .ZN(n16598) );
  NAND2_X1 U18416 ( .A1(n16604), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16597) );
  OAI211_X1 U18417 ( .C1(n16604), .C2(n16993), .A(n16598), .B(n16597), .ZN(
        P2_U2866) );
  OAI21_X1 U18418 ( .B1(n15767), .B2(n16599), .A(n15807), .ZN(n16701) );
  AND2_X1 U18419 ( .A1(n16601), .A2(n16600), .ZN(n16602) );
  OR2_X1 U18420 ( .A1(n16602), .A2(n11285), .ZN(n17017) );
  NOR2_X1 U18421 ( .A1(n17017), .A2(n16604), .ZN(n16603) );
  AOI21_X1 U18422 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16604), .A(n16603), .ZN(
        n16605) );
  OAI21_X1 U18423 ( .B1(n16701), .B2(n16606), .A(n16605), .ZN(P2_U2868) );
  OR2_X1 U18424 ( .A1(n16607), .A2(n16608), .ZN(n16609) );
  INV_X1 U18425 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16615) );
  OAI22_X1 U18426 ( .A1(n16694), .A2(n16612), .B1(n16611), .B2(n19770), .ZN(
        n16613) );
  AOI21_X1 U18427 ( .B1(n19908), .B2(BUF1_REG_29__SCAN_IN), .A(n16613), .ZN(
        n16614) );
  OAI21_X1 U18428 ( .B1(n16696), .B2(n16615), .A(n16614), .ZN(n16616) );
  AOI21_X1 U18429 ( .B1(n18956), .B2(n19822), .A(n16616), .ZN(n16617) );
  OAI21_X1 U18430 ( .B1(n16618), .B2(n19911), .A(n16617), .ZN(P2_U2890) );
  OAI22_X1 U18431 ( .A1(n16694), .A2(n16620), .B1(n16619), .B2(n19770), .ZN(
        n16622) );
  AND2_X1 U18432 ( .A1(n19908), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16621) );
  AOI211_X1 U18433 ( .C1(BUF2_REG_28__SCAN_IN), .C2(n19909), .A(n16622), .B(
        n16621), .ZN(n16626) );
  AOI21_X1 U18434 ( .B1(n16624), .B2(n16623), .A(n16607), .ZN(n18947) );
  NAND2_X1 U18435 ( .A1(n18947), .A2(n19822), .ZN(n16625) );
  OAI211_X1 U18436 ( .C1(n16627), .C2(n19911), .A(n16626), .B(n16625), .ZN(
        P2_U2891) );
  OAI21_X1 U18437 ( .B1(n16640), .B2(n16628), .A(n16623), .ZN(n16629) );
  INV_X1 U18438 ( .A(n16629), .ZN(n18936) );
  INV_X1 U18439 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n16634) );
  OAI22_X1 U18440 ( .A1(n16694), .A2(n16631), .B1(n16630), .B2(n19770), .ZN(
        n16632) );
  AOI21_X1 U18441 ( .B1(n19908), .B2(BUF1_REG_27__SCAN_IN), .A(n16632), .ZN(
        n16633) );
  OAI21_X1 U18442 ( .B1(n16696), .B2(n16634), .A(n16633), .ZN(n16635) );
  AOI21_X1 U18443 ( .B1(n18936), .B2(n19822), .A(n16635), .ZN(n16636) );
  OAI21_X1 U18444 ( .B1(n16637), .B2(n19911), .A(n16636), .ZN(P2_U2892) );
  NOR2_X1 U18445 ( .A1(n16653), .A2(n16638), .ZN(n16639) );
  OR2_X1 U18446 ( .A1(n16640), .A2(n16639), .ZN(n18923) );
  NAND2_X1 U18447 ( .A1(n16641), .A2(n19821), .ZN(n16648) );
  INV_X1 U18448 ( .A(n19908), .ZN(n16645) );
  INV_X1 U18449 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16644) );
  INV_X1 U18450 ( .A(n16694), .ZN(n19907) );
  AOI22_X1 U18451 ( .A1(n19907), .A2(n16642), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19905), .ZN(n16643) );
  OAI21_X1 U18452 ( .B1(n16645), .B2(n16644), .A(n16643), .ZN(n16646) );
  AOI21_X1 U18453 ( .B1(n19909), .B2(BUF2_REG_26__SCAN_IN), .A(n16646), .ZN(
        n16647) );
  OAI211_X1 U18454 ( .C1(n18923), .C2(n19912), .A(n16648), .B(n16647), .ZN(
        P2_U2893) );
  NAND2_X1 U18455 ( .A1(n19908), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16650) );
  NAND2_X1 U18456 ( .A1(n19905), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n16649) );
  OAI211_X1 U18457 ( .C1(n16651), .C2(n16694), .A(n16650), .B(n16649), .ZN(
        n16656) );
  AND2_X1 U18458 ( .A1(n16659), .A2(n16652), .ZN(n16654) );
  OR2_X1 U18459 ( .A1(n16654), .A2(n16653), .ZN(n18912) );
  NOR2_X1 U18460 ( .A1(n18912), .A2(n19912), .ZN(n16655) );
  AOI211_X1 U18461 ( .C1(n19909), .C2(BUF2_REG_25__SCAN_IN), .A(n16656), .B(
        n16655), .ZN(n16657) );
  OAI21_X1 U18462 ( .B1(n19911), .B2(n16658), .A(n16657), .ZN(P2_U2894) );
  INV_X1 U18463 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16667) );
  INV_X1 U18464 ( .A(n16659), .ZN(n16660) );
  AOI21_X1 U18465 ( .B1(n16661), .B2(n16673), .A(n16660), .ZN(n18898) );
  NAND2_X1 U18466 ( .A1(n18898), .A2(n19822), .ZN(n16666) );
  OAI22_X1 U18467 ( .A1(n16694), .A2(n16663), .B1(n16662), .B2(n19770), .ZN(
        n16664) );
  AOI21_X1 U18468 ( .B1(n19908), .B2(BUF1_REG_24__SCAN_IN), .A(n16664), .ZN(
        n16665) );
  OAI211_X1 U18469 ( .C1(n16696), .C2(n16667), .A(n16666), .B(n16665), .ZN(
        n16668) );
  INV_X1 U18470 ( .A(n16668), .ZN(n16669) );
  OAI21_X1 U18471 ( .B1(n19911), .B2(n16670), .A(n16669), .ZN(P2_U2895) );
  OR2_X1 U18472 ( .A1(n16976), .A2(n16671), .ZN(n16672) );
  NAND2_X1 U18473 ( .A1(n16673), .A2(n16672), .ZN(n18895) );
  OAI22_X1 U18474 ( .A1(n16694), .A2(n19527), .B1(n16674), .B2(n19770), .ZN(
        n16675) );
  AOI21_X1 U18475 ( .B1(n19908), .B2(BUF1_REG_23__SCAN_IN), .A(n16675), .ZN(
        n16677) );
  NAND2_X1 U18476 ( .A1(n19909), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16676) );
  OAI211_X1 U18477 ( .C1(n18895), .C2(n19912), .A(n16677), .B(n16676), .ZN(
        n16678) );
  AOI21_X1 U18478 ( .B1(n19821), .B2(n16679), .A(n16678), .ZN(n16680) );
  INV_X1 U18479 ( .A(n16680), .ZN(P2_U2896) );
  INV_X1 U18480 ( .A(n16977), .ZN(n16681) );
  AOI21_X1 U18481 ( .B1(n16682), .B2(n17001), .A(n16681), .ZN(n18864) );
  NAND2_X1 U18482 ( .A1(n18864), .A2(n19822), .ZN(n16689) );
  OAI22_X1 U18483 ( .A1(n16694), .A2(n19772), .B1(n16683), .B2(n19770), .ZN(
        n16684) );
  AOI21_X1 U18484 ( .B1(n19908), .B2(BUF1_REG_21__SCAN_IN), .A(n16684), .ZN(
        n16688) );
  NAND2_X1 U18485 ( .A1(n16685), .A2(n19821), .ZN(n16687) );
  NAND2_X1 U18486 ( .A1(n19909), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16686) );
  NAND4_X1 U18487 ( .A1(n16689), .A2(n16688), .A3(n16687), .A4(n16686), .ZN(
        P2_U2898) );
  XOR2_X1 U18488 ( .A(n16691), .B(n16690), .Z(n18847) );
  NAND2_X1 U18489 ( .A1(n18847), .A2(n19822), .ZN(n16700) );
  OAI22_X1 U18490 ( .A1(n16694), .A2(n16693), .B1(n16692), .B2(n19770), .ZN(
        n16698) );
  INV_X1 U18491 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16695) );
  NOR2_X1 U18492 ( .A1(n16696), .A2(n16695), .ZN(n16697) );
  AOI211_X1 U18493 ( .C1(n19908), .C2(BUF1_REG_19__SCAN_IN), .A(n16698), .B(
        n16697), .ZN(n16699) );
  OAI211_X1 U18494 ( .C1(n19911), .C2(n16701), .A(n16700), .B(n16699), .ZN(
        P2_U2900) );
  NAND2_X1 U18495 ( .A1(n11179), .A2(n11279), .ZN(n16712) );
  XNOR2_X1 U18496 ( .A(n16704), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16705) );
  XNOR2_X1 U18497 ( .A(n16706), .B(n16705), .ZN(n16913) );
  NAND2_X1 U18498 ( .A1(n11167), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16903) );
  NAND2_X1 U18499 ( .A1(n17461), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16707) );
  OAI211_X1 U18500 ( .C1(n17475), .C2(n16708), .A(n16903), .B(n16707), .ZN(
        n16710) );
  NOR2_X1 U18501 ( .A1(n16909), .A2(n17446), .ZN(n16709) );
  OAI21_X1 U18502 ( .B1(n16913), .B2(n17445), .A(n16711), .ZN(P2_U2986) );
  XNOR2_X1 U18503 ( .A(n16714), .B(n16893), .ZN(n16924) );
  INV_X1 U18504 ( .A(n16919), .ZN(n18937) );
  NOR2_X1 U18505 ( .A1(n18830), .A2(n17566), .ZN(n16915) );
  AOI21_X1 U18506 ( .B1(n17461), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16915), .ZN(n16715) );
  OAI21_X1 U18507 ( .B1(n17475), .B2(n16716), .A(n16715), .ZN(n16721) );
  NAND2_X1 U18508 ( .A1(n16717), .A2(n16893), .ZN(n16718) );
  NAND2_X1 U18509 ( .A1(n16719), .A2(n16718), .ZN(n16920) );
  NOR2_X1 U18510 ( .A1(n16920), .A2(n17446), .ZN(n16720) );
  AOI211_X1 U18511 ( .C1(n17457), .C2(n18937), .A(n16721), .B(n16720), .ZN(
        n16722) );
  OAI21_X1 U18512 ( .B1(n16924), .B2(n17445), .A(n16722), .ZN(P2_U2987) );
  OAI21_X1 U18513 ( .B1(n16723), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16717), .ZN(n16939) );
  AND2_X1 U18514 ( .A1(n16727), .A2(n16725), .ZN(n16737) );
  NAND2_X1 U18515 ( .A1(n16724), .A2(n16737), .ZN(n16736) );
  AOI21_X1 U18516 ( .B1(n16736), .B2(n16727), .A(n16726), .ZN(n16728) );
  AOI21_X1 U18517 ( .B1(n11290), .B2(n16736), .A(n16728), .ZN(n16937) );
  NAND2_X1 U18518 ( .A1(n11167), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16928) );
  OAI21_X1 U18519 ( .B1(n17452), .B2(n16729), .A(n16928), .ZN(n16730) );
  AOI21_X1 U18520 ( .B1(n17443), .B2(n11562), .A(n16730), .ZN(n16731) );
  OAI21_X1 U18521 ( .B1(n18924), .B2(n17471), .A(n16731), .ZN(n16732) );
  AOI21_X1 U18522 ( .B1(n16937), .B2(n17462), .A(n16732), .ZN(n16733) );
  OAI21_X1 U18523 ( .B1(n17446), .B2(n16939), .A(n16733), .ZN(P2_U2988) );
  INV_X1 U18524 ( .A(n16723), .ZN(n16735) );
  OAI21_X1 U18525 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16734), .A(
        n16735), .ZN(n16948) );
  OAI21_X1 U18526 ( .B1(n16724), .B2(n16737), .A(n16736), .ZN(n16946) );
  NAND2_X1 U18527 ( .A1(n16946), .A2(n17462), .ZN(n16742) );
  NAND2_X1 U18528 ( .A1(n17443), .A2(n18908), .ZN(n16738) );
  NAND2_X1 U18529 ( .A1(n11167), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16940) );
  OAI211_X1 U18530 ( .C1(n17452), .C2(n16739), .A(n16738), .B(n16940), .ZN(
        n16740) );
  AOI21_X1 U18531 ( .B1(n18914), .B2(n17457), .A(n16740), .ZN(n16741) );
  OAI211_X1 U18532 ( .C1(n16948), .C2(n17446), .A(n16742), .B(n16741), .ZN(
        P2_U2989) );
  INV_X1 U18533 ( .A(n16734), .ZN(n16744) );
  OAI21_X1 U18534 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16743), .A(
        n16744), .ZN(n16959) );
  XNOR2_X1 U18535 ( .A(n16746), .B(n16952), .ZN(n16747) );
  XNOR2_X1 U18536 ( .A(n16745), .B(n16747), .ZN(n16949) );
  NOR2_X1 U18537 ( .A1(n18897), .A2(n17471), .ZN(n16750) );
  NAND2_X1 U18538 ( .A1(n11167), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16954) );
  NAND2_X1 U18539 ( .A1(n17461), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16748) );
  OAI211_X1 U18540 ( .C1(n17475), .C2(n18901), .A(n16954), .B(n16748), .ZN(
        n16749) );
  AOI211_X1 U18541 ( .C1(n16949), .C2(n17462), .A(n16750), .B(n16749), .ZN(
        n16751) );
  OAI21_X1 U18542 ( .B1(n17446), .B2(n16959), .A(n16751), .ZN(P2_U2990) );
  INV_X1 U18543 ( .A(n16753), .ZN(n16755) );
  NAND2_X1 U18544 ( .A1(n16755), .A2(n16754), .ZN(n16756) );
  XNOR2_X1 U18545 ( .A(n16752), .B(n16756), .ZN(n16975) );
  INV_X1 U18546 ( .A(n16968), .ZN(n18889) );
  NAND2_X1 U18547 ( .A1(n17443), .A2(n16757), .ZN(n16758) );
  NAND2_X1 U18548 ( .A1(n11167), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16966) );
  OAI211_X1 U18549 ( .C1(n17452), .C2(n18885), .A(n16758), .B(n16966), .ZN(
        n16759) );
  AOI21_X1 U18550 ( .B1(n18889), .B2(n17457), .A(n16759), .ZN(n16762) );
  AOI21_X1 U18551 ( .B1(n16964), .B2(n16760), .A(n16743), .ZN(n16972) );
  NAND2_X1 U18552 ( .A1(n16972), .A2(n17467), .ZN(n16761) );
  OAI211_X1 U18553 ( .C1(n16975), .C2(n17445), .A(n16762), .B(n16761), .ZN(
        P2_U2991) );
  XNOR2_X1 U18554 ( .A(n16764), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16765) );
  XNOR2_X1 U18555 ( .A(n16763), .B(n16765), .ZN(n16988) );
  NAND2_X1 U18556 ( .A1(n11167), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16981) );
  NAND2_X1 U18557 ( .A1(n17461), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16766) );
  OAI211_X1 U18558 ( .C1(n17475), .C2(n18877), .A(n16981), .B(n16766), .ZN(
        n16767) );
  AOI21_X1 U18559 ( .B1(n18874), .B2(n17457), .A(n16767), .ZN(n16770) );
  NAND2_X1 U18560 ( .A1(n16768), .A2(n11663), .ZN(n16985) );
  NAND3_X1 U18561 ( .A1(n16760), .A2(n17467), .A3(n16985), .ZN(n16769) );
  OAI211_X1 U18562 ( .C1(n16988), .C2(n17445), .A(n16770), .B(n16769), .ZN(
        P2_U2992) );
  INV_X1 U18563 ( .A(n16772), .ZN(n16774) );
  AOI21_X1 U18564 ( .B1(n16772), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16771), .ZN(n16773) );
  INV_X1 U18565 ( .A(n16829), .ZN(n16777) );
  INV_X1 U18566 ( .A(n16820), .ZN(n16778) );
  NAND2_X1 U18567 ( .A1(n11451), .A2(n12697), .ZN(n16783) );
  NAND2_X1 U18568 ( .A1(n16781), .A2(n16780), .ZN(n16782) );
  INV_X1 U18569 ( .A(n16783), .ZN(n16784) );
  NOR2_X1 U18570 ( .A1(n16799), .A2(n16784), .ZN(n16788) );
  NAND2_X1 U18571 ( .A1(n16786), .A2(n16785), .ZN(n16787) );
  XNOR2_X1 U18572 ( .A(n16788), .B(n16787), .ZN(n16998) );
  NAND2_X1 U18573 ( .A1(n17443), .A2(n16789), .ZN(n16790) );
  NAND2_X1 U18574 ( .A1(n11167), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16991) );
  OAI211_X1 U18575 ( .C1(n17452), .C2(n16791), .A(n16790), .B(n16991), .ZN(
        n16795) );
  INV_X1 U18576 ( .A(n16792), .ZN(n16793) );
  OAI21_X1 U18577 ( .B1(n16793), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16768), .ZN(n16994) );
  NOR2_X1 U18578 ( .A1(n16994), .A2(n17446), .ZN(n16794) );
  AOI211_X1 U18579 ( .C1(n18865), .C2(n17457), .A(n16795), .B(n16794), .ZN(
        n16796) );
  OAI21_X1 U18580 ( .B1(n16998), .B2(n17445), .A(n16796), .ZN(P2_U2993) );
  INV_X1 U18581 ( .A(n16798), .ZN(n17082) );
  OAI21_X1 U18582 ( .B1(n16811), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16792), .ZN(n17016) );
  INV_X1 U18583 ( .A(n16799), .ZN(n17000) );
  NAND2_X1 U18584 ( .A1(n16800), .A2(n17012), .ZN(n16999) );
  NAND3_X1 U18585 ( .A1(n17000), .A2(n17462), .A3(n16999), .ZN(n16805) );
  INV_X1 U18586 ( .A(n16801), .ZN(n18855) );
  INV_X1 U18587 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17561) );
  NOR2_X1 U18588 ( .A1(n18830), .A2(n17561), .ZN(n17010) );
  AOI21_X1 U18589 ( .B1(n17461), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17010), .ZN(n16802) );
  OAI21_X1 U18590 ( .B1(n17475), .B2(n18858), .A(n16802), .ZN(n16803) );
  AOI21_X1 U18591 ( .B1(n18855), .B2(n17457), .A(n16803), .ZN(n16804) );
  OAI211_X1 U18592 ( .C1(n17446), .C2(n17016), .A(n16805), .B(n16804), .ZN(
        P2_U2994) );
  NAND2_X1 U18593 ( .A1(n16807), .A2(n16806), .ZN(n16810) );
  INV_X1 U18594 ( .A(n16821), .ZN(n16808) );
  NOR2_X1 U18595 ( .A1(n11258), .A2(n16808), .ZN(n16809) );
  XOR2_X1 U18596 ( .A(n16810), .B(n16809), .Z(n17029) );
  NOR2_X1 U18597 ( .A1(n18830), .A2(n17560), .ZN(n17021) );
  NOR2_X1 U18598 ( .A1(n17452), .A2(n16812), .ZN(n16813) );
  AOI211_X1 U18599 ( .C1(n16814), .C2(n17443), .A(n17021), .B(n16813), .ZN(
        n16815) );
  OAI21_X1 U18600 ( .B1(n17017), .B2(n17471), .A(n16815), .ZN(n16816) );
  AOI21_X1 U18601 ( .B1(n17027), .B2(n17467), .A(n16816), .ZN(n16817) );
  OAI21_X1 U18602 ( .B1(n16832), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n16818), .ZN(n17041) );
  NAND2_X1 U18603 ( .A1(n16821), .A2(n16820), .ZN(n16822) );
  XNOR2_X1 U18604 ( .A(n16819), .B(n16822), .ZN(n17039) );
  INV_X1 U18605 ( .A(n18840), .ZN(n16824) );
  NAND2_X1 U18606 ( .A1(n11167), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n17033) );
  OAI21_X1 U18607 ( .B1(n17452), .B2(n11565), .A(n17033), .ZN(n16823) );
  AOI21_X1 U18608 ( .B1(n17443), .B2(n16824), .A(n16823), .ZN(n16825) );
  OAI21_X1 U18609 ( .B1(n18843), .B2(n17471), .A(n16825), .ZN(n16826) );
  AOI21_X1 U18610 ( .B1(n17039), .B2(n17462), .A(n16826), .ZN(n16827) );
  OAI21_X1 U18611 ( .B1(n17446), .B2(n17041), .A(n16827), .ZN(P2_U2996) );
  NAND2_X1 U18612 ( .A1(n16829), .A2(n16828), .ZN(n16831) );
  XOR2_X1 U18613 ( .A(n16831), .B(n16830), .Z(n17046) );
  INV_X1 U18614 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17074) );
  NOR2_X2 U18615 ( .A1(n16860), .A2(n17074), .ZN(n17052) );
  NAND2_X1 U18616 ( .A1(n11167), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17042) );
  OAI21_X1 U18617 ( .B1(n17452), .B2(n11695), .A(n17042), .ZN(n16833) );
  AOI21_X1 U18618 ( .B1(n17443), .B2(n18821), .A(n16833), .ZN(n16834) );
  OAI21_X1 U18619 ( .B1(n17044), .B2(n17471), .A(n16834), .ZN(n16835) );
  OR2_X1 U18620 ( .A1(n16837), .A2(n16836), .ZN(n17060) );
  NAND3_X1 U18621 ( .A1(n17060), .A2(n16838), .A3(n17462), .ZN(n16844) );
  INV_X1 U18622 ( .A(n18813), .ZN(n17062) );
  INV_X1 U18623 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n18805) );
  NOR2_X1 U18624 ( .A1(n18830), .A2(n18805), .ZN(n17061) );
  AOI21_X1 U18625 ( .B1(n17461), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17061), .ZN(n16839) );
  OAI21_X1 U18626 ( .B1(n17475), .B2(n18811), .A(n16839), .ZN(n16840) );
  AOI21_X1 U18627 ( .B1(n17062), .B2(n17457), .A(n16840), .ZN(n16843) );
  OAI211_X1 U18628 ( .C1(n17052), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16841), .B(n17467), .ZN(n16842) );
  NAND3_X1 U18629 ( .A1(n16844), .A2(n16843), .A3(n16842), .ZN(P2_U2998) );
  INV_X1 U18630 ( .A(n17052), .ZN(n17054) );
  OAI21_X1 U18631 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11381), .A(
        n17054), .ZN(n17080) );
  OAI21_X1 U18632 ( .B1(n16849), .B2(n16846), .A(n11438), .ZN(n16854) );
  NOR2_X1 U18633 ( .A1(n16848), .A2(n16849), .ZN(n16870) );
  OAI21_X1 U18634 ( .B1(n16847), .B2(n16870), .A(n16868), .ZN(n16863) );
  OAI21_X1 U18635 ( .B1(n16850), .B2(n16849), .A(n16852), .ZN(n16851) );
  INV_X1 U18636 ( .A(n16851), .ZN(n16862) );
  NAND2_X1 U18637 ( .A1(n16863), .A2(n16862), .ZN(n16861) );
  NAND2_X1 U18638 ( .A1(n16861), .A2(n16852), .ZN(n16853) );
  XOR2_X1 U18639 ( .A(n16854), .B(n16853), .Z(n17078) );
  NAND2_X1 U18640 ( .A1(n11167), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17070) );
  OAI21_X1 U18641 ( .B1(n17452), .B2(n18793), .A(n17070), .ZN(n16855) );
  AOI21_X1 U18642 ( .B1(n17443), .B2(n18799), .A(n16855), .ZN(n16856) );
  OAI21_X1 U18643 ( .B1(n16857), .B2(n17471), .A(n16856), .ZN(n16858) );
  AOI21_X1 U18644 ( .B1(n17078), .B2(n17462), .A(n16858), .ZN(n16859) );
  OAI21_X1 U18645 ( .B1(n17446), .B2(n17080), .A(n16859), .ZN(P2_U2999) );
  OAI21_X1 U18646 ( .B1(n16874), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16860), .ZN(n17094) );
  OAI21_X1 U18647 ( .B1(n16863), .B2(n16862), .A(n16861), .ZN(n17081) );
  NAND2_X1 U18648 ( .A1(n17081), .A2(n17462), .ZN(n16867) );
  NAND2_X1 U18649 ( .A1(n11167), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n17087) );
  NAND2_X1 U18650 ( .A1(n17461), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16864) );
  OAI211_X1 U18651 ( .C1(n17475), .C2(n18782), .A(n17087), .B(n16864), .ZN(
        n16865) );
  AOI21_X1 U18652 ( .B1(n18788), .B2(n17457), .A(n16865), .ZN(n16866) );
  OAI211_X1 U18653 ( .C1(n17094), .C2(n17446), .A(n16867), .B(n16866), .ZN(
        P2_U3000) );
  INV_X1 U18654 ( .A(n16868), .ZN(n16869) );
  NOR2_X1 U18655 ( .A1(n16870), .A2(n16869), .ZN(n16871) );
  XNOR2_X1 U18656 ( .A(n16847), .B(n16871), .ZN(n17106) );
  NAND2_X1 U18657 ( .A1(n17443), .A2(n18775), .ZN(n16872) );
  NAND2_X1 U18658 ( .A1(n11167), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17095) );
  OAI211_X1 U18659 ( .C1(n17452), .C2(n11694), .A(n16872), .B(n17095), .ZN(
        n16873) );
  AOI21_X1 U18660 ( .B1(n18777), .B2(n17457), .A(n16873), .ZN(n16876) );
  AOI21_X1 U18661 ( .B1(n17099), .B2(n17468), .A(n16874), .ZN(n17103) );
  NAND2_X1 U18662 ( .A1(n17103), .A2(n17467), .ZN(n16875) );
  OAI211_X1 U18663 ( .C1(n17106), .C2(n17445), .A(n16876), .B(n16875), .ZN(
        P2_U3001) );
  NAND2_X1 U18664 ( .A1(n16877), .A2(n16878), .ZN(n16883) );
  INV_X1 U18665 ( .A(n16879), .ZN(n16881) );
  NOR2_X1 U18666 ( .A1(n16881), .A2(n16880), .ZN(n16882) );
  XNOR2_X1 U18667 ( .A(n16883), .B(n16882), .ZN(n17132) );
  NAND2_X1 U18668 ( .A1(n17146), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17133) );
  AOI21_X1 U18669 ( .B1(n17133), .B2(n17123), .A(n11172), .ZN(n17120) );
  NAND2_X1 U18670 ( .A1(n17120), .A2(n17467), .ZN(n16889) );
  NAND2_X1 U18671 ( .A1(n11167), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17125) );
  OAI21_X1 U18672 ( .B1(n17452), .B2(n18747), .A(n17125), .ZN(n16887) );
  NOR2_X1 U18673 ( .A1(n17471), .A2(n18758), .ZN(n16886) );
  AOI211_X1 U18674 ( .C1(n17443), .C2(n18753), .A(n16887), .B(n16886), .ZN(
        n16888) );
  OAI211_X1 U18675 ( .C1(n17132), .C2(n17445), .A(n16889), .B(n16888), .ZN(
        P2_U3003) );
  NAND2_X1 U18676 ( .A1(n18956), .A2(n19003), .ZN(n16897) );
  NAND2_X1 U18677 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16894), .ZN(
        n16904) );
  XNOR2_X1 U18678 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16891) );
  OAI21_X1 U18679 ( .B1(n16904), .B2(n16891), .A(n16890), .ZN(n16892) );
  AOI21_X1 U18680 ( .B1(n18958), .B2(n19017), .A(n16892), .ZN(n16896) );
  NAND2_X1 U18681 ( .A1(n16894), .A2(n16893), .ZN(n16917) );
  NAND2_X1 U18682 ( .A1(n16917), .A2(n16914), .ZN(n16902) );
  NAND2_X1 U18683 ( .A1(n16902), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16895) );
  NAND3_X1 U18684 ( .A1(n16897), .A2(n16896), .A3(n16895), .ZN(n16898) );
  AOI21_X1 U18685 ( .B1(n19007), .B2(n16899), .A(n16898), .ZN(n16900) );
  OAI21_X1 U18686 ( .B1(n16901), .B2(n17166), .A(n16900), .ZN(P2_U3017) );
  INV_X1 U18687 ( .A(n16902), .ZN(n16908) );
  OAI21_X1 U18688 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n16904), .A(
        n16903), .ZN(n16905) );
  AOI21_X1 U18689 ( .B1(n18948), .B2(n19017), .A(n16905), .ZN(n16906) );
  OAI21_X1 U18690 ( .B1(n16908), .B2(n16907), .A(n16906), .ZN(n16911) );
  NOR2_X1 U18691 ( .A1(n16909), .A2(n19015), .ZN(n16910) );
  OAI21_X1 U18692 ( .B1(n16913), .B2(n17166), .A(n16912), .ZN(P2_U3018) );
  INV_X1 U18693 ( .A(n16914), .ZN(n16916) );
  AOI21_X1 U18694 ( .B1(n16916), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16915), .ZN(n16918) );
  OAI211_X1 U18695 ( .C1(n16919), .C2(n18991), .A(n16918), .B(n16917), .ZN(
        n16922) );
  NOR2_X1 U18696 ( .A1(n16920), .A2(n19015), .ZN(n16921) );
  AOI211_X1 U18697 ( .C1(n19003), .C2(n18936), .A(n16922), .B(n16921), .ZN(
        n16923) );
  OAI21_X1 U18698 ( .B1(n16924), .B2(n17166), .A(n16923), .ZN(P2_U3019) );
  INV_X1 U18699 ( .A(n16925), .ZN(n16926) );
  NAND2_X1 U18700 ( .A1(n16926), .A2(n16931), .ZN(n16927) );
  OAI211_X1 U18701 ( .C1(n18924), .C2(n18991), .A(n16928), .B(n16927), .ZN(
        n16934) );
  NAND2_X1 U18702 ( .A1(n16929), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16930) );
  OR2_X1 U18703 ( .A1(n16953), .A2(n16930), .ZN(n16943) );
  NAND2_X1 U18704 ( .A1(n16950), .A2(n17122), .ZN(n16932) );
  AOI21_X1 U18705 ( .B1(n16943), .B2(n16932), .A(n16931), .ZN(n16933) );
  NOR2_X1 U18706 ( .A1(n16934), .A2(n16933), .ZN(n16935) );
  OAI21_X1 U18707 ( .B1(n18923), .B2(n19020), .A(n16935), .ZN(n16936) );
  AOI21_X1 U18708 ( .B1(n16937), .B2(n19024), .A(n16936), .ZN(n16938) );
  OAI21_X1 U18709 ( .B1(n19015), .B2(n16939), .A(n16938), .ZN(P2_U3020) );
  INV_X1 U18710 ( .A(n16940), .ZN(n16942) );
  AND3_X1 U18711 ( .A1(n16950), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17122), .ZN(n16941) );
  AOI211_X1 U18712 ( .C1(n18914), .C2(n19017), .A(n16942), .B(n16941), .ZN(
        n16944) );
  OAI211_X1 U18713 ( .C1(n18912), .C2(n19020), .A(n16944), .B(n16943), .ZN(
        n16945) );
  AOI21_X1 U18714 ( .B1(n16946), .B2(n19024), .A(n16945), .ZN(n16947) );
  OAI21_X1 U18715 ( .B1(n19015), .B2(n16948), .A(n16947), .ZN(P2_U3021) );
  NAND2_X1 U18716 ( .A1(n16949), .A2(n19024), .ZN(n16958) );
  INV_X1 U18717 ( .A(n16950), .ZN(n16951) );
  AOI21_X1 U18718 ( .B1(n16953), .B2(n16952), .A(n16951), .ZN(n16956) );
  OAI21_X1 U18719 ( .B1(n18897), .B2(n18991), .A(n16954), .ZN(n16955) );
  AOI211_X1 U18720 ( .C1(n18898), .C2(n19003), .A(n16956), .B(n16955), .ZN(
        n16957) );
  OAI211_X1 U18721 ( .C1(n16959), .C2(n19015), .A(n16958), .B(n16957), .ZN(
        P2_U3022) );
  INV_X1 U18722 ( .A(n18895), .ZN(n16971) );
  NAND2_X1 U18723 ( .A1(n17156), .A2(n17005), .ZN(n17069) );
  OR2_X1 U18724 ( .A1(n17069), .A2(n17004), .ZN(n17019) );
  NOR2_X1 U18725 ( .A1(n17019), .A2(n16960), .ZN(n16990) );
  NAND3_X1 U18726 ( .A1(n16990), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n11663), .ZN(n16979) );
  OAI211_X1 U18727 ( .C1(n19001), .C2(n16961), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17121), .ZN(n16989) );
  NAND2_X1 U18728 ( .A1(n16989), .A2(n17122), .ZN(n16962) );
  AOI21_X1 U18729 ( .B1(n16979), .B2(n16962), .A(n16964), .ZN(n16970) );
  INV_X1 U18730 ( .A(n16963), .ZN(n16965) );
  NAND3_X1 U18731 ( .A1(n16990), .A2(n16965), .A3(n16964), .ZN(n16967) );
  OAI211_X1 U18732 ( .C1(n16968), .C2(n18991), .A(n16967), .B(n16966), .ZN(
        n16969) );
  AOI211_X1 U18733 ( .C1(n16971), .C2(n19003), .A(n16970), .B(n16969), .ZN(
        n16974) );
  NAND2_X1 U18734 ( .A1(n16972), .A2(n19007), .ZN(n16973) );
  OAI211_X1 U18735 ( .C1(n16975), .C2(n17166), .A(n16974), .B(n16973), .ZN(
        P2_U3023) );
  AOI21_X1 U18736 ( .B1(n16978), .B2(n16977), .A(n16976), .ZN(n19728) );
  INV_X1 U18737 ( .A(n16979), .ZN(n16984) );
  NAND3_X1 U18738 ( .A1(n16989), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17122), .ZN(n16980) );
  OAI211_X1 U18739 ( .C1(n16982), .C2(n18991), .A(n16981), .B(n16980), .ZN(
        n16983) );
  AOI211_X1 U18740 ( .C1(n19728), .C2(n19003), .A(n16984), .B(n16983), .ZN(
        n16987) );
  NAND3_X1 U18741 ( .A1(n16760), .A2(n19007), .A3(n16985), .ZN(n16986) );
  OAI211_X1 U18742 ( .C1(n16988), .C2(n17166), .A(n16987), .B(n16986), .ZN(
        P2_U3024) );
  OAI21_X1 U18743 ( .B1(n16990), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16989), .ZN(n16992) );
  OAI211_X1 U18744 ( .C1(n18991), .C2(n16993), .A(n16992), .B(n16991), .ZN(
        n16996) );
  NOR2_X1 U18745 ( .A1(n16994), .A2(n19015), .ZN(n16995) );
  AOI211_X1 U18746 ( .C1(n19003), .C2(n18864), .A(n16996), .B(n16995), .ZN(
        n16997) );
  OAI21_X1 U18747 ( .B1(n16998), .B2(n17166), .A(n16997), .ZN(P2_U3025) );
  NAND3_X1 U18748 ( .A1(n17000), .A2(n19024), .A3(n16999), .ZN(n17015) );
  AOI21_X1 U18749 ( .B1(n17003), .B2(n17002), .A(n11458), .ZN(n19823) );
  NOR2_X1 U18750 ( .A1(n17019), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17034) );
  INV_X1 U18751 ( .A(n17004), .ZN(n17007) );
  OR2_X1 U18752 ( .A1(n19001), .A2(n17005), .ZN(n17006) );
  AND2_X1 U18753 ( .A1(n17006), .A2(n17121), .ZN(n17050) );
  OAI21_X1 U18754 ( .B1(n17007), .B2(n19001), .A(n17050), .ZN(n17036) );
  NOR2_X1 U18755 ( .A1(n17034), .A2(n17036), .ZN(n17025) );
  AOI21_X1 U18756 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17012), .A(
        n17024), .ZN(n17008) );
  AOI211_X1 U18757 ( .C1(n17024), .C2(n17012), .A(n17008), .B(n17019), .ZN(
        n17009) );
  AOI211_X1 U18758 ( .C1(n18855), .C2(n19017), .A(n17010), .B(n17009), .ZN(
        n17011) );
  OAI21_X1 U18759 ( .B1(n17025), .B2(n17012), .A(n17011), .ZN(n17013) );
  AOI21_X1 U18760 ( .B1(n19823), .B2(n19003), .A(n17013), .ZN(n17014) );
  OAI211_X1 U18761 ( .C1(n17016), .C2(n19015), .A(n17015), .B(n17014), .ZN(
        P2_U3026) );
  NAND2_X1 U18762 ( .A1(n18847), .A2(n19003), .ZN(n17023) );
  INV_X1 U18763 ( .A(n17017), .ZN(n18848) );
  NOR3_X1 U18764 ( .A1(n17019), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n17018), .ZN(n17020) );
  AOI211_X1 U18765 ( .C1(n18848), .C2(n19017), .A(n17021), .B(n17020), .ZN(
        n17022) );
  OAI211_X1 U18766 ( .C1(n17025), .C2(n17024), .A(n17023), .B(n17022), .ZN(
        n17026) );
  AOI21_X1 U18767 ( .B1(n17027), .B2(n19007), .A(n17026), .ZN(n17028) );
  NOR2_X1 U18768 ( .A1(n17031), .A2(n17030), .ZN(n17032) );
  OR2_X1 U18769 ( .A1(n16690), .A2(n17032), .ZN(n19913) );
  OAI21_X1 U18770 ( .B1(n18843), .B2(n18991), .A(n17033), .ZN(n17035) );
  AOI211_X1 U18771 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n17036), .A(
        n17035), .B(n17034), .ZN(n17037) );
  OAI21_X1 U18772 ( .B1(n19913), .B2(n19020), .A(n17037), .ZN(n17038) );
  AOI21_X1 U18773 ( .B1(n17039), .B2(n19024), .A(n17038), .ZN(n17040) );
  OAI21_X1 U18774 ( .B1(n19015), .B2(n17041), .A(n17040), .ZN(P2_U3028) );
  NAND2_X1 U18775 ( .A1(n18825), .A2(n19003), .ZN(n17043) );
  OAI211_X1 U18776 ( .C1(n18991), .C2(n17044), .A(n17043), .B(n17042), .ZN(
        n17045) );
  AOI21_X1 U18777 ( .B1(n17046), .B2(n19024), .A(n17045), .ZN(n17058) );
  NOR2_X1 U18778 ( .A1(n19007), .A2(n17047), .ZN(n17051) );
  NAND2_X1 U18779 ( .A1(n17048), .A2(n17074), .ZN(n17049) );
  AND2_X1 U18780 ( .A1(n17050), .A2(n17049), .ZN(n17072) );
  OAI21_X1 U18781 ( .B1(n17052), .B2(n17051), .A(n17072), .ZN(n17066) );
  AOI21_X1 U18782 ( .B1(n19001), .B2(n19015), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17053) );
  OAI21_X1 U18783 ( .B1(n17066), .B2(n17053), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17057) );
  NAND3_X1 U18784 ( .A1(n17055), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17059), .ZN(n17056) );
  NAND3_X1 U18785 ( .A1(n17056), .A2(n17057), .A3(n17058), .ZN(P2_U3029) );
  INV_X1 U18786 ( .A(n17059), .ZN(n17068) );
  NAND3_X1 U18787 ( .A1(n17060), .A2(n16838), .A3(n19024), .ZN(n17064) );
  AOI21_X1 U18788 ( .B1(n17062), .B2(n19017), .A(n17061), .ZN(n17063) );
  OAI211_X1 U18789 ( .C1(n19020), .C2(n18812), .A(n17064), .B(n17063), .ZN(
        n17065) );
  AOI21_X1 U18790 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17066), .A(
        n17065), .ZN(n17067) );
  OAI21_X1 U18791 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17068), .A(
        n17067), .ZN(P2_U3030) );
  INV_X1 U18792 ( .A(n17069), .ZN(n17075) );
  NAND2_X1 U18793 ( .A1(n18801), .A2(n19017), .ZN(n17071) );
  OAI211_X1 U18794 ( .C1(n17072), .C2(n17074), .A(n17071), .B(n17070), .ZN(
        n17073) );
  AOI21_X1 U18795 ( .B1(n17075), .B2(n17074), .A(n17073), .ZN(n17076) );
  OAI21_X1 U18796 ( .B1(n18804), .B2(n19020), .A(n17076), .ZN(n17077) );
  AOI21_X1 U18797 ( .B1(n17078), .B2(n19024), .A(n17077), .ZN(n17079) );
  OAI21_X1 U18798 ( .B1(n19015), .B2(n17080), .A(n17079), .ZN(P2_U3031) );
  NAND2_X1 U18799 ( .A1(n17081), .A2(n19024), .ZN(n17093) );
  NAND2_X1 U18800 ( .A1(n17156), .A2(n17082), .ZN(n17086) );
  OR2_X1 U18801 ( .A1(n17086), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17114) );
  NAND2_X1 U18802 ( .A1(n17121), .A2(n17082), .ZN(n17083) );
  NAND2_X1 U18803 ( .A1(n17122), .A2(n17083), .ZN(n17107) );
  AND2_X1 U18804 ( .A1(n17114), .A2(n17107), .ZN(n17100) );
  OR2_X1 U18805 ( .A1(n17086), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17096) );
  AOI21_X1 U18806 ( .B1(n17100), .B2(n17096), .A(n17084), .ZN(n17091) );
  NAND2_X1 U18807 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17085) );
  OR3_X1 U18808 ( .A1(n17086), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17085), .ZN(n17088) );
  OAI211_X1 U18809 ( .C1(n17089), .C2(n18991), .A(n17088), .B(n17087), .ZN(
        n17090) );
  AOI211_X1 U18810 ( .C1(n18787), .C2(n19003), .A(n17091), .B(n17090), .ZN(
        n17092) );
  OAI211_X1 U18811 ( .C1(n17094), .C2(n19015), .A(n17093), .B(n17092), .ZN(
        P2_U3032) );
  INV_X1 U18812 ( .A(n18780), .ZN(n17102) );
  OAI21_X1 U18813 ( .B1(n17096), .B2(n17464), .A(n17095), .ZN(n17097) );
  AOI21_X1 U18814 ( .B1(n18777), .B2(n19017), .A(n17097), .ZN(n17098) );
  OAI21_X1 U18815 ( .B1(n17100), .B2(n17099), .A(n17098), .ZN(n17101) );
  AOI21_X1 U18816 ( .B1(n17102), .B2(n19003), .A(n17101), .ZN(n17105) );
  NAND2_X1 U18817 ( .A1(n17103), .A2(n19007), .ZN(n17104) );
  OAI211_X1 U18818 ( .C1(n17106), .C2(n17166), .A(n17105), .B(n17104), .ZN(
        P2_U3033) );
  INV_X1 U18819 ( .A(n17107), .ZN(n17108) );
  AOI21_X1 U18820 ( .B1(n17468), .B2(n19007), .A(n17108), .ZN(n17119) );
  XNOR2_X1 U18821 ( .A(n17109), .B(n17464), .ZN(n17110) );
  XNOR2_X1 U18822 ( .A(n16772), .B(n17110), .ZN(n17463) );
  INV_X1 U18823 ( .A(n18764), .ZN(n17112) );
  INV_X1 U18824 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n17555) );
  NOR2_X1 U18825 ( .A1(n17555), .A2(n18830), .ZN(n17111) );
  AOI21_X1 U18826 ( .B1(n17112), .B2(n19017), .A(n17111), .ZN(n17113) );
  OAI211_X1 U18827 ( .C1(n18763), .C2(n19020), .A(n17114), .B(n17113), .ZN(
        n17117) );
  INV_X1 U18828 ( .A(n17468), .ZN(n17115) );
  NOR3_X1 U18829 ( .A1(n17115), .A2(n17465), .A3(n19015), .ZN(n17116) );
  AOI211_X1 U18830 ( .C1(n19024), .C2(n17463), .A(n17117), .B(n17116), .ZN(
        n17118) );
  OAI21_X1 U18831 ( .B1(n17119), .B2(n17464), .A(n17118), .ZN(P2_U3034) );
  NAND2_X1 U18832 ( .A1(n17120), .A2(n19007), .ZN(n17131) );
  NAND3_X1 U18833 ( .A1(n17156), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17140), .ZN(n17139) );
  NAND2_X1 U18834 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17121), .ZN(
        n17155) );
  NAND2_X1 U18835 ( .A1(n17122), .A2(n17155), .ZN(n17141) );
  AOI21_X1 U18836 ( .B1(n17139), .B2(n17141), .A(n17123), .ZN(n17129) );
  AND3_X1 U18837 ( .A1(n17156), .A2(n17124), .A3(n17123), .ZN(n17128) );
  NOR2_X1 U18838 ( .A1(n18991), .A2(n18758), .ZN(n17127) );
  OAI21_X1 U18839 ( .B1(n19020), .B2(n18746), .A(n17125), .ZN(n17126) );
  NOR4_X1 U18840 ( .A1(n17129), .A2(n17128), .A3(n17127), .A4(n17126), .ZN(
        n17130) );
  OAI211_X1 U18841 ( .C1(n17132), .C2(n17166), .A(n17131), .B(n17130), .ZN(
        P2_U3035) );
  OAI21_X1 U18842 ( .B1(n17146), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17133), .ZN(n17454) );
  NAND2_X1 U18843 ( .A1(n17134), .A2(n17149), .ZN(n17137) );
  NAND2_X1 U18844 ( .A1(n11312), .A2(n17135), .ZN(n17136) );
  XNOR2_X1 U18845 ( .A(n17137), .B(n17136), .ZN(n17458) );
  NAND2_X1 U18846 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n11167), .ZN(n17138) );
  OAI211_X1 U18847 ( .C1(n17141), .C2(n17140), .A(n17139), .B(n17138), .ZN(
        n17144) );
  OAI22_X1 U18848 ( .A1(n19020), .A2(n17142), .B1(n18991), .B2(n18744), .ZN(
        n17143) );
  AOI211_X1 U18849 ( .C1(n17458), .C2(n19024), .A(n17144), .B(n17143), .ZN(
        n17145) );
  OAI21_X1 U18850 ( .B1(n17454), .B2(n19015), .A(n17145), .ZN(P2_U3036) );
  INV_X1 U18851 ( .A(n17146), .ZN(n17147) );
  INV_X1 U18852 ( .A(n17149), .ZN(n17148) );
  OR2_X1 U18853 ( .A1(n17134), .A2(n17148), .ZN(n17154) );
  AND2_X1 U18854 ( .A1(n17150), .A2(n17149), .ZN(n17151) );
  OR2_X1 U18855 ( .A1(n17152), .A2(n17151), .ZN(n17153) );
  NAND2_X1 U18856 ( .A1(n17154), .A2(n17153), .ZN(n17444) );
  INV_X1 U18857 ( .A(n17444), .ZN(n17162) );
  INV_X1 U18858 ( .A(n17449), .ZN(n18727) );
  OAI21_X1 U18859 ( .B1(n17156), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17155), .ZN(n17160) );
  INV_X1 U18860 ( .A(n18728), .ZN(n17158) );
  INV_X1 U18861 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n17553) );
  NOR2_X1 U18862 ( .A1(n17553), .A2(n18830), .ZN(n17157) );
  AOI21_X1 U18863 ( .B1(n19003), .B2(n17158), .A(n17157), .ZN(n17159) );
  OAI211_X1 U18864 ( .C1(n18991), .C2(n18727), .A(n17160), .B(n17159), .ZN(
        n17161) );
  AOI21_X1 U18865 ( .B1(n17162), .B2(n19024), .A(n17161), .ZN(n17163) );
  OAI21_X1 U18866 ( .B1(n17447), .B2(n19015), .A(n17163), .ZN(P2_U3037) );
  OAI21_X1 U18867 ( .B1(n19015), .B2(n17165), .A(n17164), .ZN(n17169) );
  NOR2_X1 U18868 ( .A1(n17167), .A2(n17166), .ZN(n17168) );
  AOI211_X1 U18869 ( .C1(n17170), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17169), .B(n17168), .ZN(n17175) );
  AOI22_X1 U18870 ( .A1(n19017), .A2(n18648), .B1(n19003), .B2(n18646), .ZN(
        n17174) );
  INV_X1 U18871 ( .A(n19001), .ZN(n17172) );
  OAI211_X1 U18872 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n17172), .B(n17171), .ZN(n17173) );
  NAND3_X1 U18873 ( .A1(n17175), .A2(n17174), .A3(n17173), .ZN(P2_U3045) );
  OAI222_X1 U18874 ( .A1(n17179), .A2(n17488), .B1(n17178), .B2(n17177), .C1(
        n17176), .C2(n19034), .ZN(n17180) );
  MUX2_X1 U18875 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n17180), .S(
        n18988), .Z(P2_U3600) );
  INV_X1 U18876 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21676) );
  NOR2_X1 U18877 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21676), .ZN(
        n19086) );
  INV_X1 U18878 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21158) );
  INV_X1 U18879 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21668) );
  NOR2_X1 U18880 ( .A1(n21158), .A2(n21668), .ZN(n17960) );
  NAND2_X1 U18881 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17960), .ZN(n21675) );
  INV_X1 U18882 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20576) );
  OAI21_X1 U18883 ( .B1(n21190), .B2(n21182), .A(n20576), .ZN(n17318) );
  NOR2_X1 U18884 ( .A1(n18028), .A2(n17318), .ZN(n17961) );
  INV_X1 U18885 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21688) );
  NAND2_X1 U18886 ( .A1(n21158), .A2(n21668), .ZN(n20463) );
  INV_X1 U18887 ( .A(n20463), .ZN(n21681) );
  NOR2_X1 U18888 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21676), .ZN(
        n21680) );
  INV_X1 U18889 ( .A(n21680), .ZN(n17181) );
  OAI21_X1 U18890 ( .B1(n21681), .B2(n17960), .A(n17181), .ZN(n19087) );
  NAND2_X1 U18891 ( .A1(n21688), .A2(n19087), .ZN(n19294) );
  INV_X1 U18892 ( .A(n21675), .ZN(n17330) );
  NAND2_X1 U18893 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17330), .ZN(n17316) );
  OAI211_X1 U18894 ( .C1(n21675), .C2(n17961), .A(n19294), .B(n17316), .ZN(
        n17332) );
  INV_X1 U18895 ( .A(n17332), .ZN(n18537) );
  NOR2_X1 U18896 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17960), .ZN(n20467) );
  INV_X1 U18897 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22146) );
  NOR2_X1 U18898 ( .A1(n21158), .A2(n22146), .ZN(n18437) );
  INV_X1 U18899 ( .A(n18437), .ZN(n18488) );
  NAND2_X1 U18900 ( .A1(n20467), .A2(n18488), .ZN(n17183) );
  NOR2_X1 U18901 ( .A1(n21640), .A2(n21646), .ZN(n19085) );
  AOI21_X1 U18902 ( .B1(n21676), .B2(n17183), .A(n19085), .ZN(n17182) );
  NOR3_X1 U18903 ( .A1(n19086), .A2(n18537), .A3(n17182), .ZN(n18536) );
  NOR3_X1 U18904 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n22146), .ZN(n19107) );
  NAND2_X1 U18905 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17184) );
  AOI21_X1 U18906 ( .B1(n17184), .B2(n17183), .A(n18537), .ZN(n18538) );
  INV_X1 U18907 ( .A(n19294), .ZN(n19422) );
  NAND2_X1 U18908 ( .A1(n19422), .A2(n19107), .ZN(n19252) );
  INV_X2 U18909 ( .A(n19252), .ZN(n19421) );
  OAI22_X1 U18910 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19107), .B1(
        n18538), .B2(n19421), .ZN(n17185) );
  AOI22_X1 U18911 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18536), .B1(
        n17185), .B2(n21646), .ZN(P3_U2865) );
  NOR2_X1 U18912 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21688), .ZN(n21670) );
  NAND2_X1 U18913 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21670), .ZN(n21665) );
  AOI22_X1 U18914 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U18915 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U18916 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11212), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17187) );
  NOR2_X2 U18917 ( .A1(n21633), .A2(n21173), .ZN(n18018) );
  INV_X2 U18918 ( .A(n11218), .ZN(n18016) );
  AOI22_X1 U18919 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17186) );
  NAND4_X1 U18920 ( .A1(n17189), .A2(n17188), .A3(n17187), .A4(n17186), .ZN(
        n17198) );
  AOI22_X1 U18921 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17196) );
  NOR2_X2 U18922 ( .A1(n21194), .A2(n20541), .ZN(n17232) );
  AOI22_X1 U18923 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11208), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U18924 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U18925 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17193) );
  NAND4_X1 U18926 ( .A1(n17196), .A2(n17195), .A3(n17194), .A4(n17193), .ZN(
        n17197) );
  AOI22_X1 U18927 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17232), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U18928 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U18929 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18018), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17200) );
  BUF_X4 U18930 ( .A(n18017), .Z(n17992) );
  AOI22_X1 U18931 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17199) );
  NAND4_X1 U18932 ( .A1(n17202), .A2(n17201), .A3(n17200), .A4(n17199), .ZN(
        n17208) );
  AOI22_X1 U18933 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U18934 ( .A1(n18023), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17205) );
  BUF_X1 U18935 ( .A(n17233), .Z(n18061) );
  AOI22_X1 U18936 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U18937 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17203) );
  NAND4_X1 U18938 ( .A1(n17206), .A2(n17205), .A3(n17204), .A4(n17203), .ZN(
        n17207) );
  INV_X1 U18939 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17333) );
  OAI22_X1 U18940 ( .A1(n21191), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21646), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17214) );
  OAI22_X1 U18941 ( .A1(n21190), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n21640), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17300) );
  NAND2_X1 U18942 ( .A1(n21637), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17301) );
  NOR2_X1 U18943 ( .A1(n17300), .A2(n17301), .ZN(n17209) );
  AOI21_X1 U18944 ( .B1(n21640), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n17209), .ZN(n17215) );
  OR2_X1 U18945 ( .A1(n17214), .A2(n17215), .ZN(n17210) );
  OAI21_X1 U18946 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21191), .A(
        n17210), .ZN(n17211) );
  OAI22_X1 U18947 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17333), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17211), .ZN(n17217) );
  NOR2_X1 U18948 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17333), .ZN(
        n17212) );
  NAND2_X1 U18949 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n17211), .ZN(
        n17216) );
  AOI22_X1 U18950 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17217), .B1(
        n17212), .B2(n17216), .ZN(n17220) );
  OAI21_X1 U18951 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21637), .A(
        n17301), .ZN(n17979) );
  NOR2_X1 U18952 ( .A1(n17300), .A2(n17979), .ZN(n17219) );
  NAND2_X1 U18953 ( .A1(n17215), .A2(n17214), .ZN(n17213) );
  OAI211_X1 U18954 ( .C1(n17215), .C2(n17214), .A(n17220), .B(n17213), .ZN(
        n17980) );
  INV_X1 U18955 ( .A(n17980), .ZN(n17303) );
  AND2_X1 U18956 ( .A1(n17216), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17218) );
  OAI22_X1 U18957 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20576), .B1(
        n17218), .B2(n17217), .ZN(n17302) );
  AOI211_X1 U18958 ( .C1(n17220), .C2(n17219), .A(n17303), .B(n17302), .ZN(
        n21653) );
  NAND2_X1 U18959 ( .A1(n21214), .A2(n21653), .ZN(n21207) );
  AOI22_X1 U18960 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18014), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U18961 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17230) );
  INV_X1 U18962 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19169) );
  AOI22_X1 U18963 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17222) );
  OAI21_X1 U18964 ( .B1(n17238), .B2(n19169), .A(n17222), .ZN(n17228) );
  AOI22_X1 U18965 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U18966 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U18967 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11213), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U18968 ( .A1(n11211), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17223) );
  NAND4_X1 U18969 ( .A1(n17226), .A2(n17225), .A3(n17224), .A4(n17223), .ZN(
        n17227) );
  AOI22_X1 U18970 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U18971 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U18972 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U18973 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17234) );
  NAND4_X1 U18974 ( .A1(n17237), .A2(n17236), .A3(n17235), .A4(n17234), .ZN(
        n17244) );
  INV_X2 U18975 ( .A(n17238), .ZN(n18031) );
  AOI22_X1 U18976 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18031), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U18977 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U18978 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U18979 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17239) );
  NAND4_X1 U18980 ( .A1(n17242), .A2(n17241), .A3(n17240), .A4(n17239), .ZN(
        n17243) );
  AOI22_X1 U18981 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U18982 ( .A1(n11215), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U18983 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18018), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U18984 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17245) );
  NAND4_X1 U18985 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        n17254) );
  AOI22_X1 U18986 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U18987 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U18988 ( .A1(n17232), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U18989 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17249) );
  NAND4_X1 U18990 ( .A1(n17252), .A2(n17251), .A3(n17250), .A4(n17249), .ZN(
        n17253) );
  AOI22_X1 U18991 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U18992 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17262) );
  INV_X1 U18993 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19209) );
  AOI22_X1 U18994 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U18995 ( .B1(n17238), .B2(n19209), .A(n17255), .ZN(n17261) );
  AOI22_X1 U18996 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17232), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U18997 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U18998 ( .A1(n18023), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U18999 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17256) );
  NAND4_X1 U19000 ( .A1(n17259), .A2(n17258), .A3(n17257), .A4(n17256), .ZN(
        n17260) );
  AOI22_X1 U19001 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U19002 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17267) );
  AOI22_X1 U19003 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18018), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U19004 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17265) );
  NAND4_X1 U19005 ( .A1(n17268), .A2(n17267), .A3(n17266), .A4(n17265), .ZN(
        n17274) );
  AOI22_X1 U19006 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U19007 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18023), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U19008 ( .A1(n17232), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U19009 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17269) );
  NAND4_X1 U19010 ( .A1(n17272), .A2(n17271), .A3(n17270), .A4(n17269), .ZN(
        n17273) );
  AOI22_X1 U19011 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U19012 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17283) );
  INV_X1 U19013 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19418) );
  AOI22_X1 U19014 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U19015 ( .B1(n17238), .B2(n19418), .A(n17275), .ZN(n17281) );
  AOI22_X1 U19016 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17279) );
  AOI22_X1 U19017 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U19018 ( .A1(n18041), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U19019 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11212), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17276) );
  NAND4_X1 U19020 ( .A1(n17279), .A2(n17278), .A3(n17277), .A4(n17276), .ZN(
        n17280) );
  INV_X1 U19021 ( .A(n19295), .ZN(n17287) );
  NAND2_X1 U19022 ( .A1(n21218), .A2(n21026), .ZN(n17293) );
  NAND2_X1 U19023 ( .A1(n19425), .A2(n21063), .ZN(n17295) );
  NOR4_X2 U19024 ( .A1(n17287), .A2(n17285), .A3(n17293), .A4(n17295), .ZN(
        n21189) );
  NAND2_X1 U19025 ( .A1(n21189), .A2(n11506), .ZN(n17308) );
  NAND2_X1 U19026 ( .A1(n19211), .A2(n21218), .ZN(n17306) );
  INV_X1 U19027 ( .A(n17314), .ZN(n17286) );
  NAND2_X1 U19028 ( .A1(n21212), .A2(n21221), .ZN(n17313) );
  OAI211_X1 U19029 ( .C1(n21218), .C2(n17313), .A(n17287), .B(n17975), .ZN(
        n17288) );
  NAND2_X1 U19030 ( .A1(n17308), .A2(n17289), .ZN(n21628) );
  AOI21_X2 U19031 ( .B1(n17291), .B2(n21628), .A(n21666), .ZN(n17334) );
  INV_X1 U19032 ( .A(n21189), .ZN(n17298) );
  NAND2_X1 U19033 ( .A1(n21212), .A2(n19295), .ZN(n21165) );
  AOI21_X1 U19034 ( .B1(n21063), .B2(n17293), .A(n21221), .ZN(n17292) );
  AOI21_X1 U19035 ( .B1(n17293), .B2(n17310), .A(n17292), .ZN(n17297) );
  NOR2_X1 U19036 ( .A1(n20997), .A2(n21153), .ZN(n20974) );
  NOR3_X1 U19037 ( .A1(n21211), .A2(n19425), .A3(n20974), .ZN(n17305) );
  AOI211_X1 U19038 ( .C1(n19295), .C2(n17295), .A(n17305), .B(n17294), .ZN(
        n17296) );
  NAND2_X1 U19039 ( .A1(n17297), .A2(n17296), .ZN(n21167) );
  INV_X1 U19040 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18564) );
  INV_X2 U19041 ( .A(n22205), .ZN(n22153) );
  INV_X1 U19042 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22194) );
  NOR2_X1 U19043 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n22194), .ZN(n22199) );
  AND2_X1 U19044 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22153), .ZN(n18613) );
  INV_X2 U19045 ( .A(n18613), .ZN(n18616) );
  OAI21_X1 U19046 ( .B1(n22153), .B2(n22199), .A(n18616), .ZN(n21209) );
  XOR2_X1 U19047 ( .A(n17301), .B(n17300), .Z(n17304) );
  NAND2_X1 U19048 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22204) );
  NAND2_X1 U19049 ( .A1(n21656), .A2(n22204), .ZN(n21213) );
  AOI221_X1 U19050 ( .B1(n17334), .B2(n20972), .C1(n21209), .C2(n20972), .A(
        n21213), .ZN(n17315) );
  INV_X1 U19051 ( .A(n17305), .ZN(n17312) );
  OAI211_X1 U19052 ( .C1(n21153), .C2(n21221), .A(n17307), .B(n17306), .ZN(
        n17309) );
  OAI21_X1 U19053 ( .B1(n17310), .B2(n17309), .A(n17308), .ZN(n17311) );
  OAI211_X1 U19054 ( .C1(n17314), .C2(n17313), .A(n17312), .B(n17311), .ZN(
        n21215) );
  NOR2_X1 U19055 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21676), .ZN(n19088) );
  INV_X1 U19056 ( .A(n19088), .ZN(n17317) );
  OAI211_X1 U19057 ( .C1(n21665), .C2(n21644), .A(n17317), .B(n17316), .ZN(
        n21204) );
  NOR2_X1 U19058 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21202) );
  AND2_X1 U19059 ( .A1(n17318), .A2(n21163), .ZN(n21631) );
  NAND3_X1 U19060 ( .A1(n21204), .A2(n21202), .A3(n21631), .ZN(n17319) );
  OAI21_X1 U19061 ( .B1(n21204), .B2(n20576), .A(n17319), .ZN(P3_U3284) );
  INV_X1 U19062 ( .A(n17404), .ZN(n17324) );
  NOR2_X1 U19063 ( .A1(n17321), .A2(n17320), .ZN(n17322) );
  XNOR2_X1 U19064 ( .A(n17322), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21941) );
  INV_X1 U19065 ( .A(n21941), .ZN(n17323) );
  NAND4_X1 U19066 ( .A1(n22119), .A2(n17324), .A3(n22116), .A4(n17323), .ZN(
        n17325) );
  OAI21_X1 U19067 ( .B1(n22119), .B2(n17326), .A(n17325), .ZN(P1_U3468) );
  INV_X1 U19068 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17327) );
  INV_X1 U19069 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22196) );
  OAI221_X1 U19070 ( .B1(n22196), .B2(P3_STATE_REG_1__SCAN_IN), .C1(n22196), 
        .C2(n22194), .A(n22205), .ZN(n17328) );
  INV_X1 U19071 ( .A(n17328), .ZN(n22149) );
  INV_X1 U19072 ( .A(n22149), .ZN(n18604) );
  INV_X1 U19073 ( .A(BS16), .ZN(n17355) );
  NAND2_X1 U19074 ( .A1(n22194), .A2(n18564), .ZN(n22150) );
  AOI21_X1 U19075 ( .B1(n17355), .B2(n22150), .A(n18604), .ZN(n22145) );
  AOI21_X1 U19076 ( .B1(n17327), .B2(n18604), .A(n22145), .ZN(P3_U3280) );
  AND2_X1 U19077 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18604), .ZN(P3_U3028) );
  AND2_X1 U19078 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18604), .ZN(P3_U3027) );
  AND2_X1 U19079 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18604), .ZN(P3_U3026) );
  AND2_X1 U19080 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18604), .ZN(P3_U3025) );
  AND2_X1 U19081 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18604), .ZN(P3_U3024) );
  AND2_X1 U19082 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18604), .ZN(P3_U3023) );
  AND2_X1 U19083 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17328), .ZN(P3_U3022) );
  AND2_X1 U19084 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17328), .ZN(P3_U3021) );
  AND2_X1 U19085 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17328), .ZN(
        P3_U3020) );
  AND2_X1 U19086 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17328), .ZN(
        P3_U3019) );
  AND2_X1 U19087 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17328), .ZN(
        P3_U3018) );
  AND2_X1 U19088 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17328), .ZN(
        P3_U3017) );
  AND2_X1 U19089 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17328), .ZN(
        P3_U3016) );
  AND2_X1 U19090 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17328), .ZN(
        P3_U3015) );
  AND2_X1 U19091 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17328), .ZN(
        P3_U3014) );
  AND2_X1 U19092 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17328), .ZN(
        P3_U3013) );
  AND2_X1 U19093 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17328), .ZN(
        P3_U3012) );
  AND2_X1 U19094 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18604), .ZN(
        P3_U3011) );
  AND2_X1 U19095 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18604), .ZN(
        P3_U3010) );
  AND2_X1 U19096 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18604), .ZN(
        P3_U3009) );
  AND2_X1 U19097 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18604), .ZN(
        P3_U3008) );
  AND2_X1 U19098 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18604), .ZN(
        P3_U3007) );
  AND2_X1 U19099 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17328), .ZN(
        P3_U3006) );
  AND2_X1 U19100 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18604), .ZN(
        P3_U3005) );
  AND2_X1 U19101 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18604), .ZN(
        P3_U3004) );
  AND2_X1 U19102 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18604), .ZN(
        P3_U3003) );
  AND2_X1 U19103 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18604), .ZN(
        P3_U3002) );
  AND2_X1 U19104 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18604), .ZN(
        P3_U3001) );
  AND2_X1 U19105 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18604), .ZN(
        P3_U3000) );
  AND2_X1 U19106 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18604), .ZN(
        P3_U2999) );
  AOI21_X1 U19107 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17331)
         );
  INV_X1 U19108 ( .A(n22204), .ZN(n22206) );
  NAND4_X1 U19109 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n22206), .A4(n21668), .ZN(n21672) );
  INV_X1 U19110 ( .A(n21672), .ZN(n17329) );
  AOI211_X1 U19111 ( .C1(n18488), .C2(n17331), .A(n17330), .B(n17329), .ZN(
        P3_U2998) );
  NOR2_X1 U19112 ( .A1(n17333), .A2(n17332), .ZN(P3_U2867) );
  NOR2_X1 U19113 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21668), .ZN(n18231) );
  INV_X1 U19114 ( .A(n18231), .ZN(n18528) );
  NOR2_X1 U19115 ( .A1(n21158), .A2(n18528), .ZN(n18593) );
  INV_X1 U19116 ( .A(n21665), .ZN(n21690) );
  NOR3_X1 U19117 ( .A1(n17334), .A2(n21209), .A3(n20470), .ZN(n18584) );
  AND2_X1 U19118 ( .A1(n18597), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U19119 ( .A1(n21211), .A2(n11507), .ZN(n17583) );
  AOI21_X1 U19120 ( .B1(n21681), .B2(n21676), .A(n20530), .ZN(n17337) );
  INV_X1 U19121 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n17336) );
  AOI22_X1 U19122 ( .A1(n20462), .A2(n20530), .B1(n17337), .B2(n17336), .ZN(
        P3_U3298) );
  INV_X1 U19123 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18562) );
  NAND2_X1 U19124 ( .A1(n19425), .A2(n20530), .ZN(n20966) );
  INV_X1 U19125 ( .A(n20966), .ZN(n20554) );
  AOI21_X1 U19126 ( .B1(n17337), .B2(n18562), .A(n20554), .ZN(P3_U3299) );
  NOR2_X1 U19127 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22173), .ZN(n22183) );
  AOI21_X1 U19128 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22183), .A(n17338), 
        .ZN(n17339) );
  INV_X1 U19129 ( .A(n17339), .ZN(n22144) );
  INV_X1 U19130 ( .A(n22144), .ZN(n17507) );
  INV_X1 U19131 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17354) );
  NAND2_X1 U19132 ( .A1(n22181), .A2(n22173), .ZN(n22177) );
  AOI21_X1 U19133 ( .B1(n17355), .B2(n22177), .A(n17507), .ZN(n22140) );
  AOI21_X1 U19134 ( .B1(n17507), .B2(n17354), .A(n22140), .ZN(P2_U3591) );
  AND2_X1 U19135 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17507), .ZN(P2_U3208) );
  AND2_X1 U19136 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17339), .ZN(P2_U3207) );
  AND2_X1 U19137 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17507), .ZN(P2_U3206) );
  AND2_X1 U19138 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17507), .ZN(P2_U3205) );
  AND2_X1 U19139 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17507), .ZN(P2_U3204) );
  AND2_X1 U19140 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17507), .ZN(P2_U3203) );
  AND2_X1 U19141 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17339), .ZN(P2_U3202) );
  AND2_X1 U19142 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17339), .ZN(P2_U3201) );
  AND2_X1 U19143 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17339), .ZN(
        P2_U3200) );
  AND2_X1 U19144 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17339), .ZN(
        P2_U3199) );
  AND2_X1 U19145 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17339), .ZN(
        P2_U3198) );
  AND2_X1 U19146 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17339), .ZN(
        P2_U3197) );
  AND2_X1 U19147 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17339), .ZN(
        P2_U3196) );
  AND2_X1 U19148 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17339), .ZN(
        P2_U3195) );
  AND2_X1 U19149 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17339), .ZN(
        P2_U3194) );
  AND2_X1 U19150 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17339), .ZN(
        P2_U3193) );
  AND2_X1 U19151 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17339), .ZN(
        P2_U3192) );
  AND2_X1 U19152 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17339), .ZN(
        P2_U3191) );
  AND2_X1 U19153 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17507), .ZN(
        P2_U3190) );
  AND2_X1 U19154 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17507), .ZN(
        P2_U3189) );
  AND2_X1 U19155 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17507), .ZN(
        P2_U3188) );
  AND2_X1 U19156 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17507), .ZN(
        P2_U3187) );
  AND2_X1 U19157 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17339), .ZN(
        P2_U3186) );
  AND2_X1 U19158 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17507), .ZN(
        P2_U3185) );
  AND2_X1 U19159 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17507), .ZN(
        P2_U3184) );
  AND2_X1 U19160 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17507), .ZN(
        P2_U3183) );
  AND2_X1 U19161 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17507), .ZN(
        P2_U3182) );
  AND2_X1 U19162 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17507), .ZN(
        P2_U3181) );
  AND2_X1 U19163 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17507), .ZN(
        P2_U3180) );
  AND2_X1 U19164 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17507), .ZN(
        P2_U3179) );
  NAND2_X1 U19165 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n22174), .ZN(n19033) );
  AOI21_X1 U19166 ( .B1(n17340), .B2(n11739), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17341) );
  AOI221_X1 U19167 ( .B1(n19033), .B2(n17341), .C1(n14913), .C2(n17341), .A(
        n17342), .ZN(P2_U3178) );
  AOI221_X1 U19168 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17342), .C1(n19043), .C2(
        n17342), .A(n19715), .ZN(n17495) );
  INV_X1 U19169 ( .A(n17495), .ZN(n17493) );
  NOR2_X1 U19170 ( .A1(n17343), .A2(n17493), .ZN(P2_U3047) );
  AND2_X1 U19171 ( .A1(n17529), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19172 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17347) );
  NOR4_X1 U19173 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17346) );
  NOR4_X1 U19174 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17345) );
  NOR4_X1 U19175 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17344) );
  NAND4_X1 U19176 ( .A1(n17347), .A2(n17346), .A3(n17345), .A4(n17344), .ZN(
        n17353) );
  NOR4_X1 U19177 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17351) );
  AOI211_X1 U19178 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17350) );
  NOR4_X1 U19179 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17349) );
  NOR4_X1 U19180 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17348) );
  NAND4_X1 U19181 ( .A1(n17351), .A2(n17350), .A3(n17349), .A4(n17348), .ZN(
        n17352) );
  NOR2_X1 U19182 ( .A1(n17353), .A2(n17352), .ZN(n17503) );
  INV_X1 U19183 ( .A(n17503), .ZN(n17502) );
  NOR2_X1 U19184 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17502), .ZN(n17496) );
  INV_X1 U19185 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n17497) );
  INV_X1 U19186 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22143) );
  NAND3_X1 U19187 ( .A1(n17497), .A2(n22143), .A3(n17354), .ZN(n17501) );
  INV_X1 U19188 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17576) );
  AOI22_X1 U19189 ( .A1(n17496), .A2(n17501), .B1(n17502), .B2(n17576), .ZN(
        P2_U2821) );
  INV_X1 U19190 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U19191 ( .A1(n17496), .A2(n17497), .B1(n17502), .B2(n17574), .ZN(
        P2_U2820) );
  INV_X1 U19192 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17356) );
  INV_X1 U19193 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22169) );
  NAND2_X1 U19194 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22169), .ZN(n22749) );
  AND2_X1 U19195 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22164), .ZN(n17426) );
  NAND2_X1 U19196 ( .A1(n20212), .A2(n22169), .ZN(n22154) );
  AOI21_X1 U19197 ( .B1(n17355), .B2(n22154), .A(n17357), .ZN(n22138) );
  AOI21_X1 U19198 ( .B1(n17356), .B2(n17357), .A(n22138), .ZN(P1_U3464) );
  AND2_X1 U19199 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17357), .ZN(P1_U3193) );
  AND2_X1 U19200 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17357), .ZN(P1_U3192) );
  AND2_X1 U19201 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17357), .ZN(P1_U3191) );
  AND2_X1 U19202 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17357), .ZN(P1_U3190) );
  AND2_X1 U19203 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17357), .ZN(P1_U3189) );
  AND2_X1 U19204 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17357), .ZN(P1_U3188) );
  AND2_X1 U19205 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17357), .ZN(P1_U3187) );
  AND2_X1 U19206 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17357), .ZN(P1_U3186) );
  AND2_X1 U19207 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17357), .ZN(
        P1_U3185) );
  AND2_X1 U19208 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17357), .ZN(
        P1_U3184) );
  AND2_X1 U19209 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17357), .ZN(
        P1_U3183) );
  AND2_X1 U19210 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17357), .ZN(
        P1_U3182) );
  AND2_X1 U19211 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17357), .ZN(
        P1_U3181) );
  AND2_X1 U19212 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17357), .ZN(
        P1_U3180) );
  AND2_X1 U19213 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17357), .ZN(
        P1_U3179) );
  AND2_X1 U19214 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17357), .ZN(
        P1_U3178) );
  AND2_X1 U19215 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17357), .ZN(
        P1_U3177) );
  AND2_X1 U19216 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17357), .ZN(
        P1_U3176) );
  AND2_X1 U19217 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17357), .ZN(
        P1_U3175) );
  AND2_X1 U19218 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17357), .ZN(
        P1_U3174) );
  AND2_X1 U19219 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17357), .ZN(
        P1_U3173) );
  AND2_X1 U19220 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17357), .ZN(
        P1_U3172) );
  AND2_X1 U19221 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17357), .ZN(
        P1_U3171) );
  AND2_X1 U19222 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17357), .ZN(
        P1_U3170) );
  AND2_X1 U19223 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17357), .ZN(
        P1_U3169) );
  AND2_X1 U19224 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17357), .ZN(
        P1_U3168) );
  AND2_X1 U19225 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17357), .ZN(
        P1_U3167) );
  AND2_X1 U19226 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17357), .ZN(
        P1_U3166) );
  AND2_X1 U19227 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17357), .ZN(
        P1_U3165) );
  AND2_X1 U19228 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17357), .ZN(
        P1_U3164) );
  INV_X1 U19229 ( .A(n17358), .ZN(n17418) );
  OR2_X1 U19230 ( .A1(n17383), .A2(n13058), .ZN(n17382) );
  NAND2_X1 U19231 ( .A1(n17360), .A2(n17359), .ZN(n17380) );
  NAND2_X1 U19232 ( .A1(n17368), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n17361) );
  NAND2_X1 U19233 ( .A1(n17361), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17362) );
  NAND2_X1 U19234 ( .A1(n17363), .A2(n17362), .ZN(n22115) );
  AND2_X1 U19235 ( .A1(n17364), .A2(n22115), .ZN(n17377) );
  NAND2_X1 U19236 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17365) );
  AND2_X1 U19237 ( .A1(n17365), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17366) );
  OAI22_X1 U19238 ( .A1(n17370), .A2(n17366), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17374) );
  INV_X1 U19239 ( .A(n17367), .ZN(n17373) );
  MUX2_X1 U19240 ( .A(n17369), .B(n13058), .S(n17368), .Z(n17371) );
  NOR2_X1 U19241 ( .A1(n17371), .A2(n17370), .ZN(n17372) );
  OAI22_X1 U19242 ( .A1(n17375), .A2(n17374), .B1(n17373), .B2(n17372), .ZN(
        n17376) );
  AOI21_X1 U19243 ( .B1(n17378), .B2(n17377), .A(n17376), .ZN(n17379) );
  NAND2_X1 U19244 ( .A1(n17380), .A2(n17379), .ZN(n22117) );
  NAND2_X1 U19245 ( .A1(n17383), .A2(n22117), .ZN(n17381) );
  NAND2_X1 U19246 ( .A1(n17382), .A2(n17381), .ZN(n17396) );
  MUX2_X1 U19247 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17384), .S(
        n17383), .Z(n17391) );
  INV_X1 U19248 ( .A(n17391), .ZN(n17398) );
  NOR3_X1 U19249 ( .A1(n17386), .A2(n17385), .A3(n22251), .ZN(n17387) );
  NAND2_X1 U19250 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17387), .ZN(
        n17390) );
  OAI22_X1 U19251 ( .A1(n17405), .A2(n17388), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17387), .ZN(n17389) );
  OAI211_X1 U19252 ( .C1(n17391), .C2(n22237), .A(n17390), .B(n17389), .ZN(
        n17392) );
  OAI21_X1 U19253 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17398), .A(
        n17392), .ZN(n17393) );
  OAI21_X1 U19254 ( .B1(n13197), .B2(n17396), .A(n17393), .ZN(n17395) );
  NAND2_X1 U19255 ( .A1(n17396), .A2(n13197), .ZN(n17394) );
  AOI21_X1 U19256 ( .B1(n17395), .B2(n17394), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17410) );
  INV_X1 U19257 ( .A(n17396), .ZN(n17397) );
  NOR2_X1 U19258 ( .A1(n17398), .A2(n17397), .ZN(n17409) );
  NOR2_X1 U19259 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n17402) );
  INV_X1 U19260 ( .A(n17399), .ZN(n17401) );
  OAI211_X1 U19261 ( .C1(n17403), .C2(n17402), .A(n17401), .B(n17400), .ZN(
        n17408) );
  NOR2_X1 U19262 ( .A1(n21941), .A2(n17404), .ZN(n17406) );
  MUX2_X1 U19263 ( .A(n17406), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n17405), .Z(n17407) );
  NOR4_X1 U19264 ( .A1(n17410), .A2(n17409), .A3(n17408), .A4(n17407), .ZN(
        n22136) );
  OR2_X1 U19265 ( .A1(n17411), .A2(n21697), .ZN(n17416) );
  NAND2_X1 U19266 ( .A1(n17412), .A2(n22282), .ZN(n21699) );
  NOR3_X1 U19267 ( .A1(n17414), .A2(n17413), .A3(n21699), .ZN(n17415) );
  AOI21_X1 U19268 ( .B1(n17417), .B2(n17416), .A(n17415), .ZN(n17420) );
  OAI221_X1 U19269 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n22136), 
        .A(n17420), .ZN(n22127) );
  OAI211_X1 U19270 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21697), .A(n17418), 
        .B(n22127), .ZN(n22132) );
  NOR2_X1 U19271 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22165), .ZN(n17419) );
  OAI221_X1 U19272 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n22122), .C2(n17419), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n22123) );
  AOI21_X1 U19273 ( .B1(n22123), .B2(n17421), .A(n17420), .ZN(n17422) );
  AOI21_X1 U19274 ( .B1(n22121), .B2(n22132), .A(n17422), .ZN(P1_U3162) );
  NOR2_X1 U19275 ( .A1(n17424), .A2(n17423), .ZN(P1_U3032) );
  AND2_X1 U19276 ( .A1(n20199), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19277 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17425) );
  AOI21_X1 U19278 ( .B1(n17426), .B2(n17425), .A(n20459), .ZN(P1_U2802) );
  AOI22_X1 U19279 ( .A1(n18628), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_0__SCAN_IN), .B2(n17427), .ZN(n17428) );
  INV_X1 U19280 ( .A(n17428), .ZN(P2_U2816) );
  AOI22_X1 U19281 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n11167), .B1(n17443), 
        .B2(n18682), .ZN(n17433) );
  OAI22_X1 U19282 ( .A1(n17430), .A2(n17446), .B1(n17445), .B2(n17429), .ZN(
        n17431) );
  AOI21_X1 U19283 ( .B1(n17457), .B2(n18683), .A(n17431), .ZN(n17432) );
  OAI211_X1 U19284 ( .C1(n18676), .C2(n17452), .A(n17433), .B(n17432), .ZN(
        P2_U3009) );
  AOI22_X1 U19285 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17461), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n11167), .ZN(n17442) );
  XOR2_X1 U19286 ( .A(n17434), .B(n17435), .Z(n19008) );
  INV_X1 U19287 ( .A(n18720), .ZN(n19006) );
  INV_X1 U19288 ( .A(n17437), .ZN(n17439) );
  NOR2_X1 U19289 ( .A1(n17439), .A2(n17438), .ZN(n17440) );
  XNOR2_X1 U19290 ( .A(n17436), .B(n17440), .ZN(n19005) );
  AOI222_X1 U19291 ( .A1(n19008), .A2(n17467), .B1(n17457), .B2(n19006), .C1(
        n17462), .C2(n19005), .ZN(n17441) );
  OAI211_X1 U19292 ( .C1(n17475), .C2(n18715), .A(n17442), .B(n17441), .ZN(
        P2_U3006) );
  AOI22_X1 U19293 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n11167), .B1(n17443), 
        .B2(n18722), .ZN(n17451) );
  OAI22_X1 U19294 ( .A1(n17447), .A2(n17446), .B1(n17445), .B2(n17444), .ZN(
        n17448) );
  AOI21_X1 U19295 ( .B1(n17457), .B2(n17449), .A(n17448), .ZN(n17450) );
  OAI211_X1 U19296 ( .C1(n17453), .C2(n17452), .A(n17451), .B(n17450), .ZN(
        P2_U3005) );
  AOI22_X1 U19297 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17461), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n11167), .ZN(n17460) );
  INV_X1 U19298 ( .A(n18744), .ZN(n17456) );
  INV_X1 U19299 ( .A(n17454), .ZN(n17455) );
  AOI222_X1 U19300 ( .A1(n17458), .A2(n17462), .B1(n17457), .B2(n17456), .C1(
        n17467), .C2(n17455), .ZN(n17459) );
  OAI211_X1 U19301 ( .C1(n17475), .C2(n18738), .A(n17460), .B(n17459), .ZN(
        P2_U3004) );
  AOI22_X1 U19302 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17461), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n11167), .ZN(n17474) );
  NAND2_X1 U19303 ( .A1(n17463), .A2(n17462), .ZN(n17470) );
  NAND2_X1 U19304 ( .A1(n17465), .A2(n17464), .ZN(n17466) );
  NAND3_X1 U19305 ( .A1(n17468), .A2(n17467), .A3(n17466), .ZN(n17469) );
  OAI211_X1 U19306 ( .C1(n18764), .C2(n17471), .A(n17470), .B(n17469), .ZN(
        n17472) );
  INV_X1 U19307 ( .A(n17472), .ZN(n17473) );
  OAI211_X1 U19308 ( .C1(n17475), .C2(n18760), .A(n17474), .B(n17473), .ZN(
        P2_U3002) );
  OAI22_X1 U19309 ( .A1(n17477), .A2(n18630), .B1(n19594), .B2(n17476), .ZN(
        n17478) );
  AOI21_X1 U19310 ( .B1(n19612), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17478), 
        .ZN(n17479) );
  OAI22_X1 U19311 ( .A1(n19612), .A2(n17493), .B1(n17495), .B2(n17479), .ZN(
        P2_U3605) );
  INV_X1 U19312 ( .A(n19605), .ZN(n17480) );
  NAND2_X1 U19313 ( .A1(n17481), .A2(n17480), .ZN(n19661) );
  INV_X1 U19314 ( .A(n19661), .ZN(n17483) );
  NAND2_X1 U19315 ( .A1(n19605), .A2(n19708), .ZN(n17482) );
  NAND2_X1 U19316 ( .A1(n17482), .A2(n19034), .ZN(n17492) );
  AOI222_X1 U19317 ( .A1(n17484), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19708), 
        .B2(n17483), .C1(n17492), .C2(n19642), .ZN(n17485) );
  AOI22_X1 U19318 ( .A1(n17495), .A2(n19592), .B1(n17485), .B2(n17493), .ZN(
        P2_U3603) );
  NOR2_X1 U19319 ( .A1(n19694), .A2(n22141), .ZN(n17489) );
  OR2_X1 U19320 ( .A1(n19551), .A2(n17489), .ZN(n17486) );
  AOI22_X1 U19321 ( .A1(n17492), .A2(n17486), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n18646), .ZN(n17487) );
  AOI22_X1 U19322 ( .A1(n17495), .A2(n19689), .B1(n17487), .B2(n17493), .ZN(
        P2_U3604) );
  OAI21_X1 U19323 ( .B1(n19623), .B2(n17488), .A(n19581), .ZN(n17490) );
  AOI222_X1 U19324 ( .A1(n17492), .A2(n19660), .B1(n17491), .B2(
        P2_STATE2_REG_3__SCAN_IN), .C1(n17490), .C2(n17489), .ZN(n17494) );
  AOI22_X1 U19325 ( .A1(n17495), .A2(n19563), .B1(n17494), .B2(n17493), .ZN(
        P2_U3602) );
  NAND2_X1 U19326 ( .A1(n17496), .A2(n22143), .ZN(n17500) );
  OAI21_X1 U19327 ( .B1(n17548), .B2(n17497), .A(n17503), .ZN(n17498) );
  OAI21_X1 U19328 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17503), .A(n17498), 
        .ZN(n17499) );
  OAI221_X1 U19329 ( .B1(n17500), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17500), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17499), .ZN(P2_U2822) );
  INV_X1 U19330 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17579) );
  OAI221_X1 U19331 ( .B1(n17503), .B2(n17579), .C1(n17502), .C2(n17501), .A(
        n17500), .ZN(P2_U2823) );
  INV_X1 U19332 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n17504) );
  AOI22_X1 U19333 ( .A1(n22172), .A2(n17505), .B1(n17504), .B2(n17577), .ZN(
        P2_U3611) );
  INV_X1 U19334 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17506) );
  AOI22_X1 U19335 ( .A1(n22172), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17506), 
        .B2(n17577), .ZN(P2_U3608) );
  INV_X1 U19336 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n22191) );
  INV_X1 U19337 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17508) );
  OAI21_X1 U19338 ( .B1(n22191), .B2(n17508), .A(n17507), .ZN(P2_U2815) );
  AOI22_X1 U19339 ( .A1(n17542), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17510) );
  OAI21_X1 U19340 ( .B1(n17511), .B2(n17544), .A(n17510), .ZN(P2_U2951) );
  INV_X1 U19341 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U19342 ( .A1(n17542), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17512) );
  OAI21_X1 U19343 ( .B1(n17513), .B2(n17544), .A(n17512), .ZN(P2_U2950) );
  INV_X1 U19344 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17515) );
  AOI22_X1 U19345 ( .A1(n17542), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17514) );
  OAI21_X1 U19346 ( .B1(n17515), .B2(n17544), .A(n17514), .ZN(P2_U2949) );
  INV_X1 U19347 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U19348 ( .A1(n17530), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U19349 ( .B1(n17517), .B2(n17544), .A(n17516), .ZN(P2_U2948) );
  INV_X1 U19350 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U19351 ( .A1(n17542), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17518) );
  OAI21_X1 U19352 ( .B1(n17519), .B2(n17544), .A(n17518), .ZN(P2_U2947) );
  INV_X1 U19353 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19354 ( .A1(n17530), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17520) );
  OAI21_X1 U19355 ( .B1(n19771), .B2(n17544), .A(n17520), .ZN(P2_U2946) );
  AOI22_X1 U19356 ( .A1(n17530), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U19357 ( .B1(n17522), .B2(n17544), .A(n17521), .ZN(P2_U2945) );
  AOI22_X1 U19358 ( .A1(n17530), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17523) );
  OAI21_X1 U19359 ( .B1(n17524), .B2(n17544), .A(n17523), .ZN(P2_U2944) );
  AOI22_X1 U19360 ( .A1(n17530), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17525) );
  OAI21_X1 U19361 ( .B1(n17526), .B2(n17544), .A(n17525), .ZN(P2_U2943) );
  AOI22_X1 U19362 ( .A1(n17542), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17527) );
  OAI21_X1 U19363 ( .B1(n17528), .B2(n17544), .A(n17527), .ZN(P2_U2942) );
  AOI22_X1 U19364 ( .A1(n17530), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17529), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17531) );
  OAI21_X1 U19365 ( .B1(n17532), .B2(n17544), .A(n17531), .ZN(P2_U2941) );
  AOI22_X1 U19366 ( .A1(n17542), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17533) );
  OAI21_X1 U19367 ( .B1(n17534), .B2(n17544), .A(n17533), .ZN(P2_U2940) );
  AOI22_X1 U19368 ( .A1(n17542), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17535) );
  OAI21_X1 U19369 ( .B1(n17536), .B2(n17544), .A(n17535), .ZN(P2_U2939) );
  AOI22_X1 U19370 ( .A1(n17542), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U19371 ( .B1(n17538), .B2(n17544), .A(n17537), .ZN(P2_U2938) );
  AOI22_X1 U19372 ( .A1(n17542), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17539) );
  OAI21_X1 U19373 ( .B1(n17540), .B2(n17544), .A(n17539), .ZN(P2_U2937) );
  AOI22_X1 U19374 ( .A1(n17542), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17541), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17543) );
  OAI21_X1 U19375 ( .B1(n17545), .B2(n17544), .A(n17543), .ZN(P2_U2936) );
  AOI21_X1 U19376 ( .B1(n22191), .B2(n17546), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17547) );
  AOI21_X1 U19377 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n22172), .A(n17547), 
        .ZN(P2_U2817) );
  NAND2_X1 U19378 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22172), .ZN(n17570) );
  INV_X1 U19379 ( .A(n17570), .ZN(n22180) );
  INV_X1 U19380 ( .A(n22180), .ZN(n17571) );
  OAI222_X1 U19381 ( .A1(n17572), .A2(n17549), .B1(n20120), .B2(n22172), .C1(
        n17548), .C2(n17571), .ZN(P2_U3212) );
  INV_X1 U19382 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17550) );
  INV_X1 U19383 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20122) );
  OAI222_X1 U19384 ( .A1(n17568), .A2(n17550), .B1(n20122), .B2(n22172), .C1(
        n17549), .C2(n17570), .ZN(P2_U3213) );
  INV_X1 U19385 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20124) );
  OAI222_X1 U19386 ( .A1(n17568), .A2(n11952), .B1(n20124), .B2(n22172), .C1(
        n17550), .C2(n17571), .ZN(P2_U3214) );
  INV_X1 U19387 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20126) );
  OAI222_X1 U19388 ( .A1(n17568), .A2(n11955), .B1(n20126), .B2(n22172), .C1(
        n11952), .C2(n17570), .ZN(P2_U3215) );
  INV_X1 U19389 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20128) );
  OAI222_X1 U19390 ( .A1(n17568), .A2(n11961), .B1(n20128), .B2(n22172), .C1(
        n11955), .C2(n17570), .ZN(P2_U3216) );
  INV_X1 U19391 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20130) );
  OAI222_X1 U19392 ( .A1(n17568), .A2(n17551), .B1(n20130), .B2(n22172), .C1(
        n11961), .C2(n17571), .ZN(P2_U3217) );
  INV_X1 U19393 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17552) );
  INV_X1 U19394 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20132) );
  OAI222_X1 U19395 ( .A1(n17568), .A2(n17552), .B1(n20132), .B2(n22172), .C1(
        n17551), .C2(n17571), .ZN(P2_U3218) );
  INV_X1 U19396 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20134) );
  OAI222_X1 U19397 ( .A1(n17568), .A2(n17553), .B1(n20134), .B2(n22172), .C1(
        n17552), .C2(n17570), .ZN(P2_U3219) );
  INV_X1 U19398 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20136) );
  INV_X1 U19399 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n18735) );
  OAI222_X1 U19400 ( .A1(n17571), .A2(n17553), .B1(n20136), .B2(n22172), .C1(
        n18735), .C2(n17568), .ZN(P2_U3220) );
  INV_X1 U19401 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20138) );
  INV_X1 U19402 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17554) );
  OAI222_X1 U19403 ( .A1(n17570), .A2(n18735), .B1(n20138), .B2(n22172), .C1(
        n17554), .C2(n17568), .ZN(P2_U3221) );
  INV_X1 U19404 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20140) );
  OAI222_X1 U19405 ( .A1(n17570), .A2(n17554), .B1(n20140), .B2(n22172), .C1(
        n17555), .C2(n17568), .ZN(P2_U3222) );
  INV_X1 U19406 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20142) );
  INV_X1 U19407 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n17556) );
  OAI222_X1 U19408 ( .A1(n17571), .A2(n17555), .B1(n20142), .B2(n22172), .C1(
        n17556), .C2(n17568), .ZN(P2_U3223) );
  INV_X1 U19409 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20144) );
  INV_X1 U19410 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17557) );
  OAI222_X1 U19411 ( .A1(n17570), .A2(n17556), .B1(n20144), .B2(n22172), .C1(
        n17557), .C2(n17568), .ZN(P2_U3224) );
  INV_X1 U19412 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20146) );
  OAI222_X1 U19413 ( .A1(n17570), .A2(n17557), .B1(n20146), .B2(n22172), .C1(
        n17558), .C2(n17568), .ZN(P2_U3225) );
  INV_X1 U19414 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20148) );
  OAI222_X1 U19415 ( .A1(n17570), .A2(n17558), .B1(n20148), .B2(n22172), .C1(
        n18805), .C2(n17568), .ZN(P2_U3226) );
  INV_X1 U19416 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20150) );
  INV_X1 U19417 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17559) );
  OAI222_X1 U19418 ( .A1(n17570), .A2(n18805), .B1(n20150), .B2(n22172), .C1(
        n17559), .C2(n17568), .ZN(P2_U3227) );
  INV_X1 U19419 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20152) );
  OAI222_X1 U19420 ( .A1(n17570), .A2(n17559), .B1(n20152), .B2(n22172), .C1(
        n12400), .C2(n17568), .ZN(P2_U3228) );
  INV_X1 U19421 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20154) );
  OAI222_X1 U19422 ( .A1(n17568), .A2(n17560), .B1(n20154), .B2(n22172), .C1(
        n12400), .C2(n17571), .ZN(P2_U3229) );
  INV_X1 U19423 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20156) );
  OAI222_X1 U19424 ( .A1(n17570), .A2(n17560), .B1(n20156), .B2(n22172), .C1(
        n17561), .C2(n17568), .ZN(P2_U3230) );
  INV_X1 U19425 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17562) );
  INV_X1 U19426 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20158) );
  OAI222_X1 U19427 ( .A1(n17572), .A2(n17562), .B1(n20158), .B2(n22172), .C1(
        n17561), .C2(n17571), .ZN(P2_U3231) );
  INV_X1 U19428 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17563) );
  INV_X1 U19429 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20160) );
  OAI222_X1 U19430 ( .A1(n17572), .A2(n17563), .B1(n20160), .B2(n22172), .C1(
        n17562), .C2(n17571), .ZN(P2_U3232) );
  INV_X1 U19431 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20162) );
  OAI222_X1 U19432 ( .A1(n17572), .A2(n18882), .B1(n20162), .B2(n22172), .C1(
        n17563), .C2(n17571), .ZN(P2_U3233) );
  INV_X1 U19433 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17564) );
  INV_X1 U19434 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20164) );
  OAI222_X1 U19435 ( .A1(n17572), .A2(n17564), .B1(n20164), .B2(n22172), .C1(
        n18882), .C2(n17571), .ZN(P2_U3234) );
  INV_X1 U19436 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17565) );
  INV_X1 U19437 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20166) );
  OAI222_X1 U19438 ( .A1(n17572), .A2(n17565), .B1(n20166), .B2(n22172), .C1(
        n17564), .C2(n17571), .ZN(P2_U3235) );
  INV_X1 U19439 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20169) );
  OAI222_X1 U19440 ( .A1(n17570), .A2(n17565), .B1(n20169), .B2(n22172), .C1(
        n18921), .C2(n17568), .ZN(P2_U3236) );
  INV_X1 U19441 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20171) );
  OAI222_X1 U19442 ( .A1(n17572), .A2(n17566), .B1(n20171), .B2(n22172), .C1(
        n18921), .C2(n17571), .ZN(P2_U3237) );
  INV_X1 U19443 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20173) );
  INV_X1 U19444 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17567) );
  OAI222_X1 U19445 ( .A1(n17570), .A2(n17566), .B1(n20173), .B2(n22172), .C1(
        n17567), .C2(n17568), .ZN(P2_U3238) );
  INV_X1 U19446 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20175) );
  OAI222_X1 U19447 ( .A1(n17571), .A2(n17567), .B1(n20175), .B2(n22172), .C1(
        n17569), .C2(n17568), .ZN(P2_U3239) );
  INV_X1 U19448 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20177) );
  OAI222_X1 U19449 ( .A1(n17570), .A2(n17569), .B1(n20177), .B2(n22172), .C1(
        n15969), .C2(n17568), .ZN(P2_U3240) );
  INV_X1 U19450 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20180) );
  OAI222_X1 U19451 ( .A1(n17572), .A2(n18967), .B1(n20180), .B2(n22172), .C1(
        n15969), .C2(n17571), .ZN(P2_U3241) );
  INV_X1 U19452 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17573) );
  AOI22_X1 U19453 ( .A1(n22172), .A2(n17574), .B1(n17573), .B2(n17577), .ZN(
        P2_U3588) );
  INV_X1 U19454 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17575) );
  AOI22_X1 U19455 ( .A1(n22172), .A2(n17576), .B1(n17575), .B2(n17577), .ZN(
        P2_U3587) );
  MUX2_X1 U19456 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n22172), .Z(P2_U3586) );
  INV_X1 U19457 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U19458 ( .A1(n22172), .A2(n17579), .B1(n17578), .B2(n17577), .ZN(
        P2_U3585) );
  AND3_X1 U19459 ( .A1(n20997), .A2(n21221), .A3(n17580), .ZN(n17581) );
  AND2_X1 U19460 ( .A1(n17952), .A2(n21063), .ZN(n17954) );
  INV_X2 U19461 ( .A(n17954), .ZN(n17951) );
  INV_X1 U19462 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19291) );
  INV_X1 U19463 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20549) );
  NAND2_X1 U19464 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17589) );
  NOR2_X1 U19465 ( .A1(n20549), .A2(n17589), .ZN(n17587) );
  NAND2_X1 U19466 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17587), .ZN(n17584) );
  INV_X1 U19467 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20566) );
  OAI21_X1 U19468 ( .B1(n17953), .B2(n17584), .A(n20566), .ZN(n17585) );
  NOR2_X1 U19469 ( .A1(n20566), .A2(n17584), .ZN(n17604) );
  NAND2_X1 U19470 ( .A1(n17952), .A2(n17604), .ZN(n17614) );
  NAND3_X1 U19471 ( .A1(n17951), .A2(n17585), .A3(n17614), .ZN(n17586) );
  OAI21_X1 U19472 ( .B1(n17951), .B2(n19291), .A(n17586), .ZN(P3_U2699) );
  NAND2_X1 U19473 ( .A1(n20997), .A2(n17952), .ZN(n17956) );
  INV_X1 U19474 ( .A(n17956), .ZN(n17946) );
  NAND2_X1 U19475 ( .A1(n17946), .A2(n17587), .ZN(n17590) );
  INV_X1 U19476 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19334) );
  NAND3_X1 U19477 ( .A1(n17590), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17951), .ZN(
        n17588) );
  OAI221_X1 U19478 ( .B1(n17590), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17951), 
        .C2(n19334), .A(n17588), .ZN(P3_U2700) );
  INV_X1 U19479 ( .A(n17589), .ZN(n17950) );
  AOI21_X1 U19480 ( .B1(n17952), .B2(n17950), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17592) );
  NAND2_X1 U19481 ( .A1(n17951), .A2(n17590), .ZN(n17591) );
  INV_X1 U19482 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19374) );
  OAI22_X1 U19483 ( .A1(n17592), .A2(n17591), .B1(n19374), .B2(n17951), .ZN(
        P3_U2701) );
  AOI22_X1 U19484 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17806), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U19485 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19486 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U19487 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17594) );
  NAND4_X1 U19488 ( .A1(n17597), .A2(n17596), .A3(n17595), .A4(n17594), .ZN(
        n17603) );
  AOI22_X1 U19489 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U19490 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17600) );
  AOI22_X1 U19491 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U19492 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17598) );
  NAND4_X1 U19493 ( .A1(n17601), .A2(n17600), .A3(n17599), .A4(n17598), .ZN(
        n17602) );
  NOR2_X1 U19494 ( .A1(n17603), .A2(n17602), .ZN(n21137) );
  INV_X1 U19495 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20635) );
  INV_X1 U19496 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20601) );
  NAND2_X1 U19497 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17604), .ZN(n17611) );
  NOR2_X1 U19498 ( .A1(n20601), .A2(n17611), .ZN(n17608) );
  NAND2_X1 U19499 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17608), .ZN(n17607) );
  NOR2_X1 U19500 ( .A1(n20635), .A2(n17607), .ZN(n17725) );
  AOI211_X1 U19501 ( .C1(n20635), .C2(n17607), .A(n17725), .B(n17956), .ZN(
        n17605) );
  AOI21_X1 U19502 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17953), .A(n17605), .ZN(
        n17606) );
  OAI21_X1 U19503 ( .B1(n21137), .B2(n17951), .A(n17606), .ZN(P3_U2695) );
  AOI22_X1 U19504 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17954), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17953), .ZN(n17610) );
  OAI211_X1 U19505 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17608), .A(n17946), .B(
        n17607), .ZN(n17609) );
  NAND2_X1 U19506 ( .A1(n17610), .A2(n17609), .ZN(P3_U2696) );
  INV_X1 U19507 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U19508 ( .B1(n17615), .B2(n17614), .A(n17951), .ZN(n17617) );
  NOR3_X1 U19509 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17956), .A3(n17611), .ZN(
        n17612) );
  AOI21_X1 U19510 ( .B1(n17954), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17612), .ZN(n17613) );
  OAI21_X1 U19511 ( .B1(n17617), .B2(n20601), .A(n17613), .ZN(P3_U2697) );
  AND2_X1 U19512 ( .A1(n17615), .A2(n17614), .ZN(n17616) );
  INV_X1 U19513 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19250) );
  OAI22_X1 U19514 ( .A1(n17617), .A2(n17616), .B1(n19250), .B2(n17951), .ZN(
        P3_U2698) );
  AOI22_X1 U19515 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U19516 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U19517 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U19518 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17618) );
  NAND4_X1 U19519 ( .A1(n17621), .A2(n17620), .A3(n17619), .A4(n17618), .ZN(
        n17627) );
  AOI22_X1 U19520 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17625) );
  AOI22_X1 U19521 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17624) );
  AOI22_X1 U19522 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U19523 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17622) );
  NAND4_X1 U19524 ( .A1(n17625), .A2(n17624), .A3(n17623), .A4(n17622), .ZN(
        n17626) );
  NOR2_X1 U19525 ( .A1(n17627), .A2(n17626), .ZN(n21117) );
  NAND3_X1 U19526 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n17727) );
  NAND3_X1 U19527 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .ZN(n17728) );
  NAND2_X1 U19528 ( .A1(n17952), .A2(n17725), .ZN(n17721) );
  NOR2_X1 U19529 ( .A1(n17728), .A2(n17721), .ZN(n17682) );
  INV_X1 U19530 ( .A(n17682), .ZN(n17696) );
  NOR2_X1 U19531 ( .A1(n17727), .A2(n17696), .ZN(n17641) );
  NAND2_X1 U19532 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17641), .ZN(n17640) );
  INV_X1 U19533 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n20738) );
  OAI21_X1 U19534 ( .B1(n17954), .B2(n20738), .A(n17640), .ZN(n17628) );
  OAI221_X1 U19535 ( .B1(n20997), .B2(n17640), .C1(n17640), .C2(n20738), .A(
        n17628), .ZN(n17629) );
  OAI21_X1 U19536 ( .B1(n21117), .B2(n17951), .A(n17629), .ZN(P3_U2687) );
  AOI22_X1 U19537 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17639) );
  AOI22_X1 U19538 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U19539 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17630) );
  OAI21_X1 U19540 ( .B1(n17686), .B2(n19169), .A(n17630), .ZN(n17636) );
  AOI22_X1 U19541 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U19542 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17633) );
  AOI22_X1 U19543 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U19544 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17631) );
  NAND4_X1 U19545 ( .A1(n17634), .A2(n17633), .A3(n17632), .A4(n17631), .ZN(
        n17635) );
  AOI211_X1 U19546 ( .C1(n11169), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17636), .B(n17635), .ZN(n17637) );
  NAND3_X1 U19547 ( .A1(n17639), .A2(n17638), .A3(n17637), .ZN(n21127) );
  INV_X1 U19548 ( .A(n21127), .ZN(n17643) );
  OAI211_X1 U19549 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17641), .A(n17640), .B(
        n17951), .ZN(n17642) );
  OAI21_X1 U19550 ( .B1(n17643), .B2(n17951), .A(n17642), .ZN(P3_U2688) );
  AOI22_X1 U19551 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17653) );
  AOI22_X1 U19552 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17652) );
  AOI22_X1 U19553 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17644) );
  OAI21_X1 U19554 ( .B1(n17686), .B2(n19250), .A(n17644), .ZN(n17650) );
  AOI22_X1 U19555 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U19556 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U19557 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19558 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17645) );
  NAND4_X1 U19559 ( .A1(n17648), .A2(n17647), .A3(n17646), .A4(n17645), .ZN(
        n17649) );
  AOI211_X1 U19560 ( .C1(n18043), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n17650), .B(n17649), .ZN(n17651) );
  NAND3_X1 U19561 ( .A1(n17653), .A2(n17652), .A3(n17651), .ZN(n20975) );
  INV_X1 U19562 ( .A(n20975), .ZN(n17656) );
  INV_X1 U19563 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n20686) );
  NOR3_X1 U19564 ( .A1(n21063), .A2(n20686), .A3(n17696), .ZN(n17684) );
  NOR2_X1 U19565 ( .A1(n20686), .A2(n17696), .ZN(n17654) );
  OAI21_X1 U19566 ( .B1(n17954), .B2(n17654), .A(P3_EBX_REG_13__SCAN_IN), .ZN(
        n17657) );
  OAI21_X1 U19567 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17684), .A(n17657), .ZN(
        n17655) );
  OAI21_X1 U19568 ( .B1(n17656), .B2(n17951), .A(n17655), .ZN(P3_U2690) );
  NAND2_X1 U19569 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17657), .ZN(n17670) );
  AOI22_X1 U19570 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17667) );
  AOI22_X1 U19571 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17666) );
  AOI22_X1 U19572 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17658) );
  OAI21_X1 U19573 ( .B1(n17686), .B2(n19209), .A(n17658), .ZN(n17664) );
  AOI22_X1 U19574 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17662) );
  AOI22_X1 U19575 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17661) );
  AOI22_X1 U19576 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U19577 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17659) );
  NAND4_X1 U19578 ( .A1(n17662), .A2(n17661), .A3(n17660), .A4(n17659), .ZN(
        n17663) );
  AOI211_X1 U19579 ( .C1(n17934), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n17664), .B(n17663), .ZN(n17665) );
  NAND3_X1 U19580 ( .A1(n17667), .A2(n17666), .A3(n17665), .ZN(n21121) );
  INV_X1 U19581 ( .A(n21121), .ZN(n17669) );
  INV_X1 U19582 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20718) );
  NAND3_X1 U19583 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17684), .A3(n20718), 
        .ZN(n17668) );
  OAI221_X1 U19584 ( .B1(n17954), .B2(n17670), .C1(n17951), .C2(n17669), .A(
        n17668), .ZN(P3_U2689) );
  AOI22_X1 U19585 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U19586 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19587 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U19588 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17671), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17672) );
  NAND4_X1 U19589 ( .A1(n17675), .A2(n17674), .A3(n17673), .A4(n17672), .ZN(
        n17681) );
  AOI22_X1 U19590 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17679) );
  AOI22_X1 U19591 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U19592 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U19593 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17676) );
  NAND4_X1 U19594 ( .A1(n17679), .A2(n17678), .A3(n17677), .A4(n17676), .ZN(
        n17680) );
  NOR2_X1 U19595 ( .A1(n17681), .A2(n17680), .ZN(n20980) );
  OAI21_X1 U19596 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17682), .A(n17951), .ZN(
        n17683) );
  OAI22_X1 U19597 ( .A1(n20980), .A2(n17951), .B1(n17684), .B2(n17683), .ZN(
        P3_U2691) );
  AOI22_X1 U19598 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U19599 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17694) );
  AOI22_X1 U19600 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U19601 ( .B1(n17686), .B2(n19334), .A(n17685), .ZN(n17692) );
  AOI22_X1 U19602 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U19603 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17689) );
  AOI22_X1 U19604 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17688) );
  AOI22_X1 U19605 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11212), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17687) );
  NAND4_X1 U19606 ( .A1(n17690), .A2(n17689), .A3(n17688), .A4(n17687), .ZN(
        n17691) );
  AOI211_X1 U19607 ( .C1(n11169), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17692), .B(n17691), .ZN(n17693) );
  NAND3_X1 U19608 ( .A1(n17695), .A2(n17694), .A3(n17693), .ZN(n20983) );
  INV_X1 U19609 ( .A(n20983), .ZN(n17698) );
  INV_X1 U19610 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n20660) );
  INV_X1 U19611 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20637) );
  NOR3_X1 U19612 ( .A1(n20660), .A2(n20637), .A3(n17721), .ZN(n17710) );
  OAI21_X1 U19613 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17710), .A(n17696), .ZN(
        n17697) );
  AOI22_X1 U19614 ( .A1(n17954), .A2(n17698), .B1(n17697), .B2(n17951), .ZN(
        P3_U2692) );
  AOI22_X1 U19615 ( .A1(n17901), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U19616 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17701) );
  AOI22_X1 U19617 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U19618 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17699) );
  NAND4_X1 U19619 ( .A1(n17702), .A2(n17701), .A3(n17700), .A4(n17699), .ZN(
        n17708) );
  AOI22_X1 U19620 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U19621 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19622 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U19623 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17703) );
  NAND4_X1 U19624 ( .A1(n17706), .A2(n17705), .A3(n17704), .A4(n17703), .ZN(
        n17707) );
  NOR2_X1 U19625 ( .A1(n17708), .A2(n17707), .ZN(n20987) );
  NOR2_X1 U19626 ( .A1(n20637), .A2(n17721), .ZN(n17724) );
  OAI21_X1 U19627 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17724), .A(n17951), .ZN(
        n17709) );
  OAI22_X1 U19628 ( .A1(n20987), .A2(n17951), .B1(n17710), .B2(n17709), .ZN(
        P3_U2693) );
  AOI22_X1 U19629 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18043), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17714) );
  AOI22_X1 U19630 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11170), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17713) );
  AOI22_X1 U19631 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17992), .ZN(n17712) );
  AOI22_X1 U19632 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18016), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17934), .ZN(n17711) );
  NAND4_X1 U19633 ( .A1(n17714), .A2(n17713), .A3(n17712), .A4(n17711), .ZN(
        n17720) );
  AOI22_X1 U19634 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U19635 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n18044), .ZN(n17717) );
  AOI22_X1 U19636 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11177), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18041), .ZN(n17716) );
  AOI22_X1 U19637 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18029), .ZN(n17715) );
  NAND4_X1 U19638 ( .A1(n17718), .A2(n17717), .A3(n17716), .A4(n17715), .ZN(
        n17719) );
  NOR2_X1 U19639 ( .A1(n17720), .A2(n17719), .ZN(n20992) );
  INV_X1 U19640 ( .A(n17721), .ZN(n17722) );
  OAI21_X1 U19641 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17722), .A(n17951), .ZN(
        n17723) );
  OAI22_X1 U19642 ( .A1(n20992), .A2(n17951), .B1(n17724), .B2(n17723), .ZN(
        P3_U2694) );
  INV_X1 U19643 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20944) );
  AND4_X1 U19644 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .A4(P3_EBX_REG_25__SCAN_IN), .ZN(n17850)
         );
  INV_X1 U19645 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20835) );
  INV_X1 U19646 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n20823) );
  INV_X1 U19647 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20804) );
  INV_X1 U19648 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20779) );
  NAND3_X1 U19649 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(n17725), .ZN(n17726) );
  NOR3_X1 U19650 ( .A1(n17728), .A2(n17727), .A3(n17726), .ZN(n17947) );
  NAND2_X1 U19651 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17947), .ZN(n17945) );
  NOR2_X1 U19652 ( .A1(n17953), .A2(n17945), .ZN(n17918) );
  NAND2_X1 U19653 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17918), .ZN(n17920) );
  NOR2_X1 U19654 ( .A1(n20779), .A2(n17920), .ZN(n17933) );
  NAND2_X1 U19655 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17933), .ZN(n17840) );
  NOR4_X1 U19656 ( .A1(n20835), .A2(n20823), .A3(n20804), .A4(n17840), .ZN(
        n17729) );
  NAND4_X1 U19657 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n17850), .A4(n17729), .ZN(n17732) );
  NOR2_X1 U19658 ( .A1(n20944), .A2(n17732), .ZN(n17829) );
  NAND2_X1 U19659 ( .A1(n17951), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17731) );
  NAND2_X1 U19660 ( .A1(n17829), .A2(n20997), .ZN(n17730) );
  OAI22_X1 U19661 ( .A1(n17829), .A2(n17731), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17730), .ZN(P3_U2672) );
  NAND2_X1 U19662 ( .A1(n20944), .A2(n17732), .ZN(n17733) );
  NAND2_X1 U19663 ( .A1(n17733), .A2(n17951), .ZN(n17828) );
  AOI22_X1 U19664 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17737) );
  AOI22_X1 U19665 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U19666 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U19667 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17734) );
  NAND4_X1 U19668 ( .A1(n17737), .A2(n17736), .A3(n17735), .A4(n17734), .ZN(
        n17743) );
  AOI22_X1 U19669 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U19670 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U19671 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U19672 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17738) );
  NAND4_X1 U19673 ( .A1(n17741), .A2(n17740), .A3(n17739), .A4(n17738), .ZN(
        n17742) );
  NOR2_X1 U19674 ( .A1(n17743), .A2(n17742), .ZN(n17827) );
  AOI22_X1 U19675 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U19676 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19677 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17745) );
  AOI22_X1 U19678 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17744) );
  NAND4_X1 U19679 ( .A1(n17747), .A2(n17746), .A3(n17745), .A4(n17744), .ZN(
        n17753) );
  AOI22_X1 U19680 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U19681 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U19682 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U19683 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17748) );
  NAND4_X1 U19684 ( .A1(n17751), .A2(n17750), .A3(n17749), .A4(n17748), .ZN(
        n17752) );
  NOR2_X1 U19685 ( .A1(n17753), .A2(n17752), .ZN(n17855) );
  AOI22_X1 U19686 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U19687 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17756) );
  AOI22_X1 U19688 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U19689 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17754) );
  NAND4_X1 U19690 ( .A1(n17757), .A2(n17756), .A3(n17755), .A4(n17754), .ZN(
        n17763) );
  AOI22_X1 U19691 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U19692 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17760) );
  AOI22_X1 U19693 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17759) );
  AOI22_X1 U19694 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17758) );
  NAND4_X1 U19695 ( .A1(n17761), .A2(n17760), .A3(n17759), .A4(n17758), .ZN(
        n17762) );
  NOR2_X1 U19696 ( .A1(n17763), .A2(n17762), .ZN(n17861) );
  AOI22_X1 U19697 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11168), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n18041), .ZN(n17767) );
  AOI22_X1 U19698 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17766) );
  AOI22_X1 U19699 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11170), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18016), .ZN(n17765) );
  AOI22_X1 U19700 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11212), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17764) );
  NAND4_X1 U19701 ( .A1(n17767), .A2(n17766), .A3(n17765), .A4(n17764), .ZN(
        n17773) );
  AOI22_X1 U19702 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18029), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17771) );
  AOI22_X1 U19703 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18028), .ZN(n17770) );
  AOI22_X1 U19704 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n11177), .ZN(n17769) );
  AOI22_X1 U19705 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17768) );
  NAND4_X1 U19706 ( .A1(n17771), .A2(n17770), .A3(n17769), .A4(n17768), .ZN(
        n17772) );
  NOR2_X1 U19707 ( .A1(n17773), .A2(n17772), .ZN(n17870) );
  AOI22_X1 U19708 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17784) );
  AOI22_X1 U19709 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17783) );
  INV_X1 U19710 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U19711 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17774) );
  OAI21_X1 U19712 ( .B1(n17238), .B2(n17775), .A(n17774), .ZN(n17781) );
  AOI22_X1 U19713 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17779) );
  AOI22_X1 U19714 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U19715 ( .A1(n11203), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U19716 ( .A1(n11213), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17776) );
  NAND4_X1 U19717 ( .A1(n17779), .A2(n17778), .A3(n17777), .A4(n17776), .ZN(
        n17780) );
  AOI211_X1 U19718 ( .C1(n11169), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17781), .B(n17780), .ZN(n17782) );
  NAND3_X1 U19719 ( .A1(n17784), .A2(n17783), .A3(n17782), .ZN(n17875) );
  AOI22_X1 U19720 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U19721 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U19722 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17785) );
  OAI21_X1 U19723 ( .B1(n11245), .B2(n19169), .A(n17785), .ZN(n17791) );
  AOI22_X1 U19724 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U19725 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17788) );
  AOI22_X1 U19726 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U19727 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17786) );
  NAND4_X1 U19728 ( .A1(n17789), .A2(n17788), .A3(n17787), .A4(n17786), .ZN(
        n17790) );
  AOI211_X1 U19729 ( .C1(n18043), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n17791), .B(n17790), .ZN(n17792) );
  NAND3_X1 U19730 ( .A1(n17794), .A2(n17793), .A3(n17792), .ZN(n17876) );
  NAND2_X1 U19731 ( .A1(n17875), .A2(n17876), .ZN(n17874) );
  NOR2_X1 U19732 ( .A1(n17870), .A2(n17874), .ZN(n17869) );
  AOI22_X1 U19733 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U19734 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17804) );
  INV_X1 U19735 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17796) );
  AOI22_X1 U19736 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18029), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17795) );
  OAI21_X1 U19737 ( .B1(n17238), .B2(n17796), .A(n17795), .ZN(n17802) );
  AOI22_X1 U19738 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17800) );
  AOI22_X1 U19739 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U19740 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U19741 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17797) );
  NAND4_X1 U19742 ( .A1(n17800), .A2(n17799), .A3(n17798), .A4(n17797), .ZN(
        n17801) );
  AOI211_X1 U19743 ( .C1(n17901), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17802), .B(n17801), .ZN(n17803) );
  NAND3_X1 U19744 ( .A1(n17805), .A2(n17804), .A3(n17803), .ZN(n17866) );
  NAND2_X1 U19745 ( .A1(n17869), .A2(n17866), .ZN(n17865) );
  NOR2_X1 U19746 ( .A1(n17861), .A2(n17865), .ZN(n17860) );
  AOI22_X1 U19747 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17816) );
  AOI22_X1 U19748 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U19749 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17807) );
  OAI21_X1 U19750 ( .B1(n11246), .B2(n19291), .A(n17807), .ZN(n17813) );
  AOI22_X1 U19751 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U19752 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17810) );
  AOI22_X1 U19753 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U19754 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17808) );
  NAND4_X1 U19755 ( .A1(n17811), .A2(n17810), .A3(n17809), .A4(n17808), .ZN(
        n17812) );
  AOI211_X1 U19756 ( .C1(n11170), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17813), .B(n17812), .ZN(n17814) );
  NAND3_X1 U19757 ( .A1(n17816), .A2(n17815), .A3(n17814), .ZN(n17843) );
  NAND2_X1 U19758 ( .A1(n17860), .A2(n17843), .ZN(n17854) );
  NOR2_X1 U19759 ( .A1(n17855), .A2(n17854), .ZN(n17853) );
  AOI22_X1 U19760 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17826) );
  AOI22_X1 U19761 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U19762 ( .A1(n11215), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17817) );
  OAI21_X1 U19763 ( .B1(n11246), .B2(n19209), .A(n17817), .ZN(n17823) );
  AOI22_X1 U19764 ( .A1(n17806), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U19765 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U19766 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U19767 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17818) );
  NAND4_X1 U19768 ( .A1(n17821), .A2(n17820), .A3(n17819), .A4(n17818), .ZN(
        n17822) );
  AOI211_X1 U19769 ( .C1(n17221), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17823), .B(n17822), .ZN(n17824) );
  NAND3_X1 U19770 ( .A1(n17826), .A2(n17825), .A3(n17824), .ZN(n17846) );
  NAND2_X1 U19771 ( .A1(n17853), .A2(n17846), .ZN(n17845) );
  XNOR2_X1 U19772 ( .A(n17827), .B(n17845), .ZN(n21081) );
  OAI22_X1 U19773 ( .A1(n17829), .A2(n17828), .B1(n21081), .B2(n17951), .ZN(
        P3_U2673) );
  AOI22_X1 U19774 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U19775 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U19776 ( .A1(n11215), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17831) );
  AOI22_X1 U19777 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17830) );
  NAND4_X1 U19778 ( .A1(n17833), .A2(n17832), .A3(n17831), .A4(n17830), .ZN(
        n17839) );
  AOI22_X1 U19779 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U19780 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U19781 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U19782 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17834) );
  NAND4_X1 U19783 ( .A1(n17837), .A2(n17836), .A3(n17835), .A4(n17834), .ZN(
        n17838) );
  NOR2_X1 U19784 ( .A1(n17839), .A2(n17838), .ZN(n21029) );
  AND2_X1 U19785 ( .A1(n17951), .A2(n17840), .ZN(n17905) );
  NOR2_X1 U19786 ( .A1(n21063), .A2(n17840), .ZN(n17842) );
  AOI22_X1 U19787 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17905), .B1(n17842), 
        .B2(n20804), .ZN(n17841) );
  OAI21_X1 U19788 ( .B1(n21029), .B2(n17951), .A(n17841), .ZN(P3_U2682) );
  INV_X1 U19789 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20858) );
  NAND2_X1 U19790 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17842), .ZN(n17879) );
  NOR3_X1 U19791 ( .A1(n20835), .A2(n20823), .A3(n17879), .ZN(n17878) );
  NAND2_X1 U19792 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17878), .ZN(n17848) );
  NOR2_X1 U19793 ( .A1(n20858), .A2(n17848), .ZN(n17868) );
  NAND2_X1 U19794 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17868), .ZN(n17859) );
  OAI21_X1 U19795 ( .B1(n17860), .B2(n17843), .A(n17854), .ZN(n21098) );
  NAND3_X1 U19796 ( .A1(n17859), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17951), 
        .ZN(n17844) );
  OAI221_X1 U19797 ( .B1(n17859), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17951), 
        .C2(n21098), .A(n17844), .ZN(P3_U2676) );
  OAI21_X1 U19798 ( .B1(n17853), .B2(n17846), .A(n17845), .ZN(n21085) );
  NAND2_X1 U19799 ( .A1(n17951), .A2(n17859), .ZN(n17847) );
  OAI21_X1 U19800 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17956), .A(n17847), .ZN(
        n17856) );
  INV_X1 U19801 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20902) );
  OAI221_X1 U19802 ( .B1(n17856), .B2(n17946), .C1(n17856), .C2(n20902), .A(
        P3_EBX_REG_29__SCAN_IN), .ZN(n17852) );
  INV_X1 U19803 ( .A(n17848), .ZN(n17873) );
  INV_X1 U19804 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17849) );
  NAND3_X1 U19805 ( .A1(n17873), .A2(n17850), .A3(n17849), .ZN(n17851) );
  OAI211_X1 U19806 ( .C1(n17951), .C2(n21085), .A(n17852), .B(n17851), .ZN(
        P3_U2674) );
  AOI21_X1 U19807 ( .B1(n17855), .B2(n17854), .A(n17853), .ZN(n21086) );
  AOI22_X1 U19808 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17856), .B1(n21086), 
        .B2(n17954), .ZN(n17858) );
  NAND4_X1 U19809 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n17868), .A4(n20902), .ZN(n17857) );
  NAND2_X1 U19810 ( .A1(n17858), .A2(n17857), .ZN(P3_U2675) );
  INV_X1 U19811 ( .A(n17859), .ZN(n17864) );
  AOI21_X1 U19812 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17951), .A(n17868), .ZN(
        n17863) );
  AOI21_X1 U19813 ( .B1(n17861), .B2(n17865), .A(n17860), .ZN(n21068) );
  INV_X1 U19814 ( .A(n21068), .ZN(n17862) );
  OAI22_X1 U19815 ( .A1(n17864), .A2(n17863), .B1(n17862), .B2(n17951), .ZN(
        P3_U2677) );
  AOI21_X1 U19816 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17951), .A(n17873), .ZN(
        n17867) );
  OAI21_X1 U19817 ( .B1(n17869), .B2(n17866), .A(n17865), .ZN(n21067) );
  OAI22_X1 U19818 ( .A1(n17868), .A2(n17867), .B1(n21067), .B2(n17951), .ZN(
        P3_U2678) );
  AOI21_X1 U19819 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17951), .A(n17878), .ZN(
        n17872) );
  AOI21_X1 U19820 ( .B1(n17870), .B2(n17874), .A(n17869), .ZN(n21099) );
  INV_X1 U19821 ( .A(n21099), .ZN(n17871) );
  OAI22_X1 U19822 ( .A1(n17873), .A2(n17872), .B1(n17871), .B2(n17951), .ZN(
        P3_U2679) );
  NOR2_X1 U19823 ( .A1(n20823), .A2(n17879), .ZN(n17893) );
  AOI21_X1 U19824 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17951), .A(n17893), .ZN(
        n17877) );
  OAI21_X1 U19825 ( .B1(n17876), .B2(n17875), .A(n17874), .ZN(n21110) );
  OAI22_X1 U19826 ( .A1(n17878), .A2(n17877), .B1(n17951), .B2(n21110), .ZN(
        P3_U2680) );
  OAI21_X1 U19827 ( .B1(n20823), .B2(n17954), .A(n17879), .ZN(n17880) );
  INV_X1 U19828 ( .A(n17880), .ZN(n17892) );
  AOI22_X1 U19829 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17890) );
  AOI22_X1 U19830 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17889) );
  AOI22_X1 U19831 ( .A1(n11215), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17881) );
  OAI21_X1 U19832 ( .B1(n11245), .B2(n19209), .A(n17881), .ZN(n17887) );
  AOI22_X1 U19833 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17885) );
  AOI22_X1 U19834 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17884) );
  AOI22_X1 U19835 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17934), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17883) );
  AOI22_X1 U19836 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17882) );
  NAND4_X1 U19837 ( .A1(n17885), .A2(n17884), .A3(n17883), .A4(n17882), .ZN(
        n17886) );
  AOI211_X1 U19838 ( .C1(n11169), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17887), .B(n17886), .ZN(n17888) );
  NAND3_X1 U19839 ( .A1(n17890), .A2(n17889), .A3(n17888), .ZN(n21037) );
  INV_X1 U19840 ( .A(n21037), .ZN(n17891) );
  OAI22_X1 U19841 ( .A1(n17893), .A2(n17892), .B1(n17891), .B2(n17951), .ZN(
        P3_U2681) );
  AOI22_X1 U19842 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U19843 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U19844 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17894) );
  OAI21_X1 U19845 ( .B1(n11245), .B2(n19291), .A(n17894), .ZN(n17900) );
  AOI22_X1 U19846 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11203), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U19847 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U19848 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17896) );
  AOI22_X1 U19849 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17895) );
  NAND4_X1 U19850 ( .A1(n17898), .A2(n17897), .A3(n17896), .A4(n17895), .ZN(
        n17899) );
  AOI211_X1 U19851 ( .C1(n17901), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17900), .B(n17899), .ZN(n17902) );
  NAND3_X1 U19852 ( .A1(n17904), .A2(n17903), .A3(n17902), .ZN(n21033) );
  INV_X1 U19853 ( .A(n21033), .ZN(n17907) );
  OAI21_X1 U19854 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17933), .A(n17905), .ZN(
        n17906) );
  OAI21_X1 U19855 ( .B1(n17907), .B2(n17951), .A(n17906), .ZN(P3_U2683) );
  AOI22_X1 U19856 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17911) );
  AOI22_X1 U19857 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17910) );
  AOI22_X1 U19858 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U19859 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11212), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17908) );
  NAND4_X1 U19860 ( .A1(n17911), .A2(n17910), .A3(n17909), .A4(n17908), .ZN(
        n17917) );
  AOI22_X1 U19861 ( .A1(n11215), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17915) );
  AOI22_X1 U19862 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17914) );
  AOI22_X1 U19863 ( .A1(n18028), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U19864 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17912) );
  NAND4_X1 U19865 ( .A1(n17915), .A2(n17914), .A3(n17913), .A4(n17912), .ZN(
        n17916) );
  NOR2_X1 U19866 ( .A1(n17917), .A2(n17916), .ZN(n21055) );
  OAI21_X1 U19867 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17918), .A(n17920), .ZN(
        n17919) );
  AOI22_X1 U19868 ( .A1(n17954), .A2(n21055), .B1(n17919), .B2(n17951), .ZN(
        P3_U2685) );
  INV_X1 U19869 ( .A(n17920), .ZN(n17921) );
  OAI21_X1 U19870 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17921), .A(n17951), .ZN(
        n17932) );
  AOI22_X1 U19871 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U19872 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11215), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19873 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17923) );
  AOI22_X1 U19874 ( .A1(n17934), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17922) );
  NAND4_X1 U19875 ( .A1(n17925), .A2(n17924), .A3(n17923), .A4(n17922), .ZN(
        n17931) );
  AOI22_X1 U19876 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U19877 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U19878 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17927) );
  AOI22_X1 U19879 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17926) );
  NAND4_X1 U19880 ( .A1(n17929), .A2(n17928), .A3(n17927), .A4(n17926), .ZN(
        n17930) );
  NOR2_X1 U19881 ( .A1(n17931), .A2(n17930), .ZN(n21050) );
  OAI22_X1 U19882 ( .A1(n17933), .A2(n17932), .B1(n21050), .B2(n17951), .ZN(
        P3_U2684) );
  AOI22_X1 U19883 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17938) );
  AOI22_X1 U19884 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U19885 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17992), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n18028), .ZN(n17936) );
  AOI22_X1 U19886 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17934), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18016), .ZN(n17935) );
  NAND4_X1 U19887 ( .A1(n17938), .A2(n17937), .A3(n17936), .A4(n17935), .ZN(
        n17944) );
  AOI22_X1 U19888 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18041), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n11177), .ZN(n17942) );
  AOI22_X1 U19889 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17941) );
  AOI22_X1 U19890 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18044), .ZN(n17940) );
  AOI22_X1 U19891 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17939) );
  NAND4_X1 U19892 ( .A1(n17942), .A2(n17941), .A3(n17940), .A4(n17939), .ZN(
        n17943) );
  NOR2_X1 U19893 ( .A1(n17944), .A2(n17943), .ZN(n21060) );
  OAI211_X1 U19894 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n17947), .A(n17946), .B(
        n17945), .ZN(n17949) );
  NAND2_X1 U19895 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17953), .ZN(n17948) );
  OAI211_X1 U19896 ( .C1(n21060), .C2(n17951), .A(n17949), .B(n17948), .ZN(
        P3_U2686) );
  NOR2_X1 U19897 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20550) );
  OR2_X1 U19898 ( .A1(n20550), .A2(n17950), .ZN(n20536) );
  INV_X1 U19899 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20532) );
  OAI222_X1 U19900 ( .A1(n20536), .A2(n17956), .B1(n20532), .B2(n17952), .C1(
        n19418), .C2(n17951), .ZN(P3_U2702) );
  AOI22_X1 U19901 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17954), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17953), .ZN(n17955) );
  OAI21_X1 U19902 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17956), .A(n17955), .ZN(
        P3_U2703) );
  NAND2_X1 U19903 ( .A1(n21668), .A2(n21676), .ZN(n17959) );
  INV_X1 U19904 ( .A(n21670), .ZN(n20528) );
  INV_X1 U19905 ( .A(n21628), .ZN(n17957) );
  OAI21_X1 U19906 ( .B1(n17957), .B2(n20470), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17958) );
  OAI21_X1 U19907 ( .B1(n17959), .B2(n20528), .A(n17958), .ZN(P3_U2634) );
  OAI21_X1 U19908 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n17961), .A(n17960), .ZN(
        n21686) );
  INV_X1 U19909 ( .A(n19086), .ZN(n17963) );
  OAI21_X1 U19910 ( .B1(n20467), .B2(n18537), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17962) );
  OAI221_X1 U19911 ( .B1(n18537), .B2(n21686), .C1(n18537), .C2(n17963), .A(
        n17962), .ZN(P3_U2863) );
  AOI22_X1 U19912 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U19913 ( .A1(n11207), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17973) );
  AOI22_X1 U19914 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17964) );
  OAI21_X1 U19915 ( .B1(n11218), .B2(n19169), .A(n17964), .ZN(n17970) );
  AOI22_X1 U19916 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U19917 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17967) );
  AOI22_X1 U19918 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17966) );
  AOI22_X1 U19919 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17965) );
  NAND4_X1 U19920 ( .A1(n17968), .A2(n17967), .A3(n17966), .A4(n17965), .ZN(
        n17969) );
  AOI211_X1 U19921 ( .C1(n17971), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n17970), .B(n17969), .ZN(n17972) );
  NAND3_X1 U19922 ( .A1(n17974), .A2(n17973), .A3(n17972), .ZN(n21225) );
  INV_X1 U19923 ( .A(n21653), .ZN(n21219) );
  NAND2_X1 U19924 ( .A1(n21211), .A2(n17977), .ZN(n21164) );
  NAND2_X1 U19925 ( .A1(n21165), .A2(n21164), .ZN(n21155) );
  OAI21_X1 U19926 ( .B1(n17980), .B2(n17979), .A(n21656), .ZN(n21650) );
  INV_X1 U19927 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18133) );
  AOI22_X1 U19928 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U19929 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U19930 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U19931 ( .A1(n11213), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17981) );
  NAND4_X1 U19932 ( .A1(n17984), .A2(n17983), .A3(n17982), .A4(n17981), .ZN(
        n17990) );
  AOI22_X1 U19933 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17988) );
  AOI22_X1 U19934 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U19935 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19936 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11168), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17985) );
  NAND4_X1 U19937 ( .A1(n17988), .A2(n17987), .A3(n17986), .A4(n17985), .ZN(
        n17989) );
  AOI22_X1 U19938 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19939 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U19940 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U19941 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17993) );
  NAND4_X1 U19942 ( .A1(n17996), .A2(n17995), .A3(n17994), .A4(n17993), .ZN(
        n18003) );
  AOI22_X1 U19943 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U19944 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18000) );
  AOI22_X1 U19945 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U19946 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17998) );
  NAND4_X1 U19947 ( .A1(n18001), .A2(n18000), .A3(n17999), .A4(n17998), .ZN(
        n18002) );
  INV_X1 U19948 ( .A(n21012), .ZN(n18099) );
  AOI22_X1 U19949 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18007) );
  AOI22_X1 U19950 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18006) );
  AOI22_X1 U19951 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18018), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U19952 ( .A1(n11212), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18004) );
  NAND4_X1 U19953 ( .A1(n18007), .A2(n18006), .A3(n18005), .A4(n18004), .ZN(
        n18013) );
  AOI22_X1 U19954 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11170), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18011) );
  AOI22_X1 U19955 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18015), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18010) );
  AOI22_X1 U19956 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18014), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18009) );
  AOI22_X1 U19957 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17991), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18008) );
  NAND4_X1 U19958 ( .A1(n18011), .A2(n18010), .A3(n18009), .A4(n18008), .ZN(
        n18012) );
  AOI22_X1 U19959 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18028), .B1(
        n11203), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U19960 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n18014), .ZN(n18021) );
  AOI22_X1 U19961 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18016), .B1(
        n18015), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18020) );
  AOI22_X1 U19962 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18018), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17992), .ZN(n18019) );
  AOI22_X1 U19963 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n18044), .ZN(n18027) );
  AOI22_X1 U19964 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U19965 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11207), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18025) );
  AOI22_X1 U19966 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17997), .ZN(n18024) );
  AOI22_X1 U19967 ( .A1(n17806), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18040) );
  AOI22_X1 U19968 ( .A1(n18029), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18039) );
  AOI22_X1 U19969 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17992), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18030) );
  OAI21_X1 U19970 ( .B1(n11218), .B2(n19334), .A(n18030), .ZN(n18037) );
  AOI22_X1 U19971 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18031), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18035) );
  AOI22_X1 U19972 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U19973 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U19974 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18032) );
  NAND4_X1 U19975 ( .A1(n18035), .A2(n18034), .A3(n18033), .A4(n18032), .ZN(
        n18036) );
  AOI211_X1 U19976 ( .C1(n17997), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n18037), .B(n18036), .ZN(n18038) );
  NAND3_X1 U19977 ( .A1(n18040), .A2(n18039), .A3(n18038), .ZN(n18098) );
  AOI22_X1 U19978 ( .A1(n11170), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17997), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18053) );
  AOI22_X1 U19979 ( .A1(n17221), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18052) );
  AOI22_X1 U19980 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11212), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18042) );
  OAI21_X1 U19981 ( .B1(n11218), .B2(n19250), .A(n18042), .ZN(n18050) );
  AOI22_X1 U19982 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U19983 ( .A1(n11177), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U19984 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18046) );
  AOI22_X1 U19985 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11169), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18045) );
  NAND4_X1 U19986 ( .A1(n18048), .A2(n18047), .A3(n18046), .A4(n18045), .ZN(
        n18049) );
  AOI211_X1 U19987 ( .C1(n11168), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n18050), .B(n18049), .ZN(n18051) );
  NAND3_X1 U19988 ( .A1(n18053), .A2(n18052), .A3(n18051), .ZN(n18074) );
  NOR2_X1 U19989 ( .A1(n18329), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18208) );
  INV_X1 U19990 ( .A(n18208), .ZN(n18131) );
  OAI21_X1 U19991 ( .B1(n18133), .B2(n21505), .A(n18131), .ZN(n18093) );
  INV_X1 U19992 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21584) );
  NAND2_X1 U19993 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21505), .ZN(
        n18086) );
  XNOR2_X1 U19994 ( .A(n21012), .B(n18054), .ZN(n18055) );
  NAND2_X1 U19995 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18055), .ZN(
        n18073) );
  XOR2_X1 U19996 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18055), .Z(
        n18483) );
  NAND2_X1 U19997 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18056), .ZN(
        n18069) );
  NAND2_X1 U19998 ( .A1(n21145), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18068) );
  AOI22_X1 U19999 ( .A1(n11169), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11203), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U20000 ( .A1(n18031), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17971), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18059) );
  AOI22_X1 U20001 ( .A1(n11168), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18018), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U20002 ( .A1(n17992), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18016), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18057) );
  NAND4_X1 U20003 ( .A1(n18060), .A2(n18059), .A3(n18058), .A4(n18057), .ZN(
        n18067) );
  AOI22_X1 U20004 ( .A1(n17991), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18028), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18065) );
  AOI22_X1 U20005 ( .A1(n17997), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11177), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18064) );
  AOI22_X1 U20006 ( .A1(n11171), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18061), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U20007 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18041), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18062) );
  NAND4_X1 U20008 ( .A1(n18065), .A2(n18064), .A3(n18063), .A4(n18062), .ZN(
        n18066) );
  INV_X1 U20009 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21427) );
  NOR2_X1 U20010 ( .A1(n18526), .A2(n21427), .ZN(n18525) );
  NAND2_X1 U20011 ( .A1(n18068), .A2(n18517), .ZN(n18511) );
  NAND2_X1 U20012 ( .A1(n18069), .A2(n18510), .ZN(n18070) );
  NAND2_X1 U20013 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18070), .ZN(
        n18072) );
  XNOR2_X1 U20014 ( .A(n21015), .B(n18071), .ZN(n18499) );
  INV_X1 U20015 ( .A(n18074), .ZN(n21007) );
  XNOR2_X1 U20016 ( .A(n21007), .B(n18075), .ZN(n18077) );
  NAND2_X1 U20017 ( .A1(n18077), .A2(n18076), .ZN(n18078) );
  XOR2_X1 U20018 ( .A(n21002), .B(n18079), .Z(n18080) );
  XOR2_X1 U20019 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18080), .Z(
        n18462) );
  NAND2_X1 U20020 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18080), .ZN(
        n18081) );
  AOI21_X1 U20021 ( .B1(n21492), .B2(n18082), .A(n18329), .ZN(n18084) );
  NAND2_X1 U20022 ( .A1(n18084), .A2(n18148), .ZN(n18085) );
  INV_X1 U20023 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21329) );
  AOI22_X1 U20024 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21505), .B1(
        n18329), .B2(n21329), .ZN(n18442) );
  INV_X1 U20025 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21616) );
  INV_X1 U20026 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21597) );
  NOR2_X1 U20027 ( .A1(n21616), .A2(n21597), .ZN(n18397) );
  INV_X1 U20028 ( .A(n18397), .ZN(n21333) );
  INV_X1 U20029 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21341) );
  NOR2_X1 U20030 ( .A1(n21333), .A2(n21341), .ZN(n21349) );
  AND2_X1 U20031 ( .A1(n21349), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n21356) );
  NAND2_X1 U20032 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21356), .ZN(
        n21360) );
  INV_X1 U20033 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21372) );
  NOR2_X1 U20034 ( .A1(n21360), .A2(n21372), .ZN(n21379) );
  NAND2_X1 U20035 ( .A1(n21379), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21552) );
  INV_X1 U20036 ( .A(n21552), .ZN(n21222) );
  NAND2_X1 U20037 ( .A1(n18403), .A2(n21222), .ZN(n18091) );
  NOR2_X1 U20038 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18377) );
  NAND2_X1 U20039 ( .A1(n21616), .A2(n21597), .ZN(n18418) );
  INV_X1 U20040 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21347) );
  NAND2_X1 U20041 ( .A1(n21341), .A2(n21347), .ZN(n18169) );
  NOR3_X1 U20042 ( .A1(n18088), .A2(n18418), .A3(n18169), .ZN(n18089) );
  INV_X1 U20043 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21576) );
  NAND2_X1 U20044 ( .A1(n18370), .A2(n21576), .ZN(n18369) );
  NOR2_X1 U20045 ( .A1(n21584), .A2(n21576), .ZN(n21564) );
  INV_X1 U20046 ( .A(n18090), .ZN(n18092) );
  NAND2_X1 U20047 ( .A1(n18092), .A2(n18091), .ZN(n18253) );
  NAND2_X1 U20048 ( .A1(n21564), .A2(n18253), .ZN(n18132) );
  XNOR2_X1 U20049 ( .A(n18093), .B(n18186), .ZN(n21570) );
  NAND3_X1 U20050 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18410) );
  NAND2_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20701) );
  NAND2_X1 U20052 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20758) );
  INV_X1 U20053 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20543) );
  NOR2_X1 U20054 ( .A1(n18096), .A2(n20543), .ZN(n18361) );
  AOI21_X1 U20055 ( .B1(n18437), .B2(n18096), .A(n18515), .ZN(n18364) );
  OAI21_X1 U20056 ( .B1(n18361), .B2(n18528), .A(n18364), .ZN(n18139) );
  NOR3_X1 U20057 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18319), .A3(
        n18096), .ZN(n18140) );
  INV_X1 U20058 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20775) );
  INV_X1 U20059 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20764) );
  NAND2_X1 U20060 ( .A1(n18135), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18136) );
  OAI21_X1 U20061 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18361), .A(
        n18136), .ZN(n20771) );
  OAI22_X1 U20062 ( .A1(n21620), .A2(n20775), .B1(n20771), .B2(n18310), .ZN(
        n18097) );
  AOI211_X1 U20063 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18139), .A(
        n18140), .B(n18097), .ZN(n18128) );
  OAI21_X1 U20064 ( .B1(n21145), .B2(n18526), .A(n21020), .ZN(n18107) );
  AND2_X1 U20065 ( .A1(n18098), .A2(n18107), .ZN(n18105) );
  NAND2_X1 U20066 ( .A1(n18105), .A2(n18099), .ZN(n18103) );
  NOR2_X1 U20067 ( .A1(n21007), .A2(n18103), .ZN(n18102) );
  INV_X1 U20068 ( .A(n21002), .ZN(n18100) );
  NAND2_X1 U20069 ( .A1(n18102), .A2(n18100), .ZN(n18101) );
  NOR2_X1 U20070 ( .A1(n21492), .A2(n18101), .ZN(n18124) );
  XNOR2_X1 U20071 ( .A(n21225), .B(n18101), .ZN(n18452) );
  XNOR2_X1 U20072 ( .A(n21002), .B(n18102), .ZN(n18118) );
  XOR2_X1 U20073 ( .A(n21007), .B(n18103), .Z(n18104) );
  NAND2_X1 U20074 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18104), .ZN(
        n18117) );
  INV_X1 U20075 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21293) );
  XNOR2_X1 U20076 ( .A(n21293), .B(n18104), .ZN(n18476) );
  XNOR2_X1 U20077 ( .A(n21012), .B(n18105), .ZN(n18114) );
  XNOR2_X1 U20078 ( .A(n21015), .B(n18107), .ZN(n18106) );
  NAND2_X1 U20079 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18106), .ZN(
        n18113) );
  INV_X1 U20080 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21274) );
  XNOR2_X1 U20081 ( .A(n21274), .B(n18106), .ZN(n18497) );
  OAI21_X1 U20082 ( .B1(n18526), .B2(n18108), .A(n18107), .ZN(n18109) );
  NAND2_X1 U20083 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18109), .ZN(
        n18112) );
  XOR2_X1 U20084 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n18109), .Z(
        n18509) );
  INV_X1 U20085 ( .A(n18526), .ZN(n21146) );
  AOI21_X1 U20086 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11389), .A(
        n21146), .ZN(n18111) );
  NOR2_X1 U20087 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n11389), .ZN(
        n18110) );
  AOI221_X1 U20088 ( .B1(n21146), .B2(n11389), .C1(n18111), .C2(n21427), .A(
        n18110), .ZN(n18508) );
  NAND2_X1 U20089 ( .A1(n18509), .A2(n18508), .ZN(n18507) );
  NAND2_X1 U20090 ( .A1(n18114), .A2(n18115), .ZN(n18116) );
  NAND2_X1 U20091 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18485), .ZN(
        n18484) );
  NAND2_X1 U20092 ( .A1(n18116), .A2(n18484), .ZN(n18475) );
  NAND2_X1 U20093 ( .A1(n18476), .A2(n18475), .ZN(n18474) );
  NAND2_X1 U20094 ( .A1(n18118), .A2(n18119), .ZN(n18120) );
  INV_X1 U20095 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21316) );
  NAND2_X1 U20096 ( .A1(n18124), .A2(n18121), .ZN(n18125) );
  INV_X1 U20097 ( .A(n18121), .ZN(n18123) );
  NAND2_X1 U20098 ( .A1(n18124), .A2(n18123), .ZN(n18122) );
  INV_X1 U20099 ( .A(n18432), .ZN(n18417) );
  NAND2_X1 U20100 ( .A1(n21222), .A2(n18417), .ZN(n18164) );
  NOR2_X1 U20101 ( .A1(n21373), .A2(n18389), .ZN(n18151) );
  AOI21_X1 U20102 ( .B1(n18520), .B2(n21377), .A(n18151), .ZN(n18163) );
  OAI21_X1 U20103 ( .B1(n21564), .B2(n18164), .A(n18163), .ZN(n18368) );
  INV_X1 U20104 ( .A(n21564), .ZN(n18126) );
  NOR2_X1 U20105 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18126), .ZN(
        n21553) );
  INV_X1 U20106 ( .A(n18164), .ZN(n18371) );
  AOI22_X1 U20107 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18368), .B1(
        n21553), .B2(n18371), .ZN(n18127) );
  OAI211_X1 U20108 ( .C1(n18388), .C2(n21570), .A(n18128), .B(n18127), .ZN(
        P3_U2812) );
  NAND2_X1 U20109 ( .A1(n21564), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21223) );
  INV_X1 U20110 ( .A(n21223), .ZN(n18129) );
  NAND2_X1 U20111 ( .A1(n21222), .A2(n18129), .ZN(n21224) );
  INV_X1 U20112 ( .A(n18202), .ZN(n18223) );
  INV_X1 U20113 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21543) );
  NAND3_X1 U20114 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21373), .ZN(n21535) );
  NOR3_X1 U20115 ( .A1(n21223), .A2(n21543), .A3(n21377), .ZN(n21538) );
  INV_X1 U20116 ( .A(n21538), .ZN(n18130) );
  AOI22_X1 U20117 ( .A1(n18443), .A2(n21535), .B1(n18520), .B2(n18130), .ZN(
        n18220) );
  NOR2_X1 U20118 ( .A1(n18131), .A2(n18186), .ZN(n18198) );
  NOR3_X1 U20119 ( .A1(n21505), .A2(n18133), .A3(n18132), .ZN(n18207) );
  NOR2_X1 U20120 ( .A1(n18198), .A2(n18207), .ZN(n18134) );
  XNOR2_X1 U20121 ( .A(n18134), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21540) );
  INV_X1 U20122 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18137) );
  AND3_X1 U20123 ( .A1(n18137), .A2(n18280), .A3(n18135), .ZN(n18144) );
  NOR2_X1 U20124 ( .A1(n18214), .A2(n20543), .ZN(n18211) );
  AOI21_X1 U20125 ( .B1(n18137), .B2(n18136), .A(n18211), .ZN(n18138) );
  INV_X1 U20126 ( .A(n18138), .ZN(n20784) );
  NAND2_X1 U20127 ( .A1(n11176), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18142) );
  OAI21_X1 U20128 ( .B1(n18140), .B2(n18139), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18141) );
  OAI211_X1 U20129 ( .C1(n18310), .C2(n20784), .A(n18142), .B(n18141), .ZN(
        n18143) );
  AOI211_X1 U20130 ( .C1(n18444), .C2(n21540), .A(n18144), .B(n18143), .ZN(
        n18145) );
  OAI221_X1 U20131 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18223), 
        .C1(n21543), .C2(n18220), .A(n18145), .ZN(P3_U2811) );
  NOR2_X1 U20132 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21378), .ZN(
        n18155) );
  NAND2_X1 U20133 ( .A1(n18520), .A2(n21377), .ZN(n18154) );
  NOR2_X1 U20134 ( .A1(n18319), .A2(n18146), .ZN(n18158) );
  INV_X1 U20135 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20729) );
  NOR2_X1 U20136 ( .A1(n18146), .A2(n20543), .ZN(n20724) );
  AOI21_X1 U20137 ( .B1(n18437), .B2(n18146), .A(n18515), .ZN(n18380) );
  OAI21_X1 U20138 ( .B1(n20724), .B2(n18528), .A(n18380), .ZN(n18157) );
  NAND2_X1 U20139 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20724), .ZN(
        n20735) );
  OAI21_X1 U20140 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20724), .A(
        n20735), .ZN(n20725) );
  NAND2_X1 U20141 ( .A1(n11176), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21386) );
  OAI21_X1 U20142 ( .B1(n18310), .B2(n20725), .A(n21386), .ZN(n18147) );
  AOI221_X1 U20143 ( .B1(n18158), .B2(n20729), .C1(n18157), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18147), .ZN(n18153) );
  NAND4_X1 U20144 ( .A1(n18148), .A2(n18329), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18421) );
  INV_X1 U20145 ( .A(n18421), .ZN(n18404) );
  INV_X1 U20146 ( .A(n18418), .ZN(n18407) );
  NAND3_X1 U20147 ( .A1(n18401), .A2(n18407), .A3(n21329), .ZN(n18394) );
  NOR2_X1 U20148 ( .A1(n18169), .A2(n18394), .ZN(n18376) );
  AOI22_X1 U20149 ( .A1(n21379), .A2(n18404), .B1(n18377), .B2(n18376), .ZN(
        n18149) );
  XNOR2_X1 U20150 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18149), .ZN(
        n21384) );
  NAND2_X1 U20151 ( .A1(n18087), .A2(n21383), .ZN(n18150) );
  AOI22_X1 U20152 ( .A1(n18444), .A2(n21384), .B1(n18151), .B2(n18150), .ZN(
        n18152) );
  OAI211_X1 U20153 ( .C1(n18155), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        P3_U2815) );
  AOI22_X1 U20154 ( .A1(n18329), .A2(n21584), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21505), .ZN(n18156) );
  XOR2_X1 U20155 ( .A(n18253), .B(n18156), .Z(n21586) );
  INV_X1 U20156 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21588) );
  INV_X1 U20157 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20741) );
  AND2_X1 U20158 ( .A1(n11305), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18363) );
  AOI21_X1 U20159 ( .B1(n20741), .B2(n20735), .A(n18363), .ZN(n20736) );
  AOI22_X1 U20160 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18157), .B1(
        n18360), .B2(n20736), .ZN(n18160) );
  OAI211_X1 U20161 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18158), .B(n20758), .ZN(n18159) );
  OAI211_X1 U20162 ( .C1(n21588), .C2(n21620), .A(n18160), .B(n18159), .ZN(
        n18161) );
  AOI21_X1 U20163 ( .B1(n18444), .B2(n21586), .A(n18161), .ZN(n18162) );
  OAI221_X1 U20164 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18164), 
        .C1(n21584), .C2(n18163), .A(n18162), .ZN(P3_U2814) );
  NOR2_X1 U20165 ( .A1(n18166), .A2(n20543), .ZN(n18391) );
  AOI21_X1 U20166 ( .B1(n18437), .B2(n18166), .A(n18231), .ZN(n18165) );
  OAI21_X1 U20167 ( .B1(n18391), .B2(n18165), .A(n18527), .ZN(n18179) );
  OR2_X1 U20168 ( .A1(n18166), .A2(n18319), .ZN(n18176) );
  NAND2_X1 U20169 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18391), .ZN(
        n20698) );
  OAI21_X1 U20170 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18391), .A(
        n20698), .ZN(n20683) );
  OAI22_X1 U20171 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18176), .B1(
        n20683), .B2(n18310), .ZN(n18167) );
  AOI21_X1 U20172 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18179), .A(
        n18167), .ZN(n18173) );
  OAI22_X1 U20173 ( .A1(n21346), .A2(n18532), .B1(n18168), .B2(n18389), .ZN(
        n18183) );
  NAND2_X1 U20174 ( .A1(n21356), .A2(n18404), .ZN(n18181) );
  OAI211_X1 U20175 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n18394), .A(
        n18181), .B(n18169), .ZN(n18170) );
  NAND2_X1 U20176 ( .A1(n18397), .A2(n18404), .ZN(n18395) );
  INV_X1 U20177 ( .A(n18376), .ZN(n18180) );
  OAI221_X1 U20178 ( .B1(n18170), .B2(n21347), .C1(n18170), .C2(n18395), .A(
        n18180), .ZN(n21350) );
  AOI22_X1 U20179 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18183), .B1(
        n18444), .B2(n21350), .ZN(n18172) );
  NAND2_X1 U20180 ( .A1(n11176), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21351) );
  NAND3_X1 U20181 ( .A1(n21349), .A2(n21347), .A3(n18417), .ZN(n18171) );
  NAND4_X1 U20182 ( .A1(n18173), .A2(n18172), .A3(n21351), .A4(n18171), .ZN(
        P3_U2818) );
  INV_X1 U20183 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21359) );
  NAND2_X1 U20184 ( .A1(n21356), .A2(n21359), .ZN(n21596) );
  INV_X1 U20185 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20712) );
  NOR2_X1 U20186 ( .A1(n21620), .A2(n20712), .ZN(n18178) );
  INV_X1 U20187 ( .A(n20698), .ZN(n18174) );
  NAND2_X1 U20188 ( .A1(n18379), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18378) );
  OAI21_X1 U20189 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18174), .A(
        n18378), .ZN(n20699) );
  OAI21_X1 U20190 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n20701), .ZN(n18175) );
  OAI22_X1 U20191 ( .A1(n18310), .A2(n20699), .B1(n18176), .B2(n18175), .ZN(
        n18177) );
  AOI211_X1 U20192 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18179), .A(
        n18178), .B(n18177), .ZN(n18185) );
  NAND2_X1 U20193 ( .A1(n18181), .A2(n18180), .ZN(n18182) );
  XNOR2_X1 U20194 ( .A(n18182), .B(n21359), .ZN(n21590) );
  AOI22_X1 U20195 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18183), .B1(
        n18444), .B2(n21590), .ZN(n18184) );
  OAI211_X1 U20196 ( .C1(n18432), .C2(n21596), .A(n18185), .B(n18184), .ZN(
        P3_U2817) );
  INV_X1 U20197 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18219) );
  NOR2_X1 U20198 ( .A1(n18219), .A2(n21543), .ZN(n21237) );
  NAND2_X1 U20199 ( .A1(n21237), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21526) );
  INV_X1 U20200 ( .A(n21526), .ZN(n21390) );
  INV_X1 U20201 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21513) );
  NOR2_X1 U20202 ( .A1(n21223), .A2(n21526), .ZN(n18252) );
  AOI22_X1 U20203 ( .A1(n18520), .A2(n21233), .B1(n18443), .B2(n21236), .ZN(
        n18206) );
  INV_X1 U20204 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18205) );
  NAND4_X1 U20205 ( .A1(n18208), .A2(n18219), .A3(n21543), .A4(n18205), .ZN(
        n18224) );
  INV_X1 U20206 ( .A(n18258), .ZN(n18187) );
  AOI21_X1 U20207 ( .B1(n18224), .B2(n18259), .A(n18187), .ZN(n18225) );
  XNOR2_X1 U20208 ( .A(n18225), .B(n21513), .ZN(n21396) );
  INV_X1 U20209 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20816) );
  INV_X1 U20210 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20806) );
  INV_X1 U20211 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18213) );
  NAND2_X1 U20212 ( .A1(n18188), .A2(n18280), .ZN(n18195) );
  AOI221_X1 U20213 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n20816), .C2(n20806), .A(
        n18195), .ZN(n18193) );
  NAND2_X1 U20214 ( .A1(n18188), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18210) );
  NOR2_X1 U20215 ( .A1(n20806), .A2(n18210), .ZN(n18189) );
  NOR2_X1 U20216 ( .A1(n18227), .A2(n20543), .ZN(n18236) );
  INV_X1 U20217 ( .A(n18236), .ZN(n18230) );
  OAI21_X1 U20218 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18189), .A(
        n18230), .ZN(n20822) );
  OAI22_X1 U20219 ( .A1(n18211), .A2(n18528), .B1(n18188), .B2(n18488), .ZN(
        n18190) );
  NOR2_X1 U20220 ( .A1(n18515), .A2(n18190), .ZN(n18212) );
  OAI21_X1 U20221 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18320), .A(
        n18212), .ZN(n18197) );
  AOI22_X1 U20222 ( .A1(n11176), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18197), .ZN(n18191) );
  OAI21_X1 U20223 ( .B1(n20822), .B2(n18310), .A(n18191), .ZN(n18192) );
  AOI211_X1 U20224 ( .C1(n21396), .C2(n18444), .A(n18193), .B(n18192), .ZN(
        n18194) );
  OAI221_X1 U20225 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18278), 
        .C1(n21513), .C2(n18206), .A(n18194), .ZN(P3_U2808) );
  INV_X1 U20226 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20814) );
  NOR2_X1 U20227 ( .A1(n21620), .A2(n20814), .ZN(n21226) );
  XNOR2_X1 U20228 ( .A(n20806), .B(n18210), .ZN(n20811) );
  OAI22_X1 U20229 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18195), .B1(
        n18310), .B2(n20811), .ZN(n18196) );
  AOI211_X1 U20230 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18197), .A(
        n21226), .B(n18196), .ZN(n18204) );
  NOR2_X1 U20231 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U20232 ( .A1(n21237), .A2(n18207), .B1(n18199), .B2(n18198), .ZN(
        n18200) );
  XNOR2_X1 U20233 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18200), .ZN(
        n21227) );
  NAND2_X1 U20234 ( .A1(n18205), .A2(n21237), .ZN(n21241) );
  INV_X1 U20235 ( .A(n21241), .ZN(n18201) );
  AOI22_X1 U20236 ( .A1(n18444), .A2(n21227), .B1(n18202), .B2(n18201), .ZN(
        n18203) );
  OAI211_X1 U20237 ( .C1(n18206), .C2(n18205), .A(n18204), .B(n18203), .ZN(
        P3_U2809) );
  NAND2_X1 U20238 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18219), .ZN(
        n21551) );
  OAI221_X1 U20239 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18208), 
        .C1(n21543), .C2(n18207), .A(n18258), .ZN(n18209) );
  XNOR2_X1 U20240 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18209), .ZN(
        n21546) );
  OAI21_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18211), .A(
        n18210), .ZN(n20794) );
  INV_X1 U20242 ( .A(n20794), .ZN(n18217) );
  INV_X1 U20243 ( .A(n18320), .ZN(n18216) );
  AOI221_X1 U20244 ( .B1(n18214), .B2(n18213), .C1(n19252), .C2(n18213), .A(
        n18212), .ZN(n18215) );
  AOI221_X1 U20245 ( .B1(n18360), .B2(n18217), .C1(n18216), .C2(n18217), .A(
        n18215), .ZN(n18218) );
  NAND2_X1 U20246 ( .A1(n11176), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21548) );
  OAI211_X1 U20247 ( .C1(n18220), .C2(n18219), .A(n18218), .B(n21548), .ZN(
        n18221) );
  AOI21_X1 U20248 ( .B1(n18444), .B2(n21546), .A(n18221), .ZN(n18222) );
  OAI21_X1 U20249 ( .B1(n18223), .B2(n21551), .A(n18222), .ZN(P3_U2810) );
  NOR2_X1 U20250 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18224), .ZN(
        n18255) );
  OAI221_X1 U20251 ( .B1(n18255), .B2(n18329), .C1(n18255), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18225), .ZN(n18226) );
  XOR2_X1 U20252 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18226), .Z(
        n21524) );
  NOR2_X1 U20253 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18320), .ZN(
        n18235) );
  INV_X1 U20254 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18232) );
  NOR2_X1 U20255 ( .A1(n18246), .A2(n19252), .ZN(n18229) );
  INV_X1 U20256 ( .A(n18229), .ZN(n18228) );
  NAND2_X1 U20257 ( .A1(n11176), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21522) );
  OAI21_X1 U20258 ( .B1(n18228), .B2(n18227), .A(n21522), .ZN(n18234) );
  AOI211_X1 U20259 ( .C1(n18231), .C2(n18230), .A(n18229), .B(n18515), .ZN(
        n18244) );
  NAND2_X1 U20260 ( .A1(n18246), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18265) );
  OAI21_X1 U20261 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18236), .A(
        n18265), .ZN(n20840) );
  OAI22_X1 U20262 ( .A1(n18244), .A2(n18232), .B1(n20840), .B2(n18310), .ZN(
        n18233) );
  AOI211_X1 U20263 ( .C1(n18236), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        n18241) );
  NAND2_X1 U20264 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21525) );
  NOR2_X1 U20265 ( .A1(n21525), .A2(n21236), .ZN(n21517) );
  OR2_X1 U20266 ( .A1(n21517), .A2(n18389), .ZN(n18237) );
  OR2_X1 U20267 ( .A1(n21525), .A2(n21233), .ZN(n21514) );
  NAND2_X1 U20268 ( .A1(n18520), .A2(n21514), .ZN(n18238) );
  OAI22_X1 U20269 ( .A1(n21236), .A2(n18237), .B1(n21233), .B2(n18238), .ZN(
        n18239) );
  OAI21_X1 U20270 ( .B1(n21517), .B2(n18389), .A(n18238), .ZN(n18272) );
  AOI22_X1 U20271 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18239), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18272), .ZN(n18240) );
  OAI211_X1 U20272 ( .C1(n18388), .C2(n21524), .A(n18241), .B(n18240), .ZN(
        P3_U2807) );
  INV_X1 U20273 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21417) );
  INV_X1 U20274 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18242) );
  NOR2_X1 U20275 ( .A1(n18242), .A2(n21525), .ZN(n18277) );
  INV_X1 U20276 ( .A(n18277), .ZN(n18251) );
  NAND2_X1 U20277 ( .A1(n21417), .A2(n18277), .ZN(n21399) );
  OAI22_X1 U20278 ( .A1(n21417), .A2(n18275), .B1(n21233), .B2(n21399), .ZN(
        n18243) );
  INV_X1 U20279 ( .A(n18243), .ZN(n21405) );
  OAI21_X1 U20280 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18320), .A(
        n18244), .ZN(n18269) );
  INV_X1 U20281 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18245) );
  INV_X1 U20282 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20846) );
  NAND2_X1 U20283 ( .A1(n18246), .A2(n18280), .ZN(n18266) );
  AOI221_X1 U20284 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n18245), .C2(n20846), .A(
        n18266), .ZN(n18250) );
  INV_X1 U20285 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20868) );
  NOR2_X1 U20286 ( .A1(n20846), .A2(n18265), .ZN(n18248) );
  NOR2_X1 U20287 ( .A1(n11321), .A2(n20543), .ZN(n18309) );
  INV_X1 U20288 ( .A(n18309), .ZN(n18247) );
  OAI21_X1 U20289 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18248), .A(
        n18247), .ZN(n20865) );
  OAI22_X1 U20290 ( .A1(n21620), .A2(n20868), .B1(n20865), .B2(n18310), .ZN(
        n18249) );
  AOI211_X1 U20291 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18269), .A(
        n18250), .B(n18249), .ZN(n18262) );
  NOR2_X1 U20292 ( .A1(n18251), .A2(n21236), .ZN(n18276) );
  OAI22_X1 U20293 ( .A1(n18276), .A2(n21417), .B1(n21236), .B2(n21399), .ZN(
        n21408) );
  AND2_X1 U20294 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18252), .ZN(
        n21403) );
  INV_X1 U20295 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21518) );
  AOI21_X1 U20296 ( .B1(n18253), .B2(n21403), .A(n21518), .ZN(n18254) );
  INV_X1 U20297 ( .A(n18254), .ZN(n18256) );
  OAI21_X1 U20298 ( .B1(n21505), .B2(n18306), .A(n11693), .ZN(n18260) );
  XNOR2_X1 U20299 ( .A(n18260), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21409) );
  AOI22_X1 U20300 ( .A1(n18443), .A2(n21408), .B1(n18444), .B2(n21409), .ZN(
        n18261) );
  OAI211_X1 U20301 ( .C1(n21405), .C2(n18532), .A(n18262), .B(n18261), .ZN(
        P3_U2805) );
  AOI21_X1 U20302 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18264), .A(
        n18263), .ZN(n21532) );
  INV_X1 U20303 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20867) );
  NOR2_X1 U20304 ( .A1(n21620), .A2(n20867), .ZN(n18268) );
  XOR2_X1 U20305 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n18265), .Z(
        n20853) );
  OAI22_X1 U20306 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18266), .B1(
        n18310), .B2(n20853), .ZN(n18267) );
  AOI211_X1 U20307 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18269), .A(
        n18268), .B(n18267), .ZN(n18274) );
  INV_X1 U20308 ( .A(n18278), .ZN(n18271) );
  NOR2_X1 U20309 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21525), .ZN(
        n18270) );
  AOI22_X1 U20310 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18272), .B1(
        n18271), .B2(n18270), .ZN(n18273) );
  OAI211_X1 U20311 ( .C1(n21532), .C2(n18388), .A(n18274), .B(n18273), .ZN(
        P3_U2806) );
  INV_X1 U20312 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21502) );
  INV_X1 U20313 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21415) );
  NOR2_X1 U20314 ( .A1(n21415), .A2(n21417), .ZN(n21425) );
  NAND2_X1 U20315 ( .A1(n21425), .A2(n18275), .ZN(n21447) );
  INV_X1 U20316 ( .A(n21447), .ZN(n18340) );
  INV_X1 U20317 ( .A(n21418), .ZN(n18338) );
  OAI22_X1 U20318 ( .A1(n18340), .A2(n18532), .B1(n18338), .B2(n18389), .ZN(
        n18314) );
  NOR2_X1 U20319 ( .A1(n21502), .A2(n18314), .ZN(n18297) );
  OAI21_X1 U20320 ( .B1(n18443), .B2(n18520), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18294) );
  NAND2_X1 U20321 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18277), .ZN(
        n21414) );
  INV_X1 U20322 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20877) );
  OAI22_X1 U20323 ( .A1(n18528), .A2(n18309), .B1(n18488), .B2(n18298), .ZN(
        n18279) );
  OR2_X1 U20324 ( .A1(n18279), .A2(n18515), .ZN(n18313) );
  AOI21_X1 U20325 ( .B1(n18216), .B2(n20877), .A(n18313), .ZN(n18305) );
  INV_X1 U20326 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20889) );
  NAND3_X1 U20327 ( .A1(n18298), .A2(n20889), .A3(n18280), .ZN(n18301) );
  INV_X1 U20328 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20901) );
  AOI21_X1 U20329 ( .B1(n18305), .B2(n18301), .A(n20901), .ZN(n18283) );
  NOR3_X1 U20330 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18319), .A3(
        n11278), .ZN(n18282) );
  INV_X1 U20331 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21511) );
  NOR2_X1 U20332 ( .A1(n11278), .A2(n20543), .ZN(n18299) );
  NAND2_X1 U20333 ( .A1(n18352), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18321) );
  OAI21_X1 U20334 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18299), .A(
        n18321), .ZN(n20908) );
  OAI22_X1 U20335 ( .A1(n21620), .A2(n21511), .B1(n20908), .B2(n18310), .ZN(
        n18281) );
  NOR4_X1 U20336 ( .A1(n18284), .A2(n18283), .A3(n18282), .A4(n18281), .ZN(
        n18293) );
  NOR2_X1 U20337 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18329), .ZN(
        n18326) );
  AOI21_X1 U20338 ( .B1(n18329), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18326), .ZN(n21509) );
  INV_X1 U20339 ( .A(n21425), .ZN(n18288) );
  AOI21_X1 U20340 ( .B1(n21415), .B2(n21417), .A(n18329), .ZN(n18285) );
  INV_X1 U20341 ( .A(n18285), .ZN(n18286) );
  OAI211_X1 U20342 ( .C1(n18288), .C2(n18287), .A(n18286), .B(n11693), .ZN(
        n18289) );
  INV_X1 U20343 ( .A(n18289), .ZN(n18290) );
  NAND2_X1 U20344 ( .A1(n18290), .A2(n21502), .ZN(n21510) );
  INV_X1 U20345 ( .A(n21510), .ZN(n18327) );
  NOR2_X1 U20346 ( .A1(n18290), .A2(n21502), .ZN(n18328) );
  NOR2_X1 U20347 ( .A1(n18327), .A2(n18328), .ZN(n18296) );
  OAI211_X1 U20348 ( .C1(n21509), .C2(n18291), .A(n18444), .B(n21490), .ZN(
        n18292) );
  OAI211_X1 U20349 ( .C1(n18297), .C2(n18294), .A(n18293), .B(n18292), .ZN(
        P3_U2802) );
  OAI21_X1 U20350 ( .B1(n18329), .B2(n18296), .A(n18295), .ZN(n21437) );
  AOI21_X1 U20351 ( .B1(n21502), .B2(n18337), .A(n18297), .ZN(n18303) );
  NAND2_X1 U20352 ( .A1(n18298), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18308) );
  AOI21_X1 U20353 ( .B1(n20889), .B2(n18308), .A(n18299), .ZN(n18300) );
  INV_X1 U20354 ( .A(n18300), .ZN(n20894) );
  NAND2_X1 U20355 ( .A1(n11176), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21438) );
  OAI211_X1 U20356 ( .C1(n18310), .C2(n20894), .A(n18301), .B(n21438), .ZN(
        n18302) );
  AOI211_X1 U20357 ( .C1(n18444), .C2(n21437), .A(n18303), .B(n18302), .ZN(
        n18304) );
  OAI21_X1 U20358 ( .B1(n18305), .B2(n20889), .A(n18304), .ZN(P3_U2803) );
  OAI221_X1 U20359 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21505), 
        .C1(n21417), .C2(n18306), .A(n11693), .ZN(n18307) );
  XNOR2_X1 U20360 ( .A(n21415), .B(n18307), .ZN(n21424) );
  OAI21_X1 U20361 ( .B1(n11321), .B2(n19252), .A(n20877), .ZN(n18312) );
  OAI21_X1 U20362 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18309), .A(
        n18308), .ZN(n20882) );
  AOI21_X1 U20363 ( .B1(n18310), .B2(n18320), .A(n20882), .ZN(n18311) );
  INV_X1 U20364 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20885) );
  NOR2_X1 U20365 ( .A1(n21620), .A2(n20885), .ZN(n21413) );
  AOI211_X1 U20366 ( .C1(n18313), .C2(n18312), .A(n18311), .B(n21413), .ZN(
        n18316) );
  AOI22_X1 U20367 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18314), .B1(
        n11228), .B2(n21415), .ZN(n18315) );
  OAI211_X1 U20368 ( .C1(n18388), .C2(n21424), .A(n18316), .B(n18315), .ZN(
        P3_U2804) );
  NAND2_X1 U20369 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21476) );
  NAND2_X1 U20370 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21441) );
  XOR2_X1 U20371 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18317), .Z(
        n21483) );
  INV_X1 U20372 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20950) );
  NOR2_X1 U20373 ( .A1(n21620), .A2(n20950), .ZN(n21486) );
  OR2_X1 U20374 ( .A1(n18322), .A2(n18319), .ZN(n18336) );
  XOR2_X1 U20375 ( .A(n18318), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n18324) );
  NOR2_X1 U20376 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18320), .ZN(
        n18348) );
  INV_X1 U20377 ( .A(n18321), .ZN(n18350) );
  NAND2_X1 U20378 ( .A1(n19421), .A2(n18322), .ZN(n18323) );
  OAI211_X1 U20379 ( .C1(n18350), .C2(n18528), .A(n18323), .B(n18527), .ZN(
        n18351) );
  NOR2_X1 U20380 ( .A1(n18348), .A2(n18351), .ZN(n18335) );
  OAI22_X1 U20381 ( .A1(n18336), .A2(n18324), .B1(n18335), .B2(n18318), .ZN(
        n18325) );
  AOI211_X1 U20382 ( .C1(n20932), .C2(n18360), .A(n21486), .B(n18325), .ZN(
        n18333) );
  NAND2_X1 U20383 ( .A1(n18327), .A2(n18326), .ZN(n18344) );
  INV_X1 U20384 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21459) );
  NAND3_X1 U20385 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18329), .A3(
        n18328), .ZN(n21494) );
  INV_X1 U20386 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21468) );
  OAI33_X1 U20387 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n18344), .B1(n21459), .B2(
        n21494), .B3(n21468), .ZN(n18330) );
  XOR2_X1 U20388 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18330), .Z(
        n21484) );
  INV_X1 U20389 ( .A(n21441), .ZN(n21452) );
  NAND2_X1 U20390 ( .A1(n21452), .A2(n18340), .ZN(n21495) );
  XOR2_X1 U20391 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n18331), .Z(
        n21479) );
  AOI22_X1 U20392 ( .A1(n18444), .A2(n21484), .B1(n18520), .B2(n21479), .ZN(
        n18332) );
  OAI211_X1 U20393 ( .C1(n21483), .C2(n18389), .A(n18333), .B(n18332), .ZN(
        P3_U2799) );
  AOI22_X1 U20394 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21494), .B1(
        n18344), .B2(n21459), .ZN(n18334) );
  XNOR2_X1 U20395 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n18334), .ZN(
        n21475) );
  XNOR2_X1 U20396 ( .A(n18349), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n20948) );
  INV_X1 U20397 ( .A(n20948), .ZN(n18343) );
  NAND2_X1 U20398 ( .A1(n11176), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21474) );
  OAI221_X1 U20399 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18336), .C1(
        n11422), .C2(n18335), .A(n21474), .ZN(n18342) );
  NAND2_X1 U20400 ( .A1(n21452), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21464) );
  NOR2_X1 U20401 ( .A1(n21464), .A2(n18337), .ZN(n18341) );
  INV_X1 U20402 ( .A(n21464), .ZN(n18339) );
  NAND2_X1 U20403 ( .A1(n18338), .A2(n18339), .ZN(n21448) );
  AOI21_X1 U20404 ( .B1(n18340), .B2(n18339), .A(n18532), .ZN(n18358) );
  AOI21_X1 U20405 ( .B1(n18443), .B2(n21448), .A(n18358), .ZN(n18346) );
  NAND2_X1 U20406 ( .A1(n18344), .A2(n21494), .ZN(n18345) );
  XNOR2_X1 U20407 ( .A(n18345), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21462) );
  INV_X1 U20408 ( .A(n21495), .ZN(n18357) );
  AOI21_X1 U20409 ( .B1(n18347), .B2(n21459), .A(n18346), .ZN(n18356) );
  NOR2_X1 U20410 ( .A1(n18348), .A2(n18360), .ZN(n18354) );
  OAI21_X1 U20411 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18350), .A(
        n11423), .ZN(n20919) );
  OAI221_X1 U20412 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18352), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n19421), .A(n18351), .ZN(
        n18353) );
  NAND2_X1 U20413 ( .A1(n11176), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21460) );
  OAI211_X1 U20414 ( .C1(n18354), .C2(n20919), .A(n18353), .B(n21460), .ZN(
        n18355) );
  AOI211_X1 U20415 ( .C1(n18358), .C2(n18357), .A(n18356), .B(n18355), .ZN(
        n18359) );
  OAI21_X1 U20416 ( .B1(n21462), .B2(n18388), .A(n18359), .ZN(P3_U2801) );
  NAND2_X1 U20417 ( .A1(n11176), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21574) );
  INV_X1 U20418 ( .A(n21574), .ZN(n18367) );
  INV_X1 U20419 ( .A(n18361), .ZN(n18362) );
  OAI21_X1 U20420 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18363), .A(
        n18362), .ZN(n20759) );
  AOI21_X1 U20421 ( .B1(n11305), .B2(n19421), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18365) );
  OAI22_X1 U20422 ( .A1(n18513), .A2(n20759), .B1(n18365), .B2(n18364), .ZN(
        n18366) );
  AOI211_X1 U20423 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18368), .A(
        n18367), .B(n18366), .ZN(n18373) );
  OAI21_X1 U20424 ( .B1(n18370), .B2(n21576), .A(n18369), .ZN(n21573) );
  NOR2_X1 U20425 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21584), .ZN(
        n21572) );
  AOI22_X1 U20426 ( .A1(n18444), .A2(n21573), .B1(n21572), .B2(n18371), .ZN(
        n18372) );
  NAND2_X1 U20427 ( .A1(n18373), .A2(n18372), .ZN(P3_U2813) );
  AOI22_X1 U20428 ( .A1(n18404), .A2(n21379), .B1(n18376), .B2(n21359), .ZN(
        n18375) );
  OAI21_X1 U20429 ( .B1(n21360), .B2(n18421), .A(n21372), .ZN(n18374) );
  AOI22_X1 U20430 ( .A1(n18377), .A2(n18376), .B1(n18375), .B2(n18374), .ZN(
        n21366) );
  AOI21_X1 U20431 ( .B1(n11408), .B2(n18378), .A(n20724), .ZN(n20714) );
  AOI21_X1 U20432 ( .B1(n18379), .B2(n19421), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18381) );
  NAND2_X1 U20433 ( .A1(n11176), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n21370) );
  OAI21_X1 U20434 ( .B1(n18381), .B2(n18380), .A(n21370), .ZN(n18382) );
  AOI21_X1 U20435 ( .B1(n20714), .B2(n18521), .A(n18382), .ZN(n18387) );
  AOI21_X1 U20436 ( .B1(n21372), .B2(n18384), .A(n18383), .ZN(n21365) );
  AOI21_X1 U20437 ( .B1(n21372), .B2(n18385), .A(n21378), .ZN(n21369) );
  AOI22_X1 U20438 ( .A1(n18443), .A2(n21365), .B1(n18520), .B2(n21369), .ZN(
        n18386) );
  OAI211_X1 U20439 ( .C1(n21366), .C2(n18388), .A(n18387), .B(n18386), .ZN(
        P3_U2816) );
  OAI22_X1 U20440 ( .A1(n18532), .A2(n21331), .B1(n18389), .B2(n21557), .ZN(
        n18390) );
  INV_X1 U20441 ( .A(n18390), .ZN(n18431) );
  NAND2_X1 U20442 ( .A1(n20680), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18411) );
  AOI21_X1 U20443 ( .B1(n11425), .B2(n18411), .A(n18391), .ZN(n20672) );
  NAND2_X1 U20444 ( .A1(n20680), .A2(n19421), .ZN(n18408) );
  NAND2_X1 U20445 ( .A1(n18408), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18392) );
  NOR2_X1 U20446 ( .A1(n18515), .A2(n18437), .ZN(n18467) );
  NAND2_X1 U20447 ( .A1(n11176), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n21338) );
  OAI221_X1 U20448 ( .B1(n18408), .B2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C1(
        n18392), .C2(n18467), .A(n21338), .ZN(n18393) );
  AOI21_X1 U20449 ( .B1(n20672), .B2(n18521), .A(n18393), .ZN(n18400) );
  NAND2_X1 U20450 ( .A1(n18395), .A2(n18394), .ZN(n18396) );
  XNOR2_X1 U20451 ( .A(n18396), .B(n21341), .ZN(n21336) );
  NAND2_X1 U20452 ( .A1(n18397), .A2(n21341), .ZN(n21340) );
  OAI21_X1 U20453 ( .B1(n18397), .B2(n21341), .A(n21340), .ZN(n18398) );
  AOI22_X1 U20454 ( .A1(n18444), .A2(n21336), .B1(n18417), .B2(n18398), .ZN(
        n18399) );
  OAI211_X1 U20455 ( .C1(n18431), .C2(n21341), .A(n18400), .B(n18399), .ZN(
        P3_U2819) );
  NAND2_X1 U20456 ( .A1(n18401), .A2(n21329), .ZN(n18422) );
  AOI21_X1 U20457 ( .B1(n21505), .B2(n21616), .A(n18404), .ZN(n18402) );
  AOI211_X1 U20458 ( .C1(n21616), .C2(n18403), .A(n18402), .B(n21597), .ZN(
        n18406) );
  NOR3_X1 U20459 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18404), .A3(
        n21616), .ZN(n18405) );
  AOI211_X1 U20460 ( .C1(n18407), .C2(n18422), .A(n18406), .B(n18405), .ZN(
        n21598) );
  INV_X1 U20461 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20667) );
  NOR2_X1 U20462 ( .A1(n21620), .A2(n20667), .ZN(n18416) );
  INV_X1 U20463 ( .A(n18408), .ZN(n18414) );
  INV_X1 U20464 ( .A(n18467), .ZN(n18522) );
  NAND3_X1 U20465 ( .A1(n18409), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n19421), .ZN(n18457) );
  NOR2_X1 U20466 ( .A1(n18410), .A2(n18457), .ZN(n18427) );
  AOI21_X1 U20467 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18522), .A(
        n18427), .ZN(n18413) );
  INV_X1 U20468 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20614) );
  NOR3_X1 U20469 ( .A1(n18454), .A2(n20614), .A3(n20543), .ZN(n20622) );
  NAND2_X1 U20470 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20622), .ZN(
        n20639) );
  INV_X1 U20471 ( .A(n20639), .ZN(n18425) );
  NAND2_X1 U20472 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18425), .ZN(
        n20649) );
  INV_X1 U20473 ( .A(n20649), .ZN(n18412) );
  OAI21_X1 U20474 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18412), .A(
        n18411), .ZN(n20652) );
  OAI22_X1 U20475 ( .A1(n18414), .A2(n18413), .B1(n18513), .B2(n20652), .ZN(
        n18415) );
  AOI211_X1 U20476 ( .C1(n21598), .C2(n18444), .A(n18416), .B(n18415), .ZN(
        n18420) );
  NAND3_X1 U20477 ( .A1(n21333), .A2(n18418), .A3(n18417), .ZN(n18419) );
  OAI211_X1 U20478 ( .C1(n18431), .C2(n21597), .A(n18420), .B(n18419), .ZN(
        P3_U2820) );
  NAND2_X1 U20479 ( .A1(n18422), .A2(n18421), .ZN(n18423) );
  XNOR2_X1 U20480 ( .A(n18423), .B(n21616), .ZN(n21622) );
  NAND2_X1 U20481 ( .A1(n11176), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n21624) );
  INV_X1 U20482 ( .A(n21624), .ZN(n18429) );
  INV_X1 U20483 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20630) );
  NOR2_X1 U20484 ( .A1(n20630), .A2(n20614), .ZN(n18435) );
  INV_X1 U20485 ( .A(n18457), .ZN(n18424) );
  AOI22_X1 U20486 ( .A1(n18435), .A2(n18424), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18522), .ZN(n18426) );
  OAI21_X1 U20487 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18425), .A(
        n20649), .ZN(n20645) );
  OAI22_X1 U20488 ( .A1(n18427), .A2(n18426), .B1(n18513), .B2(n20645), .ZN(
        n18428) );
  AOI211_X1 U20489 ( .C1(n18444), .C2(n21622), .A(n18429), .B(n18428), .ZN(
        n18430) );
  OAI221_X1 U20490 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18432), .C1(
        n21616), .C2(n18431), .A(n18430), .ZN(P3_U2821) );
  OAI21_X1 U20491 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18434), .A(
        n18433), .ZN(n21322) );
  OR2_X1 U20492 ( .A1(n18454), .A2(n20614), .ZN(n18436) );
  AOI211_X1 U20493 ( .C1(n20630), .C2(n18436), .A(n18435), .B(n19252), .ZN(
        n18439) );
  OAI21_X1 U20494 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20622), .A(
        n20639), .ZN(n20623) );
  AOI21_X1 U20495 ( .B1(n18437), .B2(n18454), .A(n18515), .ZN(n18456) );
  OAI22_X1 U20496 ( .A1(n18513), .A2(n20623), .B1(n20630), .B2(n18456), .ZN(
        n18438) );
  AOI211_X1 U20497 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n11176), .A(n18439), .B(
        n18438), .ZN(n18447) );
  OAI21_X1 U20498 ( .B1(n18442), .B2(n18441), .A(n18440), .ZN(n21325) );
  INV_X1 U20499 ( .A(n21325), .ZN(n18445) );
  AOI22_X1 U20500 ( .A1(n18445), .A2(n18444), .B1(n18443), .B2(n21325), .ZN(
        n18446) );
  OAI211_X1 U20501 ( .C1(n18532), .C2(n21322), .A(n18447), .B(n18446), .ZN(
        P3_U2822) );
  OAI21_X1 U20502 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18449), .A(
        n18448), .ZN(n21309) );
  AOI21_X1 U20503 ( .B1(n18452), .B2(n18451), .A(n18450), .ZN(n18453) );
  XNOR2_X1 U20504 ( .A(n18453), .B(n21316), .ZN(n21311) );
  NOR2_X1 U20505 ( .A1(n18454), .A2(n20543), .ZN(n20607) );
  INV_X1 U20506 ( .A(n20607), .ZN(n20596) );
  AOI21_X1 U20507 ( .B1(n20614), .B2(n20596), .A(n20622), .ZN(n20609) );
  AOI22_X1 U20508 ( .A1(n11176), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n20609), 
        .B2(n18521), .ZN(n18455) );
  OAI221_X1 U20509 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18457), .C1(
        n20614), .C2(n18456), .A(n18455), .ZN(n18458) );
  AOI21_X1 U20510 ( .B1(n18520), .B2(n21311), .A(n18458), .ZN(n18459) );
  OAI21_X1 U20511 ( .B1(n18531), .B2(n21309), .A(n18459), .ZN(P3_U2823) );
  OAI21_X1 U20512 ( .B1(n18462), .B2(n18461), .A(n18460), .ZN(n21297) );
  NAND2_X1 U20513 ( .A1(n18409), .A2(n19421), .ZN(n18465) );
  OAI21_X1 U20514 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18464), .A(
        n18463), .ZN(n21303) );
  OAI22_X1 U20515 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18465), .B1(
        n21303), .B2(n18532), .ZN(n18466) );
  AOI21_X1 U20516 ( .B1(n11176), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18466), .ZN(
        n18469) );
  AOI21_X1 U20517 ( .B1(n19421), .B2(n18409), .A(n18467), .ZN(n18479) );
  NAND2_X1 U20518 ( .A1(n18409), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18473) );
  AOI21_X1 U20519 ( .B1(n11430), .B2(n18473), .A(n20607), .ZN(n20606) );
  AOI22_X1 U20520 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18479), .B1(
        n20606), .B2(n18521), .ZN(n18468) );
  OAI211_X1 U20521 ( .C1(n18531), .C2(n21297), .A(n18469), .B(n18468), .ZN(
        P3_U2824) );
  OAI21_X1 U20522 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18471), .A(
        n18470), .ZN(n21288) );
  OAI21_X1 U20523 ( .B1(n18515), .B2(n20574), .A(n18472), .ZN(n18478) );
  NOR2_X1 U20524 ( .A1(n20574), .A2(n20543), .ZN(n18490) );
  OAI21_X1 U20525 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18490), .A(
        n18473), .ZN(n20590) );
  OAI21_X1 U20526 ( .B1(n18476), .B2(n18475), .A(n18474), .ZN(n21287) );
  OAI22_X1 U20527 ( .A1(n18513), .A2(n20590), .B1(n18532), .B2(n21287), .ZN(
        n18477) );
  AOI21_X1 U20528 ( .B1(n18479), .B2(n18478), .A(n18477), .ZN(n18480) );
  NAND2_X1 U20529 ( .A1(n11176), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21292) );
  OAI211_X1 U20530 ( .C1(n18531), .C2(n21288), .A(n18480), .B(n21292), .ZN(
        P3_U2825) );
  OAI21_X1 U20531 ( .B1(n18483), .B2(n18482), .A(n18481), .ZN(n21276) );
  NOR2_X1 U20532 ( .A1(n19252), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18487) );
  INV_X1 U20533 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20586) );
  OAI21_X1 U20534 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18485), .A(
        n18484), .ZN(n21275) );
  OAI22_X1 U20535 ( .A1(n21620), .A2(n20586), .B1(n18532), .B2(n21275), .ZN(
        n18486) );
  AOI21_X1 U20536 ( .B1(n18487), .B2(n18489), .A(n18486), .ZN(n18492) );
  OAI21_X1 U20537 ( .B1(n18489), .B2(n18488), .A(n18527), .ZN(n18505) );
  INV_X1 U20538 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20569) );
  NAND2_X1 U20539 ( .A1(n18489), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18493) );
  AOI21_X1 U20540 ( .B1(n20569), .B2(n18493), .A(n18490), .ZN(n20575) );
  AOI22_X1 U20541 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18505), .B1(
        n20575), .B2(n18521), .ZN(n18491) );
  OAI211_X1 U20542 ( .C1(n18531), .C2(n21276), .A(n18492), .B(n18491), .ZN(
        P3_U2826) );
  NOR2_X1 U20543 ( .A1(n20553), .A2(n20543), .ZN(n18494) );
  OAI21_X1 U20544 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18494), .A(
        n18493), .ZN(n20556) );
  OAI211_X1 U20545 ( .C1(n18497), .C2(n18496), .A(n21651), .B(n18495), .ZN(
        n18502) );
  OAI211_X1 U20546 ( .C1(n18500), .C2(n18499), .A(n21491), .B(n18498), .ZN(
        n18501) );
  NAND2_X1 U20547 ( .A1(n18502), .A2(n18501), .ZN(n21269) );
  OAI21_X1 U20548 ( .B1(n18515), .B2(n20553), .A(n18503), .ZN(n18504) );
  AOI22_X1 U20549 ( .A1(n21692), .A2(n21269), .B1(n18505), .B2(n18504), .ZN(
        n18506) );
  NAND2_X1 U20550 ( .A1(n11176), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21272) );
  OAI211_X1 U20551 ( .C1(n18513), .C2(n20556), .A(n18506), .B(n21272), .ZN(
        P3_U2827) );
  OAI21_X1 U20552 ( .B1(n18509), .B2(n18508), .A(n18507), .ZN(n21264) );
  AOI22_X1 U20553 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20543), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20553), .ZN(n20544) );
  OAI21_X1 U20554 ( .B1(n18512), .B2(n18511), .A(n18510), .ZN(n21260) );
  OAI22_X1 U20555 ( .A1(n18513), .A2(n20544), .B1(n18531), .B2(n21260), .ZN(
        n18514) );
  NAND2_X1 U20556 ( .A1(n11176), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21262) );
  OAI211_X1 U20557 ( .C1(n18532), .C2(n21264), .A(n18516), .B(n21262), .ZN(
        P3_U2828) );
  OAI21_X1 U20558 ( .B1(n18518), .B2(n18525), .A(n18517), .ZN(n21249) );
  NAND2_X1 U20559 ( .A1(n21427), .A2(n18526), .ZN(n18519) );
  XNOR2_X1 U20560 ( .A(n18519), .B(n18518), .ZN(n21250) );
  AOI22_X1 U20561 ( .A1(n11176), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18520), 
        .B2(n21250), .ZN(n18524) );
  AOI22_X1 U20562 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18522), .B1(
        n18521), .B2(n20543), .ZN(n18523) );
  OAI211_X1 U20563 ( .C1(n18531), .C2(n21249), .A(n18524), .B(n18523), .ZN(
        P3_U2829) );
  AOI21_X1 U20564 ( .B1(n18526), .B2(n21427), .A(n18525), .ZN(n18533) );
  INV_X1 U20565 ( .A(n18533), .ZN(n21243) );
  NAND3_X1 U20566 ( .A1(n21158), .A2(n18528), .A3(n18527), .ZN(n18529) );
  AOI22_X1 U20567 ( .A1(n11176), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18529), .ZN(n18530) );
  OAI221_X1 U20568 ( .B1(n18533), .B2(n18532), .C1(n21243), .C2(n18531), .A(
        n18530), .ZN(P3_U2830) );
  INV_X1 U20569 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19083) );
  NAND2_X1 U20570 ( .A1(n19085), .A2(n19083), .ZN(n19120) );
  INV_X1 U20571 ( .A(n19120), .ZN(n19114) );
  NAND2_X1 U20572 ( .A1(n21646), .A2(n19083), .ZN(n19150) );
  INV_X1 U20573 ( .A(n19150), .ZN(n19152) );
  AOI21_X1 U20574 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n19152), .ZN(n18534) );
  AOI22_X1 U20575 ( .A1(n19114), .A2(n18538), .B1(n19421), .B2(n18534), .ZN(
        n18535) );
  OAI21_X1 U20576 ( .B1(n18536), .B2(n19083), .A(n18535), .ZN(P3_U2866) );
  NOR3_X1 U20577 ( .A1(n19107), .A2(n19086), .A3(n18537), .ZN(n18540) );
  INV_X1 U20578 ( .A(n18538), .ZN(n18539) );
  AOI22_X1 U20579 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18540), .B1(
        n18539), .B2(n21640), .ZN(P3_U2864) );
  NOR4_X1 U20580 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18544) );
  NOR4_X1 U20581 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18543) );
  NOR4_X1 U20582 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18542) );
  NOR4_X1 U20583 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18541) );
  NAND4_X1 U20584 ( .A1(n18544), .A2(n18543), .A3(n18542), .A4(n18541), .ZN(
        n18550) );
  NOR4_X1 U20585 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18548) );
  AOI211_X1 U20586 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18547) );
  NOR4_X1 U20587 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18546) );
  NOR4_X1 U20588 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18545) );
  NAND4_X1 U20589 ( .A1(n18548), .A2(n18547), .A3(n18546), .A4(n18545), .ZN(
        n18549) );
  NOR2_X1 U20590 ( .A1(n18550), .A2(n18549), .ZN(n18561) );
  INV_X1 U20591 ( .A(n18561), .ZN(n18559) );
  NOR2_X1 U20592 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18552) );
  NAND2_X1 U20593 ( .A1(n18559), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18551) );
  OAI21_X1 U20594 ( .B1(n18559), .B2(n18552), .A(n18551), .ZN(P3_U3293) );
  AOI211_X1 U20595 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18553) );
  AOI21_X1 U20596 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18553), .ZN(n18554) );
  INV_X1 U20597 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18618) );
  AOI22_X1 U20598 ( .A1(n18561), .A2(n18554), .B1(n18618), .B2(n18559), .ZN(
        P3_U3292) );
  INV_X1 U20599 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18556) );
  NOR3_X1 U20600 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18558) );
  NOR2_X1 U20601 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18558), .ZN(n18555) );
  MUX2_X1 U20602 ( .A(n18556), .B(n18555), .S(n18561), .Z(n18557) );
  INV_X1 U20603 ( .A(n18557), .ZN(P3_U2638) );
  INV_X1 U20604 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18606) );
  INV_X1 U20605 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22148) );
  AOI21_X1 U20606 ( .B1(n18606), .B2(n22148), .A(n18558), .ZN(n18560) );
  INV_X1 U20607 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U20608 ( .A1(n18561), .A2(n18560), .B1(n18620), .B2(n18559), .ZN(
        P3_U2639) );
  INV_X1 U20609 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18621) );
  AOI22_X1 U20610 ( .A1(n22153), .A2(n18562), .B1(n18621), .B2(n22205), .ZN(
        P3_U3297) );
  INV_X1 U20611 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18563) );
  AOI22_X1 U20612 ( .A1(n22153), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18563), 
        .B2(n22205), .ZN(P3_U3294) );
  OAI21_X1 U20613 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n18564), .A(n22150), 
        .ZN(n18565) );
  AOI22_X1 U20614 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n22205), .B1(n22196), .B2(
        n18565), .ZN(n18566) );
  INV_X1 U20615 ( .A(n18566), .ZN(P3_U2635) );
  INV_X1 U20616 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21151) );
  INV_X1 U20617 ( .A(n18584), .ZN(n18583) );
  AOI22_X1 U20618 ( .A1(n21627), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18567) );
  OAI21_X1 U20619 ( .B1(n21151), .B2(n18583), .A(n18567), .ZN(P3_U2767) );
  INV_X1 U20620 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21141) );
  AOI22_X1 U20621 ( .A1(n21627), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18568) );
  OAI21_X1 U20622 ( .B1(n21141), .B2(n18583), .A(n18568), .ZN(P3_U2766) );
  INV_X1 U20623 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20503) );
  AOI22_X1 U20624 ( .A1(n21627), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18569) );
  OAI21_X1 U20625 ( .B1(n20503), .B2(n18583), .A(n18569), .ZN(P3_U2765) );
  INV_X1 U20626 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U20627 ( .A1(n21627), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18570) );
  OAI21_X1 U20628 ( .B1(n20967), .B2(n18583), .A(n18570), .ZN(P3_U2764) );
  INV_X1 U20629 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21006) );
  AOI22_X1 U20630 ( .A1(n21627), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18571) );
  OAI21_X1 U20631 ( .B1(n21006), .B2(n18583), .A(n18571), .ZN(P3_U2763) );
  INV_X1 U20632 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20968) );
  AOI22_X1 U20633 ( .A1(n21627), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18572) );
  OAI21_X1 U20634 ( .B1(n20968), .B2(n18583), .A(n18572), .ZN(P3_U2762) );
  INV_X1 U20635 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20509) );
  AOI22_X1 U20636 ( .A1(n21627), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18573) );
  OAI21_X1 U20637 ( .B1(n20509), .B2(n18583), .A(n18573), .ZN(P3_U2761) );
  INV_X1 U20638 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20511) );
  AOI22_X1 U20639 ( .A1(n21627), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18574) );
  OAI21_X1 U20640 ( .B1(n20511), .B2(n18583), .A(n18574), .ZN(P3_U2760) );
  INV_X1 U20641 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21133) );
  AOI22_X1 U20642 ( .A1(n21627), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18575) );
  OAI21_X1 U20643 ( .B1(n21133), .B2(n18583), .A(n18575), .ZN(P3_U2759) );
  INV_X1 U20644 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20973) );
  AOI22_X1 U20645 ( .A1(n18593), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18576) );
  OAI21_X1 U20646 ( .B1(n20973), .B2(n18583), .A(n18576), .ZN(P3_U2758) );
  INV_X1 U20647 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20515) );
  AOI22_X1 U20648 ( .A1(n18593), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18577) );
  OAI21_X1 U20649 ( .B1(n20515), .B2(n18583), .A(n18577), .ZN(P3_U2757) );
  INV_X1 U20650 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U20651 ( .A1(n18593), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18578) );
  OAI21_X1 U20652 ( .B1(n20985), .B2(n18583), .A(n18578), .ZN(P3_U2756) );
  INV_X1 U20653 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20518) );
  AOI22_X1 U20654 ( .A1(n18593), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18579) );
  OAI21_X1 U20655 ( .B1(n20518), .B2(n18583), .A(n18579), .ZN(P3_U2755) );
  INV_X1 U20656 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20520) );
  AOI22_X1 U20657 ( .A1(n18593), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18580) );
  OAI21_X1 U20658 ( .B1(n20520), .B2(n18583), .A(n18580), .ZN(P3_U2754) );
  INV_X1 U20659 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21123) );
  AOI22_X1 U20660 ( .A1(n18593), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18581) );
  OAI21_X1 U20661 ( .B1(n21123), .B2(n18583), .A(n18581), .ZN(P3_U2753) );
  INV_X1 U20662 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21130) );
  AOI22_X1 U20663 ( .A1(n18593), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18582) );
  OAI21_X1 U20664 ( .B1(n21130), .B2(n18583), .A(n18582), .ZN(P3_U2752) );
  INV_X1 U20665 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20474) );
  NAND2_X1 U20666 ( .A1(n18584), .A2(n11507), .ZN(n18603) );
  AOI22_X1 U20667 ( .A1(n18593), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18585) );
  OAI21_X1 U20668 ( .B1(n20474), .B2(n18603), .A(n18585), .ZN(P3_U2751) );
  INV_X1 U20669 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20476) );
  AOI22_X1 U20670 ( .A1(n18593), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18586) );
  OAI21_X1 U20671 ( .B1(n20476), .B2(n18603), .A(n18586), .ZN(P3_U2750) );
  INV_X1 U20672 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20478) );
  AOI22_X1 U20673 ( .A1(n18593), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18587) );
  OAI21_X1 U20674 ( .B1(n20478), .B2(n18603), .A(n18587), .ZN(P3_U2749) );
  INV_X1 U20675 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21046) );
  AOI22_X1 U20676 ( .A1(n21627), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18588) );
  OAI21_X1 U20677 ( .B1(n21046), .B2(n18603), .A(n18588), .ZN(P3_U2748) );
  INV_X1 U20678 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20482) );
  AOI22_X1 U20679 ( .A1(n21627), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18589) );
  OAI21_X1 U20680 ( .B1(n20482), .B2(n18603), .A(n18589), .ZN(P3_U2747) );
  INV_X1 U20681 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21032) );
  AOI22_X1 U20682 ( .A1(n21627), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18590) );
  OAI21_X1 U20683 ( .B1(n21032), .B2(n18603), .A(n18590), .ZN(P3_U2746) );
  INV_X1 U20684 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20485) );
  AOI22_X1 U20685 ( .A1(n21627), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18591) );
  OAI21_X1 U20686 ( .B1(n20485), .B2(n18603), .A(n18591), .ZN(P3_U2745) );
  INV_X1 U20687 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20487) );
  AOI22_X1 U20688 ( .A1(n21627), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18592) );
  OAI21_X1 U20689 ( .B1(n20487), .B2(n18603), .A(n18592), .ZN(P3_U2744) );
  INV_X1 U20690 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20489) );
  AOI22_X1 U20691 ( .A1(n18593), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18594) );
  OAI21_X1 U20692 ( .B1(n20489), .B2(n18603), .A(n18594), .ZN(P3_U2743) );
  INV_X1 U20693 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20491) );
  AOI22_X1 U20694 ( .A1(n21627), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18595) );
  OAI21_X1 U20695 ( .B1(n20491), .B2(n18603), .A(n18595), .ZN(P3_U2742) );
  INV_X1 U20696 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21070) );
  AOI22_X1 U20697 ( .A1(n21627), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18596) );
  OAI21_X1 U20698 ( .B1(n21070), .B2(n18603), .A(n18596), .ZN(P3_U2741) );
  INV_X1 U20699 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20494) );
  AOI22_X1 U20700 ( .A1(n21627), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18597), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18598) );
  OAI21_X1 U20701 ( .B1(n20494), .B2(n18603), .A(n18598), .ZN(P3_U2740) );
  INV_X1 U20702 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U20703 ( .A1(n21627), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18599) );
  OAI21_X1 U20704 ( .B1(n21088), .B2(n18603), .A(n18599), .ZN(P3_U2739) );
  INV_X1 U20705 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20497) );
  AOI22_X1 U20706 ( .A1(n21627), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18600) );
  OAI21_X1 U20707 ( .B1(n20497), .B2(n18603), .A(n18600), .ZN(P3_U2738) );
  INV_X1 U20708 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20499) );
  AOI22_X1 U20709 ( .A1(n21627), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18601), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18602) );
  OAI21_X1 U20710 ( .B1(n20499), .B2(n18603), .A(n18602), .ZN(P3_U2737) );
  INV_X1 U20711 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n18605) );
  OAI21_X1 U20712 ( .B1(n22153), .B2(n18605), .A(n18604), .ZN(P3_U2633) );
  AND2_X1 U20713 ( .A1(n22153), .A2(n22194), .ZN(n18611) );
  INV_X1 U20714 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20542) );
  INV_X1 U20715 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20121) );
  OAI222_X1 U20716 ( .A1(n18615), .A2(n20542), .B1(n20121), .B2(n22153), .C1(
        n18606), .C2(n18616), .ZN(P3_U3032) );
  INV_X1 U20717 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20559) );
  INV_X1 U20718 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20123) );
  OAI222_X1 U20719 ( .A1(n18615), .A2(n20559), .B1(n20123), .B2(n22153), .C1(
        n20542), .C2(n18616), .ZN(P3_U3033) );
  INV_X1 U20720 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n20125) );
  OAI222_X1 U20721 ( .A1(n18615), .A2(n20586), .B1(n20125), .B2(n22153), .C1(
        n20559), .C2(n18616), .ZN(P3_U3034) );
  AOI22_X1 U20722 ( .A1(n18611), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n22205), .ZN(n18607) );
  OAI21_X1 U20723 ( .B1(n18616), .B2(n20586), .A(n18607), .ZN(P3_U3035) );
  INV_X1 U20724 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20613) );
  AOI22_X1 U20725 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18613), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n22205), .ZN(n18608) );
  OAI21_X1 U20726 ( .B1(n20613), .B2(n18615), .A(n18608), .ZN(P3_U3036) );
  AOI22_X1 U20727 ( .A1(n18611), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n22205), .ZN(n18609) );
  OAI21_X1 U20728 ( .B1(n18616), .B2(n20613), .A(n18609), .ZN(P3_U3037) );
  INV_X1 U20729 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20627) );
  AOI22_X1 U20730 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18613), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n22205), .ZN(n18610) );
  OAI21_X1 U20731 ( .B1(n20627), .B2(n18615), .A(n18610), .ZN(P3_U3038) );
  INV_X1 U20732 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20640) );
  INV_X1 U20733 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20135) );
  OAI222_X1 U20734 ( .A1(n18615), .A2(n20640), .B1(n20135), .B2(n22153), .C1(
        n20627), .C2(n18616), .ZN(P3_U3039) );
  INV_X1 U20735 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20137) );
  OAI222_X1 U20736 ( .A1(n18615), .A2(n20667), .B1(n20137), .B2(n22153), .C1(
        n20640), .C2(n18616), .ZN(P3_U3040) );
  INV_X1 U20737 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20139) );
  INV_X1 U20738 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20666) );
  OAI222_X1 U20739 ( .A1(n20667), .A2(n18616), .B1(n20139), .B2(n22153), .C1(
        n20666), .C2(n18615), .ZN(P3_U3041) );
  INV_X1 U20740 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20691) );
  INV_X1 U20741 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20141) );
  OAI222_X1 U20742 ( .A1(n18615), .A2(n20691), .B1(n20141), .B2(n22153), .C1(
        n20666), .C2(n18616), .ZN(P3_U3042) );
  INV_X1 U20743 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20143) );
  OAI222_X1 U20744 ( .A1(n18615), .A2(n20712), .B1(n20143), .B2(n22153), .C1(
        n20691), .C2(n18616), .ZN(P3_U3043) );
  AOI22_X1 U20745 ( .A1(n18611), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n22205), .ZN(n18612) );
  OAI21_X1 U20746 ( .B1(n18616), .B2(n20712), .A(n18612), .ZN(P3_U3044) );
  INV_X1 U20747 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20750) );
  AOI22_X1 U20748 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18613), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n22205), .ZN(n18614) );
  OAI21_X1 U20749 ( .B1(n20750), .B2(n18615), .A(n18614), .ZN(P3_U3045) );
  INV_X1 U20750 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20149) );
  OAI222_X1 U20751 ( .A1(n18615), .A2(n21588), .B1(n20149), .B2(n22153), .C1(
        n20750), .C2(n18616), .ZN(P3_U3046) );
  INV_X1 U20752 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20763) );
  INV_X1 U20753 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20151) );
  OAI222_X1 U20754 ( .A1(n18615), .A2(n20763), .B1(n20151), .B2(n22153), .C1(
        n21588), .C2(n18616), .ZN(P3_U3047) );
  INV_X1 U20755 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20153) );
  OAI222_X1 U20756 ( .A1(n20763), .A2(n18616), .B1(n20153), .B2(n22153), .C1(
        n20775), .C2(n18615), .ZN(P3_U3048) );
  INV_X1 U20757 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20155) );
  INV_X1 U20758 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U20759 ( .A1(n20775), .A2(n18616), .B1(n20155), .B2(n22153), .C1(
        n20787), .C2(n18615), .ZN(P3_U3049) );
  INV_X1 U20760 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20802) );
  INV_X1 U20761 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20157) );
  OAI222_X1 U20762 ( .A1(n18615), .A2(n20802), .B1(n20157), .B2(n22153), .C1(
        n20787), .C2(n18616), .ZN(P3_U3050) );
  INV_X1 U20763 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20159) );
  OAI222_X1 U20764 ( .A1(n18615), .A2(n20814), .B1(n20159), .B2(n22153), .C1(
        n20802), .C2(n18616), .ZN(P3_U3051) );
  INV_X1 U20765 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20831) );
  INV_X1 U20766 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20161) );
  OAI222_X1 U20767 ( .A1(n18615), .A2(n20831), .B1(n20161), .B2(n22153), .C1(
        n20814), .C2(n18616), .ZN(P3_U3052) );
  INV_X1 U20768 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20843) );
  INV_X1 U20769 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20163) );
  OAI222_X1 U20770 ( .A1(n18615), .A2(n20843), .B1(n20163), .B2(n22153), .C1(
        n20831), .C2(n18616), .ZN(P3_U3053) );
  INV_X1 U20771 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20165) );
  OAI222_X1 U20772 ( .A1(n18615), .A2(n20867), .B1(n20165), .B2(n22153), .C1(
        n20843), .C2(n18616), .ZN(P3_U3054) );
  INV_X1 U20773 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20167) );
  OAI222_X1 U20774 ( .A1(n18615), .A2(n20868), .B1(n20167), .B2(n22153), .C1(
        n20867), .C2(n18616), .ZN(P3_U3055) );
  INV_X1 U20775 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20170) );
  OAI222_X1 U20776 ( .A1(n18615), .A2(n20885), .B1(n20170), .B2(n22153), .C1(
        n20868), .C2(n18616), .ZN(P3_U3056) );
  INV_X1 U20777 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20898) );
  INV_X1 U20778 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20172) );
  OAI222_X1 U20779 ( .A1(n18615), .A2(n20898), .B1(n20172), .B2(n22153), .C1(
        n20885), .C2(n18616), .ZN(P3_U3057) );
  INV_X1 U20780 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20174) );
  OAI222_X1 U20781 ( .A1(n18615), .A2(n21511), .B1(n20174), .B2(n22153), .C1(
        n20898), .C2(n18616), .ZN(P3_U3058) );
  INV_X1 U20782 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20176) );
  INV_X1 U20783 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20920) );
  OAI222_X1 U20784 ( .A1(n21511), .A2(n18616), .B1(n20176), .B2(n22153), .C1(
        n20920), .C2(n18615), .ZN(P3_U3059) );
  INV_X1 U20785 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20937) );
  INV_X1 U20786 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20178) );
  OAI222_X1 U20787 ( .A1(n18615), .A2(n20937), .B1(n20178), .B2(n22153), .C1(
        n20920), .C2(n18616), .ZN(P3_U3060) );
  INV_X1 U20788 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20181) );
  OAI222_X1 U20789 ( .A1(n20937), .A2(n18616), .B1(n20181), .B2(n22153), .C1(
        n20950), .C2(n18615), .ZN(P3_U3061) );
  MUX2_X1 U20790 ( .A(P3_BE_N_REG_0__SCAN_IN), .B(P3_BYTEENABLE_REG_0__SCAN_IN), .S(n22153), .Z(P3_U3277) );
  MUX2_X1 U20791 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n22153), .Z(P3_U3276) );
  INV_X1 U20792 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18617) );
  AOI22_X1 U20793 ( .A1(n22153), .A2(n18618), .B1(n18617), .B2(n22205), .ZN(
        P3_U3275) );
  INV_X1 U20794 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18619) );
  AOI22_X1 U20795 ( .A1(n22153), .A2(n18620), .B1(n18619), .B2(n22205), .ZN(
        P3_U3274) );
  NOR4_X1 U20796 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18623)
         );
  NOR4_X1 U20797 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18621), .ZN(n18622) );
  NAND3_X1 U20798 ( .A1(n18623), .A2(n18622), .A3(U215), .ZN(U213) );
  NOR2_X1 U20799 ( .A1(n19035), .A2(n19594), .ZN(n18627) );
  OAI21_X1 U20800 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n12069), .A(n22182), 
        .ZN(n18625) );
  NAND3_X1 U20801 ( .A1(n18625), .A2(n18624), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18626) );
  OAI21_X1 U20802 ( .B1(n18627), .B2(n19049), .A(n18626), .ZN(n18633) );
  NAND4_X1 U20803 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n11739), .A4(n22174), .ZN(n18629) );
  OAI211_X1 U20804 ( .C1(n18631), .C2(n18630), .A(n18629), .B(n18628), .ZN(
        n18632) );
  MUX2_X1 U20805 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n18633), .S(n18632), 
        .Z(P2_U3610) );
  OAI22_X1 U20806 ( .A1(n18922), .A2(n18635), .B1(n18969), .B2(n18634), .ZN(
        n18636) );
  INV_X1 U20807 ( .A(n18636), .ZN(n18641) );
  NAND2_X1 U20808 ( .A1(n18957), .A2(n18637), .ZN(n18640) );
  NAND2_X1 U20809 ( .A1(n18951), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18639) );
  NAND2_X1 U20810 ( .A1(n18954), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18638) );
  AND4_X1 U20811 ( .A1(n18641), .A2(n18640), .A3(n18639), .A4(n18638), .ZN(
        n18645) );
  AOI22_X1 U20812 ( .A1(n18980), .A2(n18642), .B1(n19550), .B2(n18653), .ZN(
        n18644) );
  NAND2_X1 U20813 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18955), .ZN(
        n18643) );
  NAND3_X1 U20814 ( .A1(n18645), .A2(n18644), .A3(n18643), .ZN(P2_U2855) );
  AOI22_X1 U20815 ( .A1(n18977), .A2(n18646), .B1(n18954), .B2(
        P2_REIP_REG_1__SCAN_IN), .ZN(n18652) );
  INV_X1 U20816 ( .A(n18969), .ZN(n18952) );
  AOI22_X1 U20817 ( .A1(n18952), .A2(n18647), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18955), .ZN(n18651) );
  NAND2_X1 U20818 ( .A1(n18648), .A2(n18957), .ZN(n18650) );
  NAND2_X1 U20819 ( .A1(n18951), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n18649) );
  AND4_X1 U20820 ( .A1(n18652), .A2(n18651), .A3(n18650), .A4(n18649), .ZN(
        n18655) );
  NOR2_X1 U20821 ( .A1(n19039), .A2(n11164), .ZN(n18751) );
  AOI22_X1 U20822 ( .A1(n18751), .A2(n14249), .B1(n19551), .B2(n18653), .ZN(
        n18654) );
  OAI211_X1 U20823 ( .C1(n19039), .C2(n18656), .A(n18655), .B(n18654), .ZN(
        P2_U2854) );
  INV_X1 U20824 ( .A(n18957), .ZN(n18983) );
  NAND2_X1 U20825 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18955), .ZN(
        n18657) );
  OAI211_X1 U20826 ( .C1(n18969), .C2(n18658), .A(n18830), .B(n18657), .ZN(
        n18661) );
  NOR2_X1 U20827 ( .A1(n18922), .A2(n18659), .ZN(n18660) );
  NOR2_X1 U20828 ( .A1(n18661), .A2(n18660), .ZN(n18665) );
  OAI22_X1 U20829 ( .A1(n18884), .A2(n18662), .B1(n11952), .B2(n18968), .ZN(
        n18663) );
  INV_X1 U20830 ( .A(n18663), .ZN(n18664) );
  OAI211_X1 U20831 ( .C1(n19775), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        n18667) );
  INV_X1 U20832 ( .A(n18667), .ZN(n18674) );
  INV_X1 U20833 ( .A(n18668), .ZN(n18672) );
  NOR2_X1 U20834 ( .A1(n18809), .A2(n18669), .ZN(n18671) );
  AOI21_X1 U20835 ( .B1(n18672), .B2(n18671), .A(n19039), .ZN(n18670) );
  OAI21_X1 U20836 ( .B1(n18672), .B2(n18671), .A(n18670), .ZN(n18673) );
  OAI211_X1 U20837 ( .C1(n18675), .C2(n18983), .A(n18674), .B(n18673), .ZN(
        P2_U2851) );
  OAI21_X1 U20838 ( .B1(n18884), .B2(n12435), .A(n18830), .ZN(n18679) );
  OAI22_X1 U20839 ( .A1(n18969), .A2(n18677), .B1(n18676), .B2(n18973), .ZN(
        n18678) );
  AOI211_X1 U20840 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18954), .A(n18679), .B(
        n18678), .ZN(n18686) );
  NAND2_X1 U20841 ( .A1(n11165), .A2(n18680), .ZN(n18681) );
  XNOR2_X1 U20842 ( .A(n18682), .B(n18681), .ZN(n18684) );
  AOI22_X1 U20843 ( .A1(n18980), .A2(n18684), .B1(n18957), .B2(n18683), .ZN(
        n18685) );
  OAI211_X1 U20844 ( .C1(n18922), .C2(n19780), .A(n18686), .B(n18685), .ZN(
        P2_U2850) );
  OAI21_X1 U20845 ( .B1(n18884), .B2(n18687), .A(n18830), .ZN(n18690) );
  OAI22_X1 U20846 ( .A1(n18968), .A2(n11961), .B1(n18688), .B2(n18969), .ZN(
        n18689) );
  AOI211_X1 U20847 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18955), .A(
        n18690), .B(n18689), .ZN(n18697) );
  NOR2_X1 U20848 ( .A1(n18809), .A2(n18691), .ZN(n18693) );
  XNOR2_X1 U20849 ( .A(n18693), .B(n18692), .ZN(n18695) );
  AOI22_X1 U20850 ( .A1(n18980), .A2(n18695), .B1(n18977), .B2(n18694), .ZN(
        n18696) );
  OAI211_X1 U20851 ( .C1(n18983), .C2(n18698), .A(n18697), .B(n18696), .ZN(
        P2_U2849) );
  NAND2_X1 U20852 ( .A1(n11165), .A2(n18699), .ZN(n18701) );
  XOR2_X1 U20853 ( .A(n18701), .B(n18700), .Z(n18709) );
  AOI22_X1 U20854 ( .A1(n18952), .A2(n18702), .B1(n18954), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n18703) );
  OAI211_X1 U20855 ( .C1(n18884), .C2(n12436), .A(n18703), .B(n18830), .ZN(
        n18707) );
  OAI22_X1 U20856 ( .A1(n18922), .A2(n18705), .B1(n18983), .B2(n18704), .ZN(
        n18706) );
  AOI211_X1 U20857 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18955), .A(
        n18707), .B(n18706), .ZN(n18708) );
  OAI21_X1 U20858 ( .B1(n18709), .B2(n19039), .A(n18708), .ZN(P2_U2848) );
  INV_X1 U20859 ( .A(n18710), .ZN(n18712) );
  AOI22_X1 U20860 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18954), .ZN(n18711) );
  OAI21_X1 U20861 ( .B1(n18712), .B2(n18969), .A(n18711), .ZN(n18713) );
  AOI211_X1 U20862 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18713), .ZN(n18719) );
  NOR2_X1 U20863 ( .A1(n18809), .A2(n18714), .ZN(n18716) );
  XNOR2_X1 U20864 ( .A(n18716), .B(n18715), .ZN(n18717) );
  AOI22_X1 U20865 ( .A1(n18980), .A2(n18717), .B1(n18977), .B2(n19002), .ZN(
        n18718) );
  OAI211_X1 U20866 ( .C1(n18983), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P2_U2847) );
  NAND2_X1 U20867 ( .A1(n11164), .A2(n18721), .ZN(n18723) );
  XOR2_X1 U20868 ( .A(n18723), .B(n18722), .Z(n18732) );
  AOI22_X1 U20869 ( .A1(n18724), .A2(n18952), .B1(n18954), .B2(
        P2_REIP_REG_9__SCAN_IN), .ZN(n18725) );
  OAI211_X1 U20870 ( .C1(n18884), .C2(n18726), .A(n18725), .B(n18830), .ZN(
        n18730) );
  OAI22_X1 U20871 ( .A1(n18922), .A2(n18728), .B1(n18983), .B2(n18727), .ZN(
        n18729) );
  AOI211_X1 U20872 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18955), .A(
        n18730), .B(n18729), .ZN(n18731) );
  OAI21_X1 U20873 ( .B1(n18732), .B2(n19039), .A(n18731), .ZN(P2_U2846) );
  AOI22_X1 U20874 ( .A1(n18733), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18734) );
  OAI21_X1 U20875 ( .B1(n18735), .B2(n18968), .A(n18734), .ZN(n18736) );
  AOI211_X1 U20876 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18736), .ZN(n18743) );
  NOR2_X1 U20877 ( .A1(n18809), .A2(n18737), .ZN(n18739) );
  XNOR2_X1 U20878 ( .A(n18739), .B(n18738), .ZN(n18740) );
  AOI22_X1 U20879 ( .A1(n18741), .A2(n18977), .B1(n18980), .B2(n18740), .ZN(
        n18742) );
  OAI211_X1 U20880 ( .C1(n18744), .C2(n18983), .A(n18743), .B(n18742), .ZN(
        P2_U2845) );
  AOI22_X1 U20881 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18954), .ZN(n18745) );
  OAI211_X1 U20882 ( .C1(n18746), .C2(n18922), .A(n18745), .B(n18830), .ZN(
        n18750) );
  OAI22_X1 U20883 ( .A1(n18748), .A2(n18969), .B1(n18747), .B2(n18973), .ZN(
        n18749) );
  AOI211_X1 U20884 ( .C1(n18753), .C2(n18751), .A(n18750), .B(n18749), .ZN(
        n18757) );
  OR2_X1 U20885 ( .A1(n18809), .A2(n18752), .ZN(n18759) );
  AOI211_X1 U20886 ( .C1(n18754), .C2(n18753), .A(n19039), .B(n18759), .ZN(
        n18755) );
  INV_X1 U20887 ( .A(n18755), .ZN(n18756) );
  OAI211_X1 U20888 ( .C1(n18983), .C2(n18758), .A(n18757), .B(n18756), .ZN(
        P2_U2844) );
  XNOR2_X1 U20889 ( .A(n18760), .B(n18759), .ZN(n18768) );
  AOI22_X1 U20890 ( .A1(n18761), .A2(n18952), .B1(n18954), .B2(
        P2_REIP_REG_12__SCAN_IN), .ZN(n18762) );
  OAI211_X1 U20891 ( .C1(n18884), .C2(n11983), .A(n18762), .B(n18830), .ZN(
        n18766) );
  OAI22_X1 U20892 ( .A1(n18764), .A2(n18983), .B1(n18763), .B2(n18922), .ZN(
        n18765) );
  AOI211_X1 U20893 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18955), .A(
        n18766), .B(n18765), .ZN(n18767) );
  OAI21_X1 U20894 ( .B1(n19039), .B2(n18768), .A(n18767), .ZN(P2_U2843) );
  OAI21_X1 U20895 ( .B1(n18884), .B2(n18769), .A(n18830), .ZN(n18772) );
  OAI22_X1 U20896 ( .A1(n18770), .A2(n18969), .B1(n11694), .B2(n18973), .ZN(
        n18771) );
  AOI211_X1 U20897 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18954), .A(n18772), 
        .B(n18771), .ZN(n18779) );
  NAND2_X1 U20898 ( .A1(n11164), .A2(n18773), .ZN(n18774) );
  XNOR2_X1 U20899 ( .A(n18775), .B(n18774), .ZN(n18776) );
  AOI22_X1 U20900 ( .A1(n18777), .A2(n18957), .B1(n18980), .B2(n18776), .ZN(
        n18778) );
  OAI211_X1 U20901 ( .C1(n18780), .C2(n18922), .A(n18779), .B(n18778), .ZN(
        P2_U2842) );
  NOR2_X1 U20902 ( .A1(n18809), .A2(n18781), .ZN(n18783) );
  XOR2_X1 U20903 ( .A(n18783), .B(n18782), .Z(n18791) );
  AOI22_X1 U20904 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18954), .ZN(n18784) );
  OAI21_X1 U20905 ( .B1(n18785), .B2(n18969), .A(n18784), .ZN(n18786) );
  AOI211_X1 U20906 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18786), .ZN(n18790) );
  AOI22_X1 U20907 ( .A1(n18788), .A2(n18957), .B1(n18787), .B2(n18977), .ZN(
        n18789) );
  OAI211_X1 U20908 ( .C1(n19039), .C2(n18791), .A(n18790), .B(n18789), .ZN(
        P2_U2841) );
  OAI21_X1 U20909 ( .B1(n18884), .B2(n12440), .A(n18830), .ZN(n18796) );
  INV_X1 U20910 ( .A(n18792), .ZN(n18794) );
  OAI22_X1 U20911 ( .A1(n18794), .A2(n18969), .B1(n18793), .B2(n18973), .ZN(
        n18795) );
  AOI211_X1 U20912 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18954), .A(n18796), 
        .B(n18795), .ZN(n18803) );
  NAND2_X1 U20913 ( .A1(n11165), .A2(n18797), .ZN(n18798) );
  XNOR2_X1 U20914 ( .A(n18799), .B(n18798), .ZN(n18800) );
  AOI22_X1 U20915 ( .A1(n18801), .A2(n18957), .B1(n18980), .B2(n18800), .ZN(
        n18802) );
  OAI211_X1 U20916 ( .C1(n18804), .C2(n18922), .A(n18803), .B(n18802), .ZN(
        P2_U2840) );
  INV_X1 U20917 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18818) );
  OAI22_X1 U20918 ( .A1(n18806), .A2(n18969), .B1(n18805), .B2(n18968), .ZN(
        n18807) );
  AOI211_X1 U20919 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18807), .ZN(n18817) );
  NOR2_X1 U20920 ( .A1(n18809), .A2(n18808), .ZN(n18810) );
  XNOR2_X1 U20921 ( .A(n18811), .B(n18810), .ZN(n18815) );
  OAI22_X1 U20922 ( .A1(n18813), .A2(n18983), .B1(n18812), .B2(n18922), .ZN(
        n18814) );
  AOI21_X1 U20923 ( .B1(n18815), .B2(n18980), .A(n18814), .ZN(n18816) );
  OAI211_X1 U20924 ( .C1(n18818), .C2(n18973), .A(n18817), .B(n18816), .ZN(
        P2_U2839) );
  NAND2_X1 U20925 ( .A1(n11165), .A2(n18819), .ZN(n18820) );
  XOR2_X1 U20926 ( .A(n18821), .B(n18820), .Z(n18829) );
  AOI22_X1 U20927 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18954), .ZN(n18822) );
  OAI21_X1 U20928 ( .B1(n18823), .B2(n18969), .A(n18822), .ZN(n18824) );
  AOI211_X1 U20929 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18824), .ZN(n18828) );
  AOI22_X1 U20930 ( .A1(n18826), .A2(n18957), .B1(n18825), .B2(n18977), .ZN(
        n18827) );
  OAI211_X1 U20931 ( .C1(n19039), .C2(n18829), .A(n18828), .B(n18827), .ZN(
        P2_U2838) );
  INV_X1 U20932 ( .A(n19913), .ZN(n18837) );
  AOI22_X1 U20933 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18954), .ZN(n18831) );
  OAI211_X1 U20934 ( .C1(n18884), .C2(n18832), .A(n18831), .B(n18830), .ZN(
        n18833) );
  AOI21_X1 U20935 ( .B1(n18834), .B2(n18952), .A(n18833), .ZN(n18835) );
  INV_X1 U20936 ( .A(n18835), .ZN(n18836) );
  AOI21_X1 U20937 ( .B1(n18837), .B2(n18977), .A(n18836), .ZN(n18842) );
  OAI211_X1 U20938 ( .C1(n18840), .C2(n18839), .A(n18980), .B(n18838), .ZN(
        n18841) );
  OAI211_X1 U20939 ( .C1(n18983), .C2(n18843), .A(n18842), .B(n18841), .ZN(
        P2_U2837) );
  AOI22_X1 U20940 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18954), .ZN(n18844) );
  OAI21_X1 U20941 ( .B1(n18845), .B2(n18969), .A(n18844), .ZN(n18846) );
  AOI211_X1 U20942 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18951), .A(n11167), .B(
        n18846), .ZN(n18853) );
  AOI22_X1 U20943 ( .A1(n18848), .A2(n18957), .B1(n18847), .B2(n18977), .ZN(
        n18852) );
  NAND3_X1 U20944 ( .A1(n18853), .A2(n18852), .A3(n18851), .ZN(P2_U2836) );
  AOI22_X1 U20945 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18954), .ZN(n18862) );
  AOI22_X1 U20946 ( .A1(n18854), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18861) );
  AOI22_X1 U20947 ( .A1(n18855), .A2(n18957), .B1(n19823), .B2(n18977), .ZN(
        n18860) );
  OAI211_X1 U20948 ( .C1(n18858), .C2(n18857), .A(n18980), .B(n18856), .ZN(
        n18859) );
  NAND4_X1 U20949 ( .A1(n18862), .A2(n18861), .A3(n18860), .A4(n18859), .ZN(
        P2_U2835) );
  AOI22_X1 U20950 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18954), .ZN(n18872) );
  AOI22_X1 U20951 ( .A1(n18863), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18871) );
  AOI22_X1 U20952 ( .A1(n18865), .A2(n18957), .B1(n18864), .B2(n18977), .ZN(
        n18870) );
  OAI211_X1 U20953 ( .C1(n18868), .C2(n18867), .A(n18980), .B(n18866), .ZN(
        n18869) );
  NAND4_X1 U20954 ( .A1(n18872), .A2(n18871), .A3(n18870), .A4(n18869), .ZN(
        P2_U2834) );
  AOI22_X1 U20955 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18954), .ZN(n18881) );
  AOI22_X1 U20956 ( .A1(n18873), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U20957 ( .A1(n18874), .A2(n18957), .B1(n19728), .B2(n18977), .ZN(
        n18879) );
  OAI211_X1 U20958 ( .C1(n18877), .C2(n18876), .A(n18980), .B(n18875), .ZN(
        n18878) );
  NAND4_X1 U20959 ( .A1(n18881), .A2(n18880), .A3(n18879), .A4(n18878), .ZN(
        P2_U2833) );
  INV_X1 U20960 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n18883) );
  OAI22_X1 U20961 ( .A1(n18884), .A2(n18883), .B1(n18882), .B2(n18968), .ZN(
        n18888) );
  OAI22_X1 U20962 ( .A1(n18886), .A2(n18969), .B1(n18885), .B2(n18973), .ZN(
        n18887) );
  AOI211_X1 U20963 ( .C1(n18889), .C2(n18957), .A(n18888), .B(n18887), .ZN(
        n18894) );
  OAI211_X1 U20964 ( .C1(n18892), .C2(n18891), .A(n18980), .B(n18890), .ZN(
        n18893) );
  OAI211_X1 U20965 ( .C1(n18922), .C2(n18895), .A(n18894), .B(n18893), .ZN(
        P2_U2832) );
  AOI22_X1 U20966 ( .A1(n18896), .A2(n18952), .B1(n18954), .B2(
        P2_REIP_REG_24__SCAN_IN), .ZN(n18905) );
  AOI22_X1 U20967 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18955), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18951), .ZN(n18904) );
  INV_X1 U20968 ( .A(n18897), .ZN(n18899) );
  AOI22_X1 U20969 ( .A1(n18899), .A2(n18957), .B1(n18898), .B2(n18977), .ZN(
        n18903) );
  OAI211_X1 U20970 ( .C1(n18901), .C2(n18900), .A(n18980), .B(n18906), .ZN(
        n18902) );
  NAND4_X1 U20971 ( .A1(n18905), .A2(n18904), .A3(n18903), .A4(n18902), .ZN(
        P2_U2831) );
  NAND2_X1 U20972 ( .A1(n18906), .A2(n11165), .ZN(n18907) );
  XOR2_X1 U20973 ( .A(n18908), .B(n18907), .Z(n18916) );
  AOI22_X1 U20974 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18954), .ZN(n18911) );
  AOI22_X1 U20975 ( .A1(n18909), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18910) );
  OAI211_X1 U20976 ( .C1(n18912), .C2(n18922), .A(n18911), .B(n18910), .ZN(
        n18913) );
  AOI21_X1 U20977 ( .B1(n18914), .B2(n18957), .A(n18913), .ZN(n18915) );
  OAI21_X1 U20978 ( .B1(n19039), .B2(n18916), .A(n18915), .ZN(P2_U2830) );
  OAI21_X1 U20979 ( .B1(n18918), .B2(n18917), .A(n18980), .ZN(n18928) );
  AOI22_X1 U20980 ( .A1(n18919), .A2(n18952), .B1(n18955), .B2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18920) );
  OAI21_X1 U20981 ( .B1(n18921), .B2(n18968), .A(n18920), .ZN(n18926) );
  OAI22_X1 U20982 ( .A1(n18924), .A2(n18983), .B1(n18923), .B2(n18922), .ZN(
        n18925) );
  AOI211_X1 U20983 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n18951), .A(n18926), .B(
        n18925), .ZN(n18927) );
  OAI21_X1 U20984 ( .B1(n18929), .B2(n18928), .A(n18927), .ZN(P2_U2829) );
  AOI211_X1 U20985 ( .C1(n18931), .C2(n11293), .A(n18930), .B(n19039), .ZN(
        n18935) );
  AOI22_X1 U20986 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18954), .ZN(n18932) );
  OAI21_X1 U20987 ( .B1(n18933), .B2(n18969), .A(n18932), .ZN(n18934) );
  AOI211_X1 U20988 ( .C1(n18955), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n18935), .B(n18934), .ZN(n18939) );
  AOI22_X1 U20989 ( .A1(n18937), .A2(n18957), .B1(n18936), .B2(n18977), .ZN(
        n18938) );
  NAND2_X1 U20990 ( .A1(n18939), .A2(n18938), .ZN(P2_U2828) );
  AOI211_X1 U20991 ( .C1(n18942), .C2(n18941), .A(n18940), .B(n19039), .ZN(
        n18946) );
  AOI22_X1 U20992 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18951), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18954), .ZN(n18943) );
  OAI21_X1 U20993 ( .B1(n18944), .B2(n18969), .A(n18943), .ZN(n18945) );
  AOI211_X1 U20994 ( .C1(n18955), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n18946), .B(n18945), .ZN(n18950) );
  AOI22_X1 U20995 ( .A1(n18948), .A2(n18957), .B1(n18947), .B2(n18977), .ZN(
        n18949) );
  NAND2_X1 U20996 ( .A1(n18950), .A2(n18949), .ZN(P2_U2827) );
  AOI22_X1 U20997 ( .A1(n18953), .A2(n18952), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18951), .ZN(n18965) );
  AOI22_X1 U20998 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18955), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18954), .ZN(n18964) );
  AOI22_X1 U20999 ( .A1(n18958), .A2(n18957), .B1(n18956), .B2(n18977), .ZN(
        n18963) );
  AOI21_X1 U21000 ( .B1(n18960), .B2(n18959), .A(n18979), .ZN(n18961) );
  NAND2_X1 U21001 ( .A1(n18980), .A2(n18961), .ZN(n18962) );
  NAND4_X1 U21002 ( .A1(n18965), .A2(n18964), .A3(n18963), .A4(n18962), .ZN(
        P2_U2826) );
  INV_X1 U21003 ( .A(n18966), .ZN(n18970) );
  OAI22_X1 U21004 ( .A1(n18970), .A2(n18969), .B1(n18968), .B2(n18967), .ZN(
        n18976) );
  OAI22_X1 U21005 ( .A1(n18974), .A2(n18973), .B1(n18972), .B2(n18971), .ZN(
        n18975) );
  AOI211_X1 U21006 ( .C1(n18977), .C2(n19524), .A(n18976), .B(n18975), .ZN(
        n18982) );
  NAND4_X1 U21007 ( .A1(n18980), .A2(n18979), .A3(n18978), .A4(n11165), .ZN(
        n18981) );
  OAI211_X1 U21008 ( .C1(n16034), .C2(n18983), .A(n18982), .B(n18981), .ZN(
        P2_U2824) );
  NOR4_X1 U21009 ( .A1(n18984), .A2(n14776), .A3(n11855), .A4(n19034), .ZN(
        n18985) );
  NAND2_X1 U21010 ( .A1(n18988), .A2(n18985), .ZN(n18986) );
  OAI21_X1 U21011 ( .B1(n18988), .B2(n18987), .A(n18986), .ZN(P2_U3595) );
  AOI22_X1 U21012 ( .A1(n19024), .A2(n18990), .B1(n19003), .B2(n18989), .ZN(
        n19000) );
  OAI22_X1 U21013 ( .A1(n18994), .A2(n18993), .B1(n18992), .B2(n18991), .ZN(
        n18998) );
  OAI21_X1 U21014 ( .B1(n19015), .B2(n18996), .A(n18995), .ZN(n18997) );
  NOR2_X1 U21015 ( .A1(n18998), .A2(n18997), .ZN(n18999) );
  OAI211_X1 U21016 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19001), .A(
        n19000), .B(n18999), .ZN(P2_U3046) );
  AOI22_X1 U21017 ( .A1(n19004), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19003), .B2(n19002), .ZN(n19014) );
  AOI222_X1 U21018 ( .A1(n19008), .A2(n19007), .B1(n19017), .B2(n19006), .C1(
        n19024), .C2(n19005), .ZN(n19013) );
  NAND2_X1 U21019 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n11167), .ZN(n19012) );
  OAI211_X1 U21020 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n19010), .B(n19009), .ZN(n19011) );
  NAND4_X1 U21021 ( .A1(n19014), .A2(n19013), .A3(n19012), .A4(n19011), .ZN(
        P2_U3038) );
  NOR2_X1 U21022 ( .A1(n19016), .A2(n19015), .ZN(n19023) );
  NAND2_X1 U21023 ( .A1(n19017), .A2(n13756), .ZN(n19018) );
  OAI211_X1 U21024 ( .C1(n19021), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        n19022) );
  AOI211_X1 U21025 ( .C1(n19025), .C2(n19024), .A(n19023), .B(n19022), .ZN(
        n19029) );
  NAND3_X1 U21026 ( .A1(n19030), .A2(n19027), .A3(n19026), .ZN(n19028) );
  OAI211_X1 U21027 ( .C1(n19031), .C2(n19030), .A(n19029), .B(n19028), .ZN(
        P2_U3043) );
  NAND2_X1 U21028 ( .A1(n19046), .A2(n19032), .ZN(n19048) );
  OAI21_X1 U21029 ( .B1(n19034), .B2(n19033), .A(n19054), .ZN(n19038) );
  NAND2_X1 U21030 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19035), .ZN(n19036) );
  AOI21_X1 U21031 ( .B1(n19041), .B2(n19048), .A(n19036), .ZN(n19037) );
  AOI21_X1 U21032 ( .B1(n19048), .B2(n19038), .A(n19037), .ZN(n19040) );
  NAND2_X1 U21033 ( .A1(n19040), .A2(n19039), .ZN(P2_U3177) );
  OAI22_X1 U21034 ( .A1(n19043), .A2(n19042), .B1(n19041), .B2(n22174), .ZN(
        n19044) );
  AOI211_X1 U21035 ( .C1(n19046), .C2(P2_STATE2_REG_0__SCAN_IN), .A(n19045), 
        .B(n19044), .ZN(n19052) );
  NOR2_X1 U21036 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19047), .ZN(n19050) );
  OAI22_X1 U21037 ( .A1(n19050), .A2(n19049), .B1(n22174), .B2(n19048), .ZN(
        n19051) );
  OAI211_X1 U21038 ( .C1(n19053), .C2(n19054), .A(n19052), .B(n19051), .ZN(
        P2_U3176) );
  NOR2_X1 U21039 ( .A1(n19055), .A2(n19054), .ZN(n19058) );
  MUX2_X1 U21040 ( .A(P2_MORE_REG_SCAN_IN), .B(n19056), .S(n19058), .Z(
        P2_U3609) );
  OAI21_X1 U21041 ( .B1(n19058), .B2(n12747), .A(n19057), .ZN(P2_U2819) );
  INV_X1 U21042 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20457) );
  INV_X1 U21043 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19084) );
  AOI22_X1 U21044 ( .A1(n19293), .A2(n20457), .B1(n19084), .B2(U215), .ZN(U282) );
  OAI22_X1 U21045 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19293), .ZN(n19059) );
  INV_X1 U21046 ( .A(n19059), .ZN(U281) );
  OAI22_X1 U21047 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19419), .ZN(n19060) );
  INV_X1 U21048 ( .A(n19060), .ZN(U280) );
  INV_X1 U21049 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n19061) );
  INV_X1 U21050 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21092) );
  AOI22_X1 U21051 ( .A1(n19293), .A2(n19061), .B1(n21092), .B2(U215), .ZN(U279) );
  OAI22_X1 U21052 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19419), .ZN(n19062) );
  INV_X1 U21053 ( .A(n19062), .ZN(U278) );
  INV_X1 U21054 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n19063) );
  INV_X1 U21055 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n21074) );
  AOI22_X1 U21056 ( .A1(n19293), .A2(n19063), .B1(n21074), .B2(U215), .ZN(U277) );
  INV_X1 U21057 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n19064) );
  INV_X1 U21058 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n19962) );
  AOI22_X1 U21059 ( .A1(n19293), .A2(n19064), .B1(n19962), .B2(U215), .ZN(U276) );
  OAI22_X1 U21060 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19293), .ZN(n19065) );
  INV_X1 U21061 ( .A(n19065), .ZN(U275) );
  INV_X1 U21062 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n19066) );
  INV_X1 U21063 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19529) );
  AOI22_X1 U21064 ( .A1(n19293), .A2(n19066), .B1(n19529), .B2(U215), .ZN(U274) );
  OAI22_X1 U21065 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19419), .ZN(n19067) );
  INV_X1 U21066 ( .A(n19067), .ZN(U273) );
  INV_X1 U21067 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n19068) );
  AOI22_X1 U21068 ( .A1(n19419), .A2(n19068), .B1(n21028), .B2(U215), .ZN(U272) );
  OAI22_X1 U21069 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19293), .ZN(n19069) );
  INV_X1 U21070 ( .A(n19069), .ZN(U271) );
  OAI22_X1 U21071 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19293), .ZN(n19070) );
  INV_X1 U21072 ( .A(n19070), .ZN(U270) );
  OAI22_X1 U21073 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19293), .ZN(n19071) );
  INV_X1 U21074 ( .A(n19071), .ZN(U269) );
  OAI22_X1 U21075 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19293), .ZN(n19072) );
  INV_X1 U21076 ( .A(n19072), .ZN(U268) );
  OAI22_X1 U21077 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19293), .ZN(n19073) );
  INV_X1 U21078 ( .A(n19073), .ZN(U267) );
  OAI22_X1 U21079 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19293), .ZN(n19074) );
  INV_X1 U21080 ( .A(n19074), .ZN(U266) );
  OAI22_X1 U21081 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19293), .ZN(n19075) );
  INV_X1 U21082 ( .A(n19075), .ZN(U265) );
  OAI22_X1 U21083 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19293), .ZN(n19076) );
  INV_X1 U21084 ( .A(n19076), .ZN(U264) );
  INV_X1 U21085 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n19077) );
  INV_X1 U21086 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20982) );
  AOI22_X1 U21087 ( .A1(n19293), .A2(n19077), .B1(n20982), .B2(U215), .ZN(U263) );
  OAI22_X1 U21088 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19293), .ZN(n19078) );
  INV_X1 U21089 ( .A(n19078), .ZN(U262) );
  INV_X1 U21090 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19079) );
  INV_X1 U21091 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U21092 ( .A1(n19419), .A2(n19079), .B1(n20990), .B2(U215), .ZN(U261) );
  INV_X1 U21093 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n19080) );
  INV_X1 U21094 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20995) );
  AOI22_X1 U21095 ( .A1(n19293), .A2(n19080), .B1(n20995), .B2(U215), .ZN(U260) );
  INV_X1 U21096 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n19081) );
  INV_X1 U21097 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n21104) );
  AOI22_X1 U21098 ( .A1(n19419), .A2(n19081), .B1(n21104), .B2(U215), .ZN(U259) );
  INV_X1 U21099 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n19082) );
  INV_X1 U21100 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21001) );
  AOI22_X1 U21101 ( .A1(n19293), .A2(n19082), .B1(n21001), .B2(U215), .ZN(U258) );
  NOR3_X1 U21102 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21646), .A3(
        n19083), .ZN(n19096) );
  NAND2_X1 U21103 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19096), .ZN(
        n19523) );
  NAND2_X1 U21104 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19421), .ZN(n19157) );
  INV_X1 U21105 ( .A(n19096), .ZN(n19095) );
  NOR2_X2 U21106 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19095), .ZN(
        n19441) );
  NOR2_X1 U21107 ( .A1(n19084), .A2(n19252), .ZN(n19164) );
  NAND2_X1 U21108 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21668), .ZN(n21669) );
  INV_X1 U21109 ( .A(n21669), .ZN(n19162) );
  NAND2_X1 U21110 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19085), .ZN(
        n19091) );
  NOR2_X1 U21111 ( .A1(n19162), .A2(n19091), .ZN(n19423) );
  NOR2_X2 U21112 ( .A1(n21001), .A2(n19294), .ZN(n19163) );
  AOI22_X1 U21113 ( .A1(n19441), .A2(n19164), .B1(n19423), .B2(n19163), .ZN(
        n19090) );
  INV_X1 U21114 ( .A(n19091), .ZN(n19154) );
  NOR2_X1 U21115 ( .A1(n19086), .A2(n19294), .ZN(n19112) );
  AOI22_X1 U21116 ( .A1(n19421), .A2(n19096), .B1(n19154), .B2(n19112), .ZN(
        n19426) );
  NOR2_X2 U21117 ( .A1(n21637), .A2(n19091), .ZN(n19506) );
  NAND2_X1 U21118 ( .A1(n19088), .A2(n19087), .ZN(n19424) );
  NOR2_X2 U21119 ( .A1(n20997), .A2(n19424), .ZN(n19165) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19165), .ZN(n19089) );
  OAI211_X1 U21121 ( .C1(n19523), .C2(n19157), .A(n19090), .B(n19089), .ZN(
        P3_U2995) );
  INV_X1 U21122 ( .A(n19164), .ZN(n19145) );
  NAND2_X1 U21123 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21646), .ZN(
        n19111) );
  NOR2_X1 U21124 ( .A1(n21640), .A2(n19111), .ZN(n19104) );
  NAND2_X1 U21125 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19104), .ZN(
        n19382) );
  INV_X1 U21126 ( .A(n19157), .ZN(n19166) );
  INV_X1 U21127 ( .A(n19523), .ZN(n19435) );
  OR2_X1 U21128 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19091), .ZN(
        n19511) );
  INV_X1 U21129 ( .A(n19511), .ZN(n19515) );
  NOR2_X1 U21130 ( .A1(n19435), .A2(n19515), .ZN(n19160) );
  NOR2_X1 U21131 ( .A1(n19162), .A2(n19160), .ZN(n19429) );
  AOI22_X1 U21132 ( .A1(n19166), .A2(n19441), .B1(n19163), .B2(n19429), .ZN(
        n19094) );
  INV_X1 U21133 ( .A(n19382), .ZN(n19447) );
  NOR2_X1 U21134 ( .A1(n19441), .A2(n19447), .ZN(n19099) );
  INV_X1 U21135 ( .A(n19107), .ZN(n19124) );
  OAI21_X1 U21136 ( .B1(n19099), .B2(n19124), .A(n19160), .ZN(n19092) );
  OAI211_X1 U21137 ( .C1(n19515), .C2(n21676), .A(n19422), .B(n19092), .ZN(
        n19430) );
  AOI22_X1 U21138 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19430), .B1(
        n19165), .B2(n19515), .ZN(n19093) );
  OAI211_X1 U21139 ( .C1(n19145), .C2(n19382), .A(n19094), .B(n19093), .ZN(
        P3_U2987) );
  NAND2_X1 U21140 ( .A1(n19104), .A2(n21637), .ZN(n19439) );
  NOR2_X1 U21141 ( .A1(n19162), .A2(n19095), .ZN(n19434) );
  AOI22_X1 U21142 ( .A1(n19166), .A2(n19447), .B1(n19163), .B2(n19434), .ZN(
        n19098) );
  AOI22_X1 U21143 ( .A1(n19421), .A2(n19104), .B1(n19112), .B2(n19096), .ZN(
        n19436) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19165), .ZN(n19097) );
  OAI211_X1 U21145 ( .C1(n19145), .C2(n19439), .A(n19098), .B(n19097), .ZN(
        P3_U2979) );
  INV_X1 U21146 ( .A(n19111), .ZN(n19113) );
  NOR2_X1 U21147 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21637), .ZN(
        n19133) );
  NAND2_X1 U21148 ( .A1(n19113), .A2(n19133), .ZN(n19445) );
  INV_X1 U21149 ( .A(n19439), .ZN(n19453) );
  NOR2_X1 U21150 ( .A1(n19162), .A2(n19099), .ZN(n19440) );
  AOI22_X1 U21151 ( .A1(n19166), .A2(n19453), .B1(n19163), .B2(n19440), .ZN(
        n19102) );
  NAND2_X1 U21152 ( .A1(n19439), .A2(n19445), .ZN(n19108) );
  AOI21_X1 U21153 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19294), .ZN(n19135) );
  INV_X1 U21154 ( .A(n19099), .ZN(n19100) );
  AOI22_X1 U21155 ( .A1(n19421), .A2(n19108), .B1(n19135), .B2(n19100), .ZN(
        n19442) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19442), .B1(
        n19165), .B2(n19441), .ZN(n19101) );
  OAI211_X1 U21157 ( .C1(n19145), .C2(n19445), .A(n19102), .B(n19101), .ZN(
        P3_U2971) );
  NAND2_X1 U21158 ( .A1(n21640), .A2(n21637), .ZN(n21642) );
  NOR2_X2 U21159 ( .A1(n21642), .A2(n19111), .ZN(n19465) );
  INV_X1 U21160 ( .A(n19104), .ZN(n19103) );
  NOR2_X1 U21161 ( .A1(n19162), .A2(n19103), .ZN(n19446) );
  AOI22_X1 U21162 ( .A1(n19164), .A2(n19465), .B1(n19163), .B2(n19446), .ZN(
        n19106) );
  AOI22_X1 U21163 ( .A1(n19421), .A2(n19113), .B1(n19112), .B2(n19104), .ZN(
        n19448) );
  AOI22_X1 U21164 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19448), .B1(
        n19165), .B2(n19447), .ZN(n19105) );
  OAI211_X1 U21165 ( .C1(n19157), .C2(n19445), .A(n19106), .B(n19105), .ZN(
        P3_U2963) );
  INV_X1 U21166 ( .A(n19465), .ZN(n19451) );
  NOR2_X2 U21167 ( .A1(n21637), .A2(n19120), .ZN(n19472) );
  AND2_X1 U21168 ( .A1(n21669), .A2(n19108), .ZN(n19452) );
  AOI22_X1 U21169 ( .A1(n19164), .A2(n19472), .B1(n19163), .B2(n19452), .ZN(
        n19110) );
  INV_X1 U21170 ( .A(n19472), .ZN(n19457) );
  NAND2_X1 U21171 ( .A1(n19451), .A2(n19457), .ZN(n19117) );
  OAI221_X1 U21172 ( .B1(n19108), .B2(n19107), .C1(n19108), .C2(n19117), .A(
        n19135), .ZN(n19454) );
  AOI22_X1 U21173 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19454), .B1(
        n19165), .B2(n19453), .ZN(n19109) );
  OAI211_X1 U21174 ( .C1(n19157), .C2(n19451), .A(n19110), .B(n19109), .ZN(
        P3_U2955) );
  NAND2_X1 U21175 ( .A1(n21640), .A2(n21669), .ZN(n19151) );
  NOR2_X1 U21176 ( .A1(n19111), .A2(n19151), .ZN(n19458) );
  AOI22_X1 U21177 ( .A1(n19164), .A2(n11155), .B1(n19163), .B2(n19458), .ZN(
        n19116) );
  AND2_X1 U21178 ( .A1(n21640), .A2(n19112), .ZN(n19153) );
  AOI22_X1 U21179 ( .A1(n19421), .A2(n19114), .B1(n19113), .B2(n19153), .ZN(
        n19460) );
  INV_X1 U21180 ( .A(n19445), .ZN(n19459) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19460), .B1(
        n19165), .B2(n19459), .ZN(n19115) );
  OAI211_X1 U21182 ( .C1(n19157), .C2(n19457), .A(n19116), .B(n19115), .ZN(
        P3_U2947) );
  NOR2_X1 U21183 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21646), .ZN(
        n19129) );
  NAND2_X1 U21184 ( .A1(n19133), .A2(n19129), .ZN(n19469) );
  AND2_X1 U21185 ( .A1(n21669), .A2(n19117), .ZN(n19464) );
  AOI22_X1 U21186 ( .A1(n19166), .A2(n11155), .B1(n19163), .B2(n19464), .ZN(
        n19119) );
  INV_X1 U21187 ( .A(n11155), .ZN(n19463) );
  NAND2_X1 U21188 ( .A1(n19463), .A2(n19469), .ZN(n19123) );
  AOI22_X1 U21189 ( .A1(n19421), .A2(n19123), .B1(n19135), .B2(n19117), .ZN(
        n19466) );
  AOI22_X1 U21190 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19466), .B1(
        n19165), .B2(n19465), .ZN(n19118) );
  OAI211_X1 U21191 ( .C1(n19145), .C2(n19469), .A(n19119), .B(n19118), .ZN(
        P3_U2939) );
  AOI21_X1 U21192 ( .B1(n21640), .B2(n19124), .A(n19294), .ZN(n19142) );
  OAI211_X1 U21193 ( .C1(n19472), .C2(n21676), .A(n19129), .B(n19142), .ZN(
        n19471) );
  NOR2_X1 U21194 ( .A1(n19162), .A2(n19120), .ZN(n19470) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19471), .B1(
        n19163), .B2(n19470), .ZN(n19122) );
  INV_X1 U21196 ( .A(n19129), .ZN(n19128) );
  NOR2_X2 U21197 ( .A1(n21642), .A2(n19128), .ZN(n19487) );
  AOI22_X1 U21198 ( .A1(n19165), .A2(n19472), .B1(n19164), .B2(n19487), .ZN(
        n19121) );
  OAI211_X1 U21199 ( .C1(n19157), .C2(n19469), .A(n19122), .B(n19121), .ZN(
        P3_U2931) );
  NOR2_X1 U21200 ( .A1(n21640), .A2(n19150), .ZN(n19130) );
  NAND2_X1 U21201 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19130), .ZN(
        n19480) );
  AND2_X1 U21202 ( .A1(n21669), .A2(n19123), .ZN(n19476) );
  AOI22_X1 U21203 ( .A1(n19166), .A2(n19487), .B1(n19163), .B2(n19476), .ZN(
        n19127) );
  INV_X1 U21204 ( .A(n19480), .ZN(n19494) );
  NOR2_X1 U21205 ( .A1(n19487), .A2(n19494), .ZN(n19136) );
  OAI22_X1 U21206 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19469), .B1(n19136), 
        .B2(n19124), .ZN(n19125) );
  OAI21_X1 U21207 ( .B1(n11155), .B2(n19125), .A(n19422), .ZN(n19477) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19477), .B1(
        n19165), .B2(n11155), .ZN(n19126) );
  OAI211_X1 U21209 ( .C1(n19145), .C2(n19480), .A(n19127), .B(n19126), .ZN(
        P3_U2923) );
  INV_X1 U21210 ( .A(n19130), .ZN(n19141) );
  NOR2_X2 U21211 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19141), .ZN(
        n19499) );
  NOR2_X1 U21212 ( .A1(n19151), .A2(n19128), .ZN(n19481) );
  AOI22_X1 U21213 ( .A1(n19164), .A2(n19499), .B1(n19163), .B2(n19481), .ZN(
        n19132) );
  AOI22_X1 U21214 ( .A1(n19421), .A2(n19130), .B1(n19153), .B2(n19129), .ZN(
        n19483) );
  INV_X1 U21215 ( .A(n19469), .ZN(n19482) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19483), .B1(
        n19165), .B2(n19482), .ZN(n19131) );
  OAI211_X1 U21217 ( .C1(n19157), .C2(n19480), .A(n19132), .B(n19131), .ZN(
        P3_U2915) );
  INV_X1 U21218 ( .A(n19499), .ZN(n19491) );
  INV_X1 U21219 ( .A(n19133), .ZN(n19134) );
  NOR2_X2 U21220 ( .A1(n19134), .A2(n19150), .ZN(n19507) );
  NOR2_X1 U21221 ( .A1(n19162), .A2(n19136), .ZN(n19486) );
  AOI22_X1 U21222 ( .A1(n19164), .A2(n19507), .B1(n19163), .B2(n19486), .ZN(
        n19139) );
  NOR2_X1 U21223 ( .A1(n19499), .A2(n19507), .ZN(n19146) );
  INV_X1 U21224 ( .A(n19135), .ZN(n19159) );
  OAI22_X1 U21225 ( .A1(n19252), .A2(n19146), .B1(n19159), .B2(n19136), .ZN(
        n19137) );
  INV_X1 U21226 ( .A(n19137), .ZN(n19488) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19488), .B1(
        n19165), .B2(n19487), .ZN(n19138) );
  OAI211_X1 U21228 ( .C1(n19157), .C2(n19491), .A(n19139), .B(n19138), .ZN(
        P3_U2907) );
  INV_X1 U21229 ( .A(n21642), .ZN(n19140) );
  NAND2_X1 U21230 ( .A1(n19140), .A2(n19152), .ZN(n19504) );
  NOR2_X1 U21231 ( .A1(n19162), .A2(n19141), .ZN(n19492) );
  AOI22_X1 U21232 ( .A1(n19166), .A2(n19507), .B1(n19163), .B2(n19492), .ZN(
        n19144) );
  OAI211_X1 U21233 ( .C1(n19494), .C2(n21676), .A(n19152), .B(n19142), .ZN(
        n19493) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19493), .B1(
        n19165), .B2(n19494), .ZN(n19143) );
  OAI211_X1 U21235 ( .C1(n19145), .C2(n19504), .A(n19144), .B(n19143), .ZN(
        P3_U2899) );
  NOR2_X1 U21236 ( .A1(n19162), .A2(n19146), .ZN(n19497) );
  AOI22_X1 U21237 ( .A1(n19506), .A2(n19164), .B1(n19163), .B2(n19497), .ZN(
        n19149) );
  INV_X1 U21238 ( .A(n19507), .ZN(n19404) );
  OAI21_X1 U21239 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19404), .A(n19491), 
        .ZN(n19147) );
  INV_X1 U21240 ( .A(n19506), .ZN(n19411) );
  NAND2_X1 U21241 ( .A1(n19411), .A2(n19504), .ZN(n19158) );
  AOI22_X1 U21242 ( .A1(n19422), .A2(n19147), .B1(n19421), .B2(n19158), .ZN(
        n19500) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19500), .B1(
        n19165), .B2(n19499), .ZN(n19148) );
  OAI211_X1 U21244 ( .C1(n19157), .C2(n19504), .A(n19149), .B(n19148), .ZN(
        P3_U2891) );
  NOR2_X1 U21245 ( .A1(n19151), .A2(n19150), .ZN(n19505) );
  AOI22_X1 U21246 ( .A1(n19164), .A2(n19515), .B1(n19163), .B2(n19505), .ZN(
        n19156) );
  AOI22_X1 U21247 ( .A1(n19421), .A2(n19154), .B1(n19153), .B2(n19152), .ZN(
        n19508) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19508), .B1(
        n19165), .B2(n19507), .ZN(n19155) );
  OAI211_X1 U21249 ( .C1(n19157), .C2(n19411), .A(n19156), .B(n19155), .ZN(
        P3_U2883) );
  INV_X1 U21250 ( .A(n19158), .ZN(n19161) );
  OAI22_X1 U21251 ( .A1(n19160), .A2(n19252), .B1(n19161), .B2(n19159), .ZN(
        n19516) );
  NOR2_X1 U21252 ( .A1(n19162), .A2(n19161), .ZN(n19513) );
  AOI22_X1 U21253 ( .A1(n19435), .A2(n19164), .B1(n19163), .B2(n19513), .ZN(
        n19168) );
  INV_X1 U21254 ( .A(n19504), .ZN(n19518) );
  AOI22_X1 U21255 ( .A1(n19166), .A2(n19515), .B1(n19165), .B2(n19518), .ZN(
        n19167) );
  OAI211_X1 U21256 ( .C1(n19169), .C2(n19516), .A(n19168), .B(n19167), .ZN(
        P3_U2875) );
  INV_X1 U21257 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19170) );
  INV_X1 U21258 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21044) );
  AOI22_X1 U21259 ( .A1(n19419), .A2(n19170), .B1(n21044), .B2(U215), .ZN(U257) );
  NAND2_X1 U21260 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19421), .ZN(n19199) );
  NAND2_X1 U21261 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19421), .ZN(n19202) );
  INV_X1 U21262 ( .A(n19202), .ZN(n19204) );
  NOR2_X2 U21263 ( .A1(n21044), .A2(n19294), .ZN(n19203) );
  AOI22_X1 U21264 ( .A1(n19441), .A2(n19204), .B1(n19423), .B2(n19203), .ZN(
        n19172) );
  NOR2_X2 U21265 ( .A1(n21027), .A2(n19424), .ZN(n19205) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19205), .ZN(n19171) );
  OAI211_X1 U21267 ( .C1(n19523), .C2(n19199), .A(n19172), .B(n19171), .ZN(
        P3_U2994) );
  INV_X1 U21268 ( .A(n19199), .ZN(n19206) );
  AOI22_X1 U21269 ( .A1(n19441), .A2(n19206), .B1(n19429), .B2(n19203), .ZN(
        n19174) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19205), .ZN(n19173) );
  OAI211_X1 U21271 ( .C1(n19382), .C2(n19202), .A(n19174), .B(n19173), .ZN(
        P3_U2986) );
  AOI22_X1 U21272 ( .A1(n19453), .A2(n19204), .B1(n19434), .B2(n19203), .ZN(
        n19176) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19205), .ZN(n19175) );
  OAI211_X1 U21274 ( .C1(n19382), .C2(n19199), .A(n19176), .B(n19175), .ZN(
        P3_U2978) );
  AOI22_X1 U21275 ( .A1(n19453), .A2(n19206), .B1(n19440), .B2(n19203), .ZN(
        n19178) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19205), .ZN(n19177) );
  OAI211_X1 U21277 ( .C1(n19445), .C2(n19202), .A(n19178), .B(n19177), .ZN(
        P3_U2970) );
  AOI22_X1 U21278 ( .A1(n19459), .A2(n19206), .B1(n19446), .B2(n19203), .ZN(
        n19180) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19205), .ZN(n19179) );
  OAI211_X1 U21280 ( .C1(n19451), .C2(n19202), .A(n19180), .B(n19179), .ZN(
        P3_U2962) );
  AOI22_X1 U21281 ( .A1(n19472), .A2(n19204), .B1(n19452), .B2(n19203), .ZN(
        n19182) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19205), .ZN(n19181) );
  OAI211_X1 U21283 ( .C1(n19451), .C2(n19199), .A(n19182), .B(n19181), .ZN(
        P3_U2954) );
  AOI22_X1 U21284 ( .A1(n19472), .A2(n19206), .B1(n19458), .B2(n19203), .ZN(
        n19184) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19205), .ZN(n19183) );
  OAI211_X1 U21286 ( .C1(n19463), .C2(n19202), .A(n19184), .B(n19183), .ZN(
        P3_U2946) );
  AOI22_X1 U21287 ( .A1(n11155), .A2(n19206), .B1(n19464), .B2(n19203), .ZN(
        n19186) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19205), .ZN(n19185) );
  OAI211_X1 U21289 ( .C1(n19469), .C2(n19202), .A(n19186), .B(n19185), .ZN(
        P3_U2938) );
  AOI22_X1 U21290 ( .A1(n19487), .A2(n19204), .B1(n19470), .B2(n19203), .ZN(
        n19188) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19471), .B1(
        n19472), .B2(n19205), .ZN(n19187) );
  OAI211_X1 U21292 ( .C1(n19469), .C2(n19199), .A(n19188), .B(n19187), .ZN(
        P3_U2930) );
  INV_X1 U21293 ( .A(n19487), .ZN(n19475) );
  AOI22_X1 U21294 ( .A1(n19494), .A2(n19204), .B1(n19476), .B2(n19203), .ZN(
        n19190) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19205), .ZN(n19189) );
  OAI211_X1 U21296 ( .C1(n19475), .C2(n19199), .A(n19190), .B(n19189), .ZN(
        P3_U2922) );
  AOI22_X1 U21297 ( .A1(n19494), .A2(n19206), .B1(n19481), .B2(n19203), .ZN(
        n19192) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19205), .ZN(n19191) );
  OAI211_X1 U21299 ( .C1(n19491), .C2(n19202), .A(n19192), .B(n19191), .ZN(
        P3_U2914) );
  AOI22_X1 U21300 ( .A1(n19499), .A2(n19206), .B1(n19486), .B2(n19203), .ZN(
        n19194) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19205), .ZN(n19193) );
  OAI211_X1 U21302 ( .C1(n19404), .C2(n19202), .A(n19194), .B(n19193), .ZN(
        P3_U2906) );
  AOI22_X1 U21303 ( .A1(n19507), .A2(n19206), .B1(n19492), .B2(n19203), .ZN(
        n19196) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19493), .B1(
        n19494), .B2(n19205), .ZN(n19195) );
  OAI211_X1 U21305 ( .C1(n19504), .C2(n19202), .A(n19196), .B(n19195), .ZN(
        P3_U2898) );
  AOI22_X1 U21306 ( .A1(n19506), .A2(n19204), .B1(n19497), .B2(n19203), .ZN(
        n19198) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19205), .ZN(n19197) );
  OAI211_X1 U21308 ( .C1(n19504), .C2(n19199), .A(n19198), .B(n19197), .ZN(
        P3_U2890) );
  AOI22_X1 U21309 ( .A1(n19506), .A2(n19206), .B1(n19505), .B2(n19203), .ZN(
        n19201) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19205), .ZN(n19200) );
  OAI211_X1 U21311 ( .C1(n19511), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        P3_U2882) );
  AOI22_X1 U21312 ( .A1(n19435), .A2(n19204), .B1(n19513), .B2(n19203), .ZN(
        n19208) );
  AOI22_X1 U21313 ( .A1(n19515), .A2(n19206), .B1(n19518), .B2(n19205), .ZN(
        n19207) );
  OAI211_X1 U21314 ( .C1(n19209), .C2(n19516), .A(n19208), .B(n19207), .ZN(
        P3_U2874) );
  INV_X1 U21315 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n19210) );
  INV_X1 U21316 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U21317 ( .A1(n19293), .A2(n19210), .B1(n21010), .B2(U215), .ZN(U256) );
  NAND2_X1 U21318 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n19421), .ZN(n19243) );
  NAND2_X1 U21319 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19421), .ZN(n19228) );
  INV_X1 U21320 ( .A(n19228), .ZN(n19245) );
  NOR2_X2 U21321 ( .A1(n21010), .A2(n19294), .ZN(n19244) );
  AOI22_X1 U21322 ( .A1(n19441), .A2(n19245), .B1(n19423), .B2(n19244), .ZN(
        n19213) );
  NOR2_X2 U21323 ( .A1(n19211), .A2(n19424), .ZN(n19246) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19246), .ZN(n19212) );
  OAI211_X1 U21325 ( .C1(n19523), .C2(n19243), .A(n19213), .B(n19212), .ZN(
        P3_U2993) );
  INV_X1 U21326 ( .A(n19243), .ZN(n19247) );
  AOI22_X1 U21327 ( .A1(n19441), .A2(n19247), .B1(n19429), .B2(n19244), .ZN(
        n19215) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19246), .ZN(n19214) );
  OAI211_X1 U21329 ( .C1(n19382), .C2(n19228), .A(n19215), .B(n19214), .ZN(
        P3_U2985) );
  AOI22_X1 U21330 ( .A1(n19453), .A2(n19245), .B1(n19434), .B2(n19244), .ZN(
        n19217) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19246), .ZN(n19216) );
  OAI211_X1 U21332 ( .C1(n19382), .C2(n19243), .A(n19217), .B(n19216), .ZN(
        P3_U2977) );
  AOI22_X1 U21333 ( .A1(n19453), .A2(n19247), .B1(n19440), .B2(n19244), .ZN(
        n19219) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19246), .ZN(n19218) );
  OAI211_X1 U21335 ( .C1(n19445), .C2(n19228), .A(n19219), .B(n19218), .ZN(
        P3_U2969) );
  AOI22_X1 U21336 ( .A1(n19459), .A2(n19247), .B1(n19446), .B2(n19244), .ZN(
        n19221) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19246), .ZN(n19220) );
  OAI211_X1 U21338 ( .C1(n19451), .C2(n19228), .A(n19221), .B(n19220), .ZN(
        P3_U2961) );
  AOI22_X1 U21339 ( .A1(n19472), .A2(n19245), .B1(n19452), .B2(n19244), .ZN(
        n19223) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19246), .ZN(n19222) );
  OAI211_X1 U21341 ( .C1(n19451), .C2(n19243), .A(n19223), .B(n19222), .ZN(
        P3_U2953) );
  AOI22_X1 U21342 ( .A1(n19458), .A2(n19244), .B1(n11155), .B2(n19245), .ZN(
        n19225) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19246), .ZN(n19224) );
  OAI211_X1 U21344 ( .C1(n19457), .C2(n19243), .A(n19225), .B(n19224), .ZN(
        P3_U2945) );
  AOI22_X1 U21345 ( .A1(n11155), .A2(n19247), .B1(n19464), .B2(n19244), .ZN(
        n19227) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19246), .ZN(n19226) );
  OAI211_X1 U21347 ( .C1(n19469), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        P3_U2937) );
  AOI22_X1 U21348 ( .A1(n19487), .A2(n19245), .B1(n19470), .B2(n19244), .ZN(
        n19230) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19471), .B1(
        n19472), .B2(n19246), .ZN(n19229) );
  OAI211_X1 U21350 ( .C1(n19469), .C2(n19243), .A(n19230), .B(n19229), .ZN(
        P3_U2929) );
  AOI22_X1 U21351 ( .A1(n19494), .A2(n19245), .B1(n19476), .B2(n19244), .ZN(
        n19232) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19246), .ZN(n19231) );
  OAI211_X1 U21353 ( .C1(n19475), .C2(n19243), .A(n19232), .B(n19231), .ZN(
        P3_U2921) );
  AOI22_X1 U21354 ( .A1(n19499), .A2(n19245), .B1(n19481), .B2(n19244), .ZN(
        n19234) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19246), .ZN(n19233) );
  OAI211_X1 U21356 ( .C1(n19480), .C2(n19243), .A(n19234), .B(n19233), .ZN(
        P3_U2913) );
  AOI22_X1 U21357 ( .A1(n19507), .A2(n19245), .B1(n19486), .B2(n19244), .ZN(
        n19236) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19246), .ZN(n19235) );
  OAI211_X1 U21359 ( .C1(n19491), .C2(n19243), .A(n19236), .B(n19235), .ZN(
        P3_U2905) );
  AOI22_X1 U21360 ( .A1(n19518), .A2(n19245), .B1(n19492), .B2(n19244), .ZN(
        n19238) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19493), .B1(
        n19494), .B2(n19246), .ZN(n19237) );
  OAI211_X1 U21362 ( .C1(n19404), .C2(n19243), .A(n19238), .B(n19237), .ZN(
        P3_U2897) );
  AOI22_X1 U21363 ( .A1(n19506), .A2(n19245), .B1(n19497), .B2(n19244), .ZN(
        n19240) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19246), .ZN(n19239) );
  OAI211_X1 U21365 ( .C1(n19504), .C2(n19243), .A(n19240), .B(n19239), .ZN(
        P3_U2889) );
  AOI22_X1 U21366 ( .A1(n19515), .A2(n19245), .B1(n19505), .B2(n19244), .ZN(
        n19242) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19246), .ZN(n19241) );
  OAI211_X1 U21368 ( .C1(n19411), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P3_U2881) );
  AOI22_X1 U21369 ( .A1(n19435), .A2(n19245), .B1(n19513), .B2(n19244), .ZN(
        n19249) );
  AOI22_X1 U21370 ( .A1(n19515), .A2(n19247), .B1(n19518), .B2(n19246), .ZN(
        n19248) );
  OAI211_X1 U21371 ( .C1(n19250), .C2(n19516), .A(n19249), .B(n19248), .ZN(
        P3_U2873) );
  INV_X1 U21372 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19251) );
  INV_X1 U21373 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21036) );
  AOI22_X1 U21374 ( .A1(n19293), .A2(n19251), .B1(n21036), .B2(U215), .ZN(U255) );
  NAND2_X1 U21375 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19421), .ZN(n19284) );
  NOR2_X1 U21376 ( .A1(n21092), .A2(n19252), .ZN(n19288) );
  NOR2_X2 U21377 ( .A1(n21036), .A2(n19294), .ZN(n19285) );
  AOI22_X1 U21378 ( .A1(n19441), .A2(n19288), .B1(n19423), .B2(n19285), .ZN(
        n19254) );
  NOR2_X2 U21379 ( .A1(n21221), .A2(n19424), .ZN(n19287) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19287), .ZN(n19253) );
  OAI211_X1 U21381 ( .C1(n19523), .C2(n19284), .A(n19254), .B(n19253), .ZN(
        P3_U2992) );
  INV_X1 U21382 ( .A(n19441), .ZN(n19433) );
  AOI22_X1 U21383 ( .A1(n19447), .A2(n19288), .B1(n19429), .B2(n19285), .ZN(
        n19256) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19287), .ZN(n19255) );
  OAI211_X1 U21385 ( .C1(n19433), .C2(n19284), .A(n19256), .B(n19255), .ZN(
        P3_U2984) );
  AOI22_X1 U21386 ( .A1(n19453), .A2(n19288), .B1(n19434), .B2(n19285), .ZN(
        n19258) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19287), .ZN(n19257) );
  OAI211_X1 U21388 ( .C1(n19382), .C2(n19284), .A(n19258), .B(n19257), .ZN(
        P3_U2976) );
  AOI22_X1 U21389 ( .A1(n19459), .A2(n19288), .B1(n19440), .B2(n19285), .ZN(
        n19260) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19287), .ZN(n19259) );
  OAI211_X1 U21391 ( .C1(n19439), .C2(n19284), .A(n19260), .B(n19259), .ZN(
        P3_U2968) );
  AOI22_X1 U21392 ( .A1(n19465), .A2(n19288), .B1(n19446), .B2(n19285), .ZN(
        n19262) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19287), .ZN(n19261) );
  OAI211_X1 U21394 ( .C1(n19445), .C2(n19284), .A(n19262), .B(n19261), .ZN(
        P3_U2960) );
  INV_X1 U21395 ( .A(n19288), .ZN(n19281) );
  INV_X1 U21396 ( .A(n19284), .ZN(n19286) );
  AOI22_X1 U21397 ( .A1(n19465), .A2(n19286), .B1(n19452), .B2(n19285), .ZN(
        n19264) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19287), .ZN(n19263) );
  OAI211_X1 U21399 ( .C1(n19457), .C2(n19281), .A(n19264), .B(n19263), .ZN(
        P3_U2952) );
  AOI22_X1 U21400 ( .A1(n19458), .A2(n19285), .B1(n19288), .B2(n11155), .ZN(
        n19266) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19287), .ZN(n19265) );
  OAI211_X1 U21402 ( .C1(n19457), .C2(n19284), .A(n19266), .B(n19265), .ZN(
        P3_U2944) );
  AOI22_X1 U21403 ( .A1(n19482), .A2(n19288), .B1(n19464), .B2(n19285), .ZN(
        n19268) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19287), .ZN(n19267) );
  OAI211_X1 U21405 ( .C1(n19463), .C2(n19284), .A(n19268), .B(n19267), .ZN(
        P3_U2936) );
  AOI22_X1 U21406 ( .A1(n19482), .A2(n19286), .B1(n19470), .B2(n19285), .ZN(
        n19270) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19471), .B1(
        n19472), .B2(n19287), .ZN(n19269) );
  OAI211_X1 U21408 ( .C1(n19475), .C2(n19281), .A(n19270), .B(n19269), .ZN(
        P3_U2928) );
  AOI22_X1 U21409 ( .A1(n19487), .A2(n19286), .B1(n19476), .B2(n19285), .ZN(
        n19272) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19287), .ZN(n19271) );
  OAI211_X1 U21411 ( .C1(n19480), .C2(n19281), .A(n19272), .B(n19271), .ZN(
        P3_U2920) );
  AOI22_X1 U21412 ( .A1(n19494), .A2(n19286), .B1(n19481), .B2(n19285), .ZN(
        n19274) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19287), .ZN(n19273) );
  OAI211_X1 U21414 ( .C1(n19491), .C2(n19281), .A(n19274), .B(n19273), .ZN(
        P3_U2912) );
  AOI22_X1 U21415 ( .A1(n19507), .A2(n19288), .B1(n19486), .B2(n19285), .ZN(
        n19276) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19287), .ZN(n19275) );
  OAI211_X1 U21417 ( .C1(n19491), .C2(n19284), .A(n19276), .B(n19275), .ZN(
        P3_U2904) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19285), .ZN(n19278) );
  AOI22_X1 U21419 ( .A1(n19494), .A2(n19287), .B1(n19518), .B2(n19288), .ZN(
        n19277) );
  OAI211_X1 U21420 ( .C1(n19404), .C2(n19284), .A(n19278), .B(n19277), .ZN(
        P3_U2896) );
  AOI22_X1 U21421 ( .A1(n19518), .A2(n19286), .B1(n19497), .B2(n19285), .ZN(
        n19280) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19287), .ZN(n19279) );
  OAI211_X1 U21423 ( .C1(n19411), .C2(n19281), .A(n19280), .B(n19279), .ZN(
        P3_U2888) );
  AOI22_X1 U21424 ( .A1(n19515), .A2(n19288), .B1(n19505), .B2(n19285), .ZN(
        n19283) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19287), .ZN(n19282) );
  OAI211_X1 U21426 ( .C1(n19411), .C2(n19284), .A(n19283), .B(n19282), .ZN(
        P3_U2880) );
  AOI22_X1 U21427 ( .A1(n19515), .A2(n19286), .B1(n19513), .B2(n19285), .ZN(
        n19290) );
  AOI22_X1 U21428 ( .A1(n19435), .A2(n19288), .B1(n19518), .B2(n19287), .ZN(
        n19289) );
  OAI211_X1 U21429 ( .C1(n19291), .C2(n19516), .A(n19290), .B(n19289), .ZN(
        P3_U2872) );
  INV_X1 U21430 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n19292) );
  INV_X1 U21431 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21019) );
  AOI22_X1 U21432 ( .A1(n19293), .A2(n19292), .B1(n21019), .B2(U215), .ZN(U254) );
  NAND2_X1 U21433 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19421), .ZN(n19327) );
  NAND2_X1 U21434 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19421), .ZN(n19322) );
  INV_X1 U21435 ( .A(n19322), .ZN(n19329) );
  NOR2_X2 U21436 ( .A1(n21019), .A2(n19294), .ZN(n19328) );
  AOI22_X1 U21437 ( .A1(n19435), .A2(n19329), .B1(n19423), .B2(n19328), .ZN(
        n19297) );
  NOR2_X2 U21438 ( .A1(n19295), .A2(n19424), .ZN(n19330) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19330), .ZN(n19296) );
  OAI211_X1 U21440 ( .C1(n19433), .C2(n19327), .A(n19297), .B(n19296), .ZN(
        P3_U2991) );
  AOI22_X1 U21441 ( .A1(n19441), .A2(n19329), .B1(n19429), .B2(n19328), .ZN(
        n19299) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19330), .ZN(n19298) );
  OAI211_X1 U21443 ( .C1(n19382), .C2(n19327), .A(n19299), .B(n19298), .ZN(
        P3_U2983) );
  INV_X1 U21444 ( .A(n19327), .ZN(n19331) );
  AOI22_X1 U21445 ( .A1(n19453), .A2(n19331), .B1(n19434), .B2(n19328), .ZN(
        n19301) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19330), .ZN(n19300) );
  OAI211_X1 U21447 ( .C1(n19382), .C2(n19322), .A(n19301), .B(n19300), .ZN(
        P3_U2975) );
  AOI22_X1 U21448 ( .A1(n19459), .A2(n19331), .B1(n19440), .B2(n19328), .ZN(
        n19303) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19330), .ZN(n19302) );
  OAI211_X1 U21450 ( .C1(n19439), .C2(n19322), .A(n19303), .B(n19302), .ZN(
        P3_U2967) );
  AOI22_X1 U21451 ( .A1(n19459), .A2(n19329), .B1(n19446), .B2(n19328), .ZN(
        n19305) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19330), .ZN(n19304) );
  OAI211_X1 U21453 ( .C1(n19451), .C2(n19327), .A(n19305), .B(n19304), .ZN(
        P3_U2959) );
  AOI22_X1 U21454 ( .A1(n19465), .A2(n19329), .B1(n19452), .B2(n19328), .ZN(
        n19307) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19330), .ZN(n19306) );
  OAI211_X1 U21456 ( .C1(n19457), .C2(n19327), .A(n19307), .B(n19306), .ZN(
        P3_U2951) );
  AOI22_X1 U21457 ( .A1(n19458), .A2(n19328), .B1(n11155), .B2(n19331), .ZN(
        n19309) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19330), .ZN(n19308) );
  OAI211_X1 U21459 ( .C1(n19457), .C2(n19322), .A(n19309), .B(n19308), .ZN(
        P3_U2943) );
  AOI22_X1 U21460 ( .A1(n11155), .A2(n19329), .B1(n19464), .B2(n19328), .ZN(
        n19311) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19330), .ZN(n19310) );
  OAI211_X1 U21462 ( .C1(n19469), .C2(n19327), .A(n19311), .B(n19310), .ZN(
        P3_U2935) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19328), .ZN(n19313) );
  AOI22_X1 U21464 ( .A1(n19472), .A2(n19330), .B1(n19482), .B2(n19329), .ZN(
        n19312) );
  OAI211_X1 U21465 ( .C1(n19475), .C2(n19327), .A(n19313), .B(n19312), .ZN(
        P3_U2927) );
  AOI22_X1 U21466 ( .A1(n19494), .A2(n19331), .B1(n19476), .B2(n19328), .ZN(
        n19315) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19330), .ZN(n19314) );
  OAI211_X1 U21468 ( .C1(n19475), .C2(n19322), .A(n19315), .B(n19314), .ZN(
        P3_U2919) );
  AOI22_X1 U21469 ( .A1(n19499), .A2(n19331), .B1(n19481), .B2(n19328), .ZN(
        n19317) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19330), .ZN(n19316) );
  OAI211_X1 U21471 ( .C1(n19480), .C2(n19322), .A(n19317), .B(n19316), .ZN(
        P3_U2911) );
  AOI22_X1 U21472 ( .A1(n19499), .A2(n19329), .B1(n19486), .B2(n19328), .ZN(
        n19319) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19330), .ZN(n19318) );
  OAI211_X1 U21474 ( .C1(n19404), .C2(n19327), .A(n19319), .B(n19318), .ZN(
        P3_U2903) );
  AOI22_X1 U21475 ( .A1(n19518), .A2(n19331), .B1(n19492), .B2(n19328), .ZN(
        n19321) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19493), .B1(
        n19494), .B2(n19330), .ZN(n19320) );
  OAI211_X1 U21477 ( .C1(n19404), .C2(n19322), .A(n19321), .B(n19320), .ZN(
        P3_U2895) );
  AOI22_X1 U21478 ( .A1(n19518), .A2(n19329), .B1(n19497), .B2(n19328), .ZN(
        n19324) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19330), .ZN(n19323) );
  OAI211_X1 U21480 ( .C1(n19411), .C2(n19327), .A(n19324), .B(n19323), .ZN(
        P3_U2887) );
  AOI22_X1 U21481 ( .A1(n19506), .A2(n19329), .B1(n19505), .B2(n19328), .ZN(
        n19326) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19330), .ZN(n19325) );
  OAI211_X1 U21483 ( .C1(n19511), .C2(n19327), .A(n19326), .B(n19325), .ZN(
        P3_U2879) );
  AOI22_X1 U21484 ( .A1(n19515), .A2(n19329), .B1(n19513), .B2(n19328), .ZN(
        n19333) );
  AOI22_X1 U21485 ( .A1(n19435), .A2(n19331), .B1(n19518), .B2(n19330), .ZN(
        n19332) );
  OAI211_X1 U21486 ( .C1(n19334), .C2(n19516), .A(n19333), .B(n19332), .ZN(
        P3_U2871) );
  OAI22_X1 U21487 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19419), .ZN(n19335) );
  INV_X1 U21488 ( .A(n19335), .ZN(U253) );
  NAND2_X1 U21489 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19421), .ZN(n19364) );
  NAND2_X1 U21490 ( .A1(n19421), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19367) );
  INV_X1 U21491 ( .A(n19367), .ZN(n19371) );
  AND2_X1 U21492 ( .A1(n19422), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19368) );
  AOI22_X1 U21493 ( .A1(n19435), .A2(n19371), .B1(n19423), .B2(n19368), .ZN(
        n19337) );
  NOR2_X2 U21494 ( .A1(n21212), .A2(n19424), .ZN(n19370) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19370), .ZN(n19336) );
  OAI211_X1 U21496 ( .C1(n19433), .C2(n19364), .A(n19337), .B(n19336), .ZN(
        P3_U2990) );
  INV_X1 U21497 ( .A(n19364), .ZN(n19369) );
  AOI22_X1 U21498 ( .A1(n19447), .A2(n19369), .B1(n19429), .B2(n19368), .ZN(
        n19339) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19370), .ZN(n19338) );
  OAI211_X1 U21500 ( .C1(n19433), .C2(n19367), .A(n19339), .B(n19338), .ZN(
        P3_U2982) );
  AOI22_X1 U21501 ( .A1(n19453), .A2(n19369), .B1(n19434), .B2(n19368), .ZN(
        n19341) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19370), .ZN(n19340) );
  OAI211_X1 U21503 ( .C1(n19382), .C2(n19367), .A(n19341), .B(n19340), .ZN(
        P3_U2974) );
  AOI22_X1 U21504 ( .A1(n19459), .A2(n19369), .B1(n19440), .B2(n19368), .ZN(
        n19343) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19370), .ZN(n19342) );
  OAI211_X1 U21506 ( .C1(n19439), .C2(n19367), .A(n19343), .B(n19342), .ZN(
        P3_U2966) );
  AOI22_X1 U21507 ( .A1(n19465), .A2(n19369), .B1(n19446), .B2(n19368), .ZN(
        n19345) );
  AOI22_X1 U21508 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19370), .ZN(n19344) );
  OAI211_X1 U21509 ( .C1(n19445), .C2(n19367), .A(n19345), .B(n19344), .ZN(
        P3_U2958) );
  AOI22_X1 U21510 ( .A1(n19472), .A2(n19369), .B1(n19452), .B2(n19368), .ZN(
        n19347) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19370), .ZN(n19346) );
  OAI211_X1 U21512 ( .C1(n19451), .C2(n19367), .A(n19347), .B(n19346), .ZN(
        P3_U2950) );
  AOI22_X1 U21513 ( .A1(n19458), .A2(n19368), .B1(n11155), .B2(n19369), .ZN(
        n19349) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19370), .ZN(n19348) );
  OAI211_X1 U21515 ( .C1(n19457), .C2(n19367), .A(n19349), .B(n19348), .ZN(
        P3_U2942) );
  AOI22_X1 U21516 ( .A1(n11155), .A2(n19371), .B1(n19464), .B2(n19368), .ZN(
        n19351) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19370), .ZN(n19350) );
  OAI211_X1 U21518 ( .C1(n19469), .C2(n19364), .A(n19351), .B(n19350), .ZN(
        P3_U2934) );
  AOI22_X1 U21519 ( .A1(n19482), .A2(n19371), .B1(n19470), .B2(n19368), .ZN(
        n19353) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19471), .B1(
        n19472), .B2(n19370), .ZN(n19352) );
  OAI211_X1 U21521 ( .C1(n19475), .C2(n19364), .A(n19353), .B(n19352), .ZN(
        P3_U2926) );
  AOI22_X1 U21522 ( .A1(n19487), .A2(n19371), .B1(n19476), .B2(n19368), .ZN(
        n19355) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19370), .ZN(n19354) );
  OAI211_X1 U21524 ( .C1(n19480), .C2(n19364), .A(n19355), .B(n19354), .ZN(
        P3_U2918) );
  AOI22_X1 U21525 ( .A1(n19499), .A2(n19369), .B1(n19481), .B2(n19368), .ZN(
        n19357) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19370), .ZN(n19356) );
  OAI211_X1 U21527 ( .C1(n19480), .C2(n19367), .A(n19357), .B(n19356), .ZN(
        P3_U2910) );
  AOI22_X1 U21528 ( .A1(n19507), .A2(n19369), .B1(n19486), .B2(n19368), .ZN(
        n19359) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19370), .ZN(n19358) );
  OAI211_X1 U21530 ( .C1(n19491), .C2(n19367), .A(n19359), .B(n19358), .ZN(
        P3_U2902) );
  AOI22_X1 U21531 ( .A1(n19518), .A2(n19369), .B1(n19492), .B2(n19368), .ZN(
        n19361) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19493), .B1(
        n19494), .B2(n19370), .ZN(n19360) );
  OAI211_X1 U21533 ( .C1(n19404), .C2(n19367), .A(n19361), .B(n19360), .ZN(
        P3_U2894) );
  AOI22_X1 U21534 ( .A1(n19518), .A2(n19371), .B1(n19497), .B2(n19368), .ZN(
        n19363) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19370), .ZN(n19362) );
  OAI211_X1 U21536 ( .C1(n19411), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P3_U2886) );
  AOI22_X1 U21537 ( .A1(n19515), .A2(n19369), .B1(n19505), .B2(n19368), .ZN(
        n19366) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19370), .ZN(n19365) );
  OAI211_X1 U21539 ( .C1(n19411), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P3_U2878) );
  AOI22_X1 U21540 ( .A1(n19435), .A2(n19369), .B1(n19513), .B2(n19368), .ZN(
        n19373) );
  AOI22_X1 U21541 ( .A1(n19515), .A2(n19371), .B1(n19518), .B2(n19370), .ZN(
        n19372) );
  OAI211_X1 U21542 ( .C1(n19374), .C2(n19516), .A(n19373), .B(n19372), .ZN(
        P3_U2870) );
  OAI22_X1 U21543 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19419), .ZN(n19375) );
  INV_X1 U21544 ( .A(n19375), .ZN(U252) );
  NAND2_X1 U21545 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19421), .ZN(n19407) );
  NAND2_X1 U21546 ( .A1(n19421), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19410) );
  INV_X1 U21547 ( .A(n19410), .ZN(n19413) );
  AND2_X1 U21548 ( .A1(n19422), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19412) );
  AOI22_X1 U21549 ( .A1(n19435), .A2(n19413), .B1(n19423), .B2(n19412), .ZN(
        n19377) );
  NOR2_X2 U21550 ( .A1(n20529), .A2(n19424), .ZN(n19414) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19414), .ZN(n19376) );
  OAI211_X1 U21552 ( .C1(n19433), .C2(n19407), .A(n19377), .B(n19376), .ZN(
        P3_U2989) );
  INV_X1 U21553 ( .A(n19407), .ZN(n19415) );
  AOI22_X1 U21554 ( .A1(n19447), .A2(n19415), .B1(n19429), .B2(n19412), .ZN(
        n19379) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19414), .ZN(n19378) );
  OAI211_X1 U21556 ( .C1(n19433), .C2(n19410), .A(n19379), .B(n19378), .ZN(
        P3_U2981) );
  AOI22_X1 U21557 ( .A1(n19453), .A2(n19415), .B1(n19434), .B2(n19412), .ZN(
        n19381) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19414), .ZN(n19380) );
  OAI211_X1 U21559 ( .C1(n19382), .C2(n19410), .A(n19381), .B(n19380), .ZN(
        P3_U2973) );
  AOI22_X1 U21560 ( .A1(n19459), .A2(n19415), .B1(n19440), .B2(n19412), .ZN(
        n19384) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19414), .ZN(n19383) );
  OAI211_X1 U21562 ( .C1(n19439), .C2(n19410), .A(n19384), .B(n19383), .ZN(
        P3_U2965) );
  AOI22_X1 U21563 ( .A1(n19465), .A2(n19415), .B1(n19446), .B2(n19412), .ZN(
        n19386) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19414), .ZN(n19385) );
  OAI211_X1 U21565 ( .C1(n19445), .C2(n19410), .A(n19386), .B(n19385), .ZN(
        P3_U2957) );
  AOI22_X1 U21566 ( .A1(n19472), .A2(n19415), .B1(n19452), .B2(n19412), .ZN(
        n19388) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19414), .ZN(n19387) );
  OAI211_X1 U21568 ( .C1(n19451), .C2(n19410), .A(n19388), .B(n19387), .ZN(
        P3_U2949) );
  AOI22_X1 U21569 ( .A1(n19458), .A2(n19412), .B1(n11155), .B2(n19415), .ZN(
        n19391) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19414), .ZN(n19390) );
  OAI211_X1 U21571 ( .C1(n19457), .C2(n19410), .A(n19391), .B(n19390), .ZN(
        P3_U2941) );
  AOI22_X1 U21572 ( .A1(n19482), .A2(n19415), .B1(n19464), .B2(n19412), .ZN(
        n19393) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19414), .ZN(n19392) );
  OAI211_X1 U21574 ( .C1(n19463), .C2(n19410), .A(n19393), .B(n19392), .ZN(
        P3_U2933) );
  AOI22_X1 U21575 ( .A1(n19482), .A2(n19413), .B1(n19470), .B2(n19412), .ZN(
        n19395) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19471), .B1(
        n19472), .B2(n19414), .ZN(n19394) );
  OAI211_X1 U21577 ( .C1(n19475), .C2(n19407), .A(n19395), .B(n19394), .ZN(
        P3_U2925) );
  AOI22_X1 U21578 ( .A1(n19494), .A2(n19415), .B1(n19476), .B2(n19412), .ZN(
        n19397) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19414), .ZN(n19396) );
  OAI211_X1 U21580 ( .C1(n19475), .C2(n19410), .A(n19397), .B(n19396), .ZN(
        P3_U2917) );
  AOI22_X1 U21581 ( .A1(n19494), .A2(n19413), .B1(n19481), .B2(n19412), .ZN(
        n19399) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19414), .ZN(n19398) );
  OAI211_X1 U21583 ( .C1(n19491), .C2(n19407), .A(n19399), .B(n19398), .ZN(
        P3_U2909) );
  AOI22_X1 U21584 ( .A1(n19499), .A2(n19413), .B1(n19486), .B2(n19412), .ZN(
        n19401) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19414), .ZN(n19400) );
  OAI211_X1 U21586 ( .C1(n19404), .C2(n19407), .A(n19401), .B(n19400), .ZN(
        P3_U2901) );
  AOI22_X1 U21587 ( .A1(n19518), .A2(n19415), .B1(n19492), .B2(n19412), .ZN(
        n19403) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19493), .B1(
        n19494), .B2(n19414), .ZN(n19402) );
  OAI211_X1 U21589 ( .C1(n19404), .C2(n19410), .A(n19403), .B(n19402), .ZN(
        P3_U2893) );
  AOI22_X1 U21590 ( .A1(n19518), .A2(n19413), .B1(n19497), .B2(n19412), .ZN(
        n19406) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19414), .ZN(n19405) );
  OAI211_X1 U21592 ( .C1(n19411), .C2(n19407), .A(n19406), .B(n19405), .ZN(
        P3_U2885) );
  AOI22_X1 U21593 ( .A1(n19515), .A2(n19415), .B1(n19505), .B2(n19412), .ZN(
        n19409) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19414), .ZN(n19408) );
  OAI211_X1 U21595 ( .C1(n19411), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P3_U2877) );
  AOI22_X1 U21596 ( .A1(n19515), .A2(n19413), .B1(n19513), .B2(n19412), .ZN(
        n19417) );
  AOI22_X1 U21597 ( .A1(n19435), .A2(n19415), .B1(n19518), .B2(n19414), .ZN(
        n19416) );
  OAI211_X1 U21598 ( .C1(n19418), .C2(n19516), .A(n19417), .B(n19416), .ZN(
        P3_U2869) );
  OAI22_X1 U21599 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19419), .ZN(n19420) );
  INV_X1 U21600 ( .A(n19420), .ZN(U251) );
  NAND2_X1 U21601 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19421), .ZN(n19522) );
  NAND2_X1 U21602 ( .A1(n19421), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19503) );
  INV_X1 U21603 ( .A(n19503), .ZN(n19514) );
  AND2_X1 U21604 ( .A1(n19422), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19512) );
  AOI22_X1 U21605 ( .A1(n19435), .A2(n19514), .B1(n19423), .B2(n19512), .ZN(
        n19428) );
  NOR2_X2 U21606 ( .A1(n19425), .A2(n19424), .ZN(n19517) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19426), .B1(
        n19506), .B2(n19517), .ZN(n19427) );
  OAI211_X1 U21608 ( .C1(n19433), .C2(n19522), .A(n19428), .B(n19427), .ZN(
        P3_U2988) );
  INV_X1 U21609 ( .A(n19522), .ZN(n19498) );
  AOI22_X1 U21610 ( .A1(n19447), .A2(n19498), .B1(n19429), .B2(n19512), .ZN(
        n19432) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19430), .B1(
        n19515), .B2(n19517), .ZN(n19431) );
  OAI211_X1 U21612 ( .C1(n19433), .C2(n19503), .A(n19432), .B(n19431), .ZN(
        P3_U2980) );
  AOI22_X1 U21613 ( .A1(n19447), .A2(n19514), .B1(n19434), .B2(n19512), .ZN(
        n19438) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19436), .B1(
        n19435), .B2(n19517), .ZN(n19437) );
  OAI211_X1 U21615 ( .C1(n19439), .C2(n19522), .A(n19438), .B(n19437), .ZN(
        P3_U2972) );
  AOI22_X1 U21616 ( .A1(n19453), .A2(n19514), .B1(n19440), .B2(n19512), .ZN(
        n19444) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19517), .ZN(n19443) );
  OAI211_X1 U21618 ( .C1(n19445), .C2(n19522), .A(n19444), .B(n19443), .ZN(
        P3_U2964) );
  AOI22_X1 U21619 ( .A1(n19459), .A2(n19514), .B1(n19446), .B2(n19512), .ZN(
        n19450) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19517), .ZN(n19449) );
  OAI211_X1 U21621 ( .C1(n19451), .C2(n19522), .A(n19450), .B(n19449), .ZN(
        P3_U2956) );
  AOI22_X1 U21622 ( .A1(n19465), .A2(n19514), .B1(n19452), .B2(n19512), .ZN(
        n19456) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19454), .B1(
        n19453), .B2(n19517), .ZN(n19455) );
  OAI211_X1 U21624 ( .C1(n19457), .C2(n19522), .A(n19456), .B(n19455), .ZN(
        P3_U2948) );
  AOI22_X1 U21625 ( .A1(n19472), .A2(n19514), .B1(n19458), .B2(n19512), .ZN(
        n19462) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19517), .ZN(n19461) );
  OAI211_X1 U21627 ( .C1(n19463), .C2(n19522), .A(n19462), .B(n19461), .ZN(
        P3_U2940) );
  AOI22_X1 U21628 ( .A1(n11155), .A2(n19514), .B1(n19464), .B2(n19512), .ZN(
        n19468) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19466), .B1(
        n19465), .B2(n19517), .ZN(n19467) );
  OAI211_X1 U21630 ( .C1(n19469), .C2(n19522), .A(n19468), .B(n19467), .ZN(
        P3_U2932) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19471), .B1(
        n19470), .B2(n19512), .ZN(n19474) );
  AOI22_X1 U21632 ( .A1(n19472), .A2(n19517), .B1(n19482), .B2(n19514), .ZN(
        n19473) );
  OAI211_X1 U21633 ( .C1(n19475), .C2(n19522), .A(n19474), .B(n19473), .ZN(
        P3_U2924) );
  AOI22_X1 U21634 ( .A1(n19487), .A2(n19514), .B1(n19476), .B2(n19512), .ZN(
        n19479) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19477), .B1(
        n11155), .B2(n19517), .ZN(n19478) );
  OAI211_X1 U21636 ( .C1(n19480), .C2(n19522), .A(n19479), .B(n19478), .ZN(
        P3_U2916) );
  AOI22_X1 U21637 ( .A1(n19494), .A2(n19514), .B1(n19481), .B2(n19512), .ZN(
        n19485) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19483), .B1(
        n19482), .B2(n19517), .ZN(n19484) );
  OAI211_X1 U21639 ( .C1(n19491), .C2(n19522), .A(n19485), .B(n19484), .ZN(
        P3_U2908) );
  AOI22_X1 U21640 ( .A1(n19507), .A2(n19498), .B1(n19486), .B2(n19512), .ZN(
        n19490) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19517), .ZN(n19489) );
  OAI211_X1 U21642 ( .C1(n19491), .C2(n19503), .A(n19490), .B(n19489), .ZN(
        P3_U2900) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19512), .ZN(n19496) );
  AOI22_X1 U21644 ( .A1(n19494), .A2(n19517), .B1(n19507), .B2(n19514), .ZN(
        n19495) );
  OAI211_X1 U21645 ( .C1(n19504), .C2(n19522), .A(n19496), .B(n19495), .ZN(
        P3_U2892) );
  AOI22_X1 U21646 ( .A1(n19506), .A2(n19498), .B1(n19497), .B2(n19512), .ZN(
        n19502) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19517), .ZN(n19501) );
  OAI211_X1 U21648 ( .C1(n19504), .C2(n19503), .A(n19502), .B(n19501), .ZN(
        P3_U2884) );
  AOI22_X1 U21649 ( .A1(n19506), .A2(n19514), .B1(n19505), .B2(n19512), .ZN(
        n19510) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19508), .B1(
        n19507), .B2(n19517), .ZN(n19509) );
  OAI211_X1 U21651 ( .C1(n19511), .C2(n19522), .A(n19510), .B(n19509), .ZN(
        P3_U2876) );
  AOI22_X1 U21652 ( .A1(n19515), .A2(n19514), .B1(n19513), .B2(n19512), .ZN(
        n19521) );
  INV_X1 U21653 ( .A(n19516), .ZN(n19519) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19519), .B1(
        n19518), .B2(n19517), .ZN(n19520) );
  OAI211_X1 U21655 ( .C1(n19523), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P3_U2868) );
  AOI22_X1 U21656 ( .A1(n19524), .A2(n19822), .B1(BUF2_REG_31__SCAN_IN), .B2(
        n19909), .ZN(n19526) );
  AOI22_X1 U21657 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19905), .B1(n19908), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19525) );
  NAND2_X1 U21658 ( .A1(n19526), .A2(n19525), .ZN(P2_U2888) );
  NOR2_X2 U21659 ( .A1(n19527), .A2(n20005), .ZN(n19720) );
  NOR2_X2 U21660 ( .A1(n19528), .A2(n20007), .ZN(n19706) );
  AOI22_X1 U21661 ( .A1(n20009), .A2(n19720), .B1(n20008), .B2(n19706), .ZN(
        n19531) );
  INV_X1 U21662 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22638) );
  OAI22_X2 U21663 ( .A1(n19529), .A2(n19961), .B1(n22638), .B2(n19960), .ZN(
        n19707) );
  AOI22_X1 U21664 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20010), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20011), .ZN(n19723) );
  INV_X1 U21665 ( .A(n19723), .ZN(n19684) );
  AOI22_X1 U21666 ( .A1(n20109), .A2(n19707), .B1(n19966), .B2(n19684), .ZN(
        n19530) );
  OAI211_X1 U21667 ( .C1(n19533), .C2(n19532), .A(n19531), .B(n19530), .ZN(
        P2_U3175) );
  INV_X1 U21668 ( .A(n19707), .ZN(n19687) );
  NOR2_X1 U21669 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19534), .ZN(
        n20015) );
  AOI22_X1 U21670 ( .A1(n19684), .A2(n20016), .B1(n19706), .B2(n20015), .ZN(
        n19543) );
  NAND2_X1 U21671 ( .A1(n20021), .A2(n19708), .ZN(n19535) );
  OAI21_X1 U21672 ( .B1(n19535), .B2(n20016), .A(n19709), .ZN(n19539) );
  NOR3_X1 U21673 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19592), .A3(
        n19563), .ZN(n19548) );
  NAND2_X1 U21674 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19548), .ZN(
        n19538) );
  INV_X1 U21675 ( .A(n19648), .ZN(n19711) );
  AOI21_X1 U21676 ( .B1(n12549), .B2(n19712), .A(n19711), .ZN(n19536) );
  AOI21_X1 U21677 ( .B1(n19539), .B2(n19538), .A(n19536), .ZN(n19537) );
  INV_X1 U21678 ( .A(n19538), .ZN(n20022) );
  OAI21_X1 U21679 ( .B1(n20015), .B2(n20022), .A(n19539), .ZN(n19541) );
  OAI21_X1 U21680 ( .B1(n12549), .B2(n20015), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19540) );
  NAND2_X1 U21681 ( .A1(n19541), .A2(n19540), .ZN(n20017) );
  AOI22_X1 U21682 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20018), .B1(
        n19720), .B2(n20017), .ZN(n19542) );
  OAI211_X1 U21683 ( .C1(n19687), .C2(n20021), .A(n19543), .B(n19542), .ZN(
        P2_U3167) );
  INV_X1 U21684 ( .A(n19548), .ZN(n19558) );
  INV_X1 U21685 ( .A(n12550), .ZN(n19544) );
  OAI21_X1 U21686 ( .B1(n19544), .B2(n20022), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19545) );
  OAI21_X1 U21687 ( .B1(n19558), .B2(n19694), .A(n19545), .ZN(n20023) );
  AOI22_X1 U21688 ( .A1(n20023), .A2(n19720), .B1(n19706), .B2(n20022), .ZN(
        n19554) );
  OR2_X1 U21689 ( .A1(n19551), .A2(n22141), .ZN(n19696) );
  NOR2_X1 U21690 ( .A1(n19552), .A2(n19696), .ZN(n19549) );
  OAI21_X1 U21691 ( .B1(n19708), .B2(n20022), .A(n19715), .ZN(n19546) );
  OAI21_X1 U21692 ( .B1(n12550), .B2(n19699), .A(n19546), .ZN(n19547) );
  OAI21_X1 U21693 ( .B1(n19549), .B2(n19548), .A(n19547), .ZN(n20024) );
  NOR2_X2 U21694 ( .A1(n19552), .A2(n19633), .ZN(n20030) );
  AOI22_X1 U21695 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19684), .ZN(n19553) );
  OAI211_X1 U21696 ( .C1(n19687), .C2(n20027), .A(n19554), .B(n19553), .ZN(
        P2_U3159) );
  NOR2_X1 U21697 ( .A1(n19643), .A2(n19581), .ZN(n19561) );
  INV_X1 U21698 ( .A(n19555), .ZN(n19560) );
  INV_X1 U21699 ( .A(n19556), .ZN(n19557) );
  NAND2_X1 U21700 ( .A1(n19557), .A2(n19614), .ZN(n19647) );
  NOR2_X1 U21701 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19558), .ZN(
        n20028) );
  OAI21_X1 U21702 ( .B1(n12538), .B2(n20028), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19559) );
  OAI21_X1 U21703 ( .B1(n19560), .B2(n19647), .A(n19559), .ZN(n20029) );
  AOI22_X1 U21704 ( .A1(n20029), .A2(n19720), .B1(n19706), .B2(n20028), .ZN(
        n19569) );
  OAI21_X1 U21705 ( .B1(n19561), .B2(n20030), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19562) );
  OAI21_X1 U21706 ( .B1(n19647), .B2(n19563), .A(n19562), .ZN(n19567) );
  INV_X1 U21707 ( .A(n12538), .ZN(n19565) );
  OAI21_X1 U21708 ( .B1(n19708), .B2(n20028), .A(n19715), .ZN(n19564) );
  OAI21_X1 U21709 ( .B1(n19565), .B2(n19699), .A(n19564), .ZN(n19566) );
  NAND2_X1 U21710 ( .A1(n19567), .A2(n19566), .ZN(n20031) );
  AOI22_X1 U21711 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20030), .B2(n19707), .ZN(n19568) );
  OAI211_X1 U21712 ( .C1(n19723), .C2(n20039), .A(n19569), .B(n19568), .ZN(
        P2_U3151) );
  NOR2_X1 U21713 ( .A1(n19612), .A2(n19572), .ZN(n20034) );
  NOR2_X1 U21714 ( .A1(n12539), .A2(n20034), .ZN(n19571) );
  OAI22_X1 U21715 ( .A1(n19571), .A2(n19594), .B1(n19572), .B2(n19694), .ZN(
        n20035) );
  AOI22_X1 U21716 ( .A1(n20035), .A2(n19720), .B1(n19706), .B2(n20034), .ZN(
        n19577) );
  INV_X1 U21717 ( .A(n20034), .ZN(n19570) );
  OAI22_X1 U21718 ( .A1(n19571), .A2(n19699), .B1(n20005), .B2(n19570), .ZN(
        n19575) );
  OAI21_X1 U21719 ( .B1(n19573), .B2(n19661), .A(n19572), .ZN(n19574) );
  OAI21_X1 U21720 ( .B1(n19711), .B2(n19575), .A(n19574), .ZN(n20036) );
  AOI22_X1 U21721 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19684), .ZN(n19576) );
  OAI211_X1 U21722 ( .C1(n19687), .C2(n20039), .A(n19577), .B(n19576), .ZN(
        P2_U3143) );
  INV_X1 U21723 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U21724 ( .A1(n19707), .A2(n20041), .B1(n20040), .B2(n19706), .ZN(
        n19579) );
  AOI22_X1 U21725 ( .A1(n19720), .A2(n20042), .B1(n20048), .B2(n19684), .ZN(
        n19578) );
  OAI211_X1 U21726 ( .C1(n20046), .C2(n19580), .A(n19579), .B(n19578), .ZN(
        P2_U3135) );
  INV_X1 U21727 ( .A(n20055), .ZN(n20053) );
  AOI22_X1 U21728 ( .A1(n19707), .A2(n20048), .B1(n20047), .B2(n19706), .ZN(
        n19589) );
  OAI21_X1 U21729 ( .B1(n19581), .B2(n19696), .A(n19708), .ZN(n19587) );
  INV_X1 U21730 ( .A(n19590), .ZN(n19584) );
  AOI21_X1 U21731 ( .B1(n20047), .B2(n19715), .A(n19711), .ZN(n19582) );
  OAI21_X1 U21732 ( .B1(n12551), .B2(n19699), .A(n19582), .ZN(n19583) );
  OAI21_X1 U21733 ( .B1(n19587), .B2(n19584), .A(n19583), .ZN(n20050) );
  OAI21_X1 U21734 ( .B1(n11183), .B2(n20047), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19586) );
  OAI21_X1 U21735 ( .B1(n19587), .B2(n19590), .A(n19586), .ZN(n20049) );
  AOI22_X1 U21736 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20050), .B1(
        n19720), .B2(n20049), .ZN(n19588) );
  OAI211_X1 U21737 ( .C1(n19723), .C2(n20053), .A(n19589), .B(n19588), .ZN(
        P2_U3127) );
  NOR2_X1 U21738 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19590), .ZN(
        n20054) );
  AOI22_X1 U21739 ( .A1(n19707), .A2(n20055), .B1(n20054), .B2(n19706), .ZN(
        n19602) );
  NAND2_X1 U21740 ( .A1(n20066), .A2(n19708), .ZN(n19591) );
  OAI21_X1 U21741 ( .B1(n19591), .B2(n20055), .A(n19709), .ZN(n19597) );
  NOR2_X1 U21742 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19592), .ZN(
        n19625) );
  INV_X1 U21743 ( .A(n19625), .ZN(n19626) );
  NOR2_X1 U21744 ( .A1(n19626), .A2(n19659), .ZN(n20060) );
  INV_X1 U21745 ( .A(n20060), .ZN(n19606) );
  INV_X1 U21746 ( .A(n12535), .ZN(n19598) );
  OAI21_X1 U21747 ( .B1(n19598), .B2(n19594), .A(n19593), .ZN(n19595) );
  AOI21_X1 U21748 ( .B1(n19597), .B2(n19606), .A(n19595), .ZN(n19596) );
  OAI21_X1 U21749 ( .B1(n20054), .B2(n19596), .A(n19715), .ZN(n20057) );
  OAI21_X1 U21750 ( .B1(n20060), .B2(n20054), .A(n19597), .ZN(n19600) );
  OAI21_X1 U21751 ( .B1(n19598), .B2(n20054), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19599) );
  NAND2_X1 U21752 ( .A1(n19600), .A2(n19599), .ZN(n20056) );
  AOI22_X1 U21753 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19720), .ZN(n19601) );
  OAI211_X1 U21754 ( .C1(n19723), .C2(n20066), .A(n19602), .B(n19601), .ZN(
        P2_U3119) );
  NAND2_X1 U21755 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19625), .ZN(
        n19604) );
  OAI21_X1 U21756 ( .B1(n12546), .B2(n20060), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19603) );
  OAI21_X1 U21757 ( .B1(n19604), .B2(n19694), .A(n19603), .ZN(n20061) );
  AOI22_X1 U21758 ( .A1(n20061), .A2(n19720), .B1(n20060), .B2(n19706), .ZN(
        n19611) );
  OAI22_X1 U21759 ( .A1(n19623), .A2(n19605), .B1(n19626), .B2(n19689), .ZN(
        n19609) );
  INV_X1 U21760 ( .A(n12546), .ZN(n19607) );
  OAI211_X1 U21761 ( .C1(n19607), .C2(n19699), .A(n19606), .B(n19694), .ZN(
        n19608) );
  NAND3_X1 U21762 ( .A1(n19609), .A2(n19715), .A3(n19608), .ZN(n20063) );
  AOI22_X1 U21763 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20063), .B1(
        n19980), .B2(n19707), .ZN(n19610) );
  OAI211_X1 U21764 ( .C1(n19723), .C2(n20073), .A(n19611), .B(n19610), .ZN(
        P2_U3111) );
  NAND2_X1 U21765 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19612), .ZN(
        n19671) );
  NOR2_X1 U21766 ( .A1(n19671), .A2(n19626), .ZN(n20067) );
  OAI21_X1 U21767 ( .B1(n19615), .B2(n20067), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19613) );
  OAI21_X1 U21768 ( .B1(n19626), .B2(n19672), .A(n19613), .ZN(n20068) );
  AOI22_X1 U21769 ( .A1(n20068), .A2(n19720), .B1(n19706), .B2(n20067), .ZN(
        n19622) );
  AOI21_X1 U21770 ( .B1(n20079), .B2(n20073), .A(n22141), .ZN(n19620) );
  NOR2_X1 U21771 ( .A1(n19626), .A2(n19614), .ZN(n19619) );
  INV_X1 U21772 ( .A(n20067), .ZN(n19617) );
  NAND2_X1 U21773 ( .A1(n19615), .A2(n19712), .ZN(n19616) );
  OAI211_X1 U21774 ( .C1(n20005), .C2(n19617), .A(n19616), .B(n19648), .ZN(
        n19618) );
  AOI22_X1 U21775 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n19684), .ZN(n19621) );
  OAI211_X1 U21776 ( .C1(n19687), .C2(n20073), .A(n19622), .B(n19621), .ZN(
        P2_U3103) );
  INV_X1 U21777 ( .A(n19623), .ZN(n19634) );
  INV_X1 U21778 ( .A(n19696), .ZN(n19624) );
  NAND2_X1 U21779 ( .A1(n19634), .A2(n19624), .ZN(n19636) );
  NAND2_X1 U21780 ( .A1(n19625), .A2(n19689), .ZN(n19645) );
  NAND2_X1 U21781 ( .A1(n19636), .A2(n19645), .ZN(n19632) );
  NAND2_X1 U21782 ( .A1(n12531), .A2(n19712), .ZN(n19630) );
  NAND2_X1 U21783 ( .A1(n19689), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19692) );
  NOR2_X1 U21784 ( .A1(n19692), .A2(n19626), .ZN(n20074) );
  INV_X1 U21785 ( .A(n20074), .ZN(n19627) );
  NAND2_X1 U21786 ( .A1(n19694), .A2(n19627), .ZN(n19628) );
  NAND2_X1 U21787 ( .A1(n19715), .A2(n19628), .ZN(n19629) );
  NAND2_X1 U21788 ( .A1(n19630), .A2(n19629), .ZN(n19631) );
  INV_X1 U21789 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19641) );
  INV_X1 U21790 ( .A(n19633), .ZN(n19688) );
  NAND2_X1 U21791 ( .A1(n19634), .A2(n19688), .ZN(n19943) );
  AOI22_X1 U21792 ( .A1(n19684), .A2(n20081), .B1(n19706), .B2(n20074), .ZN(
        n19640) );
  INV_X1 U21793 ( .A(n19645), .ZN(n19635) );
  NAND3_X1 U21794 ( .A1(n19636), .A2(n19708), .A3(n19635), .ZN(n19638) );
  OAI21_X1 U21795 ( .B1(n12531), .B2(n20074), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19637) );
  NAND2_X1 U21796 ( .A1(n19638), .A2(n19637), .ZN(n20075) );
  AOI22_X1 U21797 ( .A1(n19720), .A2(n20075), .B1(n20069), .B2(n19707), .ZN(
        n19639) );
  OAI211_X1 U21798 ( .C1(n19751), .C2(n19641), .A(n19640), .B(n19639), .ZN(
        P2_U3095) );
  INV_X1 U21799 ( .A(n19643), .ZN(n19644) );
  NOR2_X1 U21800 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19645), .ZN(
        n20080) );
  AOI22_X1 U21801 ( .A1(n19707), .A2(n20081), .B1(n20080), .B2(n19706), .ZN(
        n19656) );
  NOR2_X1 U21802 ( .A1(n20081), .A2(n20088), .ZN(n19646) );
  OAI21_X1 U21803 ( .B1(n19646), .B2(n22141), .A(n19708), .ZN(n19654) );
  NOR2_X1 U21804 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19647), .ZN(
        n19651) );
  AOI21_X1 U21805 ( .B1(n12545), .B2(n19712), .A(n20080), .ZN(n19649) );
  OAI21_X1 U21806 ( .B1(n19649), .B2(n20005), .A(n19648), .ZN(n19650) );
  INV_X1 U21807 ( .A(n19651), .ZN(n19653) );
  OAI21_X1 U21808 ( .B1(n12545), .B2(n20080), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19652) );
  AOI22_X1 U21809 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20083), .B1(
        n19720), .B2(n20082), .ZN(n19655) );
  OAI211_X1 U21810 ( .C1(n19723), .C2(n20086), .A(n19656), .B(n19655), .ZN(
        P2_U3087) );
  INV_X1 U21811 ( .A(n19657), .ZN(n19658) );
  INV_X1 U21812 ( .A(n20098), .ZN(n19889) );
  NOR2_X1 U21813 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19690) );
  INV_X1 U21814 ( .A(n19690), .ZN(n19691) );
  NOR2_X1 U21815 ( .A1(n19659), .A2(n19691), .ZN(n20087) );
  AOI22_X1 U21816 ( .A1(n19684), .A2(n19889), .B1(n20087), .B2(n19706), .ZN(
        n19670) );
  OAI21_X1 U21817 ( .B1(n19661), .B2(n19660), .A(n19708), .ZN(n19668) );
  NOR2_X1 U21818 ( .A1(n19689), .A2(n19691), .ZN(n19665) );
  INV_X1 U21819 ( .A(n12547), .ZN(n19663) );
  OAI21_X1 U21820 ( .B1(n19708), .B2(n20087), .A(n19715), .ZN(n19662) );
  OAI21_X1 U21821 ( .B1(n19663), .B2(n19699), .A(n19662), .ZN(n19664) );
  OAI21_X1 U21822 ( .B1(n19668), .B2(n19665), .A(n19664), .ZN(n20090) );
  INV_X1 U21823 ( .A(n19665), .ZN(n19667) );
  OAI21_X1 U21824 ( .B1(n12547), .B2(n20087), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19666) );
  OAI21_X1 U21825 ( .B1(n19668), .B2(n19667), .A(n19666), .ZN(n20089) );
  AOI22_X1 U21826 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20090), .B1(
        n19720), .B2(n20089), .ZN(n19669) );
  OAI211_X1 U21827 ( .C1(n19687), .C2(n20086), .A(n19670), .B(n19669), .ZN(
        P2_U3079) );
  NOR2_X1 U21828 ( .A1(n19671), .A2(n19691), .ZN(n20093) );
  OAI21_X1 U21829 ( .B1(n19678), .B2(n20093), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19674) );
  INV_X1 U21830 ( .A(n19672), .ZN(n19673) );
  NAND2_X1 U21831 ( .A1(n19673), .A2(n19690), .ZN(n19677) );
  NAND2_X1 U21832 ( .A1(n19674), .A2(n19677), .ZN(n20094) );
  AOI22_X1 U21833 ( .A1(n20094), .A2(n19720), .B1(n19706), .B2(n20093), .ZN(
        n19686) );
  INV_X1 U21834 ( .A(n19675), .ZN(n19676) );
  INV_X1 U21835 ( .A(n20102), .ZN(n19811) );
  OAI221_X1 U21836 ( .B1(n22141), .B2(n20098), .C1(n22141), .C2(n19811), .A(
        n19677), .ZN(n19682) );
  INV_X1 U21837 ( .A(n19678), .ZN(n19680) );
  INV_X1 U21838 ( .A(n20093), .ZN(n19679) );
  OAI21_X1 U21839 ( .B1(n19680), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19679), 
        .ZN(n19681) );
  MUX2_X1 U21840 ( .A(n19682), .B(n19681), .S(n19694), .Z(n19683) );
  NAND2_X1 U21841 ( .A1(n19683), .A2(n19715), .ZN(n20095) );
  AOI22_X1 U21842 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19684), .ZN(n19685) );
  OAI211_X1 U21843 ( .C1(n19687), .C2(n20098), .A(n19686), .B(n19685), .ZN(
        P2_U3071) );
  NAND2_X1 U21844 ( .A1(n19690), .A2(n19689), .ZN(n19705) );
  NOR2_X1 U21845 ( .A1(n19692), .A2(n19691), .ZN(n20099) );
  OAI21_X1 U21846 ( .B1(n12532), .B2(n20099), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19693) );
  OAI21_X1 U21847 ( .B1(n19705), .B2(n19694), .A(n19693), .ZN(n20100) );
  AOI22_X1 U21848 ( .A1(n20100), .A2(n19720), .B1(n19706), .B2(n20099), .ZN(
        n19704) );
  INV_X1 U21849 ( .A(n19695), .ZN(n19697) );
  OAI21_X1 U21850 ( .B1(n19697), .B2(n19696), .A(n19705), .ZN(n19702) );
  INV_X1 U21851 ( .A(n12532), .ZN(n19700) );
  OAI21_X1 U21852 ( .B1(n19708), .B2(n20099), .A(n19715), .ZN(n19698) );
  OAI21_X1 U21853 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19701) );
  NAND2_X1 U21854 ( .A1(n19702), .A2(n19701), .ZN(n20101) );
  AOI22_X1 U21855 ( .A1(n19707), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n20101), .ZN(n19703) );
  OAI211_X1 U21856 ( .C1(n19723), .C2(n20116), .A(n19704), .B(n19703), .ZN(
        P2_U3063) );
  INV_X1 U21857 ( .A(n20109), .ZN(n19921) );
  NOR2_X1 U21858 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19705), .ZN(
        n20108) );
  AOI22_X1 U21859 ( .A1(n19707), .A2(n19899), .B1(n20108), .B2(n19706), .ZN(
        n19722) );
  NAND2_X1 U21860 ( .A1(n20116), .A2(n19708), .ZN(n19710) );
  OAI21_X1 U21861 ( .B1(n19710), .B2(n20109), .A(n19709), .ZN(n19717) );
  AOI21_X1 U21862 ( .B1(n12544), .B2(n19712), .A(n19711), .ZN(n19713) );
  AOI21_X1 U21863 ( .B1(n19717), .B2(n19714), .A(n19713), .ZN(n19716) );
  OAI21_X1 U21864 ( .B1(n20108), .B2(n19716), .A(n19715), .ZN(n20113) );
  OAI21_X1 U21865 ( .B1(n20008), .B2(n20108), .A(n19717), .ZN(n19719) );
  OAI21_X1 U21866 ( .B1(n12544), .B2(n20108), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19718) );
  NAND2_X1 U21867 ( .A1(n19719), .A2(n19718), .ZN(n20112) );
  AOI22_X1 U21868 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20113), .B1(
        n19720), .B2(n20112), .ZN(n19721) );
  OAI211_X1 U21869 ( .C1(n19723), .C2(n19921), .A(n19722), .B(n19721), .ZN(
        P2_U3055) );
  INV_X1 U21870 ( .A(n19724), .ZN(n19725) );
  AOI22_X1 U21871 ( .A1(n19907), .A2(n19725), .B1(n19905), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U21872 ( .A1(n19909), .A2(BUF2_REG_22__SCAN_IN), .B1(n19908), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19730) );
  INV_X1 U21873 ( .A(n19726), .ZN(n19727) );
  AOI22_X1 U21874 ( .A1(n19728), .A2(n19822), .B1(n19821), .B2(n19727), .ZN(
        n19729) );
  NAND3_X1 U21875 ( .A1(n19731), .A2(n19730), .A3(n19729), .ZN(P2_U2897) );
  AOI22_X1 U21876 ( .A1(n20009), .A2(n19766), .B1(n20008), .B2(n19764), .ZN(
        n19734) );
  INV_X1 U21877 ( .A(n19769), .ZN(n19758) );
  AOI22_X1 U21878 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20012), .B1(
        n19966), .B2(n19758), .ZN(n19733) );
  OAI211_X1 U21879 ( .C1(n19761), .C2(n19921), .A(n19734), .B(n19733), .ZN(
        P2_U3174) );
  AOI22_X1 U21880 ( .A1(n19765), .A2(n19966), .B1(n19764), .B2(n20015), .ZN(
        n19736) );
  AOI22_X1 U21881 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20018), .B1(
        n19766), .B2(n20017), .ZN(n19735) );
  OAI211_X1 U21882 ( .C1(n19769), .C2(n20027), .A(n19736), .B(n19735), .ZN(
        P2_U3166) );
  AOI22_X1 U21883 ( .A1(n20023), .A2(n19766), .B1(n19764), .B2(n20022), .ZN(
        n19738) );
  AOI22_X1 U21884 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19758), .ZN(n19737) );
  OAI211_X1 U21885 ( .C1(n19761), .C2(n20027), .A(n19738), .B(n19737), .ZN(
        P2_U3158) );
  AOI22_X1 U21886 ( .A1(n20029), .A2(n19766), .B1(n19764), .B2(n20028), .ZN(
        n19740) );
  AOI22_X1 U21887 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20030), .B2(n19765), .ZN(n19739) );
  OAI211_X1 U21888 ( .C1(n19769), .C2(n20039), .A(n19740), .B(n19739), .ZN(
        P2_U3150) );
  AOI22_X1 U21889 ( .A1(n20035), .A2(n19766), .B1(n19764), .B2(n20034), .ZN(
        n19742) );
  AOI22_X1 U21890 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19758), .ZN(n19741) );
  OAI211_X1 U21891 ( .C1(n19761), .C2(n20039), .A(n19742), .B(n19741), .ZN(
        P2_U3142) );
  AOI22_X1 U21892 ( .A1(n19758), .A2(n20055), .B1(n19764), .B2(n20047), .ZN(
        n19744) );
  AOI22_X1 U21893 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20050), .B1(
        n19766), .B2(n20049), .ZN(n19743) );
  OAI211_X1 U21894 ( .C1(n19761), .C2(n19979), .A(n19744), .B(n19743), .ZN(
        P2_U3126) );
  AOI22_X1 U21895 ( .A1(n19758), .A2(n19980), .B1(n19764), .B2(n20054), .ZN(
        n19746) );
  AOI22_X1 U21896 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19766), .ZN(n19745) );
  OAI211_X1 U21897 ( .C1(n19761), .C2(n20053), .A(n19746), .B(n19745), .ZN(
        P2_U3118) );
  AOI22_X1 U21898 ( .A1(n20061), .A2(n19766), .B1(n19764), .B2(n20060), .ZN(
        n19748) );
  AOI22_X1 U21899 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20063), .B1(
        n19980), .B2(n19765), .ZN(n19747) );
  OAI211_X1 U21900 ( .C1(n19769), .C2(n20073), .A(n19748), .B(n19747), .ZN(
        P2_U3110) );
  AOI22_X1 U21901 ( .A1(n20068), .A2(n19766), .B1(n19764), .B2(n20067), .ZN(
        n19750) );
  AOI22_X1 U21902 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n19758), .ZN(n19749) );
  OAI211_X1 U21903 ( .C1(n19761), .C2(n20073), .A(n19750), .B(n19749), .ZN(
        P2_U3102) );
  AOI22_X1 U21904 ( .A1(n19765), .A2(n20069), .B1(n19764), .B2(n20074), .ZN(
        n19753) );
  AOI22_X1 U21905 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20076), .B1(
        n19766), .B2(n20075), .ZN(n19752) );
  OAI211_X1 U21906 ( .C1(n19769), .C2(n19943), .A(n19753), .B(n19752), .ZN(
        P2_U3094) );
  AOI22_X1 U21907 ( .A1(n19765), .A2(n20081), .B1(n19764), .B2(n20080), .ZN(
        n19755) );
  AOI22_X1 U21908 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20083), .B1(
        n19766), .B2(n20082), .ZN(n19754) );
  OAI211_X1 U21909 ( .C1(n19769), .C2(n20086), .A(n19755), .B(n19754), .ZN(
        P2_U3086) );
  AOI22_X1 U21910 ( .A1(n19758), .A2(n19889), .B1(n19764), .B2(n20087), .ZN(
        n19757) );
  AOI22_X1 U21911 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20090), .B1(
        n19766), .B2(n20089), .ZN(n19756) );
  OAI211_X1 U21912 ( .C1(n19761), .C2(n20086), .A(n19757), .B(n19756), .ZN(
        P2_U3078) );
  AOI22_X1 U21913 ( .A1(n20094), .A2(n19766), .B1(n19764), .B2(n20093), .ZN(
        n19760) );
  AOI22_X1 U21914 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19758), .ZN(n19759) );
  OAI211_X1 U21915 ( .C1(n19761), .C2(n20098), .A(n19760), .B(n19759), .ZN(
        P2_U3070) );
  AOI22_X1 U21916 ( .A1(n20100), .A2(n19766), .B1(n19764), .B2(n20099), .ZN(
        n19763) );
  AOI22_X1 U21917 ( .A1(n19765), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n20101), .ZN(n19762) );
  OAI211_X1 U21918 ( .C1(n19769), .C2(n20116), .A(n19763), .B(n19762), .ZN(
        P2_U3062) );
  AOI22_X1 U21919 ( .A1(n19765), .A2(n19899), .B1(n19764), .B2(n20108), .ZN(
        n19768) );
  AOI22_X1 U21920 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n19766), .ZN(n19767) );
  OAI211_X1 U21921 ( .C1(n19769), .C2(n19921), .A(n19768), .B(n19767), .ZN(
        P2_U3054) );
  OAI22_X1 U21922 ( .A1(n19773), .A2(n19772), .B1(n19771), .B2(n19770), .ZN(
        n19774) );
  INV_X1 U21923 ( .A(n19774), .ZN(n19779) );
  INV_X1 U21924 ( .A(n19775), .ZN(n19776) );
  NAND3_X1 U21925 ( .A1(n19777), .A2(n19776), .A3(n19821), .ZN(n19778) );
  OAI211_X1 U21926 ( .C1(n19781), .C2(n19780), .A(n19779), .B(n19778), .ZN(
        P2_U2914) );
  AOI22_X1 U21927 ( .A1(n19808), .A2(n20016), .B1(n19813), .B2(n20015), .ZN(
        n19783) );
  AOI22_X1 U21928 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20018), .B1(
        n19815), .B2(n20017), .ZN(n19782) );
  OAI211_X1 U21929 ( .C1(n19812), .C2(n20021), .A(n19783), .B(n19782), .ZN(
        P2_U3165) );
  AOI22_X1 U21930 ( .A1(n20023), .A2(n19815), .B1(n19813), .B2(n20022), .ZN(
        n19785) );
  AOI22_X1 U21931 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19808), .ZN(n19784) );
  OAI211_X1 U21932 ( .C1(n19812), .C2(n20027), .A(n19785), .B(n19784), .ZN(
        P2_U3157) );
  AOI22_X1 U21933 ( .A1(n20029), .A2(n19815), .B1(n19813), .B2(n20028), .ZN(
        n19787) );
  AOI22_X1 U21934 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20030), .B2(n19814), .ZN(n19786) );
  OAI211_X1 U21935 ( .C1(n19818), .C2(n20039), .A(n19787), .B(n19786), .ZN(
        P2_U3149) );
  AOI22_X1 U21936 ( .A1(n20035), .A2(n19815), .B1(n19813), .B2(n20034), .ZN(
        n19789) );
  AOI22_X1 U21937 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19808), .ZN(n19788) );
  OAI211_X1 U21938 ( .C1(n19812), .C2(n20039), .A(n19789), .B(n19788), .ZN(
        P2_U3141) );
  AOI22_X1 U21939 ( .A1(n19808), .A2(n20048), .B1(n20040), .B2(n19813), .ZN(
        n19791) );
  AOI22_X1 U21940 ( .A1(n19815), .A2(n20042), .B1(n20041), .B2(n19814), .ZN(
        n19790) );
  OAI211_X1 U21941 ( .C1(n20046), .C2(n12536), .A(n19791), .B(n19790), .ZN(
        P2_U3133) );
  AOI22_X1 U21942 ( .A1(n19808), .A2(n20055), .B1(n19813), .B2(n20047), .ZN(
        n19793) );
  AOI22_X1 U21943 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20050), .B1(
        n19815), .B2(n20049), .ZN(n19792) );
  OAI211_X1 U21944 ( .C1(n19812), .C2(n19979), .A(n19793), .B(n19792), .ZN(
        P2_U3125) );
  AOI22_X1 U21945 ( .A1(n19814), .A2(n20055), .B1(n19813), .B2(n20054), .ZN(
        n19795) );
  AOI22_X1 U21946 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19815), .ZN(n19794) );
  OAI211_X1 U21947 ( .C1(n19818), .C2(n20066), .A(n19795), .B(n19794), .ZN(
        P2_U3117) );
  AOI22_X1 U21948 ( .A1(n20061), .A2(n19815), .B1(n20060), .B2(n19813), .ZN(
        n19797) );
  AOI22_X1 U21949 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20063), .B1(
        n20062), .B2(n19808), .ZN(n19796) );
  OAI211_X1 U21950 ( .C1(n19812), .C2(n20066), .A(n19797), .B(n19796), .ZN(
        P2_U3109) );
  AOI22_X1 U21951 ( .A1(n20068), .A2(n19815), .B1(n19813), .B2(n20067), .ZN(
        n19799) );
  AOI22_X1 U21952 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n19808), .ZN(n19798) );
  OAI211_X1 U21953 ( .C1(n19812), .C2(n20073), .A(n19799), .B(n19798), .ZN(
        P2_U3101) );
  AOI22_X1 U21954 ( .A1(n19808), .A2(n20081), .B1(n19813), .B2(n20074), .ZN(
        n19801) );
  AOI22_X1 U21955 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20076), .B1(
        n19815), .B2(n20075), .ZN(n19800) );
  OAI211_X1 U21956 ( .C1(n19812), .C2(n20079), .A(n19801), .B(n19800), .ZN(
        P2_U3093) );
  AOI22_X1 U21957 ( .A1(n19814), .A2(n20081), .B1(n19813), .B2(n20080), .ZN(
        n19803) );
  AOI22_X1 U21958 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20083), .B1(
        n19815), .B2(n20082), .ZN(n19802) );
  OAI211_X1 U21959 ( .C1(n19818), .C2(n20086), .A(n19803), .B(n19802), .ZN(
        P2_U3085) );
  AOI22_X1 U21960 ( .A1(n19814), .A2(n20088), .B1(n19813), .B2(n20087), .ZN(
        n19805) );
  AOI22_X1 U21961 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20090), .B1(
        n19815), .B2(n20089), .ZN(n19804) );
  OAI211_X1 U21962 ( .C1(n19818), .C2(n20098), .A(n19805), .B(n19804), .ZN(
        P2_U3077) );
  AOI22_X1 U21963 ( .A1(n20094), .A2(n19815), .B1(n19813), .B2(n20093), .ZN(
        n19807) );
  AOI22_X1 U21964 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19808), .ZN(n19806) );
  OAI211_X1 U21965 ( .C1(n19812), .C2(n20098), .A(n19807), .B(n19806), .ZN(
        P2_U3069) );
  AOI22_X1 U21966 ( .A1(n20100), .A2(n19815), .B1(n19813), .B2(n20099), .ZN(
        n19810) );
  AOI22_X1 U21967 ( .A1(n19808), .A2(n19899), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n20101), .ZN(n19809) );
  OAI211_X1 U21968 ( .C1(n19812), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        P2_U3061) );
  AOI22_X1 U21969 ( .A1(n19814), .A2(n19899), .B1(n19813), .B2(n20108), .ZN(
        n19817) );
  AOI22_X1 U21970 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n19815), .ZN(n19816) );
  OAI211_X1 U21971 ( .C1(n19818), .C2(n19921), .A(n19817), .B(n19816), .ZN(
        P2_U3053) );
  INV_X1 U21972 ( .A(n19827), .ZN(n19819) );
  AOI22_X1 U21973 ( .A1(n19907), .A2(n19819), .B1(n19905), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U21974 ( .A1(n19909), .A2(BUF2_REG_20__SCAN_IN), .B1(n19908), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U21975 ( .A1(n19823), .A2(n19822), .B1(n19821), .B2(n19820), .ZN(
        n19824) );
  NAND3_X1 U21976 ( .A1(n19826), .A2(n19825), .A3(n19824), .ZN(P2_U2899) );
  AOI22_X1 U21977 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_20__SCAN_IN), .B2(n20010), .ZN(n19866) );
  NOR2_X2 U21978 ( .A1(n19827), .A2(n20005), .ZN(n19863) );
  NOR2_X2 U21979 ( .A1(n19828), .A2(n20007), .ZN(n19861) );
  AOI22_X1 U21980 ( .A1(n20009), .A2(n19863), .B1(n20008), .B2(n19861), .ZN(
        n19830) );
  INV_X1 U21981 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20450) );
  OAI22_X1 U21982 ( .A1(n21092), .A2(n19961), .B1(n20450), .B2(n19960), .ZN(
        n19862) );
  AOI22_X1 U21983 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20012), .B1(
        n19966), .B2(n19862), .ZN(n19829) );
  OAI211_X1 U21984 ( .C1(n19866), .C2(n19921), .A(n19830), .B(n19829), .ZN(
        P2_U3172) );
  INV_X1 U21985 ( .A(n19862), .ZN(n19860) );
  INV_X1 U21986 ( .A(n19866), .ZN(n19857) );
  AOI22_X1 U21987 ( .A1(n19857), .A2(n19966), .B1(n19861), .B2(n20015), .ZN(
        n19832) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20018), .B1(
        n19863), .B2(n20017), .ZN(n19831) );
  OAI211_X1 U21989 ( .C1(n19860), .C2(n20027), .A(n19832), .B(n19831), .ZN(
        P2_U3164) );
  AOI22_X1 U21990 ( .A1(n20023), .A2(n19863), .B1(n19861), .B2(n20022), .ZN(
        n19834) );
  AOI22_X1 U21991 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19862), .ZN(n19833) );
  OAI211_X1 U21992 ( .C1(n19866), .C2(n20027), .A(n19834), .B(n19833), .ZN(
        P2_U3156) );
  AOI22_X1 U21993 ( .A1(n20029), .A2(n19863), .B1(n19861), .B2(n20028), .ZN(
        n19836) );
  AOI22_X1 U21994 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20030), .B2(n19857), .ZN(n19835) );
  OAI211_X1 U21995 ( .C1(n19860), .C2(n20039), .A(n19836), .B(n19835), .ZN(
        P2_U3148) );
  AOI22_X1 U21996 ( .A1(n20035), .A2(n19863), .B1(n19861), .B2(n20034), .ZN(
        n19838) );
  AOI22_X1 U21997 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19862), .ZN(n19837) );
  OAI211_X1 U21998 ( .C1(n19866), .C2(n20039), .A(n19838), .B(n19837), .ZN(
        P2_U3140) );
  AOI22_X1 U21999 ( .A1(n19857), .A2(n20041), .B1(n20040), .B2(n19861), .ZN(
        n19840) );
  AOI22_X1 U22000 ( .A1(n19863), .A2(n20042), .B1(n20048), .B2(n19862), .ZN(
        n19839) );
  OAI211_X1 U22001 ( .C1(n20046), .C2(n12189), .A(n19840), .B(n19839), .ZN(
        P2_U3132) );
  AOI22_X1 U22002 ( .A1(n19862), .A2(n20055), .B1(n19861), .B2(n20047), .ZN(
        n19842) );
  AOI22_X1 U22003 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20050), .B1(
        n19863), .B2(n20049), .ZN(n19841) );
  OAI211_X1 U22004 ( .C1(n19866), .C2(n19979), .A(n19842), .B(n19841), .ZN(
        P2_U3124) );
  AOI22_X1 U22005 ( .A1(n19862), .A2(n19980), .B1(n20054), .B2(n19861), .ZN(
        n19844) );
  AOI22_X1 U22006 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19863), .ZN(n19843) );
  OAI211_X1 U22007 ( .C1(n19866), .C2(n20053), .A(n19844), .B(n19843), .ZN(
        P2_U3116) );
  AOI22_X1 U22008 ( .A1(n20061), .A2(n19863), .B1(n20060), .B2(n19861), .ZN(
        n19846) );
  AOI22_X1 U22009 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20063), .B1(
        n19980), .B2(n19857), .ZN(n19845) );
  OAI211_X1 U22010 ( .C1(n19860), .C2(n20073), .A(n19846), .B(n19845), .ZN(
        P2_U3108) );
  AOI22_X1 U22011 ( .A1(n20068), .A2(n19863), .B1(n19861), .B2(n20067), .ZN(
        n19848) );
  AOI22_X1 U22012 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n19862), .ZN(n19847) );
  OAI211_X1 U22013 ( .C1(n19866), .C2(n20073), .A(n19848), .B(n19847), .ZN(
        P2_U3100) );
  AOI22_X1 U22014 ( .A1(n19857), .A2(n20069), .B1(n19861), .B2(n20074), .ZN(
        n19850) );
  AOI22_X1 U22015 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20076), .B1(
        n19863), .B2(n20075), .ZN(n19849) );
  OAI211_X1 U22016 ( .C1(n19860), .C2(n19943), .A(n19850), .B(n19849), .ZN(
        P2_U3092) );
  AOI22_X1 U22017 ( .A1(n19857), .A2(n20081), .B1(n20080), .B2(n19861), .ZN(
        n19852) );
  AOI22_X1 U22018 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20083), .B1(
        n19863), .B2(n20082), .ZN(n19851) );
  OAI211_X1 U22019 ( .C1(n19860), .C2(n20086), .A(n19852), .B(n19851), .ZN(
        P2_U3084) );
  AOI22_X1 U22020 ( .A1(n19857), .A2(n20088), .B1(n20087), .B2(n19861), .ZN(
        n19854) );
  AOI22_X1 U22021 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20090), .B1(
        n19863), .B2(n20089), .ZN(n19853) );
  OAI211_X1 U22022 ( .C1(n19860), .C2(n20098), .A(n19854), .B(n19853), .ZN(
        P2_U3076) );
  AOI22_X1 U22023 ( .A1(n20094), .A2(n19863), .B1(n19861), .B2(n20093), .ZN(
        n19856) );
  AOI22_X1 U22024 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19862), .ZN(n19855) );
  OAI211_X1 U22025 ( .C1(n19866), .C2(n20098), .A(n19856), .B(n19855), .ZN(
        P2_U3068) );
  AOI22_X1 U22026 ( .A1(n20100), .A2(n19863), .B1(n19861), .B2(n20099), .ZN(
        n19859) );
  AOI22_X1 U22027 ( .A1(n19857), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n20101), .ZN(n19858) );
  OAI211_X1 U22028 ( .C1(n19860), .C2(n20116), .A(n19859), .B(n19858), .ZN(
        P2_U3060) );
  AOI22_X1 U22029 ( .A1(n19862), .A2(n20109), .B1(n20108), .B2(n19861), .ZN(
        n19865) );
  AOI22_X1 U22030 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n19863), .ZN(n19864) );
  OAI211_X1 U22031 ( .C1(n19866), .C2(n20116), .A(n19865), .B(n19864), .ZN(
        P2_U3052) );
  AOI22_X1 U22032 ( .A1(n19900), .A2(n19966), .B1(n20015), .B2(n19898), .ZN(
        n19868) );
  AOI22_X1 U22033 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20018), .B1(
        n19901), .B2(n20017), .ZN(n19867) );
  OAI211_X1 U22034 ( .C1(n19904), .C2(n20027), .A(n19868), .B(n19867), .ZN(
        P2_U3163) );
  AOI22_X1 U22035 ( .A1(n20023), .A2(n19901), .B1(n19898), .B2(n20022), .ZN(
        n19870) );
  AOI22_X1 U22036 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19892), .ZN(n19869) );
  OAI211_X1 U22037 ( .C1(n19895), .C2(n20027), .A(n19870), .B(n19869), .ZN(
        P2_U3155) );
  AOI22_X1 U22038 ( .A1(n20029), .A2(n19901), .B1(n19898), .B2(n20028), .ZN(
        n19872) );
  AOI22_X1 U22039 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20030), .B2(n19900), .ZN(n19871) );
  OAI211_X1 U22040 ( .C1(n19904), .C2(n20039), .A(n19872), .B(n19871), .ZN(
        P2_U3147) );
  AOI22_X1 U22041 ( .A1(n20035), .A2(n19901), .B1(n19898), .B2(n20034), .ZN(
        n19874) );
  AOI22_X1 U22042 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19892), .ZN(n19873) );
  OAI211_X1 U22043 ( .C1(n19895), .C2(n20039), .A(n19874), .B(n19873), .ZN(
        P2_U3139) );
  AOI22_X1 U22044 ( .A1(n19900), .A2(n20041), .B1(n20040), .B2(n19898), .ZN(
        n19876) );
  AOI22_X1 U22045 ( .A1(n19901), .A2(n20042), .B1(n20048), .B2(n19892), .ZN(
        n19875) );
  OAI211_X1 U22046 ( .C1(n20046), .C2(n12480), .A(n19876), .B(n19875), .ZN(
        P2_U3131) );
  AOI22_X1 U22047 ( .A1(n19892), .A2(n20055), .B1(n20047), .B2(n19898), .ZN(
        n19878) );
  AOI22_X1 U22048 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20050), .B1(
        n19901), .B2(n20049), .ZN(n19877) );
  OAI211_X1 U22049 ( .C1(n19895), .C2(n19979), .A(n19878), .B(n19877), .ZN(
        P2_U3123) );
  AOI22_X1 U22050 ( .A1(n19900), .A2(n20055), .B1(n20054), .B2(n19898), .ZN(
        n19880) );
  AOI22_X1 U22051 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19901), .ZN(n19879) );
  OAI211_X1 U22052 ( .C1(n19904), .C2(n20066), .A(n19880), .B(n19879), .ZN(
        P2_U3115) );
  AOI22_X1 U22053 ( .A1(n20061), .A2(n19901), .B1(n20060), .B2(n19898), .ZN(
        n19882) );
  AOI22_X1 U22054 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20063), .B1(
        n20062), .B2(n19892), .ZN(n19881) );
  OAI211_X1 U22055 ( .C1(n19895), .C2(n20066), .A(n19882), .B(n19881), .ZN(
        P2_U3107) );
  AOI22_X1 U22056 ( .A1(n20068), .A2(n19901), .B1(n19898), .B2(n20067), .ZN(
        n19884) );
  AOI22_X1 U22057 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20070), .B1(
        n20062), .B2(n19900), .ZN(n19883) );
  OAI211_X1 U22058 ( .C1(n19904), .C2(n20079), .A(n19884), .B(n19883), .ZN(
        P2_U3099) );
  AOI22_X1 U22059 ( .A1(n19892), .A2(n20081), .B1(n20074), .B2(n19898), .ZN(
        n19886) );
  AOI22_X1 U22060 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20076), .B1(
        n19901), .B2(n20075), .ZN(n19885) );
  OAI211_X1 U22061 ( .C1(n19895), .C2(n20079), .A(n19886), .B(n19885), .ZN(
        P2_U3091) );
  AOI22_X1 U22062 ( .A1(n19900), .A2(n20081), .B1(n20080), .B2(n19898), .ZN(
        n19888) );
  AOI22_X1 U22063 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20083), .B1(
        n19901), .B2(n20082), .ZN(n19887) );
  OAI211_X1 U22064 ( .C1(n19904), .C2(n20086), .A(n19888), .B(n19887), .ZN(
        P2_U3083) );
  AOI22_X1 U22065 ( .A1(n19892), .A2(n19889), .B1(n20087), .B2(n19898), .ZN(
        n19891) );
  AOI22_X1 U22066 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20090), .B1(
        n19901), .B2(n20089), .ZN(n19890) );
  OAI211_X1 U22067 ( .C1(n19895), .C2(n20086), .A(n19891), .B(n19890), .ZN(
        P2_U3075) );
  AOI22_X1 U22068 ( .A1(n20094), .A2(n19901), .B1(n19898), .B2(n20093), .ZN(
        n19894) );
  AOI22_X1 U22069 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19892), .ZN(n19893) );
  OAI211_X1 U22070 ( .C1(n19895), .C2(n20098), .A(n19894), .B(n19893), .ZN(
        P2_U3067) );
  AOI22_X1 U22071 ( .A1(n20100), .A2(n19901), .B1(n19898), .B2(n20099), .ZN(
        n19897) );
  AOI22_X1 U22072 ( .A1(n19900), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n20101), .ZN(n19896) );
  OAI211_X1 U22073 ( .C1(n19904), .C2(n20116), .A(n19897), .B(n19896), .ZN(
        P2_U3059) );
  AOI22_X1 U22074 ( .A1(n19900), .A2(n19899), .B1(n20108), .B2(n19898), .ZN(
        n19903) );
  AOI22_X1 U22075 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n19901), .ZN(n19902) );
  OAI211_X1 U22076 ( .C1(n19904), .C2(n19921), .A(n19903), .B(n19902), .ZN(
        P2_U3051) );
  INV_X1 U22077 ( .A(n19918), .ZN(n19906) );
  AOI22_X1 U22078 ( .A1(n19907), .A2(n19906), .B1(n19905), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U22079 ( .A1(n19909), .A2(BUF2_REG_18__SCAN_IN), .B1(n19908), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n19916) );
  OAI22_X1 U22080 ( .A1(n19913), .A2(n19912), .B1(n19911), .B2(n19910), .ZN(
        n19914) );
  INV_X1 U22081 ( .A(n19914), .ZN(n19915) );
  NAND3_X1 U22082 ( .A1(n19917), .A2(n19916), .A3(n19915), .ZN(P2_U2901) );
  AOI22_X1 U22083 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_18__SCAN_IN), .B2(n20010), .ZN(n19959) );
  NOR2_X2 U22084 ( .A1(n19918), .A2(n20005), .ZN(n19956) );
  NOR2_X2 U22085 ( .A1(n11877), .A2(n20007), .ZN(n19954) );
  AOI22_X1 U22086 ( .A1(n20009), .A2(n19956), .B1(n20008), .B2(n19954), .ZN(
        n19920) );
  OAI22_X1 U22087 ( .A1(n21074), .A2(n19961), .B1(n16644), .B2(n19960), .ZN(
        n19955) );
  AOI22_X1 U22088 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20012), .B1(
        n19966), .B2(n19955), .ZN(n19919) );
  OAI211_X1 U22089 ( .C1(n19959), .C2(n19921), .A(n19920), .B(n19919), .ZN(
        P2_U3170) );
  AOI22_X1 U22090 ( .A1(n19950), .A2(n19966), .B1(n19954), .B2(n20015), .ZN(
        n19923) );
  AOI22_X1 U22091 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20018), .B1(
        n19956), .B2(n20017), .ZN(n19922) );
  OAI211_X1 U22092 ( .C1(n19953), .C2(n20027), .A(n19923), .B(n19922), .ZN(
        P2_U3162) );
  AOI22_X1 U22093 ( .A1(n20023), .A2(n19956), .B1(n19954), .B2(n20022), .ZN(
        n19925) );
  AOI22_X1 U22094 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n19955), .ZN(n19924) );
  OAI211_X1 U22095 ( .C1(n19959), .C2(n20027), .A(n19925), .B(n19924), .ZN(
        P2_U3154) );
  AOI22_X1 U22096 ( .A1(n20029), .A2(n19956), .B1(n19954), .B2(n20028), .ZN(
        n19927) );
  AOI22_X1 U22097 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20030), .B2(n19950), .ZN(n19926) );
  OAI211_X1 U22098 ( .C1(n19953), .C2(n20039), .A(n19927), .B(n19926), .ZN(
        P2_U3146) );
  AOI22_X1 U22099 ( .A1(n20035), .A2(n19956), .B1(n19954), .B2(n20034), .ZN(
        n19929) );
  AOI22_X1 U22100 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n19955), .ZN(n19928) );
  OAI211_X1 U22101 ( .C1(n19959), .C2(n20039), .A(n19929), .B(n19928), .ZN(
        P2_U3138) );
  INV_X1 U22102 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U22103 ( .A1(n19955), .A2(n20048), .B1(n20040), .B2(n19954), .ZN(
        n19931) );
  AOI22_X1 U22104 ( .A1(n19956), .A2(n20042), .B1(n20041), .B2(n19950), .ZN(
        n19930) );
  OAI211_X1 U22105 ( .C1(n20046), .C2(n19932), .A(n19931), .B(n19930), .ZN(
        P2_U3130) );
  AOI22_X1 U22106 ( .A1(n19950), .A2(n20048), .B1(n19954), .B2(n20047), .ZN(
        n19934) );
  AOI22_X1 U22107 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20050), .B1(
        n19956), .B2(n20049), .ZN(n19933) );
  OAI211_X1 U22108 ( .C1(n19953), .C2(n20053), .A(n19934), .B(n19933), .ZN(
        P2_U3122) );
  AOI22_X1 U22109 ( .A1(n19955), .A2(n19980), .B1(n19954), .B2(n20054), .ZN(
        n19936) );
  AOI22_X1 U22110 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n19956), .ZN(n19935) );
  OAI211_X1 U22111 ( .C1(n19959), .C2(n20053), .A(n19936), .B(n19935), .ZN(
        P2_U3114) );
  AOI22_X1 U22112 ( .A1(n20061), .A2(n19956), .B1(n20060), .B2(n19954), .ZN(
        n19938) );
  AOI22_X1 U22113 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20063), .B1(
        n19980), .B2(n19950), .ZN(n19937) );
  OAI211_X1 U22114 ( .C1(n19953), .C2(n20073), .A(n19938), .B(n19937), .ZN(
        P2_U3106) );
  AOI22_X1 U22115 ( .A1(n20068), .A2(n19956), .B1(n19954), .B2(n20067), .ZN(
        n19940) );
  AOI22_X1 U22116 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20070), .B1(
        n20062), .B2(n19950), .ZN(n19939) );
  OAI211_X1 U22117 ( .C1(n19953), .C2(n20079), .A(n19940), .B(n19939), .ZN(
        P2_U3098) );
  AOI22_X1 U22118 ( .A1(n19950), .A2(n20069), .B1(n19954), .B2(n20074), .ZN(
        n19942) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20076), .B1(
        n19956), .B2(n20075), .ZN(n19941) );
  OAI211_X1 U22120 ( .C1(n19953), .C2(n19943), .A(n19942), .B(n19941), .ZN(
        P2_U3090) );
  AOI22_X1 U22121 ( .A1(n19950), .A2(n20081), .B1(n20080), .B2(n19954), .ZN(
        n19945) );
  AOI22_X1 U22122 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20083), .B1(
        n19956), .B2(n20082), .ZN(n19944) );
  OAI211_X1 U22123 ( .C1(n19953), .C2(n20086), .A(n19945), .B(n19944), .ZN(
        P2_U3082) );
  AOI22_X1 U22124 ( .A1(n19950), .A2(n20088), .B1(n20087), .B2(n19954), .ZN(
        n19947) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20090), .B1(
        n19956), .B2(n20089), .ZN(n19946) );
  OAI211_X1 U22126 ( .C1(n19953), .C2(n20098), .A(n19947), .B(n19946), .ZN(
        P2_U3074) );
  AOI22_X1 U22127 ( .A1(n20094), .A2(n19956), .B1(n19954), .B2(n20093), .ZN(
        n19949) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n19955), .ZN(n19948) );
  OAI211_X1 U22129 ( .C1(n19959), .C2(n20098), .A(n19949), .B(n19948), .ZN(
        P2_U3066) );
  AOI22_X1 U22130 ( .A1(n20100), .A2(n19956), .B1(n19954), .B2(n20099), .ZN(
        n19952) );
  AOI22_X1 U22131 ( .A1(n19950), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n20101), .ZN(n19951) );
  OAI211_X1 U22132 ( .C1(n19953), .C2(n20116), .A(n19952), .B(n19951), .ZN(
        P2_U3058) );
  AOI22_X1 U22133 ( .A1(n19955), .A2(n20109), .B1(n20108), .B2(n19954), .ZN(
        n19958) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n19956), .ZN(n19957) );
  OAI211_X1 U22135 ( .C1(n19959), .C2(n20116), .A(n19958), .B(n19957), .ZN(
        P2_U3050) );
  INV_X1 U22136 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n22387) );
  OAI22_X2 U22137 ( .A1(n19962), .A2(n19961), .B1(n22387), .B2(n19960), .ZN(
        n20000) );
  INV_X1 U22138 ( .A(n20000), .ZN(n19998) );
  NOR2_X2 U22139 ( .A1(n19963), .A2(n20005), .ZN(n20001) );
  NOR2_X2 U22140 ( .A1(n12609), .A2(n20007), .ZN(n19999) );
  AOI22_X1 U22141 ( .A1(n20009), .A2(n20001), .B1(n20008), .B2(n19999), .ZN(
        n19965) );
  AOI22_X1 U22142 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n20010), .ZN(n20004) );
  INV_X1 U22143 ( .A(n20004), .ZN(n19995) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20012), .B1(
        n20109), .B2(n19995), .ZN(n19964) );
  OAI211_X1 U22145 ( .C1(n19998), .C2(n20021), .A(n19965), .B(n19964), .ZN(
        P2_U3169) );
  AOI22_X1 U22146 ( .A1(n19995), .A2(n19966), .B1(n19999), .B2(n20015), .ZN(
        n19968) );
  AOI22_X1 U22147 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20018), .B1(
        n20001), .B2(n20017), .ZN(n19967) );
  OAI211_X1 U22148 ( .C1(n19998), .C2(n20027), .A(n19968), .B(n19967), .ZN(
        P2_U3161) );
  AOI22_X1 U22149 ( .A1(n20023), .A2(n20001), .B1(n19999), .B2(n20022), .ZN(
        n19970) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n20000), .ZN(n19969) );
  OAI211_X1 U22151 ( .C1(n20004), .C2(n20027), .A(n19970), .B(n19969), .ZN(
        P2_U3153) );
  AOI22_X1 U22152 ( .A1(n20029), .A2(n20001), .B1(n19999), .B2(n20028), .ZN(
        n19972) );
  AOI22_X1 U22153 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20030), .B2(n19995), .ZN(n19971) );
  OAI211_X1 U22154 ( .C1(n19998), .C2(n20039), .A(n19972), .B(n19971), .ZN(
        P2_U3145) );
  AOI22_X1 U22155 ( .A1(n20035), .A2(n20001), .B1(n19999), .B2(n20034), .ZN(
        n19974) );
  AOI22_X1 U22156 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n20000), .ZN(n19973) );
  OAI211_X1 U22157 ( .C1(n20004), .C2(n20039), .A(n19974), .B(n19973), .ZN(
        P2_U3137) );
  AOI22_X1 U22158 ( .A1(n20000), .A2(n20048), .B1(n20040), .B2(n19999), .ZN(
        n19976) );
  AOI22_X1 U22159 ( .A1(n20001), .A2(n20042), .B1(n20041), .B2(n19995), .ZN(
        n19975) );
  OAI211_X1 U22160 ( .C1(n20046), .C2(n12515), .A(n19976), .B(n19975), .ZN(
        P2_U3129) );
  AOI22_X1 U22161 ( .A1(n20000), .A2(n20055), .B1(n20047), .B2(n19999), .ZN(
        n19978) );
  AOI22_X1 U22162 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20050), .B1(
        n20001), .B2(n20049), .ZN(n19977) );
  OAI211_X1 U22163 ( .C1(n20004), .C2(n19979), .A(n19978), .B(n19977), .ZN(
        P2_U3121) );
  AOI22_X1 U22164 ( .A1(n20000), .A2(n19980), .B1(n20054), .B2(n19999), .ZN(
        n19982) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n20001), .ZN(n19981) );
  OAI211_X1 U22166 ( .C1(n20004), .C2(n20053), .A(n19982), .B(n19981), .ZN(
        P2_U3113) );
  AOI22_X1 U22167 ( .A1(n20061), .A2(n20001), .B1(n20060), .B2(n19999), .ZN(
        n19984) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20063), .B1(
        n20062), .B2(n20000), .ZN(n19983) );
  OAI211_X1 U22169 ( .C1(n20004), .C2(n20066), .A(n19984), .B(n19983), .ZN(
        P2_U3105) );
  AOI22_X1 U22170 ( .A1(n20068), .A2(n20001), .B1(n19999), .B2(n20067), .ZN(
        n19986) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n20000), .ZN(n19985) );
  OAI211_X1 U22172 ( .C1(n20004), .C2(n20073), .A(n19986), .B(n19985), .ZN(
        P2_U3097) );
  AOI22_X1 U22173 ( .A1(n20000), .A2(n20081), .B1(n19999), .B2(n20074), .ZN(
        n19988) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20076), .B1(
        n20001), .B2(n20075), .ZN(n19987) );
  OAI211_X1 U22175 ( .C1(n20004), .C2(n20079), .A(n19988), .B(n19987), .ZN(
        P2_U3089) );
  AOI22_X1 U22176 ( .A1(n19995), .A2(n20081), .B1(n20080), .B2(n19999), .ZN(
        n19990) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20083), .B1(
        n20001), .B2(n20082), .ZN(n19989) );
  OAI211_X1 U22178 ( .C1(n19998), .C2(n20086), .A(n19990), .B(n19989), .ZN(
        P2_U3081) );
  AOI22_X1 U22179 ( .A1(n19995), .A2(n20088), .B1(n20087), .B2(n19999), .ZN(
        n19992) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20090), .B1(
        n20001), .B2(n20089), .ZN(n19991) );
  OAI211_X1 U22181 ( .C1(n19998), .C2(n20098), .A(n19992), .B(n19991), .ZN(
        P2_U3073) );
  AOI22_X1 U22182 ( .A1(n20094), .A2(n20001), .B1(n19999), .B2(n20093), .ZN(
        n19994) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n20000), .ZN(n19993) );
  OAI211_X1 U22184 ( .C1(n20004), .C2(n20098), .A(n19994), .B(n19993), .ZN(
        P2_U3065) );
  AOI22_X1 U22185 ( .A1(n20100), .A2(n20001), .B1(n19999), .B2(n20099), .ZN(
        n19997) );
  AOI22_X1 U22186 ( .A1(n19995), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n20101), .ZN(n19996) );
  OAI211_X1 U22187 ( .C1(n19998), .C2(n20116), .A(n19997), .B(n19996), .ZN(
        P2_U3057) );
  AOI22_X1 U22188 ( .A1(n20000), .A2(n20109), .B1(n20108), .B2(n19999), .ZN(
        n20003) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20001), .ZN(n20002) );
  OAI211_X1 U22190 ( .C1(n20004), .C2(n20116), .A(n20003), .B(n20002), .ZN(
        P2_U3049) );
  AOI22_X1 U22191 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20010), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20011), .ZN(n20106) );
  NOR2_X2 U22192 ( .A1(n20006), .A2(n20005), .ZN(n20111) );
  NOR2_X2 U22193 ( .A1(n11861), .A2(n20007), .ZN(n20107) );
  AOI22_X1 U22194 ( .A1(n20009), .A2(n20111), .B1(n20008), .B2(n20107), .ZN(
        n20014) );
  AOI22_X1 U22195 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n20011), .B1(
        BUF1_REG_16__SCAN_IN), .B2(n20010), .ZN(n20117) );
  INV_X1 U22196 ( .A(n20117), .ZN(n20103) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20012), .B1(
        n20109), .B2(n20103), .ZN(n20013) );
  OAI211_X1 U22198 ( .C1(n20106), .C2(n20021), .A(n20014), .B(n20013), .ZN(
        P2_U3168) );
  INV_X1 U22199 ( .A(n20106), .ZN(n20110) );
  AOI22_X1 U22200 ( .A1(n20110), .A2(n20016), .B1(n20015), .B2(n20107), .ZN(
        n20020) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20018), .B1(
        n20111), .B2(n20017), .ZN(n20019) );
  OAI211_X1 U22202 ( .C1(n20117), .C2(n20021), .A(n20020), .B(n20019), .ZN(
        P2_U3160) );
  AOI22_X1 U22203 ( .A1(n20023), .A2(n20111), .B1(n20107), .B2(n20022), .ZN(
        n20026) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20024), .B1(
        n20030), .B2(n20110), .ZN(n20025) );
  OAI211_X1 U22205 ( .C1(n20117), .C2(n20027), .A(n20026), .B(n20025), .ZN(
        P2_U3152) );
  AOI22_X1 U22206 ( .A1(n20029), .A2(n20111), .B1(n20107), .B2(n20028), .ZN(
        n20033) );
  AOI22_X1 U22207 ( .A1(n20031), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20030), .B2(n20103), .ZN(n20032) );
  OAI211_X1 U22208 ( .C1(n20106), .C2(n20039), .A(n20033), .B(n20032), .ZN(
        P2_U3144) );
  AOI22_X1 U22209 ( .A1(n20035), .A2(n20111), .B1(n20107), .B2(n20034), .ZN(
        n20038) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20036), .B1(
        n20041), .B2(n20110), .ZN(n20037) );
  OAI211_X1 U22211 ( .C1(n20117), .C2(n20039), .A(n20038), .B(n20037), .ZN(
        P2_U3136) );
  INV_X1 U22212 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U22213 ( .A1(n20103), .A2(n20041), .B1(n20040), .B2(n20107), .ZN(
        n20044) );
  AOI22_X1 U22214 ( .A1(n20111), .A2(n20042), .B1(n20048), .B2(n20110), .ZN(
        n20043) );
  OAI211_X1 U22215 ( .C1(n20046), .C2(n20045), .A(n20044), .B(n20043), .ZN(
        P2_U3128) );
  AOI22_X1 U22216 ( .A1(n20103), .A2(n20048), .B1(n20047), .B2(n20107), .ZN(
        n20052) );
  AOI22_X1 U22217 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20050), .B1(
        n20111), .B2(n20049), .ZN(n20051) );
  OAI211_X1 U22218 ( .C1(n20106), .C2(n20053), .A(n20052), .B(n20051), .ZN(
        P2_U3120) );
  AOI22_X1 U22219 ( .A1(n20103), .A2(n20055), .B1(n20054), .B2(n20107), .ZN(
        n20059) );
  AOI22_X1 U22220 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20057), .B1(
        n20056), .B2(n20111), .ZN(n20058) );
  OAI211_X1 U22221 ( .C1(n20106), .C2(n20066), .A(n20059), .B(n20058), .ZN(
        P2_U3112) );
  AOI22_X1 U22222 ( .A1(n20061), .A2(n20111), .B1(n20060), .B2(n20107), .ZN(
        n20065) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20063), .B1(
        n20062), .B2(n20110), .ZN(n20064) );
  OAI211_X1 U22224 ( .C1(n20117), .C2(n20066), .A(n20065), .B(n20064), .ZN(
        P2_U3104) );
  AOI22_X1 U22225 ( .A1(n20068), .A2(n20111), .B1(n20107), .B2(n20067), .ZN(
        n20072) );
  AOI22_X1 U22226 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20070), .B1(
        n20069), .B2(n20110), .ZN(n20071) );
  OAI211_X1 U22227 ( .C1(n20117), .C2(n20073), .A(n20072), .B(n20071), .ZN(
        P2_U3096) );
  AOI22_X1 U22228 ( .A1(n20110), .A2(n20081), .B1(n20074), .B2(n20107), .ZN(
        n20078) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20076), .B1(
        n20111), .B2(n20075), .ZN(n20077) );
  OAI211_X1 U22230 ( .C1(n20117), .C2(n20079), .A(n20078), .B(n20077), .ZN(
        P2_U3088) );
  AOI22_X1 U22231 ( .A1(n20103), .A2(n20081), .B1(n20080), .B2(n20107), .ZN(
        n20085) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20083), .B1(
        n20111), .B2(n20082), .ZN(n20084) );
  OAI211_X1 U22233 ( .C1(n20106), .C2(n20086), .A(n20085), .B(n20084), .ZN(
        P2_U3080) );
  AOI22_X1 U22234 ( .A1(n20103), .A2(n20088), .B1(n20087), .B2(n20107), .ZN(
        n20092) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20090), .B1(
        n20111), .B2(n20089), .ZN(n20091) );
  OAI211_X1 U22236 ( .C1(n20106), .C2(n20098), .A(n20092), .B(n20091), .ZN(
        P2_U3072) );
  AOI22_X1 U22237 ( .A1(n20094), .A2(n20111), .B1(n20107), .B2(n20093), .ZN(
        n20097) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20095), .B1(
        n20102), .B2(n20110), .ZN(n20096) );
  OAI211_X1 U22239 ( .C1(n20117), .C2(n20098), .A(n20097), .B(n20096), .ZN(
        P2_U3064) );
  AOI22_X1 U22240 ( .A1(n20100), .A2(n20111), .B1(n20107), .B2(n20099), .ZN(
        n20105) );
  AOI22_X1 U22241 ( .A1(n20103), .A2(n20102), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n20101), .ZN(n20104) );
  OAI211_X1 U22242 ( .C1(n20106), .C2(n20116), .A(n20105), .B(n20104), .ZN(
        P2_U3056) );
  AOI22_X1 U22243 ( .A1(n20110), .A2(n20109), .B1(n20108), .B2(n20107), .ZN(
        n20115) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20113), .B1(
        n20112), .B2(n20111), .ZN(n20114) );
  OAI211_X1 U22245 ( .C1(n20117), .C2(n20116), .A(n20115), .B(n20114), .ZN(
        P2_U3048) );
  INV_X1 U22246 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20454) );
  INV_X1 U22247 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20118) );
  AOI222_X1 U22248 ( .A1(n20454), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20457), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n20118), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20119) );
  INV_X1 U22249 ( .A(n20179), .ZN(n20168) );
  AOI22_X1 U22250 ( .A1(n20168), .A2(n20121), .B1(n20120), .B2(n20179), .ZN(
        U376) );
  INV_X1 U22251 ( .A(n20179), .ZN(n20182) );
  AOI22_X1 U22252 ( .A1(n20182), .A2(n20123), .B1(n20122), .B2(n20179), .ZN(
        U365) );
  AOI22_X1 U22253 ( .A1(n20168), .A2(n20125), .B1(n20124), .B2(n20179), .ZN(
        U354) );
  INV_X1 U22254 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20127) );
  AOI22_X1 U22255 ( .A1(n20168), .A2(n20127), .B1(n20126), .B2(n20179), .ZN(
        U353) );
  INV_X1 U22256 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20129) );
  AOI22_X1 U22257 ( .A1(n20168), .A2(n20129), .B1(n20128), .B2(n20179), .ZN(
        U352) );
  INV_X1 U22258 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U22259 ( .A1(n20168), .A2(n20131), .B1(n20130), .B2(n20179), .ZN(
        U351) );
  INV_X1 U22260 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U22261 ( .A1(n20182), .A2(n20133), .B1(n20132), .B2(n20179), .ZN(
        U350) );
  AOI22_X1 U22262 ( .A1(n20168), .A2(n20135), .B1(n20134), .B2(n20179), .ZN(
        U349) );
  AOI22_X1 U22263 ( .A1(n20168), .A2(n20137), .B1(n20136), .B2(n20179), .ZN(
        U348) );
  AOI22_X1 U22264 ( .A1(n20168), .A2(n20139), .B1(n20138), .B2(n20179), .ZN(
        U347) );
  AOI22_X1 U22265 ( .A1(n20168), .A2(n20141), .B1(n20140), .B2(n20179), .ZN(
        U375) );
  AOI22_X1 U22266 ( .A1(n20168), .A2(n20143), .B1(n20142), .B2(n20179), .ZN(
        U374) );
  INV_X1 U22267 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U22268 ( .A1(n20168), .A2(n20145), .B1(n20144), .B2(n20179), .ZN(
        U373) );
  INV_X1 U22269 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U22270 ( .A1(n20168), .A2(n20147), .B1(n20146), .B2(n20179), .ZN(
        U372) );
  AOI22_X1 U22271 ( .A1(n20168), .A2(n20149), .B1(n20148), .B2(n20179), .ZN(
        U371) );
  AOI22_X1 U22272 ( .A1(n20168), .A2(n20151), .B1(n20150), .B2(n20179), .ZN(
        U370) );
  AOI22_X1 U22273 ( .A1(n20168), .A2(n20153), .B1(n20152), .B2(n20179), .ZN(
        U369) );
  AOI22_X1 U22274 ( .A1(n20168), .A2(n20155), .B1(n20154), .B2(n20179), .ZN(
        U368) );
  AOI22_X1 U22275 ( .A1(n20168), .A2(n20157), .B1(n20156), .B2(n20179), .ZN(
        U367) );
  AOI22_X1 U22276 ( .A1(n20168), .A2(n20159), .B1(n20158), .B2(n20179), .ZN(
        U366) );
  AOI22_X1 U22277 ( .A1(n20168), .A2(n20161), .B1(n20160), .B2(n20179), .ZN(
        U364) );
  AOI22_X1 U22278 ( .A1(n20168), .A2(n20163), .B1(n20162), .B2(n20179), .ZN(
        U363) );
  AOI22_X1 U22279 ( .A1(n20168), .A2(n20165), .B1(n20164), .B2(n20179), .ZN(
        U362) );
  AOI22_X1 U22280 ( .A1(n20168), .A2(n20167), .B1(n20166), .B2(n20179), .ZN(
        U361) );
  AOI22_X1 U22281 ( .A1(n20182), .A2(n20170), .B1(n20169), .B2(n20179), .ZN(
        U360) );
  AOI22_X1 U22282 ( .A1(n20182), .A2(n20172), .B1(n20171), .B2(n20179), .ZN(
        U359) );
  AOI22_X1 U22283 ( .A1(n20182), .A2(n20174), .B1(n20173), .B2(n20179), .ZN(
        U358) );
  AOI22_X1 U22284 ( .A1(n20182), .A2(n20176), .B1(n20175), .B2(n20179), .ZN(
        U357) );
  AOI22_X1 U22285 ( .A1(n20182), .A2(n20178), .B1(n20177), .B2(n20179), .ZN(
        U356) );
  AOI22_X1 U22286 ( .A1(n20182), .A2(n20181), .B1(n20180), .B2(n20179), .ZN(
        U355) );
  AOI22_X1 U22287 ( .A1(n21698), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20184) );
  OAI21_X1 U22288 ( .B1(n13256), .B2(n20210), .A(n20184), .ZN(P1_U2936) );
  AOI22_X1 U22289 ( .A1(n20194), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20185) );
  OAI21_X1 U22290 ( .B1(n13267), .B2(n20210), .A(n20185), .ZN(P1_U2935) );
  AOI22_X1 U22291 ( .A1(n20194), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20186) );
  OAI21_X1 U22292 ( .B1(n13250), .B2(n20210), .A(n20186), .ZN(P1_U2934) );
  AOI22_X1 U22293 ( .A1(n20194), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20187) );
  OAI21_X1 U22294 ( .B1(n14822), .B2(n20210), .A(n20187), .ZN(P1_U2933) );
  AOI22_X1 U22295 ( .A1(n20194), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20188) );
  OAI21_X1 U22296 ( .B1(n20189), .B2(n20210), .A(n20188), .ZN(P1_U2932) );
  AOI22_X1 U22297 ( .A1(n20194), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20190) );
  OAI21_X1 U22298 ( .B1(n20191), .B2(n20210), .A(n20190), .ZN(P1_U2931) );
  AOI22_X1 U22299 ( .A1(n20194), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20192) );
  OAI21_X1 U22300 ( .B1(n15092), .B2(n20210), .A(n20192), .ZN(P1_U2930) );
  AOI22_X1 U22301 ( .A1(n21698), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20193) );
  OAI21_X1 U22302 ( .B1(n15117), .B2(n20210), .A(n20193), .ZN(P1_U2929) );
  AOI22_X1 U22303 ( .A1(n20194), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20195) );
  OAI21_X1 U22304 ( .B1(n20196), .B2(n20210), .A(n20195), .ZN(P1_U2928) );
  AOI22_X1 U22305 ( .A1(n21698), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20197) );
  OAI21_X1 U22306 ( .B1(n20198), .B2(n20210), .A(n20197), .ZN(P1_U2927) );
  AOI22_X1 U22307 ( .A1(n21698), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20199), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20200) );
  OAI21_X1 U22308 ( .B1(n20201), .B2(n20210), .A(n20200), .ZN(P1_U2926) );
  AOI22_X1 U22309 ( .A1(n21698), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U22310 ( .B1(n15765), .B2(n20210), .A(n20202), .ZN(P1_U2925) );
  AOI22_X1 U22311 ( .A1(n21698), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20203) );
  OAI21_X1 U22312 ( .B1(n16280), .B2(n20210), .A(n20203), .ZN(P1_U2924) );
  AOI22_X1 U22313 ( .A1(n21698), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20204) );
  OAI21_X1 U22314 ( .B1(n20205), .B2(n20210), .A(n20204), .ZN(P1_U2923) );
  AOI22_X1 U22315 ( .A1(n21698), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20206) );
  OAI21_X1 U22316 ( .B1(n20207), .B2(n20210), .A(n20206), .ZN(P1_U2922) );
  AOI22_X1 U22317 ( .A1(n21698), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20208), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20209) );
  OAI21_X1 U22318 ( .B1(n20211), .B2(n20210), .A(n20209), .ZN(P1_U2921) );
  NAND2_X1 U22319 ( .A1(n20459), .A2(n20212), .ZN(n20251) );
  CLKBUF_X1 U22320 ( .A(n20251), .Z(n20256) );
  OAI222_X1 U22321 ( .A1(n20260), .A2(n20275), .B1(n20213), .B2(n20459), .C1(
        n20214), .C2(n20256), .ZN(P1_U3197) );
  INV_X1 U22322 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20217) );
  INV_X1 U22323 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20215) );
  OAI222_X1 U22324 ( .A1(n20251), .A2(n20217), .B1(n20215), .B2(n20459), .C1(
        n20214), .C2(n20260), .ZN(P1_U3198) );
  INV_X1 U22325 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20216) );
  INV_X1 U22326 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21943) );
  OAI222_X1 U22327 ( .A1(n20260), .A2(n20217), .B1(n20216), .B2(n20459), .C1(
        n21943), .C2(n20256), .ZN(P1_U3199) );
  INV_X1 U22328 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20218) );
  OAI222_X1 U22329 ( .A1(n20260), .A2(n21943), .B1(n20218), .B2(n20459), .C1(
        n21955), .C2(n20256), .ZN(P1_U3200) );
  INV_X1 U22330 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21971) );
  INV_X1 U22331 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20219) );
  OAI222_X1 U22332 ( .A1(n20256), .A2(n21971), .B1(n20219), .B2(n20459), .C1(
        n21955), .C2(n20260), .ZN(P1_U3201) );
  INV_X1 U22333 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20220) );
  OAI222_X1 U22334 ( .A1(n20260), .A2(n21971), .B1(n20220), .B2(n20459), .C1(
        n21977), .C2(n20256), .ZN(P1_U3202) );
  INV_X1 U22335 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20221) );
  OAI222_X1 U22336 ( .A1(n20256), .A2(n20223), .B1(n20221), .B2(n20459), .C1(
        n21977), .C2(n20260), .ZN(P1_U3203) );
  INV_X1 U22337 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20222) );
  OAI222_X1 U22338 ( .A1(n20260), .A2(n20223), .B1(n20222), .B2(n20459), .C1(
        n20225), .C2(n20251), .ZN(P1_U3204) );
  INV_X1 U22339 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20224) );
  OAI222_X1 U22340 ( .A1(n20260), .A2(n20225), .B1(n20224), .B2(n20459), .C1(
        n21813), .C2(n20251), .ZN(P1_U3205) );
  INV_X1 U22341 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20226) );
  INV_X1 U22342 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21840) );
  OAI222_X1 U22343 ( .A1(n20260), .A2(n21813), .B1(n20226), .B2(n20459), .C1(
        n21840), .C2(n20256), .ZN(P1_U3206) );
  INV_X1 U22344 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20227) );
  OAI222_X1 U22345 ( .A1(n20260), .A2(n21840), .B1(n20227), .B2(n20459), .C1(
        n21828), .C2(n20256), .ZN(P1_U3207) );
  INV_X1 U22346 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20228) );
  OAI222_X1 U22347 ( .A1(n20251), .A2(n21711), .B1(n20228), .B2(n20459), .C1(
        n21828), .C2(n20260), .ZN(P1_U3208) );
  INV_X1 U22348 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20229) );
  OAI222_X1 U22349 ( .A1(n20251), .A2(n21721), .B1(n20229), .B2(n20459), .C1(
        n21711), .C2(n20260), .ZN(P1_U3209) );
  INV_X1 U22350 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20230) );
  OAI222_X1 U22351 ( .A1(n20260), .A2(n21721), .B1(n20230), .B2(n20459), .C1(
        n20231), .C2(n20256), .ZN(P1_U3210) );
  INV_X1 U22352 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20232) );
  OAI222_X1 U22353 ( .A1(n20251), .A2(n21864), .B1(n20232), .B2(n20459), .C1(
        n20231), .C2(n20260), .ZN(P1_U3211) );
  INV_X1 U22354 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20233) );
  OAI222_X1 U22355 ( .A1(n20260), .A2(n21864), .B1(n20233), .B2(n20459), .C1(
        n20235), .C2(n20256), .ZN(P1_U3212) );
  INV_X1 U22356 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20234) );
  INV_X1 U22357 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20236) );
  OAI222_X1 U22358 ( .A1(n20260), .A2(n20235), .B1(n20234), .B2(n20459), .C1(
        n20236), .C2(n20256), .ZN(P1_U3213) );
  INV_X1 U22359 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n22038) );
  INV_X1 U22360 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20237) );
  OAI222_X1 U22361 ( .A1(n20251), .A2(n22038), .B1(n20237), .B2(n20459), .C1(
        n20236), .C2(n20260), .ZN(P1_U3214) );
  INV_X1 U22362 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20238) );
  OAI222_X1 U22363 ( .A1(n20251), .A2(n20239), .B1(n20238), .B2(n20459), .C1(
        n22038), .C2(n20260), .ZN(P1_U3215) );
  INV_X1 U22364 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20240) );
  OAI222_X1 U22365 ( .A1(n20251), .A2(n22072), .B1(n20240), .B2(n20459), .C1(
        n20239), .C2(n20260), .ZN(P1_U3216) );
  INV_X1 U22366 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20241) );
  OAI222_X1 U22367 ( .A1(n20260), .A2(n22072), .B1(n20241), .B2(n20459), .C1(
        n22075), .C2(n20256), .ZN(P1_U3217) );
  INV_X1 U22368 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20242) );
  OAI222_X1 U22369 ( .A1(n20260), .A2(n22075), .B1(n20242), .B2(n20459), .C1(
        n22086), .C2(n20256), .ZN(P1_U3218) );
  INV_X1 U22370 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20243) );
  OAI222_X1 U22371 ( .A1(n20260), .A2(n22086), .B1(n20243), .B2(n20459), .C1(
        n22103), .C2(n20256), .ZN(P1_U3219) );
  INV_X1 U22372 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20244) );
  OAI222_X1 U22373 ( .A1(n20260), .A2(n22103), .B1(n20244), .B2(n20459), .C1(
        n20246), .C2(n20256), .ZN(P1_U3220) );
  INV_X1 U22374 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20245) );
  OAI222_X1 U22375 ( .A1(n20260), .A2(n20246), .B1(n20245), .B2(n20459), .C1(
        n20248), .C2(n20256), .ZN(P1_U3221) );
  INV_X1 U22376 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20247) );
  OAI222_X1 U22377 ( .A1(n20260), .A2(n20248), .B1(n20247), .B2(n20459), .C1(
        n20249), .C2(n20256), .ZN(P1_U3222) );
  INV_X1 U22378 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20250) );
  OAI222_X1 U22379 ( .A1(n20251), .A2(n20252), .B1(n20250), .B2(n20459), .C1(
        n20249), .C2(n20260), .ZN(P1_U3223) );
  INV_X1 U22380 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20253) );
  OAI222_X1 U22381 ( .A1(n20256), .A2(n20255), .B1(n20253), .B2(n20459), .C1(
        n20252), .C2(n20260), .ZN(P1_U3224) );
  INV_X1 U22382 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20254) );
  OAI222_X1 U22383 ( .A1(n20260), .A2(n20255), .B1(n20254), .B2(n20459), .C1(
        n20259), .C2(n20256), .ZN(P1_U3225) );
  INV_X1 U22384 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20258) );
  OAI222_X1 U22385 ( .A1(n20260), .A2(n20259), .B1(n20258), .B2(n20459), .C1(
        n20257), .C2(n20256), .ZN(P1_U3226) );
  INV_X1 U22386 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20261) );
  AOI22_X1 U22387 ( .A1(n20459), .A2(n20262), .B1(n20261), .B2(n22749), .ZN(
        P1_U3458) );
  AOI221_X1 U22388 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20273) );
  NOR4_X1 U22389 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20266) );
  NOR4_X1 U22390 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20265) );
  NOR4_X1 U22391 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20264) );
  NOR4_X1 U22392 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20263) );
  NAND4_X1 U22393 ( .A1(n20266), .A2(n20265), .A3(n20264), .A4(n20263), .ZN(
        n20272) );
  NOR4_X1 U22394 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20270) );
  AOI211_X1 U22395 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20269) );
  NOR4_X1 U22396 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20268) );
  NOR4_X1 U22397 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20267) );
  NAND4_X1 U22398 ( .A1(n20270), .A2(n20269), .A3(n20268), .A4(n20267), .ZN(
        n20271) );
  NOR2_X1 U22399 ( .A1(n20272), .A2(n20271), .ZN(n20286) );
  MUX2_X1 U22400 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n20273), .S(n20286), 
        .Z(P1_U2808) );
  INV_X1 U22401 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20274) );
  AOI22_X1 U22402 ( .A1(n20459), .A2(n20278), .B1(n20274), .B2(n22749), .ZN(
        P1_U3459) );
  AOI21_X1 U22403 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20276) );
  OAI221_X1 U22404 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20276), .C1(n20275), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20286), .ZN(n20277) );
  OAI21_X1 U22405 ( .B1(n20286), .B2(n20278), .A(n20277), .ZN(P1_U3481) );
  INV_X1 U22406 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20282) );
  INV_X1 U22407 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20279) );
  AOI22_X1 U22408 ( .A1(n20459), .A2(n20282), .B1(n20279), .B2(n22749), .ZN(
        P1_U3460) );
  NOR3_X1 U22409 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20280) );
  OAI21_X1 U22410 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20280), .A(n20286), .ZN(
        n20281) );
  OAI21_X1 U22411 ( .B1(n20286), .B2(n20282), .A(n20281), .ZN(P1_U2807) );
  INV_X1 U22412 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20285) );
  INV_X1 U22413 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20283) );
  AOI22_X1 U22414 ( .A1(n20459), .A2(n20285), .B1(n20283), .B2(n22749), .ZN(
        P1_U3461) );
  OAI21_X1 U22415 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(n20286), .ZN(n20284) );
  OAI21_X1 U22416 ( .B1(n20286), .B2(n20285), .A(n20284), .ZN(P1_U3482) );
  INV_X1 U22417 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21990) );
  AOI21_X1 U22418 ( .B1(n20289), .B2(n20288), .A(n20287), .ZN(n21988) );
  AOI22_X1 U22419 ( .A1(n21992), .A2(n20323), .B1(n20322), .B2(n21988), .ZN(
        n20290) );
  OAI21_X1 U22420 ( .B1(n20326), .B2(n21990), .A(n20290), .ZN(P1_U2861) );
  AOI22_X1 U22421 ( .A1(n22214), .A2(n20323), .B1(n20322), .B2(n21859), .ZN(
        n20291) );
  OAI21_X1 U22422 ( .B1(n20326), .B2(n20292), .A(n20291), .ZN(P1_U2855) );
  AOI22_X1 U22423 ( .A1(n20367), .A2(n20323), .B1(n20322), .B2(n21843), .ZN(
        n20293) );
  OAI21_X1 U22424 ( .B1(n20326), .B2(n20294), .A(n20293), .ZN(P1_U2857) );
  AND2_X1 U22425 ( .A1(n20296), .A2(n20295), .ZN(n20298) );
  OAI21_X1 U22426 ( .B1(n16175), .B2(n20300), .A(n20299), .ZN(n20301) );
  INV_X1 U22427 ( .A(n20301), .ZN(n22092) );
  AOI22_X1 U22428 ( .A1(n11248), .A2(n20323), .B1(n20322), .B2(n22092), .ZN(
        n20302) );
  OAI21_X1 U22429 ( .B1(n20326), .B2(n22089), .A(n20302), .ZN(P1_U2849) );
  INV_X1 U22430 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n22063) );
  INV_X1 U22431 ( .A(n20303), .ZN(n22220) );
  AOI22_X1 U22432 ( .A1(n22220), .A2(n20323), .B1(n22065), .B2(n20322), .ZN(
        n20304) );
  OAI21_X1 U22433 ( .B1(n20326), .B2(n22063), .A(n20304), .ZN(P1_U2851) );
  INV_X1 U22434 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n22042) );
  AND2_X1 U22435 ( .A1(n20306), .A2(n20305), .ZN(n20307) );
  OR2_X1 U22436 ( .A1(n20309), .A2(n20308), .ZN(n20310) );
  AND2_X1 U22437 ( .A1(n20311), .A2(n20310), .ZN(n22045) );
  AOI22_X1 U22438 ( .A1(n22217), .A2(n20323), .B1(n20322), .B2(n22045), .ZN(
        n20312) );
  OAI21_X1 U22439 ( .B1(n20326), .B2(n22042), .A(n20312), .ZN(P1_U2853) );
  INV_X1 U22440 ( .A(n20321), .ZN(n20315) );
  INV_X1 U22441 ( .A(n20313), .ZN(n20314) );
  OAI21_X1 U22442 ( .B1(n14947), .B2(n20315), .A(n20314), .ZN(n20317) );
  AND2_X1 U22443 ( .A1(n20317), .A2(n20316), .ZN(n21949) );
  AOI22_X1 U22444 ( .A1(n21958), .A2(n20323), .B1(n20322), .B2(n21949), .ZN(
        n20318) );
  OAI21_X1 U22445 ( .B1(n20326), .B2(n20319), .A(n20318), .ZN(P1_U2867) );
  INV_X1 U22446 ( .A(n20320), .ZN(n21946) );
  XNOR2_X1 U22447 ( .A(n14947), .B(n20321), .ZN(n21937) );
  AOI22_X1 U22448 ( .A1(n21946), .A2(n20323), .B1(n20322), .B2(n21937), .ZN(
        n20324) );
  OAI21_X1 U22449 ( .B1(n20326), .B2(n20325), .A(n20324), .ZN(P1_U2868) );
  AOI22_X1 U22450 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20388), .ZN(n20332) );
  OAI21_X1 U22451 ( .B1(n20329), .B2(n20328), .A(n20327), .ZN(n20330) );
  INV_X1 U22452 ( .A(n20330), .ZN(n21750) );
  AOI22_X1 U22453 ( .A1(n21750), .A2(n20392), .B1(n20385), .B2(n21946), .ZN(
        n20331) );
  OAI211_X1 U22454 ( .C1(n20395), .C2(n21948), .A(n20332), .B(n20331), .ZN(
        P1_U2995) );
  AOI22_X1 U22455 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20388), .ZN(n20338) );
  OAI21_X1 U22456 ( .B1(n20335), .B2(n20334), .A(n20333), .ZN(n20336) );
  INV_X1 U22457 ( .A(n20336), .ZN(n21774) );
  AOI22_X1 U22458 ( .A1(n21774), .A2(n20392), .B1(n20385), .B2(n21958), .ZN(
        n20337) );
  OAI211_X1 U22459 ( .C1(n20395), .C2(n21960), .A(n20338), .B(n20337), .ZN(
        P1_U2994) );
  AOI22_X1 U22460 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20388), .ZN(n20345) );
  OR2_X1 U22461 ( .A1(n20340), .A2(n20339), .ZN(n20341) );
  NAND2_X1 U22462 ( .A1(n20342), .A2(n20341), .ZN(n21764) );
  INV_X1 U22463 ( .A(n21764), .ZN(n20343) );
  AOI22_X1 U22464 ( .A1(n20343), .A2(n20392), .B1(n20385), .B2(n21968), .ZN(
        n20344) );
  OAI211_X1 U22465 ( .C1(n20395), .C2(n21975), .A(n20345), .B(n20344), .ZN(
        P1_U2993) );
  AOI22_X1 U22466 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20388), .ZN(n20351) );
  OAI21_X1 U22467 ( .B1(n20348), .B2(n20347), .A(n20346), .ZN(n20349) );
  INV_X1 U22468 ( .A(n20349), .ZN(n21785) );
  AOI22_X1 U22469 ( .A1(n21785), .A2(n20392), .B1(n20385), .B2(n21983), .ZN(
        n20350) );
  OAI211_X1 U22470 ( .C1(n20395), .C2(n21986), .A(n20351), .B(n20350), .ZN(
        P1_U2992) );
  AOI22_X1 U22471 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20388), .ZN(n20358) );
  AOI21_X1 U22472 ( .B1(n20353), .B2(n16389), .A(n20352), .ZN(n20356) );
  MUX2_X1 U22473 ( .A(n20354), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .S(
        n13169), .Z(n20355) );
  XNOR2_X1 U22474 ( .A(n20356), .B(n20355), .ZN(n21834) );
  AOI22_X1 U22475 ( .A1(n20385), .A2(n21992), .B1(n20392), .B2(n21834), .ZN(
        n20357) );
  OAI211_X1 U22476 ( .C1(n20395), .C2(n21995), .A(n20358), .B(n20357), .ZN(
        P1_U2988) );
  AOI21_X1 U22477 ( .B1(n20361), .B2(n20360), .A(n20359), .ZN(n21833) );
  AOI22_X1 U22478 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20388), .ZN(n20363) );
  AOI22_X1 U22479 ( .A1(n20385), .A2(n21999), .B1(n20379), .B2(n22000), .ZN(
        n20362) );
  OAI211_X1 U22480 ( .C1(n21833), .C2(n22113), .A(n20363), .B(n20362), .ZN(
        P1_U2987) );
  XOR2_X1 U22481 ( .A(n20365), .B(n20364), .Z(n21846) );
  AOI22_X1 U22482 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20388), .ZN(n20369) );
  AOI22_X1 U22483 ( .A1(n20367), .A2(n20385), .B1(n20379), .B2(n20366), .ZN(
        n20368) );
  OAI211_X1 U22484 ( .C1(n21846), .C2(n22113), .A(n20369), .B(n20368), .ZN(
        P1_U2984) );
  INV_X1 U22485 ( .A(n20370), .ZN(n20372) );
  OAI211_X1 U22486 ( .C1(n20374), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        n20375) );
  MUX2_X1 U22487 ( .A(n20377), .B(n20376), .S(n20375), .Z(n20378) );
  XNOR2_X1 U22488 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n20378), .ZN(
        n21863) );
  AOI22_X1 U22489 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20388), .ZN(n20382) );
  AOI22_X1 U22490 ( .A1(n22214), .A2(n20385), .B1(n20380), .B2(n20379), .ZN(
        n20381) );
  OAI211_X1 U22491 ( .C1(n21863), .C2(n22113), .A(n20382), .B(n20381), .ZN(
        P1_U2982) );
  AOI22_X1 U22492 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20388), .ZN(n20387) );
  XNOR2_X1 U22493 ( .A(n13169), .B(n21874), .ZN(n20383) );
  XNOR2_X1 U22494 ( .A(n20384), .B(n20383), .ZN(n21885) );
  AOI22_X1 U22495 ( .A1(n21885), .A2(n20392), .B1(n20385), .B2(n22217), .ZN(
        n20386) );
  OAI211_X1 U22496 ( .C1(n20395), .C2(n22041), .A(n20387), .B(n20386), .ZN(
        P1_U2980) );
  AOI22_X1 U22497 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n21923), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20388), .ZN(n20394) );
  XNOR2_X1 U22498 ( .A(n13169), .B(n20389), .ZN(n20390) );
  XNOR2_X1 U22499 ( .A(n20391), .B(n20390), .ZN(n21914) );
  AOI22_X1 U22500 ( .A1(n11248), .A2(n20385), .B1(n20392), .B2(n21914), .ZN(
        n20393) );
  OAI211_X1 U22501 ( .C1(n20395), .C2(n22097), .A(n20394), .B(n20393), .ZN(
        P1_U2976) );
  INV_X1 U22502 ( .A(n20396), .ZN(n20397) );
  OAI21_X1 U22503 ( .B1(n20397), .B2(n22135), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20398) );
  OAI21_X1 U22504 ( .B1(n20399), .B2(n22122), .A(n20398), .ZN(P1_U2803) );
  OAI222_X1 U22505 ( .A1(n20459), .A2(n22154), .B1(n20459), .B2(n20400), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(n22749), .ZN(P1_U2804) );
  INV_X1 U22506 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20403) );
  AOI22_X1 U22507 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n11174), .ZN(n20402) );
  OAI21_X1 U22508 ( .B1(n20403), .B2(n20456), .A(n20402), .ZN(U247) );
  INV_X1 U22509 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20405) );
  AOI22_X1 U22510 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n11174), .ZN(n20404) );
  OAI21_X1 U22511 ( .B1(n20405), .B2(n20456), .A(n20404), .ZN(U246) );
  AOI22_X1 U22512 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n11174), .ZN(n20406) );
  OAI21_X1 U22513 ( .B1(n20407), .B2(n20456), .A(n20406), .ZN(U245) );
  AOI22_X1 U22514 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n11174), .ZN(n20408) );
  OAI21_X1 U22515 ( .B1(n20409), .B2(n20456), .A(n20408), .ZN(U244) );
  INV_X1 U22516 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20411) );
  AOI22_X1 U22517 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n11174), .ZN(n20410) );
  OAI21_X1 U22518 ( .B1(n20411), .B2(n20456), .A(n20410), .ZN(U243) );
  AOI22_X1 U22519 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n11174), .ZN(n20412) );
  OAI21_X1 U22520 ( .B1(n20413), .B2(n20456), .A(n20412), .ZN(U242) );
  INV_X1 U22521 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20415) );
  AOI22_X1 U22522 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n11174), .ZN(n20414) );
  OAI21_X1 U22523 ( .B1(n20415), .B2(n20456), .A(n20414), .ZN(U241) );
  AOI22_X1 U22524 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11174), .ZN(n20416) );
  OAI21_X1 U22525 ( .B1(n20417), .B2(n20456), .A(n20416), .ZN(U240) );
  AOI22_X1 U22526 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n11174), .ZN(n20418) );
  OAI21_X1 U22527 ( .B1(n20419), .B2(n20456), .A(n20418), .ZN(U239) );
  AOI22_X1 U22528 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n11174), .ZN(n20420) );
  OAI21_X1 U22529 ( .B1(n20421), .B2(n20456), .A(n20420), .ZN(U238) );
  AOI22_X1 U22530 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n11174), .ZN(n20422) );
  OAI21_X1 U22531 ( .B1(n14203), .B2(n20456), .A(n20422), .ZN(U237) );
  INV_X1 U22532 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20424) );
  AOI22_X1 U22533 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n11174), .ZN(n20423) );
  OAI21_X1 U22534 ( .B1(n20424), .B2(n20456), .A(n20423), .ZN(U236) );
  INV_X1 U22535 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20426) );
  AOI22_X1 U22536 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11174), .ZN(n20425) );
  OAI21_X1 U22537 ( .B1(n20426), .B2(n20456), .A(n20425), .ZN(U235) );
  INV_X1 U22538 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20428) );
  AOI22_X1 U22539 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n11174), .ZN(n20427) );
  OAI21_X1 U22540 ( .B1(n20428), .B2(n20456), .A(n20427), .ZN(U234) );
  INV_X1 U22541 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20430) );
  AOI22_X1 U22542 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n11174), .ZN(n20429) );
  OAI21_X1 U22543 ( .B1(n20430), .B2(n20456), .A(n20429), .ZN(U233) );
  INV_X1 U22544 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20432) );
  AOI22_X1 U22545 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n11174), .ZN(n20431) );
  OAI21_X1 U22546 ( .B1(n20432), .B2(n20456), .A(n20431), .ZN(U232) );
  INV_X1 U22547 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n22246) );
  AOI22_X1 U22548 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n11174), .ZN(n20433) );
  OAI21_X1 U22549 ( .B1(n22246), .B2(n20456), .A(n20433), .ZN(U231) );
  INV_X1 U22550 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n22389) );
  AOI22_X1 U22551 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n11174), .ZN(n20434) );
  OAI21_X1 U22552 ( .B1(n22389), .B2(n20456), .A(n20434), .ZN(U230) );
  INV_X1 U22553 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20436) );
  AOI22_X1 U22554 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11174), .ZN(n20435) );
  OAI21_X1 U22555 ( .B1(n20436), .B2(n20456), .A(n20435), .ZN(U229) );
  INV_X1 U22556 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n22460) );
  AOI22_X1 U22557 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n11174), .ZN(n20437) );
  OAI21_X1 U22558 ( .B1(n22460), .B2(n20456), .A(n20437), .ZN(U228) );
  AOI22_X1 U22559 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n11174), .ZN(n20438) );
  OAI21_X1 U22560 ( .B1(n20439), .B2(n20456), .A(n20438), .ZN(U227) );
  AOI22_X1 U22561 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n11174), .ZN(n20440) );
  OAI21_X1 U22562 ( .B1(n22531), .B2(n20456), .A(n20440), .ZN(U226) );
  INV_X1 U22563 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20442) );
  AOI22_X1 U22564 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n11174), .ZN(n20441) );
  OAI21_X1 U22565 ( .B1(n20442), .B2(n20456), .A(n20441), .ZN(U225) );
  AOI22_X1 U22566 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n11174), .ZN(n20443) );
  OAI21_X1 U22567 ( .B1(n22638), .B2(n20456), .A(n20443), .ZN(U224) );
  INV_X1 U22568 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n22239) );
  AOI22_X1 U22569 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n11174), .ZN(n20444) );
  OAI21_X1 U22570 ( .B1(n22239), .B2(n20456), .A(n20444), .ZN(U223) );
  AOI22_X1 U22571 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n11174), .ZN(n20445) );
  OAI21_X1 U22572 ( .B1(n22387), .B2(n20456), .A(n20445), .ZN(U222) );
  AOI22_X1 U22573 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n11174), .ZN(n20447) );
  OAI21_X1 U22574 ( .B1(n16644), .B2(n20456), .A(n20447), .ZN(U221) );
  INV_X1 U22575 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n22458) );
  AOI22_X1 U22576 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n11174), .ZN(n20448) );
  OAI21_X1 U22577 ( .B1(n22458), .B2(n20456), .A(n20448), .ZN(U220) );
  AOI22_X1 U22578 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n11174), .ZN(n20449) );
  OAI21_X1 U22579 ( .B1(n20450), .B2(n20456), .A(n20449), .ZN(U219) );
  INV_X1 U22580 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n22530) );
  AOI22_X1 U22581 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n11174), .ZN(n20451) );
  OAI21_X1 U22582 ( .B1(n22530), .B2(n20456), .A(n20451), .ZN(U218) );
  INV_X1 U22583 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20453) );
  AOI22_X1 U22584 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20446), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n11174), .ZN(n20452) );
  OAI21_X1 U22585 ( .B1(n20453), .B2(n20456), .A(n20452), .ZN(U217) );
  INV_X1 U22586 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20455) );
  OAI222_X1 U22587 ( .A1(U212), .A2(n20457), .B1(n20456), .B2(n20455), .C1(
        U214), .C2(n20454), .ZN(U216) );
  AOI22_X1 U22588 ( .A1(n20459), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20458), 
        .B2(n22749), .ZN(P1_U3483) );
  INV_X1 U22589 ( .A(n21209), .ZN(n20460) );
  OAI21_X1 U22590 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n21211), .A(n20460), 
        .ZN(n20461) );
  AOI211_X1 U22591 ( .C1(n20462), .C2(n20461), .A(n22206), .B(n21668), .ZN(
        n20464) );
  OAI21_X1 U22592 ( .B1(n20464), .B2(n21688), .A(n20463), .ZN(n20469) );
  AOI21_X1 U22593 ( .B1(n22204), .B2(n21627), .A(n20530), .ZN(n20465) );
  INV_X1 U22594 ( .A(n20465), .ZN(n20466) );
  AOI21_X1 U22595 ( .B1(n20467), .B2(n21665), .A(n20466), .ZN(n20468) );
  MUX2_X1 U22596 ( .A(n20469), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n20468), 
        .Z(P3_U3296) );
  INV_X1 U22597 ( .A(n20470), .ZN(n20471) );
  NAND2_X1 U22598 ( .A1(n21666), .A2(n20471), .ZN(n20527) );
  NAND2_X1 U22599 ( .A1(n20471), .A2(n22204), .ZN(n20971) );
  AOI22_X1 U22600 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20521), .ZN(n20473) );
  OAI21_X1 U22601 ( .B1(n20474), .B2(n20527), .A(n20473), .ZN(P3_U2768) );
  AOI22_X1 U22602 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20521), .ZN(n20475) );
  OAI21_X1 U22603 ( .B1(n20476), .B2(n20527), .A(n20475), .ZN(P3_U2769) );
  AOI22_X1 U22604 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20521), .ZN(n20477) );
  OAI21_X1 U22605 ( .B1(n20478), .B2(n20527), .A(n20477), .ZN(P3_U2770) );
  AOI22_X1 U22606 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20521), .ZN(n20480) );
  OAI21_X1 U22607 ( .B1(n21046), .B2(n20523), .A(n20480), .ZN(P3_U2771) );
  AOI22_X1 U22608 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20521), .ZN(n20481) );
  OAI21_X1 U22609 ( .B1(n20482), .B2(n20523), .A(n20481), .ZN(P3_U2772) );
  AOI22_X1 U22610 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20521), .ZN(n20483) );
  OAI21_X1 U22611 ( .B1(n21032), .B2(n20523), .A(n20483), .ZN(P3_U2773) );
  AOI22_X1 U22612 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20521), .ZN(n20484) );
  OAI21_X1 U22613 ( .B1(n20485), .B2(n20523), .A(n20484), .ZN(P3_U2774) );
  AOI22_X1 U22614 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20525), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20521), .ZN(n20486) );
  OAI21_X1 U22615 ( .B1(n20487), .B2(n20523), .A(n20486), .ZN(P3_U2775) );
  AOI22_X1 U22616 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20521), .ZN(n20488) );
  OAI21_X1 U22617 ( .B1(n20489), .B2(n20523), .A(n20488), .ZN(P3_U2776) );
  AOI22_X1 U22618 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20521), .ZN(n20490) );
  OAI21_X1 U22619 ( .B1(n20491), .B2(n20523), .A(n20490), .ZN(P3_U2777) );
  AOI22_X1 U22620 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20521), .ZN(n20492) );
  OAI21_X1 U22621 ( .B1(n21070), .B2(n20523), .A(n20492), .ZN(P3_U2778) );
  AOI22_X1 U22622 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20521), .ZN(n20493) );
  OAI21_X1 U22623 ( .B1(n20494), .B2(n20523), .A(n20493), .ZN(P3_U2779) );
  AOI22_X1 U22624 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20521), .ZN(n20495) );
  OAI21_X1 U22625 ( .B1(n21088), .B2(n20523), .A(n20495), .ZN(P3_U2780) );
  AOI22_X1 U22626 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20521), .ZN(n20496) );
  OAI21_X1 U22627 ( .B1(n20497), .B2(n20523), .A(n20496), .ZN(P3_U2781) );
  AOI22_X1 U22628 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20507), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20521), .ZN(n20498) );
  OAI21_X1 U22629 ( .B1(n20499), .B2(n20523), .A(n20498), .ZN(P3_U2782) );
  AOI22_X1 U22630 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20521), .ZN(n20500) );
  OAI21_X1 U22631 ( .B1(n21151), .B2(n20523), .A(n20500), .ZN(P3_U2783) );
  AOI22_X1 U22632 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20521), .ZN(n20501) );
  OAI21_X1 U22633 ( .B1(n21141), .B2(n20523), .A(n20501), .ZN(P3_U2784) );
  AOI22_X1 U22634 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20521), .ZN(n20502) );
  OAI21_X1 U22635 ( .B1(n20503), .B2(n20523), .A(n20502), .ZN(P3_U2785) );
  AOI22_X1 U22636 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20524), .ZN(n20504) );
  OAI21_X1 U22637 ( .B1(n20967), .B2(n20523), .A(n20504), .ZN(P3_U2786) );
  AOI22_X1 U22638 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20521), .ZN(n20505) );
  OAI21_X1 U22639 ( .B1(n21006), .B2(n20523), .A(n20505), .ZN(P3_U2787) );
  AOI22_X1 U22640 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20524), .ZN(n20506) );
  OAI21_X1 U22641 ( .B1(n20968), .B2(n20523), .A(n20506), .ZN(P3_U2788) );
  AOI22_X1 U22642 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20507), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20524), .ZN(n20508) );
  OAI21_X1 U22643 ( .B1(n20509), .B2(n20523), .A(n20508), .ZN(P3_U2789) );
  AOI22_X1 U22644 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20524), .ZN(n20510) );
  OAI21_X1 U22645 ( .B1(n20511), .B2(n20523), .A(n20510), .ZN(P3_U2790) );
  AOI22_X1 U22646 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20524), .ZN(n20512) );
  OAI21_X1 U22647 ( .B1(n21133), .B2(n20523), .A(n20512), .ZN(P3_U2791) );
  AOI22_X1 U22648 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20524), .ZN(n20513) );
  OAI21_X1 U22649 ( .B1(n20973), .B2(n20527), .A(n20513), .ZN(P3_U2792) );
  AOI22_X1 U22650 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20524), .ZN(n20514) );
  OAI21_X1 U22651 ( .B1(n20515), .B2(n20523), .A(n20514), .ZN(P3_U2793) );
  AOI22_X1 U22652 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20524), .ZN(n20516) );
  OAI21_X1 U22653 ( .B1(n20985), .B2(n20527), .A(n20516), .ZN(P3_U2794) );
  AOI22_X1 U22654 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20524), .ZN(n20517) );
  OAI21_X1 U22655 ( .B1(n20518), .B2(n20523), .A(n20517), .ZN(P3_U2795) );
  AOI22_X1 U22656 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20524), .ZN(n20519) );
  OAI21_X1 U22657 ( .B1(n20520), .B2(n20527), .A(n20519), .ZN(P3_U2796) );
  AOI22_X1 U22658 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20521), .ZN(n20522) );
  OAI21_X1 U22659 ( .B1(n21123), .B2(n20523), .A(n20522), .ZN(P3_U2797) );
  AOI22_X1 U22660 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20525), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20524), .ZN(n20526) );
  OAI21_X1 U22661 ( .B1(n21130), .B2(n20527), .A(n20526), .ZN(P3_U2798) );
  INV_X1 U22662 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20958) );
  NOR4_X1 U22663 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n21158), .ZN(n20792) );
  OAI21_X1 U22664 ( .B1(n20723), .B2(n20958), .A(n20934), .ZN(n20696) );
  INV_X1 U22665 ( .A(n20792), .ZN(n21673) );
  NOR2_X1 U22666 ( .A1(n21673), .A2(n20723), .ZN(n20949) );
  NOR2_X1 U22667 ( .A1(n20528), .A2(n21669), .ZN(n21683) );
  NOR2_X2 U22668 ( .A1(n11327), .A2(n21676), .ZN(n20941) );
  AOI21_X1 U22669 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20949), .A(
        n20941), .ZN(n20540) );
  AOI211_X1 U22670 ( .C1(n20529), .C2(n21209), .A(n22206), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n21667) );
  NAND2_X1 U22671 ( .A1(n11507), .A2(n20530), .ZN(n20531) );
  AOI211_X4 U22672 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n21211), .A(n21667), .B(
        n20531), .ZN(n20963) );
  OAI22_X1 U22673 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20957), .B1(n20903), 
        .B2(n20532), .ZN(n20538) );
  NAND2_X1 U22674 ( .A1(n22204), .A2(n22146), .ZN(n20533) );
  NAND2_X1 U22675 ( .A1(n20535), .A2(n20541), .ZN(n21157) );
  OAI22_X1 U22676 ( .A1(n20912), .A2(n20536), .B1(n21157), .B2(n20966), .ZN(
        n20537) );
  AOI211_X1 U22677 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n11327), .A(n20538), .B(
        n20537), .ZN(n20539) );
  OAI221_X1 U22678 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20696), .C1(
        n20543), .C2(n20540), .A(n20539), .ZN(P3_U2670) );
  NAND2_X1 U22679 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20541), .ZN(
        n21177) );
  NAND2_X1 U22680 ( .A1(n21173), .A2(n21177), .ZN(n21172) );
  INV_X1 U22681 ( .A(n11327), .ZN(n20956) );
  NAND2_X1 U22682 ( .A1(n20934), .A2(n20723), .ZN(n20697) );
  OAI22_X1 U22683 ( .A1(n20542), .A2(n20956), .B1(n20544), .B2(n20697), .ZN(
        n20548) );
  NOR2_X1 U22684 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20543), .ZN(
        n20679) );
  AOI21_X1 U22685 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20679), .A(
        n20723), .ZN(n20557) );
  OAI211_X1 U22686 ( .C1(n20679), .C2(n20544), .A(n20934), .B(n20557), .ZN(
        n20546) );
  NAND2_X1 U22687 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20565) );
  OAI211_X1 U22688 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20915), .B(n20565), .ZN(n20545) );
  OAI211_X1 U22689 ( .C1(n20549), .C2(n20903), .A(n20546), .B(n20545), .ZN(
        n20547) );
  AOI211_X1 U22690 ( .C1(n20554), .C2(n21172), .A(n20548), .B(n20547), .ZN(
        n20552) );
  NAND2_X1 U22691 ( .A1(n20550), .A2(n20549), .ZN(n20555) );
  OAI211_X1 U22692 ( .C1(n20550), .C2(n20549), .A(n20962), .B(n20555), .ZN(
        n20551) );
  OAI211_X1 U22693 ( .C1(n20900), .C2(n20553), .A(n20552), .B(n20551), .ZN(
        P3_U2669) );
  NAND3_X1 U22694 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20585) );
  NAND2_X1 U22695 ( .A1(n20915), .A2(n20585), .ZN(n20564) );
  NOR2_X1 U22696 ( .A1(n21191), .A2(n21190), .ZN(n21171) );
  AOI21_X1 U22697 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21171), .A(
        n21633), .ZN(n21199) );
  OR2_X1 U22698 ( .A1(n17991), .A2(n21199), .ZN(n21203) );
  AOI22_X1 U22699 ( .A1(n20963), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n20554), .B2(
        n21203), .ZN(n20563) );
  NOR2_X1 U22700 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n20555), .ZN(n20567) );
  AOI211_X1 U22701 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20555), .A(n20567), .B(
        n20912), .ZN(n20561) );
  AOI21_X1 U22702 ( .B1(n20915), .B2(n20585), .A(n11327), .ZN(n20582) );
  XOR2_X1 U22703 ( .A(n20557), .B(n20556), .Z(n20558) );
  OAI22_X1 U22704 ( .A1(n20582), .A2(n20559), .B1(n21673), .B2(n20558), .ZN(
        n20560) );
  AOI211_X1 U22705 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20561), .B(n20560), .ZN(n20562) );
  OAI211_X1 U22706 ( .C1(n20565), .C2(n20564), .A(n20563), .B(n20562), .ZN(
        P3_U2668) );
  NOR3_X1 U22707 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20957), .A3(n20585), .ZN(
        n20571) );
  NAND2_X1 U22708 ( .A1(n20567), .A2(n20566), .ZN(n20583) );
  OAI211_X1 U22709 ( .C1(n20567), .C2(n20566), .A(n20962), .B(n20583), .ZN(
        n20568) );
  OAI21_X1 U22710 ( .B1(n20900), .B2(n20569), .A(n20568), .ZN(n20570) );
  AOI211_X1 U22711 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20963), .A(n20571), .B(
        n20570), .ZN(n20581) );
  INV_X1 U22712 ( .A(n20575), .ZN(n20572) );
  AOI211_X1 U22713 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n20697), .A(
        n20696), .B(n20572), .ZN(n20579) );
  INV_X1 U22714 ( .A(n20679), .ZN(n20573) );
  OAI21_X1 U22715 ( .B1(n20574), .B2(n20573), .A(n20932), .ZN(n20589) );
  NOR3_X1 U22716 ( .A1(n20575), .A2(n21673), .A3(n20589), .ZN(n20578) );
  AOI21_X1 U22717 ( .B1(n11218), .B2(n20576), .A(n20966), .ZN(n20577) );
  NOR4_X1 U22718 ( .A1(n11176), .A2(n20579), .A3(n20578), .A4(n20577), .ZN(
        n20580) );
  OAI211_X1 U22719 ( .C1(n20582), .C2(n20586), .A(n20581), .B(n20580), .ZN(
        P3_U2667) );
  NOR2_X1 U22720 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n20583), .ZN(n20602) );
  AOI211_X1 U22721 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n20583), .A(n20602), .B(
        n20912), .ZN(n20584) );
  AOI21_X1 U22722 ( .B1(n20941), .B2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20584), .ZN(n20595) );
  NOR2_X1 U22723 ( .A1(n20586), .A2(n20585), .ZN(n20588) );
  NAND2_X1 U22724 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20588), .ZN(n20612) );
  NAND2_X1 U22725 ( .A1(n20915), .A2(n20612), .ZN(n20591) );
  INV_X1 U22726 ( .A(n20591), .ZN(n20587) );
  AOI22_X1 U22727 ( .A1(n20963), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n20588), .B2(
        n20587), .ZN(n20594) );
  XOR2_X1 U22728 ( .A(n20590), .B(n20589), .Z(n20592) );
  NAND2_X1 U22729 ( .A1(n20956), .A2(n20591), .ZN(n20617) );
  AOI22_X1 U22730 ( .A1(n20792), .A2(n20592), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n20617), .ZN(n20593) );
  NAND4_X1 U22731 ( .A1(n20595), .A2(n20594), .A3(n20593), .A4(n21620), .ZN(
        P3_U2666) );
  OAI21_X1 U22732 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20596), .A(
        n20949), .ZN(n20605) );
  NOR3_X1 U22733 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20957), .A3(n20612), .ZN(
        n20618) );
  AOI211_X1 U22734 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20941), .A(
        n11176), .B(n20618), .ZN(n20599) );
  INV_X1 U22735 ( .A(n20696), .ZN(n20597) );
  OAI211_X1 U22736 ( .C1(n20723), .C2(n11430), .A(n20606), .B(n20597), .ZN(
        n20598) );
  OAI211_X1 U22737 ( .C1(n20601), .C2(n20903), .A(n20599), .B(n20598), .ZN(
        n20600) );
  AOI21_X1 U22738 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n20617), .A(n20600), .ZN(
        n20604) );
  NAND2_X1 U22739 ( .A1(n20602), .A2(n20601), .ZN(n20610) );
  OAI211_X1 U22740 ( .C1(n20602), .C2(n20601), .A(n20962), .B(n20610), .ZN(
        n20603) );
  OAI211_X1 U22741 ( .C1(n20606), .C2(n20605), .A(n20604), .B(n20603), .ZN(
        P3_U2665) );
  AOI21_X1 U22742 ( .B1(n20607), .B2(n20958), .A(n20723), .ZN(n20608) );
  XNOR2_X1 U22743 ( .A(n20609), .B(n20608), .ZN(n20621) );
  NOR2_X1 U22744 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20610), .ZN(n20628) );
  AOI211_X1 U22745 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20610), .A(n20628), .B(
        n20912), .ZN(n20611) );
  AOI211_X1 U22746 ( .C1(n20963), .C2(P3_EBX_REG_7__SCAN_IN), .A(n11176), .B(
        n20611), .ZN(n20620) );
  NOR2_X1 U22747 ( .A1(n20613), .A2(n20612), .ZN(n20625) );
  NAND2_X1 U22748 ( .A1(n20915), .A2(n20625), .ZN(n20615) );
  OAI22_X1 U22749 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20615), .B1(n20614), 
        .B2(n20900), .ZN(n20616) );
  AOI221_X1 U22750 ( .B1(n20618), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n20617), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n20616), .ZN(n20619) );
  OAI211_X1 U22751 ( .C1(n21673), .C2(n20621), .A(n20620), .B(n20619), .ZN(
        P3_U2664) );
  AOI21_X1 U22752 ( .B1(n20622), .B2(n20958), .A(n20723), .ZN(n20624) );
  XNOR2_X1 U22753 ( .A(n20624), .B(n20623), .ZN(n20633) );
  NAND2_X1 U22754 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20625), .ZN(n20626) );
  NOR2_X1 U22755 ( .A1(n20627), .A2(n20626), .ZN(n20655) );
  OAI21_X1 U22756 ( .B1(n20655), .B2(n20957), .A(n20956), .ZN(n20644) );
  INV_X1 U22757 ( .A(n20644), .ZN(n20654) );
  AOI221_X1 U22758 ( .B1(n20957), .B2(n20627), .C1(n20626), .C2(n20627), .A(
        n20654), .ZN(n20632) );
  NAND2_X1 U22759 ( .A1(n20628), .A2(n20635), .ZN(n20636) );
  OAI211_X1 U22760 ( .C1(n20628), .C2(n20635), .A(n20962), .B(n20636), .ZN(
        n20629) );
  OAI21_X1 U22761 ( .B1(n20900), .B2(n20630), .A(n20629), .ZN(n20631) );
  AOI211_X1 U22762 ( .C1(n20792), .C2(n20633), .A(n20632), .B(n20631), .ZN(
        n20634) );
  OAI211_X1 U22763 ( .C1(n20903), .C2(n20635), .A(n20634), .B(n21620), .ZN(
        P3_U2663) );
  NOR2_X1 U22764 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20636), .ZN(n20661) );
  INV_X1 U22765 ( .A(n20636), .ZN(n20638) );
  OAI21_X1 U22766 ( .B1(n20638), .B2(n20637), .A(n20962), .ZN(n20648) );
  AOI211_X1 U22767 ( .C1(n20639), .C2(n20697), .A(n20696), .B(n20645), .ZN(
        n20643) );
  AOI22_X1 U22768 ( .A1(n20963), .A2(P3_EBX_REG_9__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20941), .ZN(n20641) );
  NAND3_X1 U22769 ( .A1(n20915), .A2(n20655), .A3(n20640), .ZN(n20653) );
  NAND3_X1 U22770 ( .A1(n20641), .A2(n21620), .A3(n20653), .ZN(n20642) );
  AOI211_X1 U22771 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n20644), .A(n20643), .B(
        n20642), .ZN(n20647) );
  OAI211_X1 U22772 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20649), .A(
        n20949), .B(n20645), .ZN(n20646) );
  OAI211_X1 U22773 ( .C1(n20661), .C2(n20648), .A(n20647), .B(n20646), .ZN(
        P3_U2662) );
  AOI21_X1 U22774 ( .B1(n20680), .B2(n20679), .A(n20723), .ZN(n20671) );
  INV_X1 U22775 ( .A(n20671), .ZN(n20669) );
  NOR2_X1 U22776 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20649), .ZN(
        n20650) );
  OAI21_X1 U22777 ( .B1(n20650), .B2(n20652), .A(n20934), .ZN(n20651) );
  AOI22_X1 U22778 ( .A1(n20652), .A2(n20669), .B1(n20697), .B2(n20651), .ZN(
        n20659) );
  AOI21_X1 U22779 ( .B1(n20654), .B2(n20653), .A(n20667), .ZN(n20658) );
  NAND2_X1 U22780 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20655), .ZN(n20665) );
  OR2_X1 U22781 ( .A1(n20957), .A2(n20665), .ZN(n20656) );
  OAI22_X1 U22782 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20656), .B1(n20903), 
        .B2(n20660), .ZN(n20657) );
  NOR4_X1 U22783 ( .A1(n11176), .A2(n20659), .A3(n20658), .A4(n20657), .ZN(
        n20663) );
  NAND2_X1 U22784 ( .A1(n20661), .A2(n20660), .ZN(n20673) );
  OAI211_X1 U22785 ( .C1(n20661), .C2(n20660), .A(n20962), .B(n20673), .ZN(
        n20662) );
  OAI211_X1 U22786 ( .C1(n20900), .C2(n20664), .A(n20663), .B(n20662), .ZN(
        P3_U2661) );
  NOR3_X1 U22787 ( .A1(n20957), .A2(n20667), .A3(n20665), .ZN(n20689) );
  NOR2_X1 U22788 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20689), .ZN(n20678) );
  NOR3_X1 U22789 ( .A1(n20667), .A2(n20666), .A3(n20665), .ZN(n20692) );
  INV_X1 U22790 ( .A(n20692), .ZN(n20668) );
  AOI21_X1 U22791 ( .B1(n20915), .B2(n20668), .A(n11327), .ZN(n20694) );
  AOI21_X1 U22792 ( .B1(n20963), .B2(P3_EBX_REG_11__SCAN_IN), .A(n11176), .ZN(
        n20677) );
  INV_X1 U22793 ( .A(n20672), .ZN(n20670) );
  AOI221_X1 U22794 ( .B1(n20672), .B2(n20671), .C1(n20670), .C2(n20669), .A(
        n21673), .ZN(n20675) );
  NOR2_X1 U22795 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n20673), .ZN(n20684) );
  AOI211_X1 U22796 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n20673), .A(n20684), .B(
        n20912), .ZN(n20674) );
  AOI211_X1 U22797 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20675), .B(n20674), .ZN(n20676) );
  OAI211_X1 U22798 ( .C1(n20678), .C2(n20694), .A(n20677), .B(n20676), .ZN(
        P3_U2660) );
  NAND3_X1 U22799 ( .A1(n20680), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n20679), .ZN(n20700) );
  NAND2_X1 U22800 ( .A1(n20932), .A2(n20700), .ZN(n20682) );
  OAI21_X1 U22801 ( .B1(n20683), .B2(n20682), .A(n20934), .ZN(n20681) );
  AOI21_X1 U22802 ( .B1(n20683), .B2(n20682), .A(n20681), .ZN(n20688) );
  NAND2_X1 U22803 ( .A1(n20684), .A2(n20686), .ZN(n20703) );
  OAI211_X1 U22804 ( .C1(n20684), .C2(n20686), .A(n20962), .B(n20703), .ZN(
        n20685) );
  OAI211_X1 U22805 ( .C1(n20903), .C2(n20686), .A(n21620), .B(n20685), .ZN(
        n20687) );
  AOI211_X1 U22806 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20688), .B(n20687), .ZN(n20690) );
  NAND3_X1 U22807 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20689), .A3(n20691), 
        .ZN(n20695) );
  OAI211_X1 U22808 ( .C1(n20691), .C2(n20694), .A(n20690), .B(n20695), .ZN(
        P3_U2659) );
  INV_X1 U22809 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20710) );
  NAND2_X1 U22810 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20692), .ZN(n20711) );
  NOR3_X1 U22811 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n20957), .A3(n20711), 
        .ZN(n20693) );
  AOI211_X1 U22812 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n20941), .A(
        n11176), .B(n20693), .ZN(n20709) );
  AOI21_X1 U22813 ( .B1(n20695), .B2(n20694), .A(n20712), .ZN(n20707) );
  AOI211_X1 U22814 ( .C1(n20698), .C2(n20697), .A(n20696), .B(n20699), .ZN(
        n20706) );
  INV_X1 U22815 ( .A(n20699), .ZN(n20702) );
  OAI21_X1 U22816 ( .B1(n20701), .B2(n20700), .A(n20932), .ZN(n20713) );
  NOR3_X1 U22817 ( .A1(n20702), .A2(n21673), .A3(n20713), .ZN(n20705) );
  NOR2_X1 U22818 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n20703), .ZN(n20719) );
  AOI211_X1 U22819 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n20703), .A(n20719), .B(
        n20912), .ZN(n20704) );
  NOR4_X1 U22820 ( .A1(n20707), .A2(n20706), .A3(n20705), .A4(n20704), .ZN(
        n20708) );
  OAI211_X1 U22821 ( .C1(n20903), .C2(n20710), .A(n20709), .B(n20708), .ZN(
        P3_U2658) );
  NOR2_X1 U22822 ( .A1(n20712), .A2(n20711), .ZN(n20722) );
  NAND2_X1 U22823 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20722), .ZN(n20749) );
  AOI21_X1 U22824 ( .B1(n20915), .B2(n20749), .A(n11327), .ZN(n20742) );
  AOI21_X1 U22825 ( .B1(n20915), .B2(n20722), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n20716) );
  XOR2_X1 U22826 ( .A(n20714), .B(n20713), .Z(n20715) );
  OAI22_X1 U22827 ( .A1(n20742), .A2(n20716), .B1(n21673), .B2(n20715), .ZN(
        n20717) );
  AOI211_X1 U22828 ( .C1(n20963), .C2(P3_EBX_REG_14__SCAN_IN), .A(n11176), .B(
        n20717), .ZN(n20721) );
  NAND2_X1 U22829 ( .A1(n20719), .A2(n20718), .ZN(n20728) );
  OAI211_X1 U22830 ( .C1(n20719), .C2(n20718), .A(n20962), .B(n20728), .ZN(
        n20720) );
  OAI211_X1 U22831 ( .C1(n20900), .C2(n11408), .A(n20721), .B(n20720), .ZN(
        P3_U2657) );
  NAND3_X1 U22832 ( .A1(n20915), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n20722), 
        .ZN(n20744) );
  AOI21_X1 U22833 ( .B1(n20724), .B2(n20958), .A(n20723), .ZN(n20757) );
  INV_X1 U22834 ( .A(n20725), .ZN(n20727) );
  INV_X1 U22835 ( .A(n20757), .ZN(n20726) );
  AOI221_X1 U22836 ( .B1(n20757), .B2(n20727), .C1(n20726), .C2(n20725), .A(
        n21673), .ZN(n20733) );
  NOR2_X1 U22837 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n20728), .ZN(n20739) );
  AOI211_X1 U22838 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20728), .A(n20739), .B(
        n20912), .ZN(n20732) );
  INV_X1 U22839 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20730) );
  OAI22_X1 U22840 ( .A1(n20903), .A2(n20730), .B1(n20729), .B2(n20900), .ZN(
        n20731) );
  NOR4_X1 U22841 ( .A1(n11176), .A2(n20733), .A3(n20732), .A4(n20731), .ZN(
        n20734) );
  OAI221_X1 U22842 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n20744), .C1(n20750), 
        .C2(n20742), .A(n20734), .ZN(P3_U2656) );
  OAI21_X1 U22843 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20735), .A(
        n20932), .ZN(n20737) );
  XOR2_X1 U22844 ( .A(n20737), .B(n20736), .Z(n20748) );
  NAND2_X1 U22845 ( .A1(n20739), .A2(n20738), .ZN(n20751) );
  OAI211_X1 U22846 ( .C1(n20739), .C2(n20738), .A(n20962), .B(n20751), .ZN(
        n20740) );
  OAI211_X1 U22847 ( .C1(n20741), .C2(n20900), .A(n21620), .B(n20740), .ZN(
        n20746) );
  XNOR2_X1 U22848 ( .A(n21588), .B(n20750), .ZN(n20743) );
  OAI22_X1 U22849 ( .A1(n20744), .A2(n20743), .B1(n21588), .B2(n20742), .ZN(
        n20745) );
  AOI211_X1 U22850 ( .C1(n20963), .C2(P3_EBX_REG_16__SCAN_IN), .A(n20746), .B(
        n20745), .ZN(n20747) );
  OAI21_X1 U22851 ( .B1(n20748), .B2(n21673), .A(n20747), .ZN(P3_U2655) );
  NOR3_X1 U22852 ( .A1(n21588), .A2(n20750), .A3(n20749), .ZN(n20752) );
  NAND2_X1 U22853 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20752), .ZN(n20790) );
  AOI21_X1 U22854 ( .B1(n20915), .B2(n20790), .A(n11327), .ZN(n20788) );
  NOR2_X1 U22855 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n20751), .ZN(n20766) );
  AOI211_X1 U22856 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n20751), .A(n20766), .B(
        n20912), .ZN(n20756) );
  INV_X1 U22857 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20754) );
  NAND3_X1 U22858 ( .A1(n20752), .A2(n20915), .A3(n20790), .ZN(n20753) );
  OAI211_X1 U22859 ( .C1(n20903), .C2(n20754), .A(n21620), .B(n20753), .ZN(
        n20755) );
  AOI211_X1 U22860 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20756), .B(n20755), .ZN(n20762) );
  NAND2_X1 U22861 ( .A1(n20760), .A2(n20759), .ZN(n20770) );
  OAI211_X1 U22862 ( .C1(n20760), .C2(n20759), .A(n20934), .B(n20770), .ZN(
        n20761) );
  OAI211_X1 U22863 ( .C1(n20788), .C2(n20763), .A(n20762), .B(n20761), .ZN(
        P3_U2654) );
  NOR2_X1 U22864 ( .A1(n20957), .A2(n20790), .ZN(n20777) );
  INV_X1 U22865 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20765) );
  OAI22_X1 U22866 ( .A1(n20903), .A2(n20765), .B1(n20764), .B2(n20900), .ZN(
        n20769) );
  NAND2_X1 U22867 ( .A1(n20766), .A2(n20765), .ZN(n20776) );
  OAI211_X1 U22868 ( .C1(n20766), .C2(n20765), .A(n20962), .B(n20776), .ZN(
        n20767) );
  NAND2_X1 U22869 ( .A1(n21620), .A2(n20767), .ZN(n20768) );
  AOI211_X1 U22870 ( .C1(n20777), .C2(n20775), .A(n20769), .B(n20768), .ZN(
        n20774) );
  OAI211_X1 U22871 ( .C1(n20772), .C2(n20771), .A(n20934), .B(n20782), .ZN(
        n20773) );
  OAI211_X1 U22872 ( .C1(n20788), .C2(n20775), .A(n20774), .B(n20773), .ZN(
        P3_U2653) );
  NOR2_X1 U22873 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n20776), .ZN(n20795) );
  AOI211_X1 U22874 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n20776), .A(n20795), .B(
        n20912), .ZN(n20781) );
  NAND2_X1 U22875 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20789) );
  OAI211_X1 U22876 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(P3_REIP_REG_19__SCAN_IN), .A(n20777), .B(n20789), .ZN(n20778) );
  OAI211_X1 U22877 ( .C1(n20903), .C2(n20779), .A(n21620), .B(n20778), .ZN(
        n20780) );
  AOI211_X1 U22878 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20781), .B(n20780), .ZN(n20786) );
  OAI211_X1 U22879 ( .C1(n20784), .C2(n20783), .A(n20934), .B(n20791), .ZN(
        n20785) );
  OAI211_X1 U22880 ( .C1(n20788), .C2(n20787), .A(n20786), .B(n20785), .ZN(
        P3_U2652) );
  NOR3_X1 U22881 ( .A1(n20802), .A2(n20790), .A3(n20789), .ZN(n20825) );
  OAI21_X1 U22882 ( .B1(n20825), .B2(n20957), .A(n20956), .ZN(n20818) );
  INV_X1 U22883 ( .A(n20818), .ZN(n20815) );
  NOR4_X1 U22884 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20957), .A3(n20790), 
        .A4(n20789), .ZN(n20800) );
  INV_X1 U22885 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20798) );
  NAND2_X1 U22886 ( .A1(n20932), .A2(n20791), .ZN(n20793) );
  NAND2_X1 U22887 ( .A1(n20793), .A2(n20794), .ZN(n20809) );
  OAI211_X1 U22888 ( .C1(n20794), .C2(n20793), .A(n20792), .B(n20809), .ZN(
        n20797) );
  NAND2_X1 U22889 ( .A1(n20795), .A2(n20798), .ZN(n20803) );
  OAI211_X1 U22890 ( .C1(n20795), .C2(n20798), .A(n20962), .B(n20803), .ZN(
        n20796) );
  OAI211_X1 U22891 ( .C1(n20798), .C2(n20903), .A(n20797), .B(n20796), .ZN(
        n20799) );
  AOI211_X1 U22892 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n20800), .B(n20799), .ZN(n20801) );
  OAI21_X1 U22893 ( .B1(n20815), .B2(n20802), .A(n20801), .ZN(P3_U2651) );
  AND3_X1 U22894 ( .A1(n20814), .A2(n20915), .A3(n20825), .ZN(n20819) );
  NOR2_X1 U22895 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n20803), .ZN(n20824) );
  INV_X1 U22896 ( .A(n20803), .ZN(n20805) );
  OAI21_X1 U22897 ( .B1(n20805), .B2(n20804), .A(n20962), .ZN(n20807) );
  OAI22_X1 U22898 ( .A1(n20824), .A2(n20807), .B1(n20900), .B2(n20806), .ZN(
        n20808) );
  AOI211_X1 U22899 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n20963), .A(n20819), .B(
        n20808), .ZN(n20813) );
  NAND2_X1 U22900 ( .A1(n20932), .A2(n20809), .ZN(n20810) );
  NAND2_X1 U22901 ( .A1(n20810), .A2(n20811), .ZN(n20820) );
  OAI211_X1 U22902 ( .C1(n20811), .C2(n20810), .A(n20934), .B(n20820), .ZN(
        n20812) );
  OAI211_X1 U22903 ( .C1(n20815), .C2(n20814), .A(n20813), .B(n20812), .ZN(
        P3_U2650) );
  OAI22_X1 U22904 ( .A1(n20903), .A2(n20823), .B1(n20816), .B2(n20900), .ZN(
        n20817) );
  AOI221_X1 U22905 ( .B1(n20819), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n20818), 
        .C2(P3_REIP_REG_22__SCAN_IN), .A(n20817), .ZN(n20829) );
  NAND2_X1 U22906 ( .A1(n20932), .A2(n20820), .ZN(n20821) );
  NAND2_X1 U22907 ( .A1(n20821), .A2(n20822), .ZN(n20838) );
  OAI211_X1 U22908 ( .C1(n20822), .C2(n20821), .A(n20934), .B(n20838), .ZN(
        n20828) );
  NAND2_X1 U22909 ( .A1(n20824), .A2(n20823), .ZN(n20832) );
  OAI211_X1 U22910 ( .C1(n20824), .C2(n20823), .A(n20962), .B(n20832), .ZN(
        n20827) );
  NAND2_X1 U22911 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20825), .ZN(n20830) );
  OR3_X1 U22912 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20957), .A3(n20830), .ZN(
        n20826) );
  NAND4_X1 U22913 ( .A1(n20829), .A2(n20828), .A3(n20827), .A4(n20826), .ZN(
        P3_U2649) );
  OR2_X1 U22914 ( .A1(n20831), .A2(n20830), .ZN(n20834) );
  NOR2_X1 U22915 ( .A1(n20843), .A2(n20834), .ZN(n20850) );
  INV_X1 U22916 ( .A(n20850), .ZN(n20866) );
  NAND2_X1 U22917 ( .A1(n20915), .A2(n20866), .ZN(n20833) );
  NAND2_X1 U22918 ( .A1(n20956), .A2(n20833), .ZN(n20861) );
  INV_X1 U22919 ( .A(n20861), .ZN(n20856) );
  NOR2_X1 U22920 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n20832), .ZN(n20844) );
  AOI211_X1 U22921 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n20832), .A(n20844), .B(
        n20912), .ZN(n20837) );
  OAI22_X1 U22922 ( .A1(n20903), .A2(n20835), .B1(n20834), .B2(n20833), .ZN(
        n20836) );
  AOI211_X1 U22923 ( .C1(n20941), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n20837), .B(n20836), .ZN(n20842) );
  NAND2_X1 U22924 ( .A1(n20932), .A2(n20838), .ZN(n20839) );
  NAND2_X1 U22925 ( .A1(n20839), .A2(n20840), .ZN(n20851) );
  OAI211_X1 U22926 ( .C1(n20840), .C2(n20839), .A(n20934), .B(n20851), .ZN(
        n20841) );
  OAI211_X1 U22927 ( .C1(n20856), .C2(n20843), .A(n20842), .B(n20841), .ZN(
        P3_U2648) );
  NOR2_X1 U22928 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20957), .ZN(n20862) );
  INV_X1 U22929 ( .A(n20844), .ZN(n20845) );
  NOR2_X1 U22930 ( .A1(n20845), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n20857) );
  AOI211_X1 U22931 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20845), .A(n20857), .B(
        n20912), .ZN(n20849) );
  INV_X1 U22932 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20847) );
  OAI22_X1 U22933 ( .A1(n20903), .A2(n20847), .B1(n20846), .B2(n20900), .ZN(
        n20848) );
  AOI211_X1 U22934 ( .C1(n20862), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        n20855) );
  NAND2_X1 U22935 ( .A1(n20932), .A2(n20851), .ZN(n20852) );
  NAND2_X1 U22936 ( .A1(n20852), .A2(n20853), .ZN(n20863) );
  OAI211_X1 U22937 ( .C1(n20853), .C2(n20852), .A(n20934), .B(n20863), .ZN(
        n20854) );
  OAI211_X1 U22938 ( .C1(n20856), .C2(n20867), .A(n20855), .B(n20854), .ZN(
        P3_U2647) );
  AOI22_X1 U22939 ( .A1(n20963), .A2(P3_EBX_REG_25__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20941), .ZN(n20872) );
  NAND2_X1 U22940 ( .A1(n20858), .A2(n20857), .ZN(n20874) );
  OAI211_X1 U22941 ( .C1(n20858), .C2(n20857), .A(n20874), .B(n20962), .ZN(
        n20859) );
  INV_X1 U22942 ( .A(n20859), .ZN(n20860) );
  AOI221_X1 U22943 ( .B1(n20862), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n20861), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n20860), .ZN(n20871) );
  NAND2_X1 U22944 ( .A1(n20932), .A2(n20863), .ZN(n20864) );
  NAND2_X1 U22945 ( .A1(n20864), .A2(n20865), .ZN(n20880) );
  OAI211_X1 U22946 ( .C1(n20865), .C2(n20864), .A(n20934), .B(n20880), .ZN(
        n20870) );
  NOR2_X1 U22947 ( .A1(n20867), .A2(n20866), .ZN(n20873) );
  NAND3_X1 U22948 ( .A1(n20915), .A2(n20873), .A3(n20868), .ZN(n20869) );
  NAND4_X1 U22949 ( .A1(n20872), .A2(n20871), .A3(n20870), .A4(n20869), .ZN(
        P3_U2646) );
  NAND2_X1 U22950 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20873), .ZN(n20876) );
  NOR2_X1 U22951 ( .A1(n20885), .A2(n20876), .ZN(n20888) );
  OR2_X1 U22952 ( .A1(n20888), .A2(n20957), .ZN(n20875) );
  NAND2_X1 U22953 ( .A1(n20956), .A2(n20875), .ZN(n20914) );
  INV_X1 U22954 ( .A(n20914), .ZN(n20899) );
  NOR2_X1 U22955 ( .A1(n20874), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n20886) );
  AOI211_X1 U22956 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20874), .A(n20886), .B(
        n20912), .ZN(n20879) );
  OAI22_X1 U22957 ( .A1(n20877), .A2(n20900), .B1(n20876), .B2(n20875), .ZN(
        n20878) );
  AOI211_X1 U22958 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20963), .A(n20879), .B(
        n20878), .ZN(n20884) );
  NAND2_X1 U22959 ( .A1(n20932), .A2(n20880), .ZN(n20881) );
  NAND2_X1 U22960 ( .A1(n20881), .A2(n20882), .ZN(n20892) );
  OAI211_X1 U22961 ( .C1(n20882), .C2(n20881), .A(n20934), .B(n20892), .ZN(
        n20883) );
  OAI211_X1 U22962 ( .C1(n20899), .C2(n20885), .A(n20884), .B(n20883), .ZN(
        P3_U2645) );
  INV_X1 U22963 ( .A(n20886), .ZN(n20887) );
  NOR2_X1 U22964 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n20887), .ZN(n20897) );
  AOI211_X1 U22965 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20887), .A(n20897), .B(
        n20912), .ZN(n20891) );
  NAND2_X1 U22966 ( .A1(n20915), .A2(n20888), .ZN(n20935) );
  OAI22_X1 U22967 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20935), .B1(n20889), 
        .B2(n20900), .ZN(n20890) );
  AOI211_X1 U22968 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n20963), .A(n20891), .B(
        n20890), .ZN(n20896) );
  NAND2_X1 U22969 ( .A1(n20932), .A2(n20892), .ZN(n20893) );
  NAND2_X1 U22970 ( .A1(n20894), .A2(n20893), .ZN(n20906) );
  OAI211_X1 U22971 ( .C1(n20894), .C2(n20893), .A(n20934), .B(n20906), .ZN(
        n20895) );
  OAI211_X1 U22972 ( .C1(n20899), .C2(n20898), .A(n20896), .B(n20895), .ZN(
        P3_U2644) );
  NAND2_X1 U22973 ( .A1(n20897), .A2(n20902), .ZN(n20913) );
  OAI21_X1 U22974 ( .B1(n20897), .B2(n20902), .A(n20913), .ZN(n20911) );
  NOR2_X1 U22975 ( .A1(n20898), .A2(n20935), .ZN(n20921) );
  OAI21_X1 U22976 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n20935), .A(n20899), 
        .ZN(n20905) );
  OAI22_X1 U22977 ( .A1(n20903), .A2(n20902), .B1(n20901), .B2(n20900), .ZN(
        n20904) );
  AOI221_X1 U22978 ( .B1(n20921), .B2(n21511), .C1(n20905), .C2(
        P3_REIP_REG_28__SCAN_IN), .A(n20904), .ZN(n20910) );
  NAND2_X1 U22979 ( .A1(n20932), .A2(n20906), .ZN(n20907) );
  OAI211_X1 U22980 ( .C1(n20908), .C2(n20907), .A(n20934), .B(n20917), .ZN(
        n20909) );
  OAI211_X1 U22981 ( .C1(n20911), .C2(n20912), .A(n20910), .B(n20909), .ZN(
        P3_U2643) );
  AOI22_X1 U22982 ( .A1(n20963), .A2(P3_EBX_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20941), .ZN(n20925) );
  NOR2_X1 U22983 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20913), .ZN(n20928) );
  NOR2_X1 U22984 ( .A1(n20928), .A2(n20912), .ZN(n20927) );
  NAND2_X1 U22985 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n20913), .ZN(n20916) );
  NAND3_X1 U22986 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n20936) );
  AOI21_X1 U22987 ( .B1(n20936), .B2(n20915), .A(n20914), .ZN(n20943) );
  INV_X1 U22988 ( .A(n20943), .ZN(n20926) );
  AOI22_X1 U22989 ( .A1(n20927), .A2(n20916), .B1(P3_REIP_REG_29__SCAN_IN), 
        .B2(n20926), .ZN(n20924) );
  OAI211_X1 U22990 ( .C1(n20919), .C2(n20918), .A(n20934), .B(n20931), .ZN(
        n20923) );
  NAND3_X1 U22991 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20921), .A3(n20920), 
        .ZN(n20922) );
  NAND4_X1 U22992 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        P3_U2642) );
  AOI22_X1 U22993 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20941), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n20926), .ZN(n20940) );
  INV_X1 U22994 ( .A(n20927), .ZN(n20930) );
  AND2_X1 U22995 ( .A1(n20962), .A2(n20928), .ZN(n20945) );
  NOR2_X1 U22996 ( .A1(n20963), .A2(n20945), .ZN(n20929) );
  MUX2_X1 U22997 ( .A(n20930), .B(n20929), .S(P3_EBX_REG_30__SCAN_IN), .Z(
        n20939) );
  NAND2_X1 U22998 ( .A1(n20947), .A2(n20948), .ZN(n20933) );
  OAI211_X1 U22999 ( .C1(n20948), .C2(n20947), .A(n20934), .B(n20933), .ZN(
        n20938) );
  NOR2_X1 U23000 ( .A1(n20936), .A2(n20935), .ZN(n20951) );
  NAND2_X1 U23001 ( .A1(n20951), .A2(n20937), .ZN(n20942) );
  NAND4_X1 U23002 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20942), .ZN(
        P3_U2641) );
  AOI22_X1 U23003 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20963), .B1(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20941), .ZN(n20955) );
  NAND2_X1 U23004 ( .A1(n20943), .A2(n20942), .ZN(n20946) );
  AOI22_X1 U23005 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20946), .B1(n20945), 
        .B2(n20944), .ZN(n20954) );
  NAND3_X1 U23006 ( .A1(n20949), .A2(n20948), .A3(n20947), .ZN(n20953) );
  NAND3_X1 U23007 ( .A1(n20951), .A2(P3_REIP_REG_30__SCAN_IN), .A3(n20950), 
        .ZN(n20952) );
  NAND4_X1 U23008 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        P3_U2640) );
  NAND2_X1 U23009 ( .A1(n20957), .A2(n20956), .ZN(n20961) );
  NOR3_X1 U23010 ( .A1(n11327), .A2(n21202), .A3(n20958), .ZN(n20960) );
  AOI21_X1 U23011 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n20961), .A(n20960), .ZN(
        n20965) );
  OAI21_X1 U23012 ( .B1(n20963), .B2(n20962), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20964) );
  OAI211_X1 U23013 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n20966), .A(
        n20965), .B(n20964), .ZN(P3_U2671) );
  NAND2_X1 U23014 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n21025) );
  NAND3_X1 U23015 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n21005) );
  NOR4_X1 U23016 ( .A1(n21005), .A2(n20968), .A3(n20967), .A4(n21006), .ZN(
        n20996) );
  NOR2_X1 U23017 ( .A1(n21063), .A2(n21134), .ZN(n21000) );
  NAND2_X1 U23018 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21000), .ZN(n20991) );
  NOR2_X1 U23019 ( .A1(n20973), .A2(n20991), .ZN(n20994) );
  NAND2_X1 U23020 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20994), .ZN(n20986) );
  NOR2_X1 U23021 ( .A1(n21025), .A2(n20986), .ZN(n21118) );
  INV_X1 U23022 ( .A(n21118), .ZN(n20978) );
  NAND2_X1 U23023 ( .A1(n20978), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U23024 ( .A1(n21150), .A2(n20974), .ZN(n21018) );
  NAND2_X1 U23025 ( .A1(n21153), .A2(n21150), .ZN(n21144) );
  AOI22_X1 U23026 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21148), .B1(n21147), .B2(
        n20975), .ZN(n20976) );
  OAI221_X1 U23027 ( .B1(n20978), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20977), 
        .C2(n21139), .A(n20976), .ZN(P3_U2722) );
  INV_X1 U23028 ( .A(n20986), .ZN(n20979) );
  AOI22_X1 U23029 ( .A1(n20979), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n21120), .ZN(n20981) );
  OAI222_X1 U23030 ( .A1(n21018), .A2(n20982), .B1(n21118), .B2(n20981), .C1(
        n21144), .C2(n20980), .ZN(P3_U2723) );
  NAND2_X1 U23031 ( .A1(n21120), .A2(n20986), .ZN(n20989) );
  AOI22_X1 U23032 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21148), .B1(n21147), .B2(
        n20983), .ZN(n20984) );
  OAI221_X1 U23033 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20986), .C1(n20985), 
        .C2(n20989), .A(n20984), .ZN(P3_U2724) );
  NOR2_X1 U23034 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20994), .ZN(n20988) );
  OAI222_X1 U23035 ( .A1(n21018), .A2(n20990), .B1(n20989), .B2(n20988), .C1(
        n21144), .C2(n20987), .ZN(P3_U2725) );
  INV_X1 U23036 ( .A(n20991), .ZN(n21125) );
  AOI21_X1 U23037 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n21120), .A(n21125), .ZN(
        n20993) );
  OAI222_X1 U23038 ( .A1(n21018), .A2(n20995), .B1(n20994), .B2(n20993), .C1(
        n21144), .C2(n20992), .ZN(P3_U2726) );
  INV_X1 U23039 ( .A(n20996), .ZN(n20998) );
  NAND2_X1 U23040 ( .A1(n20997), .A2(n21150), .ZN(n21152) );
  NOR2_X1 U23041 ( .A1(n20998), .A2(n21152), .ZN(n21009) );
  AOI22_X1 U23042 ( .A1(n21009), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n21120), .ZN(n20999) );
  OAI222_X1 U23043 ( .A1(n21018), .A2(n21001), .B1(n21000), .B2(n20999), .C1(
        n21144), .C2(n21492), .ZN(P3_U2728) );
  AND2_X1 U23044 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n21009), .ZN(n21004) );
  AOI21_X1 U23045 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21120), .A(n21009), .ZN(
        n21003) );
  OAI222_X1 U23046 ( .A1(n21044), .A2(n21018), .B1(n21004), .B2(n21003), .C1(
        n21144), .C2(n21002), .ZN(P3_U2729) );
  NOR2_X1 U23047 ( .A1(n21005), .A2(n21152), .ZN(n21023) );
  NAND2_X1 U23048 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21023), .ZN(n21011) );
  NOR2_X1 U23049 ( .A1(n21006), .A2(n21011), .ZN(n21014) );
  AOI21_X1 U23050 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21120), .A(n21014), .ZN(
        n21008) );
  OAI222_X1 U23051 ( .A1(n21010), .A2(n21018), .B1(n21009), .B2(n21008), .C1(
        n21144), .C2(n21007), .ZN(P3_U2730) );
  INV_X1 U23052 ( .A(n21011), .ZN(n21017) );
  AOI21_X1 U23053 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21120), .A(n21017), .ZN(
        n21013) );
  OAI222_X1 U23054 ( .A1(n21036), .A2(n21018), .B1(n21014), .B2(n21013), .C1(
        n21144), .C2(n21012), .ZN(P3_U2731) );
  AOI21_X1 U23055 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21120), .A(n21023), .ZN(
        n21016) );
  OAI222_X1 U23056 ( .A1(n21019), .A2(n21018), .B1(n21017), .B2(n21016), .C1(
        n21144), .C2(n21015), .ZN(P3_U2732) );
  NAND2_X1 U23057 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n21150), .ZN(n21140) );
  NOR2_X1 U23058 ( .A1(n21141), .A2(n21140), .ZN(n21138) );
  OAI21_X1 U23059 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21138), .A(n21120), .ZN(
        n21022) );
  AOI22_X1 U23060 ( .A1(n21148), .A2(BUF2_REG_2__SCAN_IN), .B1(n21147), .B2(
        n11390), .ZN(n21021) );
  OAI21_X1 U23061 ( .B1(n21023), .B2(n21022), .A(n21021), .ZN(P3_U2733) );
  NAND2_X1 U23062 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n21062) );
  NAND4_X1 U23063 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n21024)
         );
  NOR2_X1 U23064 ( .A1(n21025), .A2(n21024), .ZN(n21126) );
  NAND2_X1 U23065 ( .A1(n21132), .A2(n21126), .ZN(n21119) );
  NOR2_X1 U23066 ( .A1(n21063), .A2(n21113), .ZN(n21057) );
  NAND2_X1 U23067 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21057), .ZN(n21056) );
  NOR2_X1 U23068 ( .A1(n21062), .A2(n21056), .ZN(n21045) );
  NAND2_X1 U23069 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21045), .ZN(n21038) );
  NAND2_X1 U23070 ( .A1(n21120), .A2(n21038), .ZN(n21039) );
  NOR2_X2 U23071 ( .A1(n21026), .A2(n21120), .ZN(n21112) );
  NOR2_X2 U23072 ( .A1(n21027), .A2(n21120), .ZN(n21111) );
  INV_X1 U23073 ( .A(n21111), .ZN(n21093) );
  OAI22_X1 U23074 ( .A1(n21029), .A2(n21144), .B1(n21028), .B2(n21093), .ZN(
        n21030) );
  AOI21_X1 U23075 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21112), .A(n21030), .ZN(
        n21031) );
  OAI221_X1 U23076 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21038), .C1(n21032), 
        .C2(n21039), .A(n21031), .ZN(P3_U2714) );
  INV_X1 U23077 ( .A(n21112), .ZN(n21105) );
  AOI22_X1 U23078 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n21111), .B1(n21147), .B2(
        n21033), .ZN(n21035) );
  OAI211_X1 U23079 ( .C1(n21045), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21120), .B(
        n21038), .ZN(n21034) );
  OAI211_X1 U23080 ( .C1(n21105), .C2(n21036), .A(n21035), .B(n21034), .ZN(
        P3_U2715) );
  AOI22_X1 U23081 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n21111), .B1(n21147), .B2(
        n21037), .ZN(n21043) );
  NOR2_X1 U23082 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n21038), .ZN(n21041) );
  OAI21_X1 U23083 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21152), .A(n21039), .ZN(
        n21040) );
  AOI22_X1 U23084 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n21041), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21040), .ZN(n21042) );
  OAI211_X1 U23085 ( .C1(n21044), .C2(n21105), .A(n21043), .B(n21042), .ZN(
        P3_U2713) );
  AOI22_X1 U23086 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21111), .ZN(n21049) );
  INV_X1 U23087 ( .A(n21056), .ZN(n21052) );
  NAND2_X1 U23088 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n21052), .ZN(n21051) );
  AOI211_X1 U23089 ( .C1(n21046), .C2(n21051), .A(n21045), .B(n21139), .ZN(
        n21047) );
  INV_X1 U23090 ( .A(n21047), .ZN(n21048) );
  OAI211_X1 U23091 ( .C1(n21050), .C2(n21144), .A(n21049), .B(n21048), .ZN(
        P3_U2716) );
  AOI22_X1 U23092 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n21111), .ZN(n21054) );
  OAI211_X1 U23093 ( .C1(n21052), .C2(P3_EAX_REG_18__SCAN_IN), .A(n21120), .B(
        n21051), .ZN(n21053) );
  OAI211_X1 U23094 ( .C1(n21055), .C2(n21144), .A(n21054), .B(n21053), .ZN(
        P3_U2717) );
  AOI22_X1 U23095 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21111), .ZN(n21059) );
  OAI211_X1 U23096 ( .C1(n21057), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21120), .B(
        n21056), .ZN(n21058) );
  OAI211_X1 U23097 ( .C1(n21060), .C2(n21144), .A(n21059), .B(n21058), .ZN(
        P3_U2718) );
  AOI22_X1 U23098 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n21111), .ZN(n21066) );
  NAND4_X1 U23099 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n21061)
         );
  NAND2_X1 U23100 ( .A1(n21107), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21106) );
  NAND2_X1 U23101 ( .A1(n21101), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21100) );
  OAI211_X1 U23102 ( .C1(n21064), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21120), .B(
        n21069), .ZN(n21065) );
  OAI211_X1 U23103 ( .C1(n21067), .C2(n21144), .A(n21066), .B(n21065), .ZN(
        P3_U2710) );
  AOI22_X1 U23104 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21112), .B1(n21147), .B2(
        n21068), .ZN(n21073) );
  AOI211_X1 U23105 ( .C1(n21070), .C2(n21069), .A(n21095), .B(n21139), .ZN(
        n21071) );
  INV_X1 U23106 ( .A(n21071), .ZN(n21072) );
  OAI211_X1 U23107 ( .C1(n21093), .C2(n21074), .A(n21073), .B(n21072), .ZN(
        P3_U2709) );
  NAND2_X1 U23108 ( .A1(n21087), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n21082) );
  NAND2_X1 U23109 ( .A1(n21078), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21077) );
  OAI22_X1 U23110 ( .A1(n21139), .A2(n21078), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n21152), .ZN(n21075) );
  AOI22_X1 U23111 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21111), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n21075), .ZN(n21076) );
  OAI21_X1 U23112 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n21077), .A(n21076), .ZN(
        P3_U2704) );
  AOI22_X1 U23113 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n21111), .ZN(n21080) );
  OAI211_X1 U23114 ( .C1(n21078), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21120), .B(
        n21077), .ZN(n21079) );
  OAI211_X1 U23115 ( .C1(n21081), .C2(n21144), .A(n21080), .B(n21079), .ZN(
        P3_U2705) );
  AOI22_X1 U23116 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n21111), .ZN(n21084) );
  OAI211_X1 U23117 ( .C1(n21087), .C2(P3_EAX_REG_29__SCAN_IN), .A(n21120), .B(
        n21082), .ZN(n21083) );
  OAI211_X1 U23118 ( .C1(n21085), .C2(n21144), .A(n21084), .B(n21083), .ZN(
        P3_U2706) );
  AOI22_X1 U23119 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21112), .B1(n21147), .B2(
        n21086), .ZN(n21091) );
  AOI211_X1 U23120 ( .C1(n21088), .C2(n21094), .A(n21087), .B(n21139), .ZN(
        n21089) );
  INV_X1 U23121 ( .A(n21089), .ZN(n21090) );
  OAI211_X1 U23122 ( .C1(n21093), .C2(n21092), .A(n21091), .B(n21090), .ZN(
        P3_U2707) );
  AOI22_X1 U23123 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n21111), .ZN(n21097) );
  OAI211_X1 U23124 ( .C1(n21095), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21120), .B(
        n21094), .ZN(n21096) );
  OAI211_X1 U23125 ( .C1(n21098), .C2(n21144), .A(n21097), .B(n21096), .ZN(
        P3_U2708) );
  AOI22_X1 U23126 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n21111), .B1(n21147), .B2(
        n21099), .ZN(n21103) );
  OAI211_X1 U23127 ( .C1(n21101), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21120), .B(
        n21100), .ZN(n21102) );
  OAI211_X1 U23128 ( .C1(n21105), .C2(n21104), .A(n21103), .B(n21102), .ZN(
        P3_U2711) );
  AOI22_X1 U23129 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n21111), .ZN(n21109) );
  OAI211_X1 U23130 ( .C1(n21107), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21120), .B(
        n21106), .ZN(n21108) );
  OAI211_X1 U23131 ( .C1(n21110), .C2(n21144), .A(n21109), .B(n21108), .ZN(
        P3_U2712) );
  AOI22_X1 U23132 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21112), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21111), .ZN(n21116) );
  OAI211_X1 U23133 ( .C1(n21114), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21120), .B(
        n21113), .ZN(n21115) );
  OAI211_X1 U23134 ( .C1(n21117), .C2(n21144), .A(n21116), .B(n21115), .ZN(
        P3_U2719) );
  NAND2_X1 U23135 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21118), .ZN(n21124) );
  NAND2_X1 U23136 ( .A1(n21120), .A2(n21119), .ZN(n21129) );
  AOI22_X1 U23137 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21148), .B1(n21147), .B2(
        n21121), .ZN(n21122) );
  OAI221_X1 U23138 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n21124), .C1(n21123), 
        .C2(n21129), .A(n21122), .ZN(P3_U2721) );
  NAND2_X1 U23139 ( .A1(n21126), .A2(n21125), .ZN(n21131) );
  AOI22_X1 U23140 ( .A1(n21147), .A2(n21127), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n21148), .ZN(n21128) );
  OAI221_X1 U23141 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n21131), .C1(n21130), 
        .C2(n21129), .A(n21128), .ZN(P3_U2720) );
  AOI211_X1 U23142 ( .C1(n21134), .C2(n21133), .A(n21139), .B(n21132), .ZN(
        n21135) );
  AOI21_X1 U23143 ( .B1(n21148), .B2(BUF2_REG_8__SCAN_IN), .A(n21135), .ZN(
        n21136) );
  OAI21_X1 U23144 ( .B1(n21137), .B2(n21144), .A(n21136), .ZN(P3_U2727) );
  AOI211_X1 U23145 ( .C1(n21141), .C2(n21140), .A(n21139), .B(n21138), .ZN(
        n21142) );
  AOI21_X1 U23146 ( .B1(n21148), .B2(BUF2_REG_1__SCAN_IN), .A(n21142), .ZN(
        n21143) );
  OAI21_X1 U23147 ( .B1(n21145), .B2(n21144), .A(n21143), .ZN(P3_U2734) );
  AOI22_X1 U23148 ( .A1(n21148), .A2(BUF2_REG_0__SCAN_IN), .B1(n21147), .B2(
        n21146), .ZN(n21149) );
  OAI221_X1 U23149 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21152), .C1(n21151), 
        .C2(n21150), .A(n21149), .ZN(P3_U2735) );
  INV_X1 U23150 ( .A(n21204), .ZN(n21206) );
  INV_X1 U23151 ( .A(n21611), .ZN(n21391) );
  NOR2_X1 U23152 ( .A1(n21153), .A2(n21391), .ZN(n21156) );
  AOI22_X1 U23153 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21619), .B1(
        n21156), .B2(n21181), .ZN(n21641) );
  AOI222_X1 U23154 ( .A1(n21427), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21641), 
        .B2(n21202), .C1(n21181), .C2(n21680), .ZN(n21154) );
  AOI22_X1 U23155 ( .A1(n21206), .A2(n21181), .B1(n21154), .B2(n21204), .ZN(
        P3_U3290) );
  NOR3_X2 U23156 ( .A1(n21189), .A2(n21188), .A3(n21155), .ZN(n21610) );
  INV_X1 U23157 ( .A(n21610), .ZN(n21561) );
  OAI21_X1 U23158 ( .B1(n21600), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21561), .ZN(n21162) );
  OAI22_X1 U23159 ( .A1(n21156), .A2(n21157), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21162), .ZN(n21639) );
  INV_X1 U23160 ( .A(n21157), .ZN(n21160) );
  INV_X1 U23161 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21489) );
  AOI22_X1 U23162 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n21489), .B2(n11550), .ZN(
        n21176) );
  INV_X1 U23163 ( .A(n21176), .ZN(n21159) );
  NOR2_X1 U23164 ( .A1(n21158), .A2(n21427), .ZN(n21175) );
  AOI222_X1 U23165 ( .A1(n21639), .A2(n21202), .B1(n21160), .B2(n21680), .C1(
        n21159), .C2(n21175), .ZN(n21161) );
  AOI22_X1 U23166 ( .A1(n21206), .A2(n21190), .B1(n21161), .B2(n21204), .ZN(
        P3_U3289) );
  INV_X1 U23167 ( .A(n21652), .ZN(n21565) );
  NOR2_X1 U23168 ( .A1(n21190), .A2(n21162), .ZN(n21192) );
  AOI21_X1 U23169 ( .B1(n21163), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n21192), .ZN(n21170) );
  OAI22_X1 U23170 ( .A1(n21166), .A2(n21165), .B1(n21188), .B2(n21164), .ZN(
        n21200) );
  AOI211_X1 U23171 ( .C1(n21190), .C2(n21168), .A(n21167), .B(n21200), .ZN(
        n21169) );
  OAI222_X1 U23172 ( .A1(n21172), .A2(n21565), .B1(n21171), .B2(n21170), .C1(
        n21177), .C2(n21169), .ZN(n21635) );
  INV_X1 U23173 ( .A(n21173), .ZN(n21174) );
  AOI222_X1 U23174 ( .A1(n21635), .A2(n21202), .B1(n21176), .B2(n21175), .C1(
        n21174), .C2(n21680), .ZN(n21180) );
  INV_X1 U23175 ( .A(n21177), .ZN(n21178) );
  AOI22_X1 U23176 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21206), .B1(
        n21680), .B2(n21178), .ZN(n21179) );
  OAI21_X1 U23177 ( .B1(n21206), .B2(n21180), .A(n21179), .ZN(P3_U3288) );
  NAND2_X1 U23178 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21181), .ZN(
        n21186) );
  OAI211_X1 U23179 ( .C1(n21184), .C2(n21183), .A(n21652), .B(n21182), .ZN(
        n21185) );
  OAI22_X1 U23180 ( .A1(n21187), .A2(n21186), .B1(n18018), .B2(n21185), .ZN(
        n21198) );
  NOR2_X1 U23181 ( .A1(n21189), .A2(n21188), .ZN(n21196) );
  OAI21_X1 U23182 ( .B1(n21191), .B2(n21190), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21195) );
  INV_X1 U23183 ( .A(n21192), .ZN(n21193) );
  OAI22_X1 U23184 ( .A1(n21196), .A2(n21195), .B1(n21194), .B2(n21193), .ZN(
        n21197) );
  AOI211_X1 U23185 ( .C1(n21200), .C2(n21199), .A(n21198), .B(n21197), .ZN(
        n21632) );
  INV_X1 U23186 ( .A(n21632), .ZN(n21201) );
  AOI22_X1 U23187 ( .A1(n21680), .A2(n21203), .B1(n21202), .B2(n21201), .ZN(
        n21205) );
  AOI22_X1 U23188 ( .A1(n21206), .A2(n21633), .B1(n21205), .B2(n21204), .ZN(
        P3_U3285) );
  OAI21_X1 U23189 ( .B1(n21208), .B2(n21650), .A(n21207), .ZN(n21217) );
  OAI21_X1 U23190 ( .B1(n21212), .B2(n21211), .A(n21209), .ZN(n21210) );
  AOI21_X1 U23191 ( .B1(n21212), .B2(n21211), .A(n21210), .ZN(n21629) );
  NOR3_X1 U23192 ( .A1(n21214), .A2(n21629), .A3(n21213), .ZN(n21216) );
  AOI211_X1 U23193 ( .C1(n21218), .C2(n21217), .A(n21216), .B(n21215), .ZN(
        n21220) );
  AOI221_X4 U23194 ( .B1(n21221), .B2(n21220), .C1(n21219), .C2(n21220), .A(
        n21665), .ZN(n21602) );
  AOI22_X1 U23195 ( .A1(n21536), .A2(n21557), .B1(n21651), .B2(n21331), .ZN(
        n21330) );
  AOI21_X1 U23196 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21268) );
  NAND3_X1 U23197 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21295) );
  NOR2_X1 U23198 ( .A1(n21268), .A2(n21295), .ZN(n21283) );
  NAND2_X1 U23199 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21283), .ZN(
        n21306) );
  NOR3_X1 U23200 ( .A1(n21329), .A2(n21316), .A3(n21306), .ZN(n21355) );
  NAND2_X1 U23201 ( .A1(n21222), .A2(n21355), .ZN(n21402) );
  NOR2_X1 U23202 ( .A1(n21223), .A2(n21402), .ZN(n21231) );
  NAND2_X1 U23203 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21265) );
  NOR2_X1 U23204 ( .A1(n21295), .A2(n21265), .ZN(n21282) );
  NAND2_X1 U23205 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21282), .ZN(
        n21305) );
  NOR2_X1 U23206 ( .A1(n21316), .A2(n21305), .ZN(n21617) );
  NAND2_X1 U23207 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21617), .ZN(
        n21599) );
  NOR2_X1 U23208 ( .A1(n21224), .A2(n21599), .ZN(n21228) );
  OAI21_X1 U23209 ( .B1(n21611), .B2(n21427), .A(n21619), .ZN(n21255) );
  AOI22_X1 U23210 ( .A1(n21652), .A2(n21231), .B1(n21228), .B2(n21255), .ZN(
        n21400) );
  OAI21_X1 U23211 ( .B1(n21330), .B2(n21224), .A(n21400), .ZN(n21389) );
  NAND2_X1 U23212 ( .A1(n21602), .A2(n21389), .ZN(n21550) );
  NAND2_X1 U23213 ( .A1(n21491), .A2(n21225), .ZN(n21321) );
  AOI21_X1 U23214 ( .B1(n21623), .B2(n21227), .A(n21226), .ZN(n21240) );
  OAI221_X1 U23215 ( .B1(n21611), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21611), .C2(n21228), .A(n21602), .ZN(n21534) );
  INV_X1 U23216 ( .A(n21228), .ZN(n21229) );
  OAI21_X1 U23217 ( .B1(n21229), .B2(n21543), .A(n21600), .ZN(n21230) );
  OAI21_X1 U23218 ( .B1(n21231), .B2(n21565), .A(n21230), .ZN(n21533) );
  OAI22_X1 U23219 ( .A1(n21565), .A2(n21237), .B1(n21619), .B2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21232) );
  AOI21_X1 U23220 ( .B1(n21233), .B2(n21651), .A(n21232), .ZN(n21234) );
  INV_X1 U23221 ( .A(n21234), .ZN(n21235) );
  AOI211_X1 U23222 ( .C1(n21536), .C2(n21236), .A(n21533), .B(n21235), .ZN(
        n21393) );
  OAI21_X1 U23223 ( .B1(n21611), .B2(n21237), .A(n21393), .ZN(n21238) );
  OAI211_X1 U23224 ( .C1(n21534), .C2(n21238), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n21620), .ZN(n21239) );
  OAI211_X1 U23225 ( .C1(n21241), .C2(n21550), .A(n21240), .B(n21239), .ZN(
        P3_U2841) );
  NAND2_X1 U23226 ( .A1(n21611), .A2(n21565), .ZN(n21542) );
  OAI22_X1 U23227 ( .A1(n21619), .A2(n21427), .B1(n21243), .B2(n21658), .ZN(
        n21242) );
  AOI21_X1 U23228 ( .B1(n21427), .B2(n21542), .A(n21242), .ZN(n21246) );
  NOR2_X2 U23229 ( .A1(n11176), .A2(n21602), .ZN(n21615) );
  NOR2_X1 U23230 ( .A1(n21470), .A2(n21579), .ZN(n21419) );
  AOI22_X1 U23231 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21615), .B1(
        n21419), .B2(n21243), .ZN(n21245) );
  NAND2_X1 U23232 ( .A1(n11176), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21244) );
  OAI211_X1 U23233 ( .C1(n21246), .C2(n21470), .A(n21245), .B(n21244), .ZN(
        P3_U2862) );
  NAND3_X1 U23234 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21427), .A3(
        n21542), .ZN(n21248) );
  OAI211_X1 U23235 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n21600), .A(
        n11550), .B(n21582), .ZN(n21247) );
  OAI211_X1 U23236 ( .C1(n21249), .C2(n21658), .A(n21248), .B(n21247), .ZN(
        n21251) );
  AOI22_X1 U23237 ( .A1(n21602), .A2(n21251), .B1(n21419), .B2(n21250), .ZN(
        n21253) );
  NAND2_X1 U23238 ( .A1(n11176), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21252) );
  OAI211_X1 U23239 ( .C1(n21591), .C2(n11550), .A(n21253), .B(n21252), .ZN(
        P3_U2861) );
  INV_X1 U23240 ( .A(n21419), .ZN(n21304) );
  NOR2_X1 U23241 ( .A1(n11550), .A2(n21427), .ZN(n21254) );
  OAI221_X1 U23242 ( .B1(n21268), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n21268), .C2(n21254), .A(n21652), .ZN(n21259) );
  NOR2_X1 U23243 ( .A1(n21611), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21401) );
  INV_X1 U23244 ( .A(n21401), .ZN(n21554) );
  OAI21_X1 U23245 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21610), .A(
        n21554), .ZN(n21257) );
  INV_X1 U23246 ( .A(n21255), .ZN(n21444) );
  NOR3_X1 U23247 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21444), .A3(
        n11550), .ZN(n21256) );
  AOI21_X1 U23248 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21257), .A(
        n21256), .ZN(n21258) );
  OAI211_X1 U23249 ( .C1(n21658), .C2(n21260), .A(n21259), .B(n21258), .ZN(
        n21261) );
  AOI22_X1 U23250 ( .A1(n21602), .A2(n21261), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21615), .ZN(n21263) );
  OAI211_X1 U23251 ( .C1(n21304), .C2(n21264), .A(n21263), .B(n21262), .ZN(
        P3_U2860) );
  OAI22_X1 U23252 ( .A1(n21565), .A2(n21268), .B1(n21265), .B2(n21444), .ZN(
        n21286) );
  INV_X1 U23253 ( .A(n21286), .ZN(n21296) );
  INV_X1 U23254 ( .A(n21265), .ZN(n21266) );
  AOI21_X1 U23255 ( .B1(n21266), .B2(n21554), .A(n21610), .ZN(n21267) );
  AOI211_X1 U23256 ( .C1(n21652), .C2(n21268), .A(n21267), .B(n21274), .ZN(
        n21273) );
  AOI21_X1 U23257 ( .B1(n21296), .B2(n21274), .A(n21273), .ZN(n21270) );
  OAI21_X1 U23258 ( .B1(n21270), .B2(n21269), .A(n21602), .ZN(n21271) );
  OAI211_X1 U23259 ( .C1(n21591), .C2(n21274), .A(n21272), .B(n21271), .ZN(
        P3_U2859) );
  INV_X1 U23260 ( .A(n21582), .ZN(n21318) );
  NOR2_X1 U23261 ( .A1(n21318), .A2(n21273), .ZN(n21279) );
  NOR3_X1 U23262 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21296), .A3(
        n21274), .ZN(n21278) );
  OAI22_X1 U23263 ( .A1(n21658), .A2(n21276), .B1(n21579), .B2(n21275), .ZN(
        n21277) );
  AOI211_X1 U23264 ( .C1(n21279), .C2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n21278), .B(n21277), .ZN(n21281) );
  AOI22_X1 U23265 ( .A1(n11176), .A2(P3_REIP_REG_4__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21615), .ZN(n21280) );
  OAI21_X1 U23266 ( .B1(n21281), .B2(n21470), .A(n21280), .ZN(P3_U2858) );
  OAI22_X1 U23267 ( .A1(n21283), .A2(n21565), .B1(n21282), .B2(n21610), .ZN(
        n21284) );
  NOR2_X1 U23268 ( .A1(n21401), .A2(n21284), .ZN(n21285) );
  OAI21_X1 U23269 ( .B1(n21285), .B2(n21470), .A(n21591), .ZN(n21299) );
  INV_X1 U23270 ( .A(n21299), .ZN(n21294) );
  AND4_X1 U23271 ( .A1(n21293), .A2(n21286), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21290) );
  OAI22_X1 U23272 ( .A1(n21658), .A2(n21288), .B1(n21579), .B2(n21287), .ZN(
        n21289) );
  OAI21_X1 U23273 ( .B1(n21290), .B2(n21289), .A(n21602), .ZN(n21291) );
  OAI211_X1 U23274 ( .C1(n21294), .C2(n21293), .A(n21292), .B(n21291), .ZN(
        P3_U2857) );
  NOR2_X1 U23275 ( .A1(n21296), .A2(n21295), .ZN(n21308) );
  INV_X1 U23276 ( .A(n21308), .ZN(n21298) );
  OAI22_X1 U23277 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21298), .B1(
        n21658), .B2(n21297), .ZN(n21300) );
  AOI22_X1 U23278 ( .A1(n21602), .A2(n21300), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21299), .ZN(n21302) );
  NAND2_X1 U23279 ( .A1(n11176), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21301) );
  OAI211_X1 U23280 ( .C1(n21304), .C2(n21303), .A(n21302), .B(n21301), .ZN(
        P3_U2856) );
  AOI22_X1 U23281 ( .A1(n21652), .A2(n21306), .B1(n21305), .B2(n21561), .ZN(
        n21307) );
  AND3_X1 U23282 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n21307), .A3(
        n21554), .ZN(n21317) );
  NAND2_X1 U23283 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21308), .ZN(
        n21315) );
  AND2_X1 U23284 ( .A1(n21316), .A2(n21315), .ZN(n21310) );
  OAI22_X1 U23285 ( .A1(n21317), .A2(n21310), .B1(n21658), .B2(n21309), .ZN(
        n21312) );
  AOI22_X1 U23286 ( .A1(n21602), .A2(n21312), .B1(n21419), .B2(n21311), .ZN(
        n21314) );
  NAND2_X1 U23287 ( .A1(n11176), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21313) );
  OAI211_X1 U23288 ( .C1(n21591), .C2(n21316), .A(n21314), .B(n21313), .ZN(
        P3_U2855) );
  INV_X1 U23289 ( .A(n21328), .ZN(n21320) );
  NOR2_X1 U23290 ( .A1(n21318), .A2(n21317), .ZN(n21319) );
  MUX2_X1 U23291 ( .A(n21320), .B(n21319), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n21324) );
  OAI22_X1 U23292 ( .A1(n21579), .A2(n21322), .B1(n21321), .B2(n21325), .ZN(
        n21323) );
  AOI211_X1 U23293 ( .C1(n21536), .C2(n21325), .A(n21324), .B(n21323), .ZN(
        n21327) );
  AOI22_X1 U23294 ( .A1(n11176), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21615), .ZN(n21326) );
  OAI21_X1 U23295 ( .B1(n21327), .B2(n21470), .A(n21326), .ZN(P3_U2854) );
  NOR2_X1 U23296 ( .A1(n21329), .A2(n21328), .ZN(n21380) );
  INV_X1 U23297 ( .A(n21380), .ZN(n21354) );
  NAND2_X1 U23298 ( .A1(n21330), .A2(n21354), .ZN(n21348) );
  NAND2_X1 U23299 ( .A1(n21602), .A2(n21348), .ZN(n21626) );
  NOR2_X1 U23300 ( .A1(n21427), .A2(n21599), .ZN(n21609) );
  NAND2_X1 U23301 ( .A1(n21556), .A2(n21579), .ZN(n21559) );
  NOR2_X1 U23302 ( .A1(n21355), .A2(n21565), .ZN(n21614) );
  OAI22_X1 U23303 ( .A1(n21557), .A2(n21556), .B1(n21579), .B2(n21331), .ZN(
        n21612) );
  AOI211_X1 U23304 ( .C1(n21333), .C2(n21559), .A(n21614), .B(n21612), .ZN(
        n21332) );
  OAI221_X1 U23305 ( .B1(n21611), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n21611), .C2(n21609), .A(n21332), .ZN(n21605) );
  OAI21_X1 U23306 ( .B1(n21333), .B2(n21599), .A(n21600), .ZN(n21334) );
  OAI21_X1 U23307 ( .B1(n21349), .B2(n21565), .A(n21334), .ZN(n21342) );
  AOI211_X1 U23308 ( .C1(n21391), .C2(n21597), .A(n21605), .B(n21342), .ZN(
        n21335) );
  OAI21_X1 U23309 ( .B1(n21335), .B2(n21470), .A(n21591), .ZN(n21337) );
  AOI22_X1 U23310 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21337), .B1(
        n21623), .B2(n21336), .ZN(n21339) );
  OAI211_X1 U23311 ( .C1(n21626), .C2(n21340), .A(n21339), .B(n21338), .ZN(
        P3_U2851) );
  AOI21_X1 U23312 ( .B1(n21356), .B2(n21609), .A(n21611), .ZN(n21357) );
  AOI211_X1 U23313 ( .C1(n21600), .C2(n21341), .A(n21357), .B(n21614), .ZN(
        n21345) );
  AOI21_X1 U23314 ( .B1(n21536), .B2(n21343), .A(n21342), .ZN(n21344) );
  OAI211_X1 U23315 ( .C1(n21346), .C2(n21579), .A(n21345), .B(n21344), .ZN(
        n21593) );
  OAI222_X1 U23316 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21349), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21348), .C1(n21593), 
        .C2(n21347), .ZN(n21353) );
  AOI22_X1 U23317 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21615), .B1(
        n21623), .B2(n21350), .ZN(n21352) );
  OAI211_X1 U23318 ( .C1(n21470), .C2(n21353), .A(n21352), .B(n21351), .ZN(
        P3_U2850) );
  NOR3_X1 U23319 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21360), .A3(
        n21354), .ZN(n21364) );
  AOI21_X1 U23320 ( .B1(n21356), .B2(n21355), .A(n21565), .ZN(n21358) );
  AOI211_X1 U23321 ( .C1(n21359), .C2(n21542), .A(n21358), .B(n21357), .ZN(
        n21362) );
  OAI21_X1 U23322 ( .B1(n21360), .B2(n21599), .A(n21600), .ZN(n21361) );
  AOI21_X1 U23323 ( .B1(n21362), .B2(n21361), .A(n21372), .ZN(n21363) );
  AOI211_X1 U23324 ( .C1(n21536), .C2(n21365), .A(n21364), .B(n21363), .ZN(
        n21367) );
  OAI22_X1 U23325 ( .A1(n21367), .A2(n21470), .B1(n21366), .B2(n21569), .ZN(
        n21368) );
  AOI21_X1 U23326 ( .B1(n21419), .B2(n21369), .A(n21368), .ZN(n21371) );
  OAI211_X1 U23327 ( .C1(n21591), .C2(n21372), .A(n21371), .B(n21370), .ZN(
        P3_U2848) );
  NOR2_X1 U23328 ( .A1(n21373), .A2(n21556), .ZN(n21376) );
  INV_X1 U23329 ( .A(n21599), .ZN(n21375) );
  AOI211_X1 U23330 ( .C1(n21402), .C2(n21652), .A(n21401), .B(n18087), .ZN(
        n21374) );
  OAI221_X1 U23331 ( .B1(n21610), .B2(n21379), .C1(n21610), .C2(n21375), .A(
        n21374), .ZN(n21581) );
  AOI221_X1 U23332 ( .B1(n21376), .B2(n21602), .C1(n21581), .C2(n21602), .A(
        n21615), .ZN(n21388) );
  INV_X1 U23333 ( .A(n21376), .ZN(n21578) );
  OAI211_X1 U23334 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n21378), .A(
        n21651), .B(n21377), .ZN(n21382) );
  NAND3_X1 U23335 ( .A1(n21380), .A2(n21379), .A3(n21581), .ZN(n21381) );
  OAI211_X1 U23336 ( .C1(n21578), .C2(n21383), .A(n21382), .B(n21381), .ZN(
        n21385) );
  AOI22_X1 U23337 ( .A1(n21602), .A2(n21385), .B1(n21623), .B2(n21384), .ZN(
        n21387) );
  OAI211_X1 U23338 ( .C1(n21388), .C2(n18087), .A(n21387), .B(n21386), .ZN(
        P3_U2847) );
  NAND2_X1 U23339 ( .A1(n21390), .A2(n21389), .ZN(n21512) );
  AOI21_X1 U23340 ( .B1(n21512), .B2(n21513), .A(n21470), .ZN(n21395) );
  NOR2_X1 U23341 ( .A1(n21552), .A2(n21599), .ZN(n21555) );
  NAND2_X1 U23342 ( .A1(n21403), .A2(n21555), .ZN(n21426) );
  OAI22_X1 U23343 ( .A1(n21401), .A2(n21426), .B1(n21391), .B2(n21513), .ZN(
        n21392) );
  OAI211_X1 U23344 ( .C1(n21603), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n21393), .B(n21392), .ZN(n21394) );
  AOI22_X1 U23345 ( .A1(n21623), .A2(n21396), .B1(n21395), .B2(n21394), .ZN(
        n21398) );
  NAND2_X1 U23346 ( .A1(n11176), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21397) );
  OAI211_X1 U23347 ( .C1(n21591), .C2(n21513), .A(n21398), .B(n21397), .ZN(
        P3_U2840) );
  NOR3_X1 U23348 ( .A1(n21400), .A2(n21526), .A3(n21399), .ZN(n21407) );
  OAI21_X1 U23349 ( .B1(n21401), .B2(n21426), .A(n21561), .ZN(n21515) );
  INV_X1 U23350 ( .A(n21402), .ZN(n21563) );
  NAND2_X1 U23351 ( .A1(n21563), .A2(n21403), .ZN(n21428) );
  NAND2_X1 U23352 ( .A1(n21652), .A2(n21428), .ZN(n21519) );
  NAND4_X1 U23353 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n21515), .A4(n21519), .ZN(
        n21416) );
  NAND3_X1 U23354 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21582), .A3(
        n21416), .ZN(n21404) );
  OAI21_X1 U23355 ( .B1(n21405), .B2(n21579), .A(n21404), .ZN(n21406) );
  AOI211_X1 U23356 ( .C1(n21536), .C2(n21408), .A(n21407), .B(n21406), .ZN(
        n21412) );
  AOI22_X1 U23357 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21615), .B1(
        n21623), .B2(n21409), .ZN(n21411) );
  NAND2_X1 U23358 ( .A1(n11176), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21410) );
  OAI211_X1 U23359 ( .C1(n21412), .C2(n21470), .A(n21411), .B(n21410), .ZN(
        P3_U2837) );
  AOI21_X1 U23360 ( .B1(n21615), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21413), .ZN(n21423) );
  NOR2_X1 U23361 ( .A1(n21512), .A2(n21414), .ZN(n21433) );
  AOI221_X1 U23362 ( .B1(n21417), .B2(n21582), .C1(n21416), .C2(n21582), .A(
        n21415), .ZN(n21420) );
  NAND2_X1 U23363 ( .A1(n21536), .A2(n21418), .ZN(n21430) );
  NAND2_X1 U23364 ( .A1(n21419), .A2(n21447), .ZN(n21434) );
  OAI221_X1 U23365 ( .B1(n21470), .B2(n21420), .C1(n21470), .C2(n21430), .A(
        n21434), .ZN(n21421) );
  OAI21_X1 U23366 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21433), .A(
        n21421), .ZN(n21422) );
  OAI211_X1 U23367 ( .C1(n21424), .C2(n21569), .A(n21423), .B(n21422), .ZN(
        P3_U2836) );
  NAND3_X1 U23368 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n21425), .ZN(n21429) );
  NOR2_X1 U23369 ( .A1(n21426), .A2(n21429), .ZN(n21451) );
  INV_X1 U23370 ( .A(n21451), .ZN(n21442) );
  NOR2_X1 U23371 ( .A1(n21427), .A2(n21442), .ZN(n21453) );
  NOR2_X1 U23372 ( .A1(n21429), .A2(n21428), .ZN(n21440) );
  NOR2_X1 U23373 ( .A1(n21440), .A2(n21565), .ZN(n21463) );
  NOR2_X1 U23374 ( .A1(n21463), .A2(n21502), .ZN(n21446) );
  OAI21_X1 U23375 ( .B1(n21619), .B2(n21451), .A(n21446), .ZN(n21497) );
  INV_X1 U23376 ( .A(n21497), .ZN(n21431) );
  OAI211_X1 U23377 ( .C1(n21611), .C2(n21453), .A(n21431), .B(n21430), .ZN(
        n21432) );
  AOI22_X1 U23378 ( .A1(n21602), .A2(n21432), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21615), .ZN(n21435) );
  NAND2_X1 U23379 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21433), .ZN(
        n21503) );
  AOI22_X1 U23380 ( .A1(n21435), .A2(n21434), .B1(n21503), .B2(n21502), .ZN(
        n21436) );
  AOI21_X1 U23381 ( .B1(n21623), .B2(n21437), .A(n21436), .ZN(n21439) );
  NAND2_X1 U23382 ( .A1(n21439), .A2(n21438), .ZN(P3_U2835) );
  NAND2_X1 U23383 ( .A1(n21652), .A2(n21440), .ZN(n21443) );
  AOI221_X1 U23384 ( .B1(n21444), .B2(n21443), .C1(n21442), .C2(n21443), .A(
        n21441), .ZN(n21477) );
  AOI21_X1 U23385 ( .B1(n21536), .B2(n21499), .A(n21477), .ZN(n21445) );
  OAI21_X1 U23386 ( .B1(n21579), .B2(n21495), .A(n21445), .ZN(n21472) );
  NAND2_X1 U23387 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21446), .ZN(
        n21456) );
  NOR2_X1 U23388 ( .A1(n21447), .A2(n21464), .ZN(n21450) );
  INV_X1 U23389 ( .A(n21448), .ZN(n21449) );
  OAI22_X1 U23390 ( .A1(n21450), .A2(n21579), .B1(n21449), .B2(n21556), .ZN(
        n21467) );
  NAND2_X1 U23391 ( .A1(n21452), .A2(n21451), .ZN(n21454) );
  AOI21_X1 U23392 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21453), .A(
        n21611), .ZN(n21496) );
  AOI21_X1 U23393 ( .B1(n21600), .B2(n21454), .A(n21496), .ZN(n21466) );
  INV_X1 U23394 ( .A(n21466), .ZN(n21455) );
  AOI211_X1 U23395 ( .C1(n21542), .C2(n21456), .A(n21467), .B(n21455), .ZN(
        n21457) );
  OAI21_X1 U23396 ( .B1(n21457), .B2(n21470), .A(n21591), .ZN(n21458) );
  OAI222_X1 U23397 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21602), 
        .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21472), .C1(n21459), 
        .C2(n21458), .ZN(n21461) );
  OAI211_X1 U23398 ( .C1(n21462), .C2(n21569), .A(n21461), .B(n21460), .ZN(
        P3_U2833) );
  AOI211_X1 U23399 ( .C1(n21582), .C2(n21464), .A(n21463), .B(n21468), .ZN(
        n21465) );
  NAND2_X1 U23400 ( .A1(n21466), .A2(n21465), .ZN(n21480) );
  OAI22_X1 U23401 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n21467), .B2(n21480), .ZN(
        n21469) );
  OAI22_X1 U23402 ( .A1(n21470), .A2(n21469), .B1(n21591), .B2(n21468), .ZN(
        n21471) );
  OAI21_X1 U23403 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21472), .A(
        n21471), .ZN(n21473) );
  OAI211_X1 U23404 ( .C1(n21475), .C2(n21569), .A(n21474), .B(n21473), .ZN(
        P3_U2832) );
  NOR2_X1 U23405 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21476), .ZN(
        n21478) );
  AOI22_X1 U23406 ( .A1(n21479), .A2(n21651), .B1(n21478), .B2(n21477), .ZN(
        n21482) );
  NAND3_X1 U23407 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21582), .A3(
        n21480), .ZN(n21481) );
  OAI211_X1 U23408 ( .C1(n21483), .C2(n21556), .A(n21482), .B(n21481), .ZN(
        n21485) );
  AOI22_X1 U23409 ( .A1(n21602), .A2(n21485), .B1(n21623), .B2(n21484), .ZN(
        n21488) );
  INV_X1 U23410 ( .A(n21486), .ZN(n21487) );
  OAI211_X1 U23411 ( .C1(n21489), .C2(n21591), .A(n21488), .B(n21487), .ZN(
        P3_U2831) );
  OAI21_X1 U23412 ( .B1(n21492), .B2(n21504), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21493) );
  INV_X1 U23413 ( .A(n21603), .ZN(n21498) );
  AOI211_X1 U23414 ( .C1(n21498), .C2(n21497), .A(n21496), .B(n21615), .ZN(
        n21501) );
  OAI22_X1 U23415 ( .A1(n21505), .A2(n21504), .B1(n21503), .B2(n21502), .ZN(
        n21506) );
  NOR3_X1 U23416 ( .A1(n21615), .A2(n21513), .A3(n21512), .ZN(n21521) );
  AOI21_X1 U23417 ( .B1(n21651), .B2(n21514), .A(n21615), .ZN(n21516) );
  OAI211_X1 U23418 ( .C1(n21517), .C2(n21556), .A(n21516), .B(n21515), .ZN(
        n21529) );
  NOR2_X1 U23419 ( .A1(n21518), .A2(n21529), .ZN(n21520) );
  AOI21_X1 U23420 ( .B1(n21520), .B2(n21519), .A(n11176), .ZN(n21528) );
  OAI21_X1 U23421 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21521), .A(
        n21528), .ZN(n21523) );
  OAI211_X1 U23422 ( .C1(n21569), .C2(n21524), .A(n21523), .B(n21522), .ZN(
        P3_U2839) );
  NOR4_X1 U23423 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21526), .A3(
        n21525), .A4(n21550), .ZN(n21527) );
  AOI21_X1 U23424 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n11176), .A(n21527), 
        .ZN(n21531) );
  OAI211_X1 U23425 ( .C1(n21582), .C2(n21529), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21528), .ZN(n21530) );
  OAI211_X1 U23426 ( .C1(n21532), .C2(n21569), .A(n21531), .B(n21530), .ZN(
        P3_U2838) );
  AOI211_X1 U23427 ( .C1(n21536), .C2(n21535), .A(n21534), .B(n21533), .ZN(
        n21537) );
  OAI21_X1 U23428 ( .B1(n21579), .B2(n21538), .A(n21537), .ZN(n21539) );
  NAND2_X1 U23429 ( .A1(n21539), .A2(n21620), .ZN(n21544) );
  AOI22_X1 U23430 ( .A1(n11176), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n21623), 
        .B2(n21540), .ZN(n21541) );
  OAI221_X1 U23431 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21550), 
        .C1(n21543), .C2(n21544), .A(n21541), .ZN(P3_U2843) );
  NAND3_X1 U23432 ( .A1(n21543), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n21542), 
        .ZN(n21545) );
  NAND2_X1 U23433 ( .A1(n21545), .A2(n21544), .ZN(n21547) );
  AOI22_X1 U23434 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21547), .B1(
        n21623), .B2(n21546), .ZN(n21549) );
  OAI211_X1 U23435 ( .C1(n21551), .C2(n21550), .A(n21549), .B(n21548), .ZN(
        P3_U2842) );
  NOR2_X1 U23436 ( .A1(n21552), .A2(n21626), .ZN(n21585) );
  AOI22_X1 U23437 ( .A1(n11176), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n21585), 
        .B2(n21553), .ZN(n21568) );
  NAND3_X1 U23438 ( .A1(n21555), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n21554), .ZN(n21560) );
  OAI211_X1 U23439 ( .C1(n21557), .C2(n21556), .A(n21564), .B(n21580), .ZN(
        n21558) );
  AOI22_X1 U23440 ( .A1(n21561), .A2(n21560), .B1(n21559), .B2(n21558), .ZN(
        n21562) );
  OAI221_X1 U23441 ( .B1(n21565), .B2(n21564), .C1(n21565), .C2(n21563), .A(
        n21562), .ZN(n21571) );
  OAI21_X1 U23442 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n21610), .A(
        n21602), .ZN(n21566) );
  OAI211_X1 U23443 ( .C1(n21571), .C2(n21566), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n21620), .ZN(n21567) );
  OAI211_X1 U23444 ( .C1(n21570), .C2(n21569), .A(n21568), .B(n21567), .ZN(
        P3_U2844) );
  AOI21_X1 U23445 ( .B1(n21602), .B2(n21571), .A(n21615), .ZN(n21577) );
  AOI22_X1 U23446 ( .A1(n21623), .A2(n21573), .B1(n21585), .B2(n21572), .ZN(
        n21575) );
  OAI211_X1 U23447 ( .C1(n21577), .C2(n21576), .A(n21575), .B(n21574), .ZN(
        P3_U2845) );
  OAI211_X1 U23448 ( .C1(n21580), .C2(n21579), .A(n21602), .B(n21578), .ZN(
        n21583) );
  OAI221_X1 U23449 ( .B1(n21583), .B2(n21582), .C1(n21583), .C2(n21581), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21589) );
  AOI22_X1 U23450 ( .A1(n21586), .A2(n21623), .B1(n21585), .B2(n21584), .ZN(
        n21587) );
  OAI221_X1 U23451 ( .B1(n11176), .B2(n21589), .C1(n21620), .C2(n21588), .A(
        n21587), .ZN(P3_U2846) );
  AOI22_X1 U23452 ( .A1(n11176), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21623), 
        .B2(n21590), .ZN(n21595) );
  OAI21_X1 U23453 ( .B1(n21603), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n21591), .ZN(n21592) );
  OAI211_X1 U23454 ( .C1(n21593), .C2(n21592), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n21620), .ZN(n21594) );
  OAI211_X1 U23455 ( .C1(n21596), .C2(n21626), .A(n21595), .B(n21594), .ZN(
        P3_U2849) );
  NAND2_X1 U23456 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21597), .ZN(
        n21608) );
  AOI22_X1 U23457 ( .A1(n11176), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21623), 
        .B2(n21598), .ZN(n21607) );
  NAND2_X1 U23458 ( .A1(n21600), .A2(n21599), .ZN(n21601) );
  OAI211_X1 U23459 ( .C1(n21603), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21602), .B(n21601), .ZN(n21604) );
  OAI211_X1 U23460 ( .C1(n21605), .C2(n21604), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21620), .ZN(n21606) );
  OAI211_X1 U23461 ( .C1(n21608), .C2(n21626), .A(n21607), .B(n21606), .ZN(
        P3_U2852) );
  AOI211_X1 U23462 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n21611), .A(
        n21610), .B(n21609), .ZN(n21613) );
  NOR4_X1 U23463 ( .A1(n21615), .A2(n21614), .A3(n21613), .A4(n21612), .ZN(
        n21618) );
  AOI221_X1 U23464 ( .B1(n21619), .B2(n21618), .C1(n21617), .C2(n21618), .A(
        n21616), .ZN(n21621) );
  AOI22_X1 U23465 ( .A1(n21623), .A2(n21622), .B1(n21621), .B2(n21620), .ZN(
        n21625) );
  OAI211_X1 U23466 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21626), .A(
        n21625), .B(n21624), .ZN(P3_U2853) );
  NAND2_X1 U23467 ( .A1(n22206), .A2(n21627), .ZN(n21678) );
  NOR2_X1 U23468 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(P3_MORE_REG_SCAN_IN), .ZN(
        n21664) );
  OAI211_X1 U23469 ( .C1(n21629), .C2(n22206), .A(n21656), .B(n21628), .ZN(
        n21689) );
  AOI211_X1 U23470 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21644), .A(
        n21631), .B(n21630), .ZN(n21663) );
  INV_X1 U23471 ( .A(n21644), .ZN(n21634) );
  AOI22_X1 U23472 ( .A1(n21644), .A2(n21633), .B1(n21632), .B2(n21634), .ZN(
        n21661) );
  AOI22_X1 U23473 ( .A1(n21644), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21635), .B2(n21634), .ZN(n21636) );
  OAI21_X1 U23474 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21636), .ZN(n21660) );
  INV_X1 U23475 ( .A(n21661), .ZN(n21649) );
  INV_X1 U23476 ( .A(n21636), .ZN(n21647) );
  OR3_X1 U23477 ( .A1(n21641), .A2(n21640), .A3(n21637), .ZN(n21638) );
  AOI22_X1 U23478 ( .A1(n21641), .A2(n21640), .B1(n21639), .B2(n21638), .ZN(
        n21643) );
  OAI21_X1 U23479 ( .B1(n21644), .B2(n21643), .A(n21642), .ZN(n21645) );
  AOI222_X1 U23480 ( .A1(n21647), .A2(n21646), .B1(n21647), .B2(n21645), .C1(
        n21646), .C2(n21645), .ZN(n21648) );
  AOI211_X1 U23481 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n21649), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n21648), .ZN(n21659) );
  INV_X1 U23482 ( .A(n21650), .ZN(n21657) );
  NOR2_X1 U23483 ( .A1(n21652), .A2(n21651), .ZN(n21654) );
  OAI222_X1 U23484 ( .A1(n21658), .A2(n21657), .B1(n21656), .B2(n21655), .C1(
        n21654), .C2(n21653), .ZN(n21691) );
  AOI211_X1 U23485 ( .C1(n21661), .C2(n21660), .A(n21659), .B(n21691), .ZN(
        n21662) );
  OAI211_X1 U23486 ( .C1(n21664), .C2(n21689), .A(n21663), .B(n21662), .ZN(
        n21684) );
  AOI211_X1 U23487 ( .C1(n21667), .C2(n21666), .A(n21665), .B(n21684), .ZN(
        n21674) );
  AOI21_X1 U23488 ( .B1(n22206), .B2(n21668), .A(n21674), .ZN(n21687) );
  NAND3_X1 U23489 ( .A1(n21670), .A2(n21687), .A3(n21669), .ZN(n21671) );
  NAND4_X1 U23490 ( .A1(n21673), .A2(n21678), .A3(n21672), .A4(n21671), .ZN(
        P3_U2997) );
  NOR2_X1 U23491 ( .A1(n21674), .A2(n21688), .ZN(n21677) );
  OAI21_X1 U23492 ( .B1(n21677), .B2(n21676), .A(n21675), .ZN(P3_U3282) );
  INV_X1 U23493 ( .A(n21678), .ZN(n21679) );
  AOI211_X1 U23494 ( .C1(n21681), .C2(n21680), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n21679), .ZN(n21682) );
  AOI211_X1 U23495 ( .C1(n21690), .C2(n21684), .A(n21683), .B(n21682), .ZN(
        n21685) );
  OAI221_X1 U23496 ( .B1(n21688), .B2(n21687), .C1(n21688), .C2(n21686), .A(
        n21685), .ZN(P3_U2996) );
  NAND2_X1 U23497 ( .A1(n21690), .A2(n21689), .ZN(n21693) );
  MUX2_X1 U23498 ( .A(n21691), .B(P3_MORE_REG_SCAN_IN), .S(n21693), .Z(
        P3_U3295) );
  AOI21_X1 U23499 ( .B1(n21693), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21692), .ZN(
        n21694) );
  INV_X1 U23500 ( .A(n21694), .ZN(P3_U2637) );
  INV_X1 U23501 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22160) );
  AOI211_X1 U23502 ( .C1(n21698), .C2(n21697), .A(n21696), .B(n21695), .ZN(
        n21704) );
  NAND2_X1 U23503 ( .A1(n21699), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21700) );
  OAI21_X1 U23504 ( .B1(n21701), .B2(n21700), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21703) );
  NOR2_X1 U23505 ( .A1(n21704), .A2(n22130), .ZN(n21702) );
  AOI22_X1 U23506 ( .A1(n22160), .A2(n21704), .B1(n21703), .B2(n21702), .ZN(
        P1_U3485) );
  INV_X1 U23507 ( .A(n21878), .ZN(n21709) );
  OAI22_X1 U23508 ( .A1(n21715), .A2(n21707), .B1(n21706), .B2(n21705), .ZN(
        n21708) );
  AOI211_X1 U23509 ( .C1(n21709), .C2(n21710), .A(n21819), .B(n21708), .ZN(
        n21720) );
  AND2_X1 U23510 ( .A1(n21710), .A2(n21709), .ZN(n21714) );
  NOR2_X1 U23511 ( .A1(n21711), .A2(n21915), .ZN(n21713) );
  AND2_X1 U23512 ( .A1(n21712), .A2(n21729), .ZN(n21724) );
  AOI211_X1 U23513 ( .C1(n21715), .C2(n21714), .A(n21713), .B(n21724), .ZN(
        n21719) );
  AOI22_X1 U23514 ( .A1(n21925), .A2(n21717), .B1(n11156), .B2(n21716), .ZN(
        n21718) );
  OAI211_X1 U23515 ( .C1(n21720), .C2(n21729), .A(n21719), .B(n21718), .ZN(
        P1_U3018) );
  INV_X1 U23516 ( .A(n21720), .ZN(n21723) );
  NOR2_X1 U23517 ( .A1(n21721), .A2(n21915), .ZN(n21722) );
  AOI221_X1 U23518 ( .B1(n21724), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n21723), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n21722), .ZN(
        n21733) );
  NAND2_X1 U23519 ( .A1(n21821), .A2(n21779), .ZN(n21726) );
  NAND3_X1 U23520 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n21725), .ZN(n21763) );
  NAND2_X1 U23521 ( .A1(n21726), .A2(n21763), .ZN(n21799) );
  NAND2_X1 U23522 ( .A1(n21727), .A2(n21799), .ZN(n21835) );
  NOR3_X1 U23523 ( .A1(n21729), .A2(n21728), .A3(n21835), .ZN(n21841) );
  AOI22_X1 U23524 ( .A1(n11156), .A2(n21731), .B1(n21841), .B2(n21730), .ZN(
        n21732) );
  OAI211_X1 U23525 ( .C1(n21906), .C2(n22007), .A(n21733), .B(n21732), .ZN(
        P1_U3017) );
  NOR2_X1 U23526 ( .A1(n21743), .A2(n21936), .ZN(n21736) );
  OAI21_X1 U23527 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21826), .A(
        n21734), .ZN(n21735) );
  AOI21_X1 U23528 ( .B1(n21821), .B2(n21736), .A(n21735), .ZN(n21746) );
  INV_X1 U23529 ( .A(n21737), .ZN(n21742) );
  INV_X1 U23530 ( .A(n21779), .ZN(n21738) );
  NAND2_X1 U23531 ( .A1(n21821), .A2(n21738), .ZN(n21749) );
  OAI211_X1 U23532 ( .C1(n21906), .C2(n21740), .A(n21749), .B(n21739), .ZN(
        n21741) );
  AOI21_X1 U23533 ( .B1(n21742), .B2(n11156), .A(n21741), .ZN(n21745) );
  INV_X1 U23534 ( .A(n21826), .ZN(n21747) );
  NAND2_X1 U23535 ( .A1(n21743), .A2(n21878), .ZN(n21921) );
  NAND4_X1 U23536 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21748), .A3(
        n21747), .A4(n21921), .ZN(n21744) );
  OAI211_X1 U23537 ( .C1(n21746), .C2(n21748), .A(n21745), .B(n21744), .ZN(
        P1_U3029) );
  OAI21_X1 U23538 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21799), .ZN(n21753) );
  AOI22_X1 U23539 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21923), .B1(n21925), 
        .B2(n21937), .ZN(n21752) );
  AOI221_X1 U23540 ( .B1(n21748), .B2(n21747), .C1(n21936), .C2(n21747), .A(
        n21819), .ZN(n21780) );
  NAND2_X1 U23541 ( .A1(n21749), .A2(n21780), .ZN(n21802) );
  AOI22_X1 U23542 ( .A1(n21750), .A2(n11156), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21802), .ZN(n21751) );
  OAI211_X1 U23543 ( .C1(n21761), .C2(n21753), .A(n21752), .B(n21751), .ZN(
        P1_U3027) );
  INV_X1 U23544 ( .A(n21799), .ZN(n21766) );
  AOI22_X1 U23545 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21923), .B1(n21925), 
        .B2(n21754), .ZN(n21758) );
  INV_X1 U23546 ( .A(n21755), .ZN(n21756) );
  AOI22_X1 U23547 ( .A1(n21756), .A2(n11156), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21802), .ZN(n21757) );
  OAI211_X1 U23548 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n21766), .A(
        n21758), .B(n21757), .ZN(P1_U3028) );
  INV_X1 U23549 ( .A(n21765), .ZN(n21781) );
  NAND2_X1 U23550 ( .A1(n21781), .A2(n21779), .ZN(n21760) );
  OAI21_X1 U23551 ( .B1(n21826), .B2(n21761), .A(n21780), .ZN(n21759) );
  AOI21_X1 U23552 ( .B1(n21821), .B2(n21760), .A(n21759), .ZN(n21778) );
  NAND2_X1 U23553 ( .A1(n21761), .A2(n21777), .ZN(n21772) );
  AOI221_X1 U23554 ( .B1(n21763), .B2(n21778), .C1(n21772), .C2(n21778), .A(
        n21762), .ZN(n21769) );
  NOR2_X1 U23555 ( .A1(n21764), .A2(n21862), .ZN(n21768) );
  NOR3_X1 U23556 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21766), .A3(
        n21765), .ZN(n21767) );
  NOR3_X1 U23557 ( .A1(n21769), .A2(n21768), .A3(n21767), .ZN(n21771) );
  NAND2_X1 U23558 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21923), .ZN(n21770) );
  OAI211_X1 U23559 ( .C1(n21906), .C2(n21966), .A(n21771), .B(n21770), .ZN(
        P1_U3025) );
  AOI22_X1 U23560 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21923), .B1(n21925), 
        .B2(n21949), .ZN(n21776) );
  INV_X1 U23561 ( .A(n21772), .ZN(n21773) );
  AOI22_X1 U23562 ( .A1(n21774), .A2(n11156), .B1(n21773), .B2(n21799), .ZN(
        n21775) );
  OAI211_X1 U23563 ( .C1(n21778), .C2(n21777), .A(n21776), .B(n21775), .ZN(
        P1_U3026) );
  NAND2_X1 U23564 ( .A1(n21800), .A2(n21799), .ZN(n21788) );
  NAND4_X1 U23565 ( .A1(n21781), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n21780), .A4(n21779), .ZN(n21782) );
  NAND2_X1 U23566 ( .A1(n21783), .A2(n21782), .ZN(n21797) );
  INV_X1 U23567 ( .A(n21976), .ZN(n21784) );
  AOI222_X1 U23568 ( .A1(n21785), .A2(n11156), .B1(n21925), .B2(n21784), .C1(
        n21923), .C2(P1_REIP_REG_7__SCAN_IN), .ZN(n21786) );
  OAI221_X1 U23569 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21788), .C1(
        n21789), .C2(n21797), .A(n21786), .ZN(P1_U3024) );
  INV_X1 U23570 ( .A(n21787), .ZN(n21795) );
  AOI211_X1 U23571 ( .C1(n21798), .C2(n21789), .A(n21801), .B(n21788), .ZN(
        n21794) );
  INV_X1 U23572 ( .A(n21790), .ZN(n21791) );
  OAI21_X1 U23573 ( .B1(n21906), .B2(n21792), .A(n21791), .ZN(n21793) );
  AOI211_X1 U23574 ( .C1(n21795), .C2(n11156), .A(n21794), .B(n21793), .ZN(
        n21796) );
  OAI21_X1 U23575 ( .B1(n21798), .B2(n21797), .A(n21796), .ZN(P1_U3023) );
  NAND3_X1 U23576 ( .A1(n21801), .A2(n21800), .A3(n21799), .ZN(n21810) );
  INV_X1 U23577 ( .A(n21848), .ZN(n21922) );
  AOI21_X1 U23578 ( .B1(n21922), .B2(n21803), .A(n21802), .ZN(n21818) );
  INV_X1 U23579 ( .A(n21804), .ZN(n21808) );
  NOR2_X1 U23580 ( .A1(n21805), .A2(n21862), .ZN(n21806) );
  AOI211_X1 U23581 ( .C1(n21925), .C2(n21808), .A(n21807), .B(n21806), .ZN(
        n21809) );
  OAI221_X1 U23582 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21810), .C1(
        n21811), .C2(n21818), .A(n21809), .ZN(P1_U3022) );
  AOI221_X1 U23583 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n21811), .C2(n15685), .A(
        n21810), .ZN(n21815) );
  OAI22_X1 U23584 ( .A1(n21813), .A2(n21915), .B1(n21906), .B2(n21812), .ZN(
        n21814) );
  AOI211_X1 U23585 ( .C1(n21816), .C2(n11156), .A(n21815), .B(n21814), .ZN(
        n21817) );
  OAI21_X1 U23586 ( .B1(n21818), .B2(n15685), .A(n21817), .ZN(P1_U3021) );
  AOI21_X1 U23587 ( .B1(n21821), .B2(n21820), .A(n21819), .ZN(n21824) );
  AOI21_X1 U23588 ( .B1(n21826), .B2(n21824), .A(n21822), .ZN(n21831) );
  INV_X1 U23589 ( .A(n21823), .ZN(n21825) );
  OAI211_X1 U23590 ( .C1(n21826), .C2(n21825), .A(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n21824), .ZN(n21836) );
  NOR3_X1 U23591 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n20354), .A3(
        n21835), .ZN(n21830) );
  OAI22_X1 U23592 ( .A1(n21828), .A2(n21915), .B1(n21906), .B2(n21827), .ZN(
        n21829) );
  AOI211_X1 U23593 ( .C1(n21831), .C2(n21836), .A(n21830), .B(n21829), .ZN(
        n21832) );
  OAI21_X1 U23594 ( .B1(n21833), .B2(n21862), .A(n21832), .ZN(P1_U3019) );
  AOI22_X1 U23595 ( .A1(n21925), .A2(n21988), .B1(n11156), .B2(n21834), .ZN(
        n21839) );
  INV_X1 U23596 ( .A(n21835), .ZN(n21837) );
  OAI21_X1 U23597 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21837), .A(
        n21836), .ZN(n21838) );
  OAI211_X1 U23598 ( .C1(n21915), .C2(n21840), .A(n21839), .B(n21838), .ZN(
        P1_U3020) );
  AOI22_X1 U23599 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n21923), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21847), .ZN(n21845) );
  NAND2_X1 U23600 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21841), .ZN(
        n21856) );
  INV_X1 U23601 ( .A(n21856), .ZN(n21871) );
  AOI22_X1 U23602 ( .A1(n21843), .A2(n21925), .B1(n21871), .B2(n21842), .ZN(
        n21844) );
  OAI211_X1 U23603 ( .C1(n21846), .C2(n21862), .A(n21845), .B(n21844), .ZN(
        P1_U3016) );
  INV_X1 U23604 ( .A(n21847), .ZN(n21866) );
  OAI21_X1 U23605 ( .B1(n21848), .B2(n21850), .A(n21866), .ZN(n21858) );
  AOI22_X1 U23606 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n21923), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21858), .ZN(n21854) );
  INV_X1 U23607 ( .A(n21849), .ZN(n21852) );
  NOR2_X1 U23608 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21856), .ZN(
        n21851) );
  AOI22_X1 U23609 ( .A1(n21852), .A2(n11156), .B1(n21851), .B2(n21850), .ZN(
        n21853) );
  OAI211_X1 U23610 ( .C1(n21906), .C2(n22031), .A(n21854), .B(n21853), .ZN(
        P1_U3013) );
  OAI21_X1 U23611 ( .B1(n21870), .B2(n21856), .A(n21855), .ZN(n21857) );
  AOI22_X1 U23612 ( .A1(n21925), .A2(n21859), .B1(n21858), .B2(n21857), .ZN(
        n21861) );
  NAND2_X1 U23613 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21923), .ZN(n21860) );
  OAI211_X1 U23614 ( .C1(n21863), .C2(n21862), .A(n21861), .B(n21860), .ZN(
        P1_U3014) );
  OAI22_X1 U23615 ( .A1(n21866), .A2(n21865), .B1(n21864), .B2(n21915), .ZN(
        n21867) );
  AOI21_X1 U23616 ( .B1(n11156), .B2(n21868), .A(n21867), .ZN(n21873) );
  NAND3_X1 U23617 ( .A1(n21871), .A2(n21870), .A3(n21869), .ZN(n21872) );
  OAI211_X1 U23618 ( .C1(n22016), .C2(n21906), .A(n21873), .B(n21872), .ZN(
        P1_U3015) );
  NOR2_X1 U23619 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21874), .ZN(
        n21875) );
  AOI22_X1 U23620 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n21923), .B1(n21875), 
        .B2(n21883), .ZN(n21882) );
  OAI221_X1 U23621 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21878), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21877), .A(n21876), .ZN(
        n21880) );
  AOI22_X1 U23622 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21880), .B1(
        n11156), .B2(n21879), .ZN(n21881) );
  OAI211_X1 U23623 ( .C1(n21906), .C2(n22051), .A(n21882), .B(n21881), .ZN(
        P1_U3011) );
  INV_X1 U23624 ( .A(n21883), .ZN(n21889) );
  AOI22_X1 U23625 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n21923), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21884), .ZN(n21887) );
  AOI22_X1 U23626 ( .A1(n21885), .A2(n11156), .B1(n21925), .B2(n22045), .ZN(
        n21886) );
  OAI211_X1 U23627 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21889), .A(
        n21887), .B(n21886), .ZN(P1_U3012) );
  NOR2_X1 U23628 ( .A1(n22075), .A2(n21915), .ZN(n21891) );
  NOR3_X1 U23629 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21889), .A3(
        n21888), .ZN(n21890) );
  AOI211_X1 U23630 ( .C1(n21892), .C2(n11156), .A(n21891), .B(n21890), .ZN(
        n21897) );
  INV_X1 U23631 ( .A(n21893), .ZN(n21894) );
  OAI21_X1 U23632 ( .B1(n21895), .B2(n21894), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21896) );
  OAI211_X1 U23633 ( .C1(n21906), .C2(n22083), .A(n21897), .B(n21896), .ZN(
        P1_U3009) );
  AOI22_X1 U23634 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21923), .B1(n11156), 
        .B2(n21898), .ZN(n21904) );
  INV_X1 U23635 ( .A(n21899), .ZN(n21902) );
  AND2_X1 U23636 ( .A1(n21900), .A2(n21912), .ZN(n21907) );
  OAI22_X1 U23637 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21902), .B1(
        n21907), .B2(n21901), .ZN(n21903) );
  OAI211_X1 U23638 ( .C1(n21906), .C2(n21905), .A(n21904), .B(n21903), .ZN(
        P1_U3005) );
  AOI21_X1 U23639 ( .B1(n21923), .B2(P1_REIP_REG_25__SCAN_IN), .A(n21907), 
        .ZN(n21911) );
  AOI22_X1 U23640 ( .A1(n21925), .A2(n21909), .B1(n11156), .B2(n21908), .ZN(
        n21910) );
  OAI211_X1 U23641 ( .C1(n21913), .C2(n21912), .A(n21911), .B(n21910), .ZN(
        P1_U3006) );
  AOI22_X1 U23642 ( .A1(n21914), .A2(n11156), .B1(n21925), .B2(n22092), .ZN(
        n21920) );
  NOR2_X1 U23643 ( .A1(n22086), .A2(n21915), .ZN(n21916) );
  AOI211_X1 U23644 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21918), .A(
        n21917), .B(n21916), .ZN(n21919) );
  NAND2_X1 U23645 ( .A1(n21920), .A2(n21919), .ZN(P1_U3008) );
  NAND3_X1 U23646 ( .A1(n21936), .A2(n21922), .A3(n21921), .ZN(n21932) );
  NAND2_X1 U23647 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21923), .ZN(n21931) );
  NAND2_X1 U23648 ( .A1(n21925), .A2(n21924), .ZN(n21930) );
  NAND3_X1 U23649 ( .A1(n11156), .A2(n21927), .A3(n21926), .ZN(n21929) );
  AND4_X1 U23650 ( .A1(n21932), .A2(n21931), .A3(n21930), .A4(n21929), .ZN(
        n21933) );
  OAI221_X1 U23651 ( .B1(n21936), .B2(n21935), .C1(n21936), .C2(n21934), .A(
        n21933), .ZN(P1_U3030) );
  AOI22_X1 U23652 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(n22079), .B1(n22093), .B2(
        n21937), .ZN(n21939) );
  AOI21_X1 U23653 ( .B1(n22061), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22044), .ZN(n21938) );
  OAI211_X1 U23654 ( .C1(n21941), .C2(n21940), .A(n21939), .B(n21938), .ZN(
        n21945) );
  AOI21_X1 U23655 ( .B1(n22073), .B2(n21950), .A(n21964), .ZN(n21954) );
  AOI21_X1 U23656 ( .B1(n21943), .B2(n21942), .A(n21954), .ZN(n21944) );
  AOI211_X1 U23657 ( .C1(n21946), .C2(n21957), .A(n21945), .B(n21944), .ZN(
        n21947) );
  OAI21_X1 U23658 ( .B1(n21948), .B2(n22096), .A(n21947), .ZN(P1_U2836) );
  AOI22_X1 U23659 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n22079), .B1(n22093), .B2(
        n21949), .ZN(n21953) );
  NOR3_X1 U23660 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21950), .A3(n22069), .ZN(
        n21951) );
  AOI211_X1 U23661 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n22044), .B(n21951), .ZN(n21952) );
  OAI211_X1 U23662 ( .C1(n21955), .C2(n21954), .A(n21953), .B(n21952), .ZN(
        n21956) );
  AOI21_X1 U23663 ( .B1(n21958), .B2(n21957), .A(n21956), .ZN(n21959) );
  OAI21_X1 U23664 ( .B1(n21960), .B2(n22096), .A(n21959), .ZN(P1_U2835) );
  NOR2_X1 U23665 ( .A1(n21961), .A2(n22069), .ZN(n21962) );
  AOI22_X1 U23666 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n22079), .B1(n21963), .B2(
        n21962), .ZN(n21974) );
  AOI21_X1 U23667 ( .B1(n22073), .B2(n21965), .A(n21964), .ZN(n21978) );
  OAI21_X1 U23668 ( .B1(n21966), .B2(n22111), .A(n22023), .ZN(n21967) );
  AOI21_X1 U23669 ( .B1(n22061), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21967), .ZN(n21970) );
  NAND2_X1 U23670 ( .A1(n21968), .A2(n22108), .ZN(n21969) );
  OAI211_X1 U23671 ( .C1(n21978), .C2(n21971), .A(n21970), .B(n21969), .ZN(
        n21972) );
  INV_X1 U23672 ( .A(n21972), .ZN(n21973) );
  OAI211_X1 U23673 ( .C1(n21975), .C2(n22096), .A(n21974), .B(n21973), .ZN(
        P1_U2834) );
  OAI22_X1 U23674 ( .A1(n21978), .A2(n21977), .B1(n22111), .B2(n21976), .ZN(
        n21979) );
  AOI211_X1 U23675 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22044), .B(n21979), .ZN(n21985) );
  OAI22_X1 U23676 ( .A1(n21981), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n21980), 
        .B2(n22100), .ZN(n21982) );
  AOI21_X1 U23677 ( .B1(n22108), .B2(n21983), .A(n21982), .ZN(n21984) );
  OAI211_X1 U23678 ( .C1(n21986), .C2(n22096), .A(n21985), .B(n21984), .ZN(
        P1_U2833) );
  NOR2_X1 U23679 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22069), .ZN(n22002) );
  AOI22_X1 U23680 ( .A1(n22093), .A2(n21988), .B1(n21987), .B2(n22002), .ZN(
        n21994) );
  AOI22_X1 U23681 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22001), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n22061), .ZN(n21989) );
  OAI211_X1 U23682 ( .C1(n22100), .C2(n21990), .A(n21989), .B(n22023), .ZN(
        n21991) );
  AOI21_X1 U23683 ( .B1(n22108), .B2(n21992), .A(n21991), .ZN(n21993) );
  OAI211_X1 U23684 ( .C1(n21995), .C2(n22096), .A(n21994), .B(n21993), .ZN(
        P1_U2829) );
  AOI22_X1 U23685 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(n22079), .B1(n22093), 
        .B2(n21996), .ZN(n22006) );
  NOR3_X1 U23686 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n21997), .A3(n22069), 
        .ZN(n21998) );
  AOI211_X1 U23687 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22044), .B(n21998), .ZN(n22005) );
  AOI22_X1 U23688 ( .A1(n22000), .A2(n22107), .B1(n22108), .B2(n21999), .ZN(
        n22004) );
  OAI21_X1 U23689 ( .B1(n22002), .B2(n22001), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n22003) );
  NAND4_X1 U23690 ( .A1(n22006), .A2(n22005), .A3(n22004), .A4(n22003), .ZN(
        P1_U2828) );
  AOI22_X1 U23691 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(n22079), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n22061), .ZN(n22015) );
  OAI22_X1 U23692 ( .A1(n22008), .A2(n22052), .B1(n22111), .B2(n22007), .ZN(
        n22009) );
  AOI21_X1 U23693 ( .B1(n22010), .B2(n22107), .A(n22009), .ZN(n22014) );
  OAI211_X1 U23694 ( .C1(P1_REIP_REG_14__SCAN_IN), .C2(n22012), .A(n22011), 
        .B(n22040), .ZN(n22013) );
  NAND4_X1 U23695 ( .A1(n22015), .A2(n22014), .A3(n22023), .A4(n22013), .ZN(
        P1_U2826) );
  AOI22_X1 U23696 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n22079), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n22061), .ZN(n22025) );
  OAI22_X1 U23697 ( .A1(n22017), .A2(n22052), .B1(n22111), .B2(n22016), .ZN(
        n22018) );
  AOI21_X1 U23698 ( .B1(n22019), .B2(n22107), .A(n22018), .ZN(n22024) );
  OAI211_X1 U23699 ( .C1(n22021), .C2(P1_REIP_REG_16__SCAN_IN), .A(n22040), 
        .B(n22020), .ZN(n22022) );
  NAND4_X1 U23700 ( .A1(n22025), .A2(n22024), .A3(n22023), .A4(n22022), .ZN(
        P1_U2824) );
  NAND2_X1 U23701 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n22026), .ZN(n22037) );
  INV_X1 U23702 ( .A(n22037), .ZN(n22039) );
  AOI21_X1 U23703 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n22040), .A(n22026), 
        .ZN(n22036) );
  OAI22_X1 U23704 ( .A1(n22028), .A2(n22100), .B1(n22027), .B2(n22098), .ZN(
        n22029) );
  AOI211_X1 U23705 ( .C1(n22107), .C2(n22030), .A(n22044), .B(n22029), .ZN(
        n22035) );
  INV_X1 U23706 ( .A(n22031), .ZN(n22032) );
  AOI22_X1 U23707 ( .A1(n22033), .A2(n22108), .B1(n22093), .B2(n22032), .ZN(
        n22034) );
  OAI211_X1 U23708 ( .C1(n22039), .C2(n22036), .A(n22035), .B(n22034), .ZN(
        P1_U2822) );
  NOR2_X1 U23709 ( .A1(n22038), .A2(n22037), .ZN(n22055) );
  AOI21_X1 U23710 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n22040), .A(n22039), 
        .ZN(n22048) );
  OAI22_X1 U23711 ( .A1(n22042), .A2(n22100), .B1(n22041), .B2(n22096), .ZN(
        n22043) );
  AOI211_X1 U23712 ( .C1(n22061), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22044), .B(n22043), .ZN(n22047) );
  AOI22_X1 U23713 ( .A1(n22217), .A2(n22108), .B1(n22093), .B2(n22045), .ZN(
        n22046) );
  OAI211_X1 U23714 ( .C1(n22055), .C2(n22048), .A(n22047), .B(n22046), .ZN(
        P1_U2821) );
  AOI22_X1 U23715 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n22061), .B1(
        n22049), .B2(n22107), .ZN(n22057) );
  OAI21_X1 U23716 ( .B1(n22060), .B2(n22069), .A(n22050), .ZN(n22071) );
  OAI22_X1 U23717 ( .A1(n22053), .A2(n22052), .B1(n22111), .B2(n22051), .ZN(
        n22054) );
  AOI221_X1 U23718 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n22071), .C1(n22055), 
        .C2(n22071), .A(n22054), .ZN(n22056) );
  OAI211_X1 U23719 ( .C1(n22058), .C2(n22100), .A(n22057), .B(n22056), .ZN(
        P1_U2820) );
  NOR2_X1 U23720 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22069), .ZN(n22059) );
  AOI22_X1 U23721 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n22061), .B1(
        n22060), .B2(n22059), .ZN(n22062) );
  OAI21_X1 U23722 ( .B1(n22063), .B2(n22100), .A(n22062), .ZN(n22064) );
  AOI21_X1 U23723 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22071), .A(n22064), 
        .ZN(n22067) );
  AOI22_X1 U23724 ( .A1(n22220), .A2(n22108), .B1(n22093), .B2(n22065), .ZN(
        n22066) );
  OAI211_X1 U23725 ( .C1(n22068), .C2(n22096), .A(n22067), .B(n22066), .ZN(
        P1_U2819) );
  NOR3_X1 U23726 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n22070), .A3(n22069), 
        .ZN(n22078) );
  AOI21_X1 U23727 ( .B1(n22073), .B2(n22072), .A(n22071), .ZN(n22076) );
  OAI22_X1 U23728 ( .A1(n22076), .A2(n22075), .B1(n22074), .B2(n22098), .ZN(
        n22077) );
  AOI211_X1 U23729 ( .C1(n22079), .C2(P1_EBX_REG_22__SCAN_IN), .A(n22078), .B(
        n22077), .ZN(n22082) );
  AOI22_X1 U23730 ( .A1(n22224), .A2(n22108), .B1(n22080), .B2(n22107), .ZN(
        n22081) );
  OAI211_X1 U23731 ( .C1(n22111), .C2(n22083), .A(n22082), .B(n22081), .ZN(
        P1_U2818) );
  NOR2_X1 U23732 ( .A1(n22085), .A2(n22084), .ZN(n22105) );
  NAND2_X1 U23733 ( .A1(n22087), .A2(n22086), .ZN(n22091) );
  INV_X1 U23734 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n22088) );
  OAI22_X1 U23735 ( .A1(n22089), .A2(n22100), .B1(n22088), .B2(n22098), .ZN(
        n22090) );
  AOI21_X1 U23736 ( .B1(n22105), .B2(n22091), .A(n22090), .ZN(n22095) );
  AOI22_X1 U23737 ( .A1(n11248), .A2(n22108), .B1(n22093), .B2(n22092), .ZN(
        n22094) );
  OAI211_X1 U23738 ( .C1(n22097), .C2(n22096), .A(n22095), .B(n22094), .ZN(
        P1_U2817) );
  OAI22_X1 U23739 ( .A1(n22101), .A2(n22100), .B1(n22099), .B2(n22098), .ZN(
        n22102) );
  AOI221_X1 U23740 ( .B1(n22105), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n22104), 
        .C2(n22103), .A(n22102), .ZN(n22110) );
  AOI22_X1 U23741 ( .A1(n22380), .A2(n22108), .B1(n22107), .B2(n22106), .ZN(
        n22109) );
  OAI211_X1 U23742 ( .C1(n22112), .C2(n22111), .A(n22110), .B(n22109), .ZN(
        P1_U2816) );
  OAI21_X1 U23743 ( .B1(n22114), .B2(n14602), .A(n22113), .ZN(P1_U2806) );
  AOI22_X1 U23744 ( .A1(n22117), .A2(n22116), .B1(n22115), .B2(n22129), .ZN(
        n22118) );
  INV_X1 U23745 ( .A(n22118), .ZN(n22120) );
  MUX2_X1 U23746 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n22120), .S(
        n22119), .Z(P1_U3469) );
  NOR2_X1 U23747 ( .A1(n22122), .A2(n22121), .ZN(n22124) );
  OAI21_X1 U23748 ( .B1(n22124), .B2(n22253), .A(n22123), .ZN(P1_U3163) );
  OAI211_X1 U23749 ( .C1(n22316), .C2(n22127), .A(n22126), .B(n22125), .ZN(
        P1_U3466) );
  INV_X1 U23750 ( .A(n22127), .ZN(n22128) );
  AOI21_X1 U23751 ( .B1(n22130), .B2(n22129), .A(n22128), .ZN(n22131) );
  OAI22_X1 U23752 ( .A1(n22133), .A2(n22132), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22131), .ZN(n22134) );
  OAI21_X1 U23753 ( .B1(n22136), .B2(n22135), .A(n22134), .ZN(P1_U3161) );
  AOI21_X1 U23754 ( .B1(n17357), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n22138), 
        .ZN(n22137) );
  INV_X1 U23755 ( .A(n22137), .ZN(P1_U2805) );
  AOI21_X1 U23756 ( .B1(n17357), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n22138), 
        .ZN(n22139) );
  INV_X1 U23757 ( .A(n22139), .ZN(P1_U3465) );
  INV_X1 U23758 ( .A(n22140), .ZN(n22142) );
  OAI21_X1 U23759 ( .B1(n22144), .B2(n22141), .A(n22142), .ZN(P2_U2818) );
  OAI21_X1 U23760 ( .B1(n22144), .B2(n22143), .A(n22142), .ZN(P2_U3592) );
  INV_X1 U23761 ( .A(n22145), .ZN(n22147) );
  OAI21_X1 U23762 ( .B1(n22149), .B2(n22146), .A(n22147), .ZN(P3_U2636) );
  OAI21_X1 U23763 ( .B1(n22149), .B2(n22148), .A(n22147), .ZN(P3_U3281) );
  INV_X1 U23764 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22197) );
  AOI21_X1 U23765 ( .B1(HOLD), .B2(n22150), .A(n22197), .ZN(n22152) );
  AOI21_X1 U23766 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22206), .A(n22196), 
        .ZN(n22213) );
  OAI21_X1 U23767 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n22175), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n22212) );
  INV_X1 U23768 ( .A(n22212), .ZN(n22151) );
  OAI22_X1 U23769 ( .A1(n22153), .A2(n22152), .B1(n22213), .B2(n22151), .ZN(
        P3_U3029) );
  AOI21_X1 U23770 ( .B1(n22165), .B2(n22175), .A(n22164), .ZN(n22159) );
  OAI211_X1 U23771 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n22160), .A(HOLD), .B(
        P1_STATE_REG_0__SCAN_IN), .ZN(n22158) );
  NAND2_X1 U23772 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22165), .ZN(n22162) );
  OAI21_X1 U23773 ( .B1(n22160), .B2(n22162), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n22155) );
  NAND3_X1 U23774 ( .A1(n22155), .A2(n22175), .A3(n22154), .ZN(n22157) );
  OAI211_X1 U23775 ( .C1(n22165), .C2(n22169), .A(P1_STATE_REG_2__SCAN_IN), 
        .B(P1_STATE_REG_1__SCAN_IN), .ZN(n22156) );
  OAI211_X1 U23776 ( .C1(n22159), .C2(n22158), .A(n22157), .B(n22156), .ZN(
        P1_U3196) );
  NAND2_X1 U23777 ( .A1(HOLD), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22166) );
  AOI21_X1 U23778 ( .B1(HOLD), .B2(P1_STATE_REG_2__SCAN_IN), .A(n22160), .ZN(
        n22167) );
  AOI21_X1 U23779 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n22167), .A(n22161), 
        .ZN(n22163) );
  OAI211_X1 U23780 ( .C1(n22164), .C2(n22166), .A(n22163), .B(n22162), .ZN(
        P1_U3195) );
  AOI21_X1 U23781 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22165), .A(n22169), 
        .ZN(n22171) );
  NAND2_X1 U23782 ( .A1(n22167), .A2(n22166), .ZN(n22168) );
  AOI21_X1 U23783 ( .B1(NA), .B2(n22169), .A(n22168), .ZN(n22170) );
  OAI22_X1 U23784 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22171), .B1(n20459), 
        .B2(n22170), .ZN(P1_U3194) );
  INV_X1 U23785 ( .A(HOLD), .ZN(n22195) );
  NOR2_X1 U23786 ( .A1(n22172), .A2(n22195), .ZN(n22178) );
  NOR2_X1 U23787 ( .A1(n22174), .A2(n22173), .ZN(n22186) );
  NOR2_X1 U23788 ( .A1(n22186), .A2(n22191), .ZN(n22193) );
  INV_X1 U23789 ( .A(n22193), .ZN(n22176) );
  OAI21_X1 U23790 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n22175), .A(
        P2_STATE_REG_2__SCAN_IN), .ZN(n22192) );
  AOI22_X1 U23791 ( .A1(n22178), .A2(n22177), .B1(n22176), .B2(n22192), .ZN(
        n22179) );
  OAI21_X1 U23792 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n22180), .A(n22179), .ZN(P2_U3209) );
  NOR2_X1 U23793 ( .A1(n22181), .A2(n22195), .ZN(n22189) );
  NAND2_X1 U23794 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22185) );
  AOI211_X1 U23795 ( .C1(n22183), .C2(HOLD), .A(n22186), .B(n22182), .ZN(
        n22184) );
  OAI21_X1 U23796 ( .B1(n22189), .B2(n22185), .A(n22184), .ZN(P2_U3210) );
  INV_X1 U23797 ( .A(n22186), .ZN(n22187) );
  OAI22_X1 U23798 ( .A1(NA), .A2(n22187), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22188) );
  OAI22_X1 U23799 ( .A1(n22189), .A2(n22188), .B1(HOLD), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22190) );
  OAI22_X1 U23800 ( .A1(n22193), .A2(n22192), .B1(n22191), .B2(n22190), .ZN(
        P2_U3211) );
  NOR2_X1 U23801 ( .A1(n22195), .A2(n22194), .ZN(n22209) );
  NOR3_X1 U23802 ( .A1(n22209), .A2(n22197), .A3(n22196), .ZN(n22198) );
  NOR2_X1 U23803 ( .A1(n22199), .A2(n22198), .ZN(n22202) );
  NOR2_X1 U23804 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22211)
         );
  AOI221_X1 U23805 ( .B1(n22209), .B2(n22204), .C1(n22211), .C2(n22204), .A(
        n22199), .ZN(n22200) );
  INV_X1 U23806 ( .A(n22200), .ZN(n22201) );
  MUX2_X1 U23807 ( .A(n22202), .B(n22201), .S(P3_STATE_REG_1__SCAN_IN), .Z(
        n22203) );
  OAI221_X1 U23808 ( .B1(n22205), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n22205), 
        .C2(n22204), .A(n22203), .ZN(P3_U3030) );
  NAND2_X1 U23809 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n22206), .ZN(n22207) );
  OAI22_X1 U23810 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n22207), .ZN(n22208) );
  OAI21_X1 U23811 ( .B1(n22209), .B2(n22208), .A(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n22210) );
  OAI22_X1 U23812 ( .A1(n22213), .A2(n22212), .B1(n22211), .B2(n22210), .ZN(
        P3_U3031) );
  INV_X1 U23813 ( .A(DATAI_17_), .ZN(n22390) );
  AOI22_X1 U23814 ( .A1(n22377), .A2(n22385), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n22375), .ZN(n22216) );
  AOI22_X1 U23815 ( .A1(n22214), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n22215) );
  OAI211_X1 U23816 ( .C1(n22390), .C2(n22383), .A(n22216), .B(n22215), .ZN(
        P1_U2887) );
  INV_X1 U23817 ( .A(DATAI_19_), .ZN(n22461) );
  AOI22_X1 U23818 ( .A1(n22377), .A2(n22456), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n22375), .ZN(n22219) );
  AOI22_X1 U23819 ( .A1(n22217), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n22218) );
  OAI211_X1 U23820 ( .C1(n22461), .C2(n22383), .A(n22219), .B(n22218), .ZN(
        P1_U2885) );
  INV_X1 U23821 ( .A(DATAI_21_), .ZN(n22532) );
  AOI22_X1 U23822 ( .A1(n22377), .A2(n22527), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n22375), .ZN(n22222) );
  AOI22_X1 U23823 ( .A1(n22220), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n22221) );
  OAI211_X1 U23824 ( .C1(n22532), .C2(n22383), .A(n22222), .B(n22221), .ZN(
        P1_U2883) );
  AOI22_X1 U23825 ( .A1(n22377), .A2(n22223), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n22375), .ZN(n22226) );
  AOI22_X1 U23826 ( .A1(n22224), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n22225) );
  OAI211_X1 U23827 ( .C1(n22227), .C2(n22383), .A(n22226), .B(n22225), .ZN(
        P1_U2882) );
  INV_X1 U23828 ( .A(DATAI_23_), .ZN(n22641) );
  AOI22_X1 U23829 ( .A1(n22377), .A2(n22631), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n22375), .ZN(n22229) );
  AOI22_X1 U23830 ( .A1(n11248), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n22228) );
  OAI211_X1 U23831 ( .C1(n22641), .C2(n22383), .A(n22229), .B(n22228), .ZN(
        P1_U2881) );
  INV_X1 U23832 ( .A(n22230), .ZN(n22231) );
  NAND3_X1 U23833 ( .A1(n22232), .A2(n22292), .A3(n22245), .ZN(n22233) );
  INV_X1 U23834 ( .A(n22337), .ZN(n22293) );
  NAND2_X1 U23835 ( .A1(n22233), .A2(n22293), .ZN(n22243) );
  NOR2_X1 U23836 ( .A1(n22250), .A2(n22354), .ZN(n22240) );
  INV_X1 U23837 ( .A(n22323), .ZN(n22234) );
  NOR2_X1 U23838 ( .A1(n22309), .A2(n22234), .ZN(n22279) );
  AOI22_X1 U23839 ( .A1(n22243), .A2(n22240), .B1(n22325), .B2(n22279), .ZN(
        n22645) );
  NAND2_X1 U23840 ( .A1(n22632), .A2(n22235), .ZN(n22350) );
  NOR2_X2 U23841 ( .A1(n22634), .A2(n22236), .ZN(n22370) );
  NAND3_X1 U23842 ( .A1(n22238), .A2(n13197), .A3(n22237), .ZN(n22254) );
  NOR2_X1 U23843 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22254), .ZN(
        n22637) );
  INV_X1 U23844 ( .A(DATAI_24_), .ZN(n22384) );
  AOI22_X1 U23845 ( .A1(n22370), .A2(n22637), .B1(n22743), .B2(n22365), .ZN(
        n22249) );
  INV_X1 U23846 ( .A(n22240), .ZN(n22242) );
  INV_X1 U23847 ( .A(n22637), .ZN(n22241) );
  AOI22_X1 U23848 ( .A1(n22243), .A2(n22242), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22241), .ZN(n22244) );
  OAI211_X1 U23849 ( .C1(n22279), .C2(n22253), .A(n22314), .B(n22244), .ZN(
        n22642) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22371), .ZN(n22248) );
  OAI211_X1 U23851 ( .C1(n22645), .C2(n22350), .A(n22249), .B(n22248), .ZN(
        P1_U3033) );
  INV_X1 U23852 ( .A(n22371), .ZN(n22368) );
  INV_X1 U23853 ( .A(n22250), .ZN(n22264) );
  NOR2_X1 U23854 ( .A1(n22251), .A2(n22254), .ZN(n22646) );
  AOI21_X1 U23855 ( .B1(n22264), .B2(n22252), .A(n22646), .ZN(n22255) );
  OAI22_X1 U23856 ( .A1(n22255), .A2(n22358), .B1(n22254), .B2(n22253), .ZN(
        n22647) );
  AOI22_X1 U23857 ( .A1(n22647), .A2(n22369), .B1(n22370), .B2(n22646), .ZN(
        n22259) );
  INV_X1 U23858 ( .A(n22254), .ZN(n22257) );
  OAI211_X1 U23859 ( .C1(n22275), .C2(n22282), .A(n22292), .B(n22255), .ZN(
        n22256) );
  OAI211_X1 U23860 ( .C1(n22292), .C2(n22257), .A(n22268), .B(n22256), .ZN(
        n22649) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22365), .ZN(n22258) );
  OAI211_X1 U23862 ( .C1(n22368), .C2(n22652), .A(n22259), .B(n22258), .ZN(
        P1_U3041) );
  INV_X1 U23863 ( .A(n22260), .ZN(n22653) );
  AOI22_X1 U23864 ( .A1(n22660), .A2(n22371), .B1(n22370), .B2(n22653), .ZN(
        n22262) );
  AOI22_X1 U23865 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22655), .B1(
        n22654), .B2(n22365), .ZN(n22261) );
  OAI211_X1 U23866 ( .C1(n22658), .C2(n22350), .A(n22262), .B(n22261), .ZN(
        P1_U3049) );
  AND2_X1 U23867 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22273), .ZN(
        n22659) );
  AOI21_X1 U23868 ( .B1(n22264), .B2(n22263), .A(n22659), .ZN(n22271) );
  INV_X1 U23869 ( .A(n22271), .ZN(n22267) );
  INV_X1 U23870 ( .A(n22275), .ZN(n22266) );
  AOI21_X1 U23871 ( .B1(n22266), .B2(n22265), .A(n22358), .ZN(n22270) );
  AOI22_X1 U23872 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22273), .B1(n22267), 
        .B2(n22270), .ZN(n22664) );
  AOI22_X1 U23873 ( .A1(n22660), .A2(n22365), .B1(n22370), .B2(n22659), .ZN(
        n22277) );
  INV_X1 U23874 ( .A(n22268), .ZN(n22269) );
  AOI21_X1 U23875 ( .B1(n22271), .B2(n22270), .A(n22269), .ZN(n22272) );
  OAI21_X1 U23876 ( .B1(n22292), .B2(n22273), .A(n22272), .ZN(n22661) );
  AOI22_X1 U23877 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22661), .B1(
        n22667), .B2(n22371), .ZN(n22276) );
  OAI211_X1 U23878 ( .C1(n22664), .C2(n22350), .A(n22277), .B(n22276), .ZN(
        P1_U3057) );
  NOR2_X1 U23879 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22278), .ZN(
        n22666) );
  INV_X1 U23880 ( .A(n22279), .ZN(n22281) );
  NAND3_X1 U23881 ( .A1(n22295), .A2(n22292), .A3(n22339), .ZN(n22280) );
  OAI21_X1 U23882 ( .B1(n22356), .B2(n22281), .A(n22280), .ZN(n22665) );
  AOI22_X1 U23883 ( .A1(n22370), .A2(n22666), .B1(n22665), .B2(n22369), .ZN(
        n22288) );
  AOI21_X1 U23884 ( .B1(n22671), .B2(n22577), .A(n22282), .ZN(n22283) );
  AOI21_X1 U23885 ( .B1(n22295), .B2(n22339), .A(n22283), .ZN(n22284) );
  NOR2_X1 U23886 ( .A1(n22284), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22286) );
  AOI22_X1 U23887 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22365), .ZN(n22287) );
  OAI211_X1 U23888 ( .C1(n22368), .C2(n22671), .A(n22288), .B(n22287), .ZN(
        P1_U3065) );
  INV_X1 U23889 ( .A(n22365), .ZN(n22374) );
  AOI22_X1 U23890 ( .A1(n22370), .A2(n22673), .B1(n22672), .B2(n22369), .ZN(
        n22290) );
  AOI22_X1 U23891 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22675), .B1(
        n22583), .B2(n22371), .ZN(n22289) );
  OAI211_X1 U23892 ( .C1(n22374), .C2(n22671), .A(n22290), .B(n22289), .ZN(
        P1_U3073) );
  NOR2_X1 U23893 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22291), .ZN(
        n22678) );
  AOI22_X1 U23894 ( .A1(n22583), .A2(n22365), .B1(n22370), .B2(n22678), .ZN(
        n22304) );
  NAND3_X1 U23895 ( .A1(n22593), .A2(n22683), .A3(n22292), .ZN(n22294) );
  NAND2_X1 U23896 ( .A1(n22294), .A2(n22293), .ZN(n22299) );
  NAND2_X1 U23897 ( .A1(n22295), .A2(n22354), .ZN(n22301) );
  INV_X1 U23898 ( .A(n22678), .ZN(n22296) );
  AOI22_X1 U23899 ( .A1(n22299), .A2(n22301), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22296), .ZN(n22298) );
  NAND3_X1 U23900 ( .A1(n22362), .A2(n22298), .A3(n22297), .ZN(n22680) );
  INV_X1 U23901 ( .A(n22299), .ZN(n22302) );
  OAI22_X1 U23902 ( .A1(n22302), .A2(n22301), .B1(n22300), .B2(n22356), .ZN(
        n22679) );
  AOI22_X1 U23903 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22680), .B1(
        n22369), .B2(n22679), .ZN(n22303) );
  OAI211_X1 U23904 ( .C1(n22368), .C2(n22593), .A(n22304), .B(n22303), .ZN(
        P1_U3081) );
  INV_X1 U23905 ( .A(n22588), .ZN(n22684) );
  AOI22_X1 U23906 ( .A1(n22685), .A2(n22370), .B1(n22684), .B2(n22369), .ZN(
        n22306) );
  AOI22_X1 U23907 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22687), .B1(
        n22693), .B2(n22371), .ZN(n22305) );
  OAI211_X1 U23908 ( .C1(n22374), .C2(n22593), .A(n22306), .B(n22305), .ZN(
        P1_U3089) );
  INV_X1 U23909 ( .A(n22322), .ZN(n22308) );
  NOR2_X1 U23910 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22307), .ZN(
        n22691) );
  AOI21_X1 U23911 ( .B1(n22308), .B2(n22339), .A(n22691), .ZN(n22312) );
  INV_X1 U23912 ( .A(n22325), .ZN(n22310) );
  NAND2_X1 U23913 ( .A1(n22309), .A2(n22323), .ZN(n22344) );
  OAI22_X1 U23914 ( .A1(n22312), .A2(n22358), .B1(n22310), .B2(n22344), .ZN(
        n22692) );
  AOI22_X1 U23915 ( .A1(n22692), .A2(n22369), .B1(n22370), .B2(n22691), .ZN(
        n22318) );
  OAI21_X1 U23916 ( .B1(n22311), .B2(n22693), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22313) );
  NAND2_X1 U23917 ( .A1(n22313), .A2(n22312), .ZN(n22315) );
  AOI22_X1 U23918 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22365), .ZN(n22317) );
  OAI211_X1 U23919 ( .C1(n22368), .C2(n22702), .A(n22318), .B(n22317), .ZN(
        P1_U3097) );
  AOI22_X1 U23920 ( .A1(n22370), .A2(n22698), .B1(n22697), .B2(n22369), .ZN(
        n22320) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22371), .ZN(n22319) );
  OAI211_X1 U23922 ( .C1(n22374), .C2(n22702), .A(n22320), .B(n22319), .ZN(
        P1_U3105) );
  NOR3_X1 U23923 ( .A1(n22704), .A2(n22705), .A3(n22358), .ZN(n22321) );
  NOR2_X1 U23924 ( .A1(n22321), .A2(n22337), .ZN(n22332) );
  INV_X1 U23925 ( .A(n22332), .ZN(n22326) );
  NOR2_X1 U23926 ( .A1(n22322), .A2(n22339), .ZN(n22331) );
  OR2_X1 U23927 ( .A1(n22323), .A2(n13197), .ZN(n22357) );
  INV_X1 U23928 ( .A(n22357), .ZN(n22324) );
  NOR2_X1 U23929 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22327), .ZN(
        n22703) );
  AOI22_X1 U23930 ( .A1(n22705), .A2(n22365), .B1(n22370), .B2(n22703), .ZN(
        n22334) );
  INV_X1 U23931 ( .A(n22703), .ZN(n22598) );
  NAND2_X1 U23932 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22357), .ZN(n22363) );
  INV_X1 U23933 ( .A(n22363), .ZN(n22328) );
  AOI211_X1 U23934 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22598), .A(n22329), 
        .B(n22328), .ZN(n22330) );
  OAI21_X1 U23935 ( .B1(n22332), .B2(n22331), .A(n22330), .ZN(n22706) );
  AOI22_X1 U23936 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22706), .B1(
        n22704), .B2(n22371), .ZN(n22333) );
  OAI211_X1 U23937 ( .C1(n22709), .C2(n22350), .A(n22334), .B(n22333), .ZN(
        P1_U3113) );
  INV_X1 U23938 ( .A(n22602), .ZN(n22710) );
  AOI22_X1 U23939 ( .A1(n22370), .A2(n22711), .B1(n22710), .B2(n22369), .ZN(
        n22336) );
  AOI22_X1 U23940 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22371), .ZN(n22335) );
  OAI211_X1 U23941 ( .C1(n22374), .C2(n22715), .A(n22336), .B(n22335), .ZN(
        P1_U3121) );
  NOR3_X1 U23942 ( .A1(n22718), .A2(n22717), .A3(n22358), .ZN(n22338) );
  NOR2_X1 U23943 ( .A1(n22338), .A2(n22337), .ZN(n22347) );
  INV_X1 U23944 ( .A(n22347), .ZN(n22342) );
  AND2_X1 U23945 ( .A1(n22355), .A2(n22339), .ZN(n22346) );
  INV_X1 U23946 ( .A(n22356), .ZN(n22341) );
  INV_X1 U23947 ( .A(n22344), .ZN(n22340) );
  NOR2_X1 U23948 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22343), .ZN(
        n22716) );
  AOI22_X1 U23949 ( .A1(n22717), .A2(n22371), .B1(n22370), .B2(n22716), .ZN(
        n22349) );
  INV_X1 U23950 ( .A(n22716), .ZN(n22607) );
  AOI22_X1 U23951 ( .A1(n22344), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n22607), .ZN(n22345) );
  OAI211_X1 U23952 ( .C1(n22347), .C2(n22346), .A(n22362), .B(n22345), .ZN(
        n22719) );
  AOI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22365), .ZN(n22348) );
  OAI211_X1 U23954 ( .C1(n22723), .C2(n22350), .A(n22349), .B(n22348), .ZN(
        P1_U3129) );
  INV_X1 U23955 ( .A(n22611), .ZN(n22724) );
  AOI22_X1 U23956 ( .A1(n22370), .A2(n22725), .B1(n22724), .B2(n22369), .ZN(
        n22352) );
  AOI22_X1 U23957 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22371), .ZN(n22351) );
  OAI211_X1 U23958 ( .C1(n22374), .C2(n22729), .A(n22352), .B(n22351), .ZN(
        P1_U3137) );
  NOR2_X1 U23959 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22353), .ZN(
        n22731) );
  NAND2_X1 U23960 ( .A1(n22355), .A2(n22354), .ZN(n22360) );
  OAI22_X1 U23961 ( .A1(n22360), .A2(n22358), .B1(n22357), .B2(n22356), .ZN(
        n22730) );
  AOI22_X1 U23962 ( .A1(n22370), .A2(n22731), .B1(n22730), .B2(n22369), .ZN(
        n22367) );
  OAI21_X1 U23963 ( .B1(n22359), .B2(n22733), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n22361) );
  AOI21_X1 U23964 ( .B1(n22361), .B2(n22360), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n22364) );
  OAI211_X1 U23965 ( .C1(n22364), .C2(n22731), .A(n22363), .B(n22362), .ZN(
        n22734) );
  AOI22_X1 U23966 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22365), .ZN(n22366) );
  OAI211_X1 U23967 ( .C1(n22368), .C2(n22747), .A(n22367), .B(n22366), .ZN(
        P1_U3145) );
  INV_X1 U23968 ( .A(n22622), .ZN(n22739) );
  AOI22_X1 U23969 ( .A1(n22741), .A2(n22370), .B1(n22739), .B2(n22369), .ZN(
        n22373) );
  AOI22_X1 U23970 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22371), .ZN(n22372) );
  OAI211_X1 U23971 ( .C1(n22374), .C2(n22747), .A(n22373), .B(n22372), .ZN(
        P1_U3153) );
  AOI22_X1 U23972 ( .A1(n22377), .A2(n22376), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n22375), .ZN(n22382) );
  AOI22_X1 U23973 ( .A1(n22380), .A2(n22379), .B1(n22378), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n22381) );
  OAI211_X1 U23974 ( .C1(n22384), .C2(n22383), .A(n22382), .B(n22381), .ZN(
        P1_U2880) );
  NAND2_X1 U23975 ( .A1(n22632), .A2(n22385), .ZN(n22417) );
  NOR2_X2 U23976 ( .A1(n22634), .A2(n22386), .ZN(n22425) );
  AOI22_X1 U23977 ( .A1(n22425), .A2(n22637), .B1(n22743), .B2(n22420), .ZN(
        n22392) );
  AOI22_X1 U23978 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22426), .ZN(n22391) );
  OAI211_X1 U23979 ( .C1(n22645), .C2(n22417), .A(n22392), .B(n22391), .ZN(
        P1_U3034) );
  INV_X1 U23980 ( .A(n22426), .ZN(n22423) );
  AOI22_X1 U23981 ( .A1(n22647), .A2(n22424), .B1(n22425), .B2(n22646), .ZN(
        n22394) );
  AOI22_X1 U23982 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22420), .ZN(n22393) );
  OAI211_X1 U23983 ( .C1(n22423), .C2(n22652), .A(n22394), .B(n22393), .ZN(
        P1_U3042) );
  AOI22_X1 U23984 ( .A1(n22654), .A2(n22420), .B1(n22425), .B2(n22653), .ZN(
        n22396) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22655), .B1(
        n22660), .B2(n22426), .ZN(n22395) );
  OAI211_X1 U23986 ( .C1(n22658), .C2(n22417), .A(n22396), .B(n22395), .ZN(
        P1_U3050) );
  AOI22_X1 U23987 ( .A1(n22660), .A2(n22420), .B1(n22425), .B2(n22659), .ZN(
        n22398) );
  AOI22_X1 U23988 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22661), .B1(
        n22667), .B2(n22426), .ZN(n22397) );
  OAI211_X1 U23989 ( .C1(n22664), .C2(n22417), .A(n22398), .B(n22397), .ZN(
        P1_U3058) );
  AOI22_X1 U23990 ( .A1(n22425), .A2(n22666), .B1(n22665), .B2(n22424), .ZN(
        n22400) );
  AOI22_X1 U23991 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22420), .ZN(n22399) );
  OAI211_X1 U23992 ( .C1(n22423), .C2(n22671), .A(n22400), .B(n22399), .ZN(
        P1_U3066) );
  AOI22_X1 U23993 ( .A1(n22425), .A2(n22673), .B1(n22672), .B2(n22424), .ZN(
        n22402) );
  AOI22_X1 U23994 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22675), .B1(
        n22674), .B2(n22420), .ZN(n22401) );
  OAI211_X1 U23995 ( .C1(n22423), .C2(n22683), .A(n22402), .B(n22401), .ZN(
        P1_U3074) );
  AOI22_X1 U23996 ( .A1(n22583), .A2(n22420), .B1(n22425), .B2(n22678), .ZN(
        n22404) );
  AOI22_X1 U23997 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22680), .B1(
        n22424), .B2(n22679), .ZN(n22403) );
  OAI211_X1 U23998 ( .C1(n22423), .C2(n22593), .A(n22404), .B(n22403), .ZN(
        P1_U3082) );
  INV_X1 U23999 ( .A(n22420), .ZN(n22429) );
  AOI22_X1 U24000 ( .A1(n22685), .A2(n22425), .B1(n22684), .B2(n22424), .ZN(
        n22406) );
  AOI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22687), .B1(
        n22693), .B2(n22426), .ZN(n22405) );
  OAI211_X1 U24002 ( .C1(n22429), .C2(n22593), .A(n22406), .B(n22405), .ZN(
        P1_U3090) );
  AOI22_X1 U24003 ( .A1(n22692), .A2(n22424), .B1(n22425), .B2(n22691), .ZN(
        n22408) );
  AOI22_X1 U24004 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22420), .ZN(n22407) );
  OAI211_X1 U24005 ( .C1(n22423), .C2(n22702), .A(n22408), .B(n22407), .ZN(
        P1_U3098) );
  AOI22_X1 U24006 ( .A1(n22425), .A2(n22698), .B1(n22697), .B2(n22424), .ZN(
        n22410) );
  AOI22_X1 U24007 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22426), .ZN(n22409) );
  OAI211_X1 U24008 ( .C1(n22429), .C2(n22702), .A(n22410), .B(n22409), .ZN(
        P1_U3106) );
  AOI22_X1 U24009 ( .A1(n22704), .A2(n22426), .B1(n22425), .B2(n22703), .ZN(
        n22412) );
  AOI22_X1 U24010 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22706), .B1(
        n22705), .B2(n22420), .ZN(n22411) );
  OAI211_X1 U24011 ( .C1(n22709), .C2(n22417), .A(n22412), .B(n22411), .ZN(
        P1_U3114) );
  AOI22_X1 U24012 ( .A1(n22425), .A2(n22711), .B1(n22710), .B2(n22424), .ZN(
        n22414) );
  AOI22_X1 U24013 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22426), .ZN(n22413) );
  OAI211_X1 U24014 ( .C1(n22429), .C2(n22715), .A(n22414), .B(n22413), .ZN(
        P1_U3122) );
  AOI22_X1 U24015 ( .A1(n22717), .A2(n22426), .B1(n22425), .B2(n22716), .ZN(
        n22416) );
  AOI22_X1 U24016 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22420), .ZN(n22415) );
  OAI211_X1 U24017 ( .C1(n22723), .C2(n22417), .A(n22416), .B(n22415), .ZN(
        P1_U3130) );
  AOI22_X1 U24018 ( .A1(n22425), .A2(n22725), .B1(n22724), .B2(n22424), .ZN(
        n22419) );
  AOI22_X1 U24019 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22426), .ZN(n22418) );
  OAI211_X1 U24020 ( .C1(n22429), .C2(n22729), .A(n22419), .B(n22418), .ZN(
        P1_U3138) );
  AOI22_X1 U24021 ( .A1(n22425), .A2(n22731), .B1(n22730), .B2(n22424), .ZN(
        n22422) );
  AOI22_X1 U24022 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22420), .ZN(n22421) );
  OAI211_X1 U24023 ( .C1(n22423), .C2(n22747), .A(n22422), .B(n22421), .ZN(
        P1_U3146) );
  AOI22_X1 U24024 ( .A1(n22741), .A2(n22425), .B1(n22739), .B2(n22424), .ZN(
        n22428) );
  AOI22_X1 U24025 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22426), .ZN(n22427) );
  OAI211_X1 U24026 ( .C1(n22429), .C2(n22747), .A(n22428), .B(n22427), .ZN(
        P1_U3154) );
  AOI22_X1 U24027 ( .A1(n22637), .A2(n22451), .B1(n22743), .B2(n22452), .ZN(
        n22431) );
  AOI22_X1 U24028 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22446), .ZN(n22430) );
  OAI211_X1 U24029 ( .C1(n22645), .C2(n22449), .A(n22431), .B(n22430), .ZN(
        P1_U3035) );
  AOI22_X1 U24030 ( .A1(n22450), .A2(n22647), .B1(n22451), .B2(n22646), .ZN(
        n22433) );
  AOI22_X1 U24031 ( .A1(n22649), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n22648), .B2(n22452), .ZN(n22432) );
  OAI211_X1 U24032 ( .C1(n22455), .C2(n22652), .A(n22433), .B(n22432), .ZN(
        P1_U3043) );
  AOI22_X1 U24033 ( .A1(n22660), .A2(n22446), .B1(n22451), .B2(n22653), .ZN(
        n22435) );
  AOI22_X1 U24034 ( .A1(n22655), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22654), .B2(n22452), .ZN(n22434) );
  OAI211_X1 U24035 ( .C1(n22658), .C2(n22449), .A(n22435), .B(n22434), .ZN(
        P1_U3051) );
  AOI22_X1 U24036 ( .A1(n22660), .A2(n22452), .B1(n22451), .B2(n22659), .ZN(
        n22437) );
  AOI22_X1 U24037 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22661), .B1(
        n22667), .B2(n22446), .ZN(n22436) );
  OAI211_X1 U24038 ( .C1(n22664), .C2(n22449), .A(n22437), .B(n22436), .ZN(
        P1_U3059) );
  AOI22_X1 U24039 ( .A1(n22451), .A2(n22666), .B1(n22450), .B2(n22665), .ZN(
        n22439) );
  AOI22_X1 U24040 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n22667), .B2(n22452), .ZN(n22438) );
  OAI211_X1 U24041 ( .C1(n22455), .C2(n22671), .A(n22439), .B(n22438), .ZN(
        P1_U3067) );
  AOI22_X1 U24042 ( .A1(n22583), .A2(n22452), .B1(n22451), .B2(n22678), .ZN(
        n22441) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22680), .B1(
        n22450), .B2(n22679), .ZN(n22440) );
  OAI211_X1 U24044 ( .C1(n22455), .C2(n22593), .A(n22441), .B(n22440), .ZN(
        P1_U3083) );
  AOI22_X1 U24045 ( .A1(n22450), .A2(n22692), .B1(n22451), .B2(n22691), .ZN(
        n22443) );
  AOI22_X1 U24046 ( .A1(n22694), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22693), .B2(n22452), .ZN(n22442) );
  OAI211_X1 U24047 ( .C1(n22455), .C2(n22702), .A(n22443), .B(n22442), .ZN(
        P1_U3099) );
  AOI22_X1 U24048 ( .A1(n22705), .A2(n22452), .B1(n22703), .B2(n22451), .ZN(
        n22445) );
  AOI22_X1 U24049 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22706), .B1(
        n22704), .B2(n22446), .ZN(n22444) );
  OAI211_X1 U24050 ( .C1(n22709), .C2(n22449), .A(n22445), .B(n22444), .ZN(
        P1_U3115) );
  AOI22_X1 U24051 ( .A1(n22717), .A2(n22446), .B1(n22451), .B2(n22716), .ZN(
        n22448) );
  AOI22_X1 U24052 ( .A1(n22719), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22718), .B2(n22452), .ZN(n22447) );
  OAI211_X1 U24053 ( .C1(n22723), .C2(n22449), .A(n22448), .B(n22447), .ZN(
        P1_U3131) );
  AOI22_X1 U24054 ( .A1(n22451), .A2(n22731), .B1(n22450), .B2(n22730), .ZN(
        n22454) );
  AOI22_X1 U24055 ( .A1(n22734), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n22733), .B2(n22452), .ZN(n22453) );
  OAI211_X1 U24056 ( .C1(n22455), .C2(n22747), .A(n22454), .B(n22453), .ZN(
        P1_U3147) );
  NAND2_X1 U24057 ( .A1(n22632), .A2(n22456), .ZN(n22488) );
  NOR2_X2 U24058 ( .A1(n22634), .A2(n22457), .ZN(n22496) );
  AOI22_X1 U24059 ( .A1(n22496), .A2(n22637), .B1(n22743), .B2(n22491), .ZN(
        n22463) );
  OAI22_X1 U24060 ( .A1(n22461), .A2(n22640), .B1(n22639), .B2(n22460), .ZN(
        n22497) );
  AOI22_X1 U24061 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22497), .ZN(n22462) );
  OAI211_X1 U24062 ( .C1(n22645), .C2(n22488), .A(n22463), .B(n22462), .ZN(
        P1_U3036) );
  INV_X1 U24063 ( .A(n22497), .ZN(n22494) );
  AOI22_X1 U24064 ( .A1(n22647), .A2(n22495), .B1(n22496), .B2(n22646), .ZN(
        n22465) );
  AOI22_X1 U24065 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22491), .ZN(n22464) );
  OAI211_X1 U24066 ( .C1(n22494), .C2(n22652), .A(n22465), .B(n22464), .ZN(
        P1_U3044) );
  AOI22_X1 U24067 ( .A1(n22654), .A2(n22491), .B1(n22496), .B2(n22653), .ZN(
        n22467) );
  AOI22_X1 U24068 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22655), .B1(
        n22660), .B2(n22497), .ZN(n22466) );
  OAI211_X1 U24069 ( .C1(n22658), .C2(n22488), .A(n22467), .B(n22466), .ZN(
        P1_U3052) );
  AOI22_X1 U24070 ( .A1(n22667), .A2(n22497), .B1(n22496), .B2(n22659), .ZN(
        n22469) );
  AOI22_X1 U24071 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22661), .B1(
        n22660), .B2(n22491), .ZN(n22468) );
  OAI211_X1 U24072 ( .C1(n22664), .C2(n22488), .A(n22469), .B(n22468), .ZN(
        P1_U3060) );
  AOI22_X1 U24073 ( .A1(n22496), .A2(n22666), .B1(n22665), .B2(n22495), .ZN(
        n22471) );
  AOI22_X1 U24074 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22491), .ZN(n22470) );
  OAI211_X1 U24075 ( .C1(n22494), .C2(n22671), .A(n22471), .B(n22470), .ZN(
        P1_U3068) );
  AOI22_X1 U24076 ( .A1(n22496), .A2(n22673), .B1(n22672), .B2(n22495), .ZN(
        n22473) );
  AOI22_X1 U24077 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22675), .B1(
        n22674), .B2(n22491), .ZN(n22472) );
  OAI211_X1 U24078 ( .C1(n22494), .C2(n22683), .A(n22473), .B(n22472), .ZN(
        P1_U3076) );
  AOI22_X1 U24079 ( .A1(n22583), .A2(n22491), .B1(n22496), .B2(n22678), .ZN(
        n22475) );
  AOI22_X1 U24080 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22680), .B1(
        n22495), .B2(n22679), .ZN(n22474) );
  OAI211_X1 U24081 ( .C1(n22494), .C2(n22593), .A(n22475), .B(n22474), .ZN(
        P1_U3084) );
  AOI22_X1 U24082 ( .A1(n22685), .A2(n22496), .B1(n22684), .B2(n22495), .ZN(
        n22477) );
  AOI22_X1 U24083 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22687), .B1(
        n22686), .B2(n22491), .ZN(n22476) );
  OAI211_X1 U24084 ( .C1(n22494), .C2(n22690), .A(n22477), .B(n22476), .ZN(
        P1_U3092) );
  AOI22_X1 U24085 ( .A1(n22692), .A2(n22495), .B1(n22496), .B2(n22691), .ZN(
        n22479) );
  AOI22_X1 U24086 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22491), .ZN(n22478) );
  OAI211_X1 U24087 ( .C1(n22494), .C2(n22702), .A(n22479), .B(n22478), .ZN(
        P1_U3100) );
  INV_X1 U24088 ( .A(n22491), .ZN(n22500) );
  AOI22_X1 U24089 ( .A1(n22496), .A2(n22698), .B1(n22697), .B2(n22495), .ZN(
        n22481) );
  AOI22_X1 U24090 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22497), .ZN(n22480) );
  OAI211_X1 U24091 ( .C1(n22500), .C2(n22702), .A(n22481), .B(n22480), .ZN(
        P1_U3108) );
  AOI22_X1 U24092 ( .A1(n22704), .A2(n22497), .B1(n22496), .B2(n22703), .ZN(
        n22483) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22706), .B1(
        n22705), .B2(n22491), .ZN(n22482) );
  OAI211_X1 U24094 ( .C1(n22709), .C2(n22488), .A(n22483), .B(n22482), .ZN(
        P1_U3116) );
  AOI22_X1 U24095 ( .A1(n22496), .A2(n22711), .B1(n22710), .B2(n22495), .ZN(
        n22485) );
  AOI22_X1 U24096 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22497), .ZN(n22484) );
  OAI211_X1 U24097 ( .C1(n22500), .C2(n22715), .A(n22485), .B(n22484), .ZN(
        P1_U3124) );
  AOI22_X1 U24098 ( .A1(n22717), .A2(n22497), .B1(n22496), .B2(n22716), .ZN(
        n22487) );
  AOI22_X1 U24099 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22491), .ZN(n22486) );
  OAI211_X1 U24100 ( .C1(n22723), .C2(n22488), .A(n22487), .B(n22486), .ZN(
        P1_U3132) );
  AOI22_X1 U24101 ( .A1(n22496), .A2(n22725), .B1(n22724), .B2(n22495), .ZN(
        n22490) );
  AOI22_X1 U24102 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22497), .ZN(n22489) );
  OAI211_X1 U24103 ( .C1(n22500), .C2(n22729), .A(n22490), .B(n22489), .ZN(
        P1_U3140) );
  AOI22_X1 U24104 ( .A1(n22496), .A2(n22731), .B1(n22730), .B2(n22495), .ZN(
        n22493) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22491), .ZN(n22492) );
  OAI211_X1 U24106 ( .C1(n22494), .C2(n22747), .A(n22493), .B(n22492), .ZN(
        P1_U3148) );
  AOI22_X1 U24107 ( .A1(n22741), .A2(n22496), .B1(n22739), .B2(n22495), .ZN(
        n22499) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22497), .ZN(n22498) );
  OAI211_X1 U24109 ( .C1(n22500), .C2(n22747), .A(n22499), .B(n22498), .ZN(
        P1_U3156) );
  AOI22_X1 U24110 ( .A1(n22521), .A2(n22637), .B1(n22743), .B2(n22523), .ZN(
        n22502) );
  AOI22_X1 U24111 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22517), .ZN(n22501) );
  OAI211_X1 U24112 ( .C1(n22645), .C2(n22520), .A(n22502), .B(n22501), .ZN(
        P1_U3037) );
  AOI22_X1 U24113 ( .A1(n22522), .A2(n22647), .B1(n22521), .B2(n22646), .ZN(
        n22504) );
  AOI22_X1 U24114 ( .A1(n22649), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n22648), .B2(n22523), .ZN(n22503) );
  OAI211_X1 U24115 ( .C1(n22526), .C2(n22652), .A(n22504), .B(n22503), .ZN(
        P1_U3045) );
  AOI22_X1 U24116 ( .A1(n22654), .A2(n22523), .B1(n22521), .B2(n22653), .ZN(
        n22506) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22655), .B1(
        n22660), .B2(n22517), .ZN(n22505) );
  OAI211_X1 U24118 ( .C1(n22658), .C2(n22520), .A(n22506), .B(n22505), .ZN(
        P1_U3053) );
  AOI22_X1 U24119 ( .A1(n22517), .A2(n22667), .B1(n22521), .B2(n22659), .ZN(
        n22508) );
  AOI22_X1 U24120 ( .A1(n22661), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22660), .B2(n22523), .ZN(n22507) );
  OAI211_X1 U24121 ( .C1(n22664), .C2(n22520), .A(n22508), .B(n22507), .ZN(
        P1_U3061) );
  AOI22_X1 U24122 ( .A1(n22522), .A2(n22665), .B1(n22521), .B2(n22666), .ZN(
        n22510) );
  AOI22_X1 U24123 ( .A1(n22668), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n22667), .B2(n22523), .ZN(n22509) );
  OAI211_X1 U24124 ( .C1(n22526), .C2(n22671), .A(n22510), .B(n22509), .ZN(
        P1_U3069) );
  AOI22_X1 U24125 ( .A1(n22521), .A2(n22678), .B1(n22583), .B2(n22523), .ZN(
        n22512) );
  AOI22_X1 U24126 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22680), .B1(
        n22522), .B2(n22679), .ZN(n22511) );
  OAI211_X1 U24127 ( .C1(n22526), .C2(n22593), .A(n22512), .B(n22511), .ZN(
        P1_U3085) );
  AOI22_X1 U24128 ( .A1(n22522), .A2(n22692), .B1(n22521), .B2(n22691), .ZN(
        n22514) );
  AOI22_X1 U24129 ( .A1(n22694), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22693), .B2(n22523), .ZN(n22513) );
  OAI211_X1 U24130 ( .C1(n22526), .C2(n22702), .A(n22514), .B(n22513), .ZN(
        P1_U3101) );
  AOI22_X1 U24131 ( .A1(n22704), .A2(n22517), .B1(n22521), .B2(n22703), .ZN(
        n22516) );
  AOI22_X1 U24132 ( .A1(n22706), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22705), .B2(n22523), .ZN(n22515) );
  OAI211_X1 U24133 ( .C1(n22709), .C2(n22520), .A(n22516), .B(n22515), .ZN(
        P1_U3117) );
  AOI22_X1 U24134 ( .A1(n22521), .A2(n22716), .B1(n22717), .B2(n22517), .ZN(
        n22519) );
  AOI22_X1 U24135 ( .A1(n22719), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22718), .B2(n22523), .ZN(n22518) );
  OAI211_X1 U24136 ( .C1(n22723), .C2(n22520), .A(n22519), .B(n22518), .ZN(
        P1_U3133) );
  AOI22_X1 U24137 ( .A1(n22522), .A2(n22730), .B1(n22521), .B2(n22731), .ZN(
        n22525) );
  AOI22_X1 U24138 ( .A1(n22734), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n22733), .B2(n22523), .ZN(n22524) );
  OAI211_X1 U24139 ( .C1(n22526), .C2(n22747), .A(n22525), .B(n22524), .ZN(
        P1_U3149) );
  NAND2_X1 U24140 ( .A1(n22632), .A2(n22527), .ZN(n22559) );
  NOR2_X2 U24141 ( .A1(n22634), .A2(n22528), .ZN(n22567) );
  AOI22_X1 U24142 ( .A1(n22567), .A2(n22637), .B1(n22743), .B2(n22562), .ZN(
        n22534) );
  OAI22_X1 U24143 ( .A1(n22532), .A2(n22640), .B1(n22639), .B2(n22531), .ZN(
        n22568) );
  AOI22_X1 U24144 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22568), .ZN(n22533) );
  OAI211_X1 U24145 ( .C1(n22645), .C2(n22559), .A(n22534), .B(n22533), .ZN(
        P1_U3038) );
  INV_X1 U24146 ( .A(n22568), .ZN(n22565) );
  AOI22_X1 U24147 ( .A1(n22647), .A2(n22566), .B1(n22567), .B2(n22646), .ZN(
        n22536) );
  AOI22_X1 U24148 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22562), .ZN(n22535) );
  OAI211_X1 U24149 ( .C1(n22565), .C2(n22652), .A(n22536), .B(n22535), .ZN(
        P1_U3046) );
  AOI22_X1 U24150 ( .A1(n22654), .A2(n22562), .B1(n22567), .B2(n22653), .ZN(
        n22538) );
  AOI22_X1 U24151 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22655), .B1(
        n22660), .B2(n22568), .ZN(n22537) );
  OAI211_X1 U24152 ( .C1(n22658), .C2(n22559), .A(n22538), .B(n22537), .ZN(
        P1_U3054) );
  AOI22_X1 U24153 ( .A1(n22660), .A2(n22562), .B1(n22567), .B2(n22659), .ZN(
        n22540) );
  AOI22_X1 U24154 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22661), .B1(
        n22667), .B2(n22568), .ZN(n22539) );
  OAI211_X1 U24155 ( .C1(n22664), .C2(n22559), .A(n22540), .B(n22539), .ZN(
        P1_U3062) );
  AOI22_X1 U24156 ( .A1(n22567), .A2(n22666), .B1(n22665), .B2(n22566), .ZN(
        n22542) );
  AOI22_X1 U24157 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22562), .ZN(n22541) );
  OAI211_X1 U24158 ( .C1(n22565), .C2(n22671), .A(n22542), .B(n22541), .ZN(
        P1_U3070) );
  AOI22_X1 U24159 ( .A1(n22567), .A2(n22673), .B1(n22672), .B2(n22566), .ZN(
        n22544) );
  AOI22_X1 U24160 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22675), .B1(
        n22674), .B2(n22562), .ZN(n22543) );
  OAI211_X1 U24161 ( .C1(n22565), .C2(n22683), .A(n22544), .B(n22543), .ZN(
        P1_U3078) );
  AOI22_X1 U24162 ( .A1(n22583), .A2(n22562), .B1(n22567), .B2(n22678), .ZN(
        n22546) );
  AOI22_X1 U24163 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22680), .B1(
        n22566), .B2(n22679), .ZN(n22545) );
  OAI211_X1 U24164 ( .C1(n22565), .C2(n22593), .A(n22546), .B(n22545), .ZN(
        P1_U3086) );
  AOI22_X1 U24165 ( .A1(n22685), .A2(n22567), .B1(n22684), .B2(n22566), .ZN(
        n22548) );
  AOI22_X1 U24166 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22687), .B1(
        n22686), .B2(n22562), .ZN(n22547) );
  OAI211_X1 U24167 ( .C1(n22565), .C2(n22690), .A(n22548), .B(n22547), .ZN(
        P1_U3094) );
  AOI22_X1 U24168 ( .A1(n22692), .A2(n22566), .B1(n22567), .B2(n22691), .ZN(
        n22550) );
  AOI22_X1 U24169 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22562), .ZN(n22549) );
  OAI211_X1 U24170 ( .C1(n22565), .C2(n22702), .A(n22550), .B(n22549), .ZN(
        P1_U3102) );
  INV_X1 U24171 ( .A(n22562), .ZN(n22571) );
  AOI22_X1 U24172 ( .A1(n22567), .A2(n22698), .B1(n22697), .B2(n22566), .ZN(
        n22552) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22568), .ZN(n22551) );
  OAI211_X1 U24174 ( .C1(n22571), .C2(n22702), .A(n22552), .B(n22551), .ZN(
        P1_U3110) );
  AOI22_X1 U24175 ( .A1(n22705), .A2(n22562), .B1(n22567), .B2(n22703), .ZN(
        n22554) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22706), .B1(
        n22704), .B2(n22568), .ZN(n22553) );
  OAI211_X1 U24177 ( .C1(n22709), .C2(n22559), .A(n22554), .B(n22553), .ZN(
        P1_U3118) );
  AOI22_X1 U24178 ( .A1(n22567), .A2(n22711), .B1(n22710), .B2(n22566), .ZN(
        n22556) );
  AOI22_X1 U24179 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22568), .ZN(n22555) );
  OAI211_X1 U24180 ( .C1(n22571), .C2(n22715), .A(n22556), .B(n22555), .ZN(
        P1_U3126) );
  AOI22_X1 U24181 ( .A1(n22717), .A2(n22568), .B1(n22567), .B2(n22716), .ZN(
        n22558) );
  AOI22_X1 U24182 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22562), .ZN(n22557) );
  OAI211_X1 U24183 ( .C1(n22723), .C2(n22559), .A(n22558), .B(n22557), .ZN(
        P1_U3134) );
  AOI22_X1 U24184 ( .A1(n22567), .A2(n22725), .B1(n22724), .B2(n22566), .ZN(
        n22561) );
  AOI22_X1 U24185 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22568), .ZN(n22560) );
  OAI211_X1 U24186 ( .C1(n22571), .C2(n22729), .A(n22561), .B(n22560), .ZN(
        P1_U3142) );
  AOI22_X1 U24187 ( .A1(n22567), .A2(n22731), .B1(n22730), .B2(n22566), .ZN(
        n22564) );
  AOI22_X1 U24188 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22562), .ZN(n22563) );
  OAI211_X1 U24189 ( .C1(n22565), .C2(n22747), .A(n22564), .B(n22563), .ZN(
        P1_U3150) );
  AOI22_X1 U24190 ( .A1(n22741), .A2(n22567), .B1(n22739), .B2(n22566), .ZN(
        n22570) );
  AOI22_X1 U24191 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22568), .ZN(n22569) );
  OAI211_X1 U24192 ( .C1(n22571), .C2(n22747), .A(n22570), .B(n22569), .ZN(
        P1_U3158) );
  AOI22_X1 U24193 ( .A1(n22617), .A2(n22637), .B1(n22743), .B2(n22618), .ZN(
        n22573) );
  INV_X1 U24194 ( .A(n22621), .ZN(n22627) );
  AOI22_X1 U24195 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22627), .ZN(n22572) );
  OAI211_X1 U24196 ( .C1(n22645), .C2(n22623), .A(n22573), .B(n22572), .ZN(
        P1_U3039) );
  INV_X1 U24197 ( .A(n22623), .ZN(n22616) );
  AOI22_X1 U24198 ( .A1(n22617), .A2(n22646), .B1(n22647), .B2(n22616), .ZN(
        n22575) );
  AOI22_X1 U24199 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22618), .ZN(n22574) );
  OAI211_X1 U24200 ( .C1(n22621), .C2(n22652), .A(n22575), .B(n22574), .ZN(
        P1_U3047) );
  INV_X1 U24201 ( .A(n22659), .ZN(n22576) );
  OAI22_X1 U24202 ( .A1(n22621), .A2(n22577), .B1(n22625), .B2(n22576), .ZN(
        n22578) );
  INV_X1 U24203 ( .A(n22578), .ZN(n22580) );
  AOI22_X1 U24204 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22661), .B1(
        n22660), .B2(n22618), .ZN(n22579) );
  OAI211_X1 U24205 ( .C1(n22664), .C2(n22623), .A(n22580), .B(n22579), .ZN(
        P1_U3063) );
  AOI22_X1 U24206 ( .A1(n22617), .A2(n22666), .B1(n22616), .B2(n22665), .ZN(
        n22582) );
  AOI22_X1 U24207 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22618), .ZN(n22581) );
  OAI211_X1 U24208 ( .C1(n22621), .C2(n22671), .A(n22582), .B(n22581), .ZN(
        P1_U3071) );
  AOI22_X1 U24209 ( .A1(n22617), .A2(n22673), .B1(n22616), .B2(n22672), .ZN(
        n22585) );
  AOI22_X1 U24210 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22675), .B1(
        n22583), .B2(n22627), .ZN(n22584) );
  OAI211_X1 U24211 ( .C1(n22630), .C2(n22671), .A(n22585), .B(n22584), .ZN(
        P1_U3079) );
  AOI22_X1 U24212 ( .A1(n22617), .A2(n22678), .B1(n22686), .B2(n22627), .ZN(
        n22587) );
  AOI22_X1 U24213 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22680), .B1(
        n22616), .B2(n22679), .ZN(n22586) );
  OAI211_X1 U24214 ( .C1(n22630), .C2(n22683), .A(n22587), .B(n22586), .ZN(
        P1_U3087) );
  OAI22_X1 U24215 ( .A1(n22625), .A2(n22589), .B1(n22623), .B2(n22588), .ZN(
        n22590) );
  INV_X1 U24216 ( .A(n22590), .ZN(n22592) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22687), .B1(
        n22693), .B2(n22627), .ZN(n22591) );
  OAI211_X1 U24218 ( .C1(n22630), .C2(n22593), .A(n22592), .B(n22591), .ZN(
        P1_U3095) );
  AOI22_X1 U24219 ( .A1(n22617), .A2(n22691), .B1(n22692), .B2(n22616), .ZN(
        n22595) );
  AOI22_X1 U24220 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22618), .ZN(n22594) );
  OAI211_X1 U24221 ( .C1(n22621), .C2(n22702), .A(n22595), .B(n22594), .ZN(
        P1_U3103) );
  AOI22_X1 U24222 ( .A1(n22617), .A2(n22698), .B1(n22616), .B2(n22697), .ZN(
        n22597) );
  AOI22_X1 U24223 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22627), .ZN(n22596) );
  OAI211_X1 U24224 ( .C1(n22630), .C2(n22702), .A(n22597), .B(n22596), .ZN(
        P1_U3111) );
  OAI22_X1 U24225 ( .A1(n22715), .A2(n22621), .B1(n22598), .B2(n22625), .ZN(
        n22599) );
  INV_X1 U24226 ( .A(n22599), .ZN(n22601) );
  AOI22_X1 U24227 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22706), .B1(
        n22705), .B2(n22618), .ZN(n22600) );
  OAI211_X1 U24228 ( .C1(n22709), .C2(n22623), .A(n22601), .B(n22600), .ZN(
        P1_U3119) );
  OAI22_X1 U24229 ( .A1(n22625), .A2(n22603), .B1(n22623), .B2(n22602), .ZN(
        n22604) );
  INV_X1 U24230 ( .A(n22604), .ZN(n22606) );
  AOI22_X1 U24231 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22627), .ZN(n22605) );
  OAI211_X1 U24232 ( .C1(n22630), .C2(n22715), .A(n22606), .B(n22605), .ZN(
        P1_U3127) );
  OAI22_X1 U24233 ( .A1(n22625), .A2(n22607), .B1(n22729), .B2(n22621), .ZN(
        n22608) );
  INV_X1 U24234 ( .A(n22608), .ZN(n22610) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22618), .ZN(n22609) );
  OAI211_X1 U24236 ( .C1(n22723), .C2(n22623), .A(n22610), .B(n22609), .ZN(
        P1_U3135) );
  OAI22_X1 U24237 ( .A1(n22625), .A2(n22612), .B1(n22623), .B2(n22611), .ZN(
        n22613) );
  INV_X1 U24238 ( .A(n22613), .ZN(n22615) );
  AOI22_X1 U24239 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22627), .ZN(n22614) );
  OAI211_X1 U24240 ( .C1(n22630), .C2(n22729), .A(n22615), .B(n22614), .ZN(
        P1_U3143) );
  AOI22_X1 U24241 ( .A1(n22617), .A2(n22731), .B1(n22616), .B2(n22730), .ZN(
        n22620) );
  AOI22_X1 U24242 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22618), .ZN(n22619) );
  OAI211_X1 U24243 ( .C1(n22621), .C2(n22747), .A(n22620), .B(n22619), .ZN(
        P1_U3151) );
  OAI22_X1 U24244 ( .A1(n22625), .A2(n22624), .B1(n22623), .B2(n22622), .ZN(
        n22626) );
  INV_X1 U24245 ( .A(n22626), .ZN(n22629) );
  AOI22_X1 U24246 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22627), .ZN(n22628) );
  OAI211_X1 U24247 ( .C1(n22630), .C2(n22747), .A(n22629), .B(n22628), .ZN(
        P1_U3159) );
  NAND2_X1 U24248 ( .A1(n22632), .A2(n22631), .ZN(n22722) );
  NOR2_X2 U24249 ( .A1(n22634), .A2(n22633), .ZN(n22740) );
  AOI22_X1 U24250 ( .A1(DATAI_31_), .A2(n22636), .B1(n22635), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n22748) );
  INV_X1 U24251 ( .A(n22748), .ZN(n22732) );
  AOI22_X1 U24252 ( .A1(n22740), .A2(n22637), .B1(n22743), .B2(n22732), .ZN(
        n22644) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22642), .B1(
        n22648), .B2(n22742), .ZN(n22643) );
  OAI211_X1 U24254 ( .C1(n22645), .C2(n22722), .A(n22644), .B(n22643), .ZN(
        P1_U3040) );
  INV_X1 U24255 ( .A(n22742), .ZN(n22737) );
  AOI22_X1 U24256 ( .A1(n22647), .A2(n22738), .B1(n22740), .B2(n22646), .ZN(
        n22651) );
  AOI22_X1 U24257 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22649), .B1(
        n22648), .B2(n22732), .ZN(n22650) );
  OAI211_X1 U24258 ( .C1(n22737), .C2(n22652), .A(n22651), .B(n22650), .ZN(
        P1_U3048) );
  AOI22_X1 U24259 ( .A1(n22654), .A2(n22732), .B1(n22740), .B2(n22653), .ZN(
        n22657) );
  AOI22_X1 U24260 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22655), .B1(
        n22660), .B2(n22742), .ZN(n22656) );
  OAI211_X1 U24261 ( .C1(n22658), .C2(n22722), .A(n22657), .B(n22656), .ZN(
        P1_U3056) );
  AOI22_X1 U24262 ( .A1(n22660), .A2(n22732), .B1(n22740), .B2(n22659), .ZN(
        n22663) );
  AOI22_X1 U24263 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22661), .B1(
        n22667), .B2(n22742), .ZN(n22662) );
  OAI211_X1 U24264 ( .C1(n22664), .C2(n22722), .A(n22663), .B(n22662), .ZN(
        P1_U3064) );
  AOI22_X1 U24265 ( .A1(n22740), .A2(n22666), .B1(n22665), .B2(n22738), .ZN(
        n22670) );
  AOI22_X1 U24266 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22668), .B1(
        n22667), .B2(n22732), .ZN(n22669) );
  OAI211_X1 U24267 ( .C1(n22737), .C2(n22671), .A(n22670), .B(n22669), .ZN(
        P1_U3072) );
  AOI22_X1 U24268 ( .A1(n22740), .A2(n22673), .B1(n22672), .B2(n22738), .ZN(
        n22677) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22675), .B1(
        n22674), .B2(n22732), .ZN(n22676) );
  OAI211_X1 U24270 ( .C1(n22737), .C2(n22683), .A(n22677), .B(n22676), .ZN(
        P1_U3080) );
  AOI22_X1 U24271 ( .A1(n22686), .A2(n22742), .B1(n22740), .B2(n22678), .ZN(
        n22682) );
  AOI22_X1 U24272 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22680), .B1(
        n22738), .B2(n22679), .ZN(n22681) );
  OAI211_X1 U24273 ( .C1(n22748), .C2(n22683), .A(n22682), .B(n22681), .ZN(
        P1_U3088) );
  AOI22_X1 U24274 ( .A1(n22685), .A2(n22740), .B1(n22684), .B2(n22738), .ZN(
        n22689) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22687), .B1(
        n22686), .B2(n22732), .ZN(n22688) );
  OAI211_X1 U24276 ( .C1(n22737), .C2(n22690), .A(n22689), .B(n22688), .ZN(
        P1_U3096) );
  AOI22_X1 U24277 ( .A1(n22692), .A2(n22738), .B1(n22740), .B2(n22691), .ZN(
        n22696) );
  AOI22_X1 U24278 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22694), .B1(
        n22693), .B2(n22732), .ZN(n22695) );
  OAI211_X1 U24279 ( .C1(n22737), .C2(n22702), .A(n22696), .B(n22695), .ZN(
        P1_U3104) );
  AOI22_X1 U24280 ( .A1(n22740), .A2(n22698), .B1(n22697), .B2(n22738), .ZN(
        n22701) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22699), .B1(
        n22705), .B2(n22742), .ZN(n22700) );
  OAI211_X1 U24282 ( .C1(n22748), .C2(n22702), .A(n22701), .B(n22700), .ZN(
        P1_U3112) );
  AOI22_X1 U24283 ( .A1(n22704), .A2(n22742), .B1(n22740), .B2(n22703), .ZN(
        n22708) );
  AOI22_X1 U24284 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22706), .B1(
        n22705), .B2(n22732), .ZN(n22707) );
  OAI211_X1 U24285 ( .C1(n22709), .C2(n22722), .A(n22708), .B(n22707), .ZN(
        P1_U3120) );
  AOI22_X1 U24286 ( .A1(n22740), .A2(n22711), .B1(n22710), .B2(n22738), .ZN(
        n22714) );
  AOI22_X1 U24287 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22712), .B1(
        n22718), .B2(n22742), .ZN(n22713) );
  OAI211_X1 U24288 ( .C1(n22748), .C2(n22715), .A(n22714), .B(n22713), .ZN(
        P1_U3128) );
  AOI22_X1 U24289 ( .A1(n22717), .A2(n22742), .B1(n22740), .B2(n22716), .ZN(
        n22721) );
  AOI22_X1 U24290 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22719), .B1(
        n22718), .B2(n22732), .ZN(n22720) );
  OAI211_X1 U24291 ( .C1(n22723), .C2(n22722), .A(n22721), .B(n22720), .ZN(
        P1_U3136) );
  AOI22_X1 U24292 ( .A1(n22740), .A2(n22725), .B1(n22724), .B2(n22738), .ZN(
        n22728) );
  AOI22_X1 U24293 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22726), .B1(
        n22733), .B2(n22742), .ZN(n22727) );
  OAI211_X1 U24294 ( .C1(n22748), .C2(n22729), .A(n22728), .B(n22727), .ZN(
        P1_U3144) );
  AOI22_X1 U24295 ( .A1(n22740), .A2(n22731), .B1(n22730), .B2(n22738), .ZN(
        n22736) );
  AOI22_X1 U24296 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22734), .B1(
        n22733), .B2(n22732), .ZN(n22735) );
  OAI211_X1 U24297 ( .C1(n22737), .C2(n22747), .A(n22736), .B(n22735), .ZN(
        P1_U3152) );
  AOI22_X1 U24298 ( .A1(n22741), .A2(n22740), .B1(n22739), .B2(n22738), .ZN(
        n22746) );
  AOI22_X1 U24299 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22744), .B1(
        n22743), .B2(n22742), .ZN(n22745) );
  OAI211_X1 U24300 ( .C1(n22748), .C2(n22747), .A(n22746), .B(n22745), .ZN(
        P1_U3160) );
  INV_X1 U24301 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22751) );
  AOI22_X1 U24302 ( .A1(n20459), .A2(n22751), .B1(n22750), .B2(n22749), .ZN(
        P1_U3486) );
  AND2_X1 U11520 ( .A1(n12248), .A2(n12247), .ZN(n16849) );
  NOR2_X1 U14008 ( .A1(n12494), .A2(n12500), .ZN(n12531) );
  NOR2_X1 U12901 ( .A1(n12494), .A2(n12501), .ZN(n12545) );
  AND2_X1 U11366 ( .A1(n13796), .A2(n11317), .ZN(n15098) );
  CLKBUF_X1 U11266 ( .A(n13422), .Z(n13709) );
  CLKBUF_X1 U11276 ( .A(n11376), .Z(n11157) );
  AND2_X1 U11299 ( .A1(n13938), .A2(n14785), .ZN(n12096) );
  OR2_X1 U11315 ( .A1(n12902), .A2(n12901), .ZN(n12977) );
  CLKBUF_X1 U11316 ( .A(n11913), .Z(n12045) );
  CLKBUF_X1 U11318 ( .A(n11937), .Z(n11865) );
  CLKBUF_X1 U11331 ( .A(n12548), .Z(n19678) );
  NOR2_X1 U11353 ( .A1(n12494), .A2(n12497), .ZN(n12546) );
  CLKBUF_X1 U11354 ( .A(n11355), .Z(n16004) );
  CLKBUF_X3 U11371 ( .A(n17593), .Z(n17971) );
  CLKBUF_X2 U11392 ( .A(n15881), .Z(n11159) );
  CLKBUF_X1 U11537 ( .A(n11707), .Z(n11164) );
  CLKBUF_X2 U11543 ( .A(n11707), .Z(n11165) );
  CLKBUF_X1 U12176 ( .A(n17529), .Z(n17541) );
  INV_X1 U12292 ( .A(n20183), .ZN(n20210) );
  INV_X2 U12442 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14483) );
  NOR2_X1 U12471 ( .A1(n20183), .A2(n21698), .ZN(n20199) );
  NAND2_X1 U12719 ( .A1(n20932), .A2(n20770), .ZN(n11403) );
endmodule

